module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35074 , n35075 , n35076 , n35077 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 ;
  assign n2152 = x444 ^ x92 ;
  assign n2153 = n2152 ^ x284 ;
  assign n2154 = n2153 ^ x28 ;
  assign n2221 = n2154 ^ x187 ;
  assign n2222 = n2221 ^ x379 ;
  assign n2223 = n2222 ^ x123 ;
  assign n2302 = n2223 ^ x282 ;
  assign n2303 = n2302 ^ x474 ;
  assign n2304 = n2303 ^ x218 ;
  assign n2383 = n2304 ^ x377 ;
  assign n2272 = x474 ^ x122 ;
  assign n2273 = n2272 ^ x314 ;
  assign n2274 = n2273 ^ x58 ;
  assign n2384 = n2383 ^ n2274 ;
  assign n2385 = n2384 ^ x313 ;
  assign n20766 = n2385 ^ x472 ;
  assign n2351 = n2274 ^ x217 ;
  assign n2352 = n2351 ^ x409 ;
  assign n2353 = n2352 ^ x153 ;
  assign n20767 = n20766 ^ n2353 ;
  assign n20768 = n20767 ^ x408 ;
  assign n13647 = x472 ^ x120 ;
  assign n13648 = n13647 ^ x312 ;
  assign n13649 = n13648 ^ x56 ;
  assign n22371 = n20768 ^ n13649 ;
  assign n2434 = n2353 ^ x312 ;
  assign n2435 = n2434 ^ x504 ;
  assign n2436 = n2435 ^ x248 ;
  assign n22372 = n22371 ^ n2436 ;
  assign n22373 = n22372 ^ x503 ;
  assign n15591 = n13649 ^ x215 ;
  assign n15592 = n15591 ^ x407 ;
  assign n15593 = n15592 ^ x151 ;
  assign n24542 = n22373 ^ n15593 ;
  assign n19524 = n2436 ^ x407 ;
  assign n2904 = x504 ^ x152 ;
  assign n2905 = n2904 ^ x344 ;
  assign n2906 = n2905 ^ x88 ;
  assign n19525 = n19524 ^ n2906 ;
  assign n19526 = n19525 ^ x343 ;
  assign n24543 = n24542 ^ n19526 ;
  assign n1478 = x503 ^ x151 ;
  assign n1479 = n1478 ^ x343 ;
  assign n1480 = n1479 ^ x87 ;
  assign n24544 = n24543 ^ n1480 ;
  assign n17478 = n15593 ^ x310 ;
  assign n17479 = n17478 ^ x502 ;
  assign n17480 = n17479 ^ x246 ;
  assign n26515 = n24544 ^ n17480 ;
  assign n21157 = n19526 ^ x502 ;
  assign n2907 = n2906 ^ x247 ;
  assign n2908 = n2907 ^ x439 ;
  assign n2909 = n2908 ^ x183 ;
  assign n21158 = n21157 ^ n2909 ;
  assign n21159 = n21158 ^ x438 ;
  assign n26516 = n26515 ^ n21159 ;
  assign n1490 = n1480 ^ x246 ;
  assign n1491 = n1490 ^ x438 ;
  assign n1492 = n1491 ^ x182 ;
  assign n26517 = n26516 ^ n1492 ;
  assign n19480 = n17480 ^ x405 ;
  assign n1484 = x502 ^ x150 ;
  assign n1485 = n1484 ^ x342 ;
  assign n1486 = n1485 ^ x86 ;
  assign n19481 = n19480 ^ n1486 ;
  assign n19482 = n19481 ^ x341 ;
  assign n28627 = n26517 ^ n19482 ;
  assign n23070 = n21159 ^ n1486 ;
  assign n2922 = n2909 ^ x342 ;
  assign n513 = x439 ^ x87 ;
  assign n514 = n513 ^ x279 ;
  assign n515 = n514 ^ x23 ;
  assign n2923 = n2922 ^ n515 ;
  assign n2924 = n2923 ^ x278 ;
  assign n23071 = n23070 ^ n2924 ;
  assign n1503 = x438 ^ x86 ;
  assign n1504 = n1503 ^ x278 ;
  assign n1505 = n1504 ^ x22 ;
  assign n23072 = n23071 ^ n1505 ;
  assign n28628 = n28627 ^ n23072 ;
  assign n1502 = n1492 ^ x341 ;
  assign n1506 = n1505 ^ n1502 ;
  assign n1507 = n1506 ^ x277 ;
  assign n28629 = n28628 ^ n1507 ;
  assign n2289 = x442 ^ x90 ;
  assign n2290 = n2289 ^ x282 ;
  assign n2291 = n2290 ^ x26 ;
  assign n2370 = n2291 ^ x185 ;
  assign n2371 = n2370 ^ x377 ;
  assign n2372 = n2371 ^ x121 ;
  assign n16709 = n2372 ^ x280 ;
  assign n16710 = n16709 ^ x472 ;
  assign n16711 = n16710 ^ x216 ;
  assign n18809 = n16711 ^ x375 ;
  assign n18810 = n18809 ^ n13649 ;
  assign n18811 = n18810 ^ x311 ;
  assign n20758 = n18811 ^ x470 ;
  assign n20759 = n20758 ^ n15593 ;
  assign n20760 = n20759 ^ x406 ;
  assign n543 = x470 ^ x118 ;
  assign n544 = n543 ^ x310 ;
  assign n545 = n544 ^ x54 ;
  assign n22774 = n20760 ^ n545 ;
  assign n22775 = n22774 ^ n17480 ;
  assign n22776 = n22775 ^ x501 ;
  assign n546 = n545 ^ x213 ;
  assign n547 = n546 ^ x405 ;
  assign n548 = n547 ^ x149 ;
  assign n24535 = n22776 ^ n548 ;
  assign n24536 = n24535 ^ n19482 ;
  assign n611 = x501 ^ x149 ;
  assign n612 = n611 ^ x341 ;
  assign n613 = n612 ^ x85 ;
  assign n24537 = n24536 ^ n613 ;
  assign n34561 = n28629 ^ n24537 ;
  assign n2028 = x509 ^ x157 ;
  assign n2029 = n2028 ^ x349 ;
  assign n2030 = n2029 ^ x93 ;
  assign n2088 = n2030 ^ x252 ;
  assign n2089 = n2088 ^ x444 ;
  assign n2090 = n2089 ^ x188 ;
  assign n2157 = n2090 ^ x347 ;
  assign n2158 = n2157 ^ n2154 ;
  assign n2159 = n2158 ^ x283 ;
  assign n2226 = n2159 ^ x442 ;
  assign n2227 = n2226 ^ n2223 ;
  assign n2228 = n2227 ^ x378 ;
  assign n2307 = n2291 ^ n2228 ;
  assign n2308 = n2307 ^ n2304 ;
  assign n2309 = n2308 ^ x473 ;
  assign n2388 = n2372 ^ n2309 ;
  assign n2389 = n2388 ^ n2385 ;
  assign n1449 = x473 ^ x121 ;
  assign n1450 = n1449 ^ x313 ;
  assign n1451 = n1450 ^ x57 ;
  assign n2390 = n2389 ^ n1451 ;
  assign n25830 = n16711 ^ n2390 ;
  assign n25831 = n25830 ^ n20768 ;
  assign n1452 = n1451 ^ x216 ;
  assign n1453 = n1452 ^ x408 ;
  assign n1454 = n1453 ^ x152 ;
  assign n25832 = n25831 ^ n1454 ;
  assign n27801 = n25832 ^ n18811 ;
  assign n27802 = n27801 ^ n22373 ;
  assign n1471 = n1454 ^ x311 ;
  assign n1472 = n1471 ^ x503 ;
  assign n1473 = n1472 ^ x247 ;
  assign n27803 = n27802 ^ n1473 ;
  assign n1477 = n1473 ^ x406 ;
  assign n1481 = n1480 ^ n1477 ;
  assign n1482 = n1481 ^ x342 ;
  assign n29778 = n27803 ^ n1482 ;
  assign n29779 = n29778 ^ n24544 ;
  assign n29780 = n29779 ^ n20760 ;
  assign n32006 = n29780 ^ n22776 ;
  assign n32007 = n32006 ^ n26517 ;
  assign n1489 = n1482 ^ x501 ;
  assign n1493 = n1492 ^ n1489 ;
  assign n1494 = n1493 ^ x437 ;
  assign n32008 = n32007 ^ n1494 ;
  assign n34562 = n34561 ^ n32008 ;
  assign n1509 = x437 ^ x85 ;
  assign n1510 = n1509 ^ x277 ;
  assign n1511 = n1510 ^ x21 ;
  assign n1501 = n1494 ^ n613 ;
  assign n1508 = n1507 ^ n1501 ;
  assign n1512 = n1511 ^ n1508 ;
  assign n34563 = n34562 ^ n1512 ;
  assign n549 = n548 ^ x308 ;
  assign n550 = n549 ^ x500 ;
  assign n551 = n550 ^ x244 ;
  assign n26523 = n24537 ^ n551 ;
  assign n21150 = n19482 ^ x500 ;
  assign n1496 = n1486 ^ x245 ;
  assign n1497 = n1496 ^ x437 ;
  assign n1498 = n1497 ^ x181 ;
  assign n21151 = n21150 ^ n1498 ;
  assign n21152 = n21151 ^ x436 ;
  assign n26524 = n26523 ^ n21152 ;
  assign n624 = n613 ^ x244 ;
  assign n625 = n624 ^ x436 ;
  assign n626 = n625 ^ x180 ;
  assign n26525 = n26524 ^ n626 ;
  assign n37087 = n34563 ^ n26525 ;
  assign n30668 = n28629 ^ n21152 ;
  assign n25049 = n23072 ^ n1498 ;
  assign n2931 = n2924 ^ x437 ;
  assign n516 = n515 ^ x182 ;
  assign n517 = n516 ^ x374 ;
  assign n518 = n517 ^ x118 ;
  assign n2932 = n2931 ^ n518 ;
  assign n2933 = n2932 ^ x373 ;
  assign n25050 = n25049 ^ n2933 ;
  assign n1521 = n1505 ^ x181 ;
  assign n1522 = n1521 ^ x373 ;
  assign n1523 = n1522 ^ x117 ;
  assign n25051 = n25050 ^ n1523 ;
  assign n30669 = n30668 ^ n25051 ;
  assign n1520 = n1507 ^ x436 ;
  assign n1524 = n1523 ^ n1520 ;
  assign n1525 = n1524 ^ x372 ;
  assign n30670 = n30669 ^ n1525 ;
  assign n37088 = n37087 ^ n30670 ;
  assign n1527 = n1511 ^ x180 ;
  assign n1528 = n1527 ^ x372 ;
  assign n1529 = n1528 ^ x116 ;
  assign n1519 = n1512 ^ n626 ;
  assign n1526 = n1525 ^ n1519 ;
  assign n1530 = n1529 ^ n1526 ;
  assign n37089 = n37088 ^ n1530 ;
  assign n553 = x500 ^ x148 ;
  assign n554 = n553 ^ x340 ;
  assign n555 = n554 ^ x84 ;
  assign n552 = n551 ^ x403 ;
  assign n556 = n555 ^ n552 ;
  assign n557 = n556 ^ x339 ;
  assign n28620 = n26525 ^ n557 ;
  assign n23151 = n21152 ^ n555 ;
  assign n1514 = n1498 ^ x340 ;
  assign n1515 = n1514 ^ n1511 ;
  assign n1516 = n1515 ^ x276 ;
  assign n23152 = n23151 ^ n1516 ;
  assign n658 = x436 ^ x84 ;
  assign n659 = n658 ^ x276 ;
  assign n660 = n659 ^ x20 ;
  assign n23153 = n23152 ^ n660 ;
  assign n28621 = n28620 ^ n23153 ;
  assign n657 = n626 ^ x339 ;
  assign n661 = n660 ^ n657 ;
  assign n662 = n661 ^ x275 ;
  assign n28622 = n28621 ^ n662 ;
  assign n39232 = n37089 ^ n28622 ;
  assign n33085 = n30670 ^ n23153 ;
  assign n27193 = n25051 ^ n1516 ;
  assign n2940 = n2933 ^ n1511 ;
  assign n519 = n518 ^ x277 ;
  assign n520 = n519 ^ x469 ;
  assign n521 = n520 ^ x213 ;
  assign n2941 = n2940 ^ n521 ;
  assign n2942 = n2941 ^ x468 ;
  assign n27194 = n27193 ^ n2942 ;
  assign n1539 = n1523 ^ x276 ;
  assign n1540 = n1539 ^ x468 ;
  assign n1541 = n1540 ^ x212 ;
  assign n27195 = n27194 ^ n1541 ;
  assign n33086 = n33085 ^ n27195 ;
  assign n1538 = n1525 ^ n660 ;
  assign n1542 = n1541 ^ n1538 ;
  assign n1543 = n1542 ^ x467 ;
  assign n33087 = n33086 ^ n1543 ;
  assign n39233 = n39232 ^ n33087 ;
  assign n1545 = n1529 ^ x275 ;
  assign n1546 = n1545 ^ x467 ;
  assign n1547 = n1546 ^ x211 ;
  assign n1537 = n1530 ^ n662 ;
  assign n1544 = n1543 ^ n1537 ;
  assign n1548 = n1547 ^ n1544 ;
  assign n39234 = n39233 ^ n1548 ;
  assign n635 = n557 ^ x498 ;
  assign n630 = n555 ^ x243 ;
  assign n631 = n630 ^ x435 ;
  assign n632 = n631 ^ x179 ;
  assign n636 = n635 ^ n632 ;
  assign n637 = n636 ^ x434 ;
  assign n30662 = n28622 ^ n637 ;
  assign n24971 = n23153 ^ n632 ;
  assign n1532 = n1516 ^ x435 ;
  assign n1533 = n1532 ^ n1529 ;
  assign n1534 = n1533 ^ x371 ;
  assign n24972 = n24971 ^ n1534 ;
  assign n700 = n660 ^ x179 ;
  assign n701 = n700 ^ x371 ;
  assign n702 = n701 ^ x115 ;
  assign n24973 = n24972 ^ n702 ;
  assign n30663 = n30662 ^ n24973 ;
  assign n699 = n662 ^ x434 ;
  assign n703 = n702 ^ n699 ;
  assign n704 = n703 ^ x370 ;
  assign n30664 = n30663 ^ n704 ;
  assign n41660 = n39234 ^ n30664 ;
  assign n35561 = n33087 ^ n24973 ;
  assign n29409 = n27195 ^ n1534 ;
  assign n2949 = n2942 ^ n1529 ;
  assign n523 = x469 ^ x117 ;
  assign n524 = n523 ^ x309 ;
  assign n525 = n524 ^ x53 ;
  assign n522 = n521 ^ x372 ;
  assign n526 = n525 ^ n522 ;
  assign n527 = n526 ^ x308 ;
  assign n2950 = n2949 ^ n527 ;
  assign n1563 = x468 ^ x116 ;
  assign n1564 = n1563 ^ x308 ;
  assign n1565 = n1564 ^ x52 ;
  assign n2951 = n2950 ^ n1565 ;
  assign n29410 = n29409 ^ n2951 ;
  assign n1562 = n1541 ^ x371 ;
  assign n1566 = n1565 ^ n1562 ;
  assign n1567 = n1566 ^ x307 ;
  assign n29411 = n29410 ^ n1567 ;
  assign n35562 = n35561 ^ n29411 ;
  assign n1568 = n1567 ^ n702 ;
  assign n1569 = n1568 ^ n1543 ;
  assign n534 = x467 ^ x115 ;
  assign n535 = n534 ^ x307 ;
  assign n536 = n535 ^ x51 ;
  assign n1570 = n1569 ^ n536 ;
  assign n35563 = n35562 ^ n1570 ;
  assign n41661 = n41660 ^ n35563 ;
  assign n1561 = n1548 ^ n704 ;
  assign n1571 = n1570 ^ n1561 ;
  assign n1555 = n1547 ^ x370 ;
  assign n1556 = n1555 ^ n536 ;
  assign n1557 = n1556 ^ x306 ;
  assign n1572 = n1571 ^ n1557 ;
  assign n41662 = n41661 ^ n1572 ;
  assign n676 = x434 ^ x82 ;
  assign n677 = n676 ^ x274 ;
  assign n678 = n677 ^ x18 ;
  assign n650 = x498 ^ x146 ;
  assign n651 = n650 ^ x338 ;
  assign n652 = n651 ^ x82 ;
  assign n674 = n652 ^ n637 ;
  assign n669 = n632 ^ x338 ;
  assign n664 = x435 ^ x83 ;
  assign n665 = n664 ^ x275 ;
  assign n666 = n665 ^ x19 ;
  assign n670 = n669 ^ n666 ;
  assign n671 = n670 ^ x274 ;
  assign n675 = n674 ^ n671 ;
  assign n679 = n678 ^ n675 ;
  assign n33053 = n30664 ^ n679 ;
  assign n27186 = n24973 ^ n671 ;
  assign n1550 = n1547 ^ n666 ;
  assign n1551 = n1550 ^ n1534 ;
  assign n1552 = n1551 ^ x466 ;
  assign n27187 = n27186 ^ n1552 ;
  assign n748 = n702 ^ x274 ;
  assign n749 = n748 ^ x466 ;
  assign n750 = n749 ^ x210 ;
  assign n27188 = n27187 ^ n750 ;
  assign n33054 = n33053 ^ n27188 ;
  assign n747 = n704 ^ n678 ;
  assign n751 = n750 ^ n747 ;
  assign n752 = n751 ^ x465 ;
  assign n33055 = n33054 ^ n752 ;
  assign n43771 = n41662 ^ n33055 ;
  assign n37641 = n35563 ^ n27188 ;
  assign n31382 = n29411 ^ n1552 ;
  assign n2958 = n2951 ^ n1547 ;
  assign n529 = n525 ^ x212 ;
  assign n530 = n529 ^ x404 ;
  assign n531 = n530 ^ x148 ;
  assign n528 = n527 ^ x467 ;
  assign n532 = n531 ^ n528 ;
  assign n533 = n532 ^ x403 ;
  assign n2959 = n2958 ^ n533 ;
  assign n1579 = n1565 ^ x211 ;
  assign n1580 = n1579 ^ x403 ;
  assign n1581 = n1580 ^ x147 ;
  assign n2960 = n2959 ^ n1581 ;
  assign n31383 = n31382 ^ n2960 ;
  assign n1578 = n1567 ^ x466 ;
  assign n1582 = n1581 ^ n1578 ;
  assign n1583 = n1582 ^ x402 ;
  assign n31384 = n31383 ^ n1583 ;
  assign n37642 = n37641 ^ n31384 ;
  assign n1577 = n1570 ^ n750 ;
  assign n1584 = n1583 ^ n1577 ;
  assign n639 = n536 ^ x210 ;
  assign n640 = n639 ^ x402 ;
  assign n641 = n640 ^ x146 ;
  assign n1585 = n1584 ^ n641 ;
  assign n37643 = n37642 ^ n1585 ;
  assign n43772 = n43771 ^ n37643 ;
  assign n1587 = n1557 ^ x465 ;
  assign n1588 = n1587 ^ n641 ;
  assign n1589 = n1588 ^ x401 ;
  assign n1576 = n1572 ^ n752 ;
  assign n1586 = n1585 ^ n1576 ;
  assign n1590 = n1589 ^ n1586 ;
  assign n43773 = n43772 ^ n1590 ;
  assign n718 = n678 ^ x177 ;
  assign n719 = n718 ^ x369 ;
  assign n720 = n719 ^ x113 ;
  assign n692 = n652 ^ x241 ;
  assign n693 = n692 ^ x433 ;
  assign n694 = n693 ^ x177 ;
  assign n716 = n694 ^ n679 ;
  assign n711 = n671 ^ x433 ;
  assign n706 = n666 ^ x178 ;
  assign n707 = n706 ^ x370 ;
  assign n708 = n707 ^ x114 ;
  assign n712 = n711 ^ n708 ;
  assign n713 = n712 ^ x369 ;
  assign n717 = n716 ^ n713 ;
  assign n721 = n720 ^ n717 ;
  assign n35549 = n33055 ^ n721 ;
  assign n29401 = n27188 ^ n713 ;
  assign n1554 = n1552 ^ n708 ;
  assign n1558 = n1557 ^ n1554 ;
  assign n797 = x466 ^ x114 ;
  assign n798 = n797 ^ x306 ;
  assign n799 = n798 ^ x50 ;
  assign n1559 = n1558 ^ n799 ;
  assign n29402 = n29401 ^ n1559 ;
  assign n796 = n750 ^ x369 ;
  assign n800 = n799 ^ n796 ;
  assign n801 = n800 ^ x305 ;
  assign n29403 = n29402 ^ n801 ;
  assign n35550 = n35549 ^ n29403 ;
  assign n803 = x465 ^ x113 ;
  assign n804 = n803 ^ x305 ;
  assign n805 = n804 ^ x49 ;
  assign n795 = n752 ^ n720 ;
  assign n802 = n801 ^ n795 ;
  assign n806 = n805 ^ n802 ;
  assign n35551 = n35550 ^ n806 ;
  assign n45764 = n43773 ^ n35551 ;
  assign n40098 = n37643 ^ n29403 ;
  assign n33878 = n31384 ^ n1559 ;
  assign n2967 = n2960 ^ n1557 ;
  assign n538 = n531 ^ x307 ;
  assign n539 = n538 ^ x499 ;
  assign n540 = n539 ^ x243 ;
  assign n537 = n536 ^ n533 ;
  assign n541 = n540 ^ n537 ;
  assign n542 = n541 ^ x498 ;
  assign n2968 = n2967 ^ n542 ;
  assign n1600 = n1581 ^ x306 ;
  assign n1601 = n1600 ^ x498 ;
  assign n1602 = n1601 ^ x242 ;
  assign n2969 = n2968 ^ n1602 ;
  assign n33879 = n33878 ^ n2969 ;
  assign n1599 = n1583 ^ n799 ;
  assign n1603 = n1602 ^ n1599 ;
  assign n1604 = n1603 ^ x497 ;
  assign n33880 = n33879 ^ n1604 ;
  assign n40099 = n40098 ^ n33880 ;
  assign n1598 = n1585 ^ n801 ;
  assign n1605 = n1604 ^ n1598 ;
  assign n681 = n641 ^ x305 ;
  assign n682 = n681 ^ x497 ;
  assign n683 = n682 ^ x241 ;
  assign n1606 = n1605 ^ n683 ;
  assign n40100 = n40099 ^ n1606 ;
  assign n45765 = n45764 ^ n40100 ;
  assign n1608 = n1589 ^ n805 ;
  assign n1609 = n1608 ^ n683 ;
  assign n1610 = n1609 ^ x496 ;
  assign n1597 = n1590 ^ n806 ;
  assign n1607 = n1606 ^ n1597 ;
  assign n1611 = n1610 ^ n1607 ;
  assign n45766 = n45765 ^ n1611 ;
  assign n766 = n720 ^ x272 ;
  assign n767 = n766 ^ x464 ;
  assign n768 = n767 ^ x208 ;
  assign n740 = n694 ^ x336 ;
  assign n735 = x433 ^ x81 ;
  assign n736 = n735 ^ x273 ;
  assign n737 = n736 ^ x17 ;
  assign n741 = n740 ^ n737 ;
  assign n742 = n741 ^ x272 ;
  assign n764 = n742 ^ n721 ;
  assign n759 = n737 ^ n713 ;
  assign n754 = n708 ^ x273 ;
  assign n755 = n754 ^ x465 ;
  assign n756 = n755 ^ x209 ;
  assign n760 = n759 ^ n756 ;
  assign n761 = n760 ^ x464 ;
  assign n765 = n764 ^ n761 ;
  assign n769 = n768 ^ n765 ;
  assign n37765 = n35551 ^ n769 ;
  assign n31354 = n29403 ^ n761 ;
  assign n1592 = n1559 ^ n756 ;
  assign n1593 = n1592 ^ n1589 ;
  assign n863 = n799 ^ x209 ;
  assign n864 = n863 ^ x401 ;
  assign n865 = n864 ^ x145 ;
  assign n1594 = n1593 ^ n865 ;
  assign n31355 = n31354 ^ n1594 ;
  assign n862 = n801 ^ x464 ;
  assign n866 = n865 ^ n862 ;
  assign n867 = n866 ^ x400 ;
  assign n31356 = n31355 ^ n867 ;
  assign n37766 = n37765 ^ n31356 ;
  assign n869 = n805 ^ x208 ;
  assign n870 = n869 ^ x400 ;
  assign n871 = n870 ^ x144 ;
  assign n861 = n806 ^ n768 ;
  assign n868 = n867 ^ n861 ;
  assign n872 = n871 ^ n868 ;
  assign n37767 = n37766 ^ n872 ;
  assign n48026 = n45766 ^ n37767 ;
  assign n42481 = n40100 ^ n31356 ;
  assign n36320 = n33880 ^ n1594 ;
  assign n2976 = n2969 ^ n1589 ;
  assign n644 = x499 ^ x147 ;
  assign n645 = n644 ^ x339 ;
  assign n646 = n645 ^ x83 ;
  assign n643 = n540 ^ x402 ;
  assign n647 = n646 ^ n643 ;
  assign n648 = n647 ^ x338 ;
  assign n642 = n641 ^ n542 ;
  assign n649 = n648 ^ n642 ;
  assign n653 = n652 ^ n649 ;
  assign n2977 = n2976 ^ n653 ;
  assign n1621 = n1602 ^ x401 ;
  assign n1622 = n1621 ^ n652 ;
  assign n1623 = n1622 ^ x337 ;
  assign n2978 = n2977 ^ n1623 ;
  assign n36321 = n36320 ^ n2978 ;
  assign n1620 = n1604 ^ n865 ;
  assign n1624 = n1623 ^ n1620 ;
  assign n723 = x497 ^ x145 ;
  assign n724 = n723 ^ x337 ;
  assign n725 = n724 ^ x81 ;
  assign n1625 = n1624 ^ n725 ;
  assign n36322 = n36321 ^ n1625 ;
  assign n42482 = n42481 ^ n36322 ;
  assign n1619 = n1606 ^ n867 ;
  assign n1626 = n1625 ^ n1619 ;
  assign n726 = n683 ^ x400 ;
  assign n727 = n726 ^ n725 ;
  assign n728 = n727 ^ x336 ;
  assign n1627 = n1626 ^ n728 ;
  assign n42483 = n42482 ^ n1627 ;
  assign n48027 = n48026 ^ n42483 ;
  assign n1629 = n1610 ^ n871 ;
  assign n1630 = n1629 ^ n728 ;
  assign n1011 = x496 ^ x144 ;
  assign n1012 = n1011 ^ x336 ;
  assign n1013 = n1012 ^ x80 ;
  assign n1631 = n1630 ^ n1013 ;
  assign n1618 = n1611 ^ n872 ;
  assign n1628 = n1627 ^ n1618 ;
  assign n1632 = n1631 ^ n1628 ;
  assign n48028 = n48027 ^ n1632 ;
  assign n823 = n768 ^ x367 ;
  assign n815 = x464 ^ x112 ;
  assign n816 = n815 ^ x304 ;
  assign n817 = n816 ^ x48 ;
  assign n824 = n823 ^ n817 ;
  assign n825 = n824 ^ x303 ;
  assign n788 = n742 ^ x431 ;
  assign n783 = n737 ^ x176 ;
  assign n784 = n783 ^ x368 ;
  assign n785 = n784 ^ x112 ;
  assign n789 = n788 ^ n785 ;
  assign n790 = n789 ^ x367 ;
  assign n821 = n790 ^ n769 ;
  assign n813 = n785 ^ n761 ;
  assign n808 = n756 ^ x368 ;
  assign n809 = n808 ^ n805 ;
  assign n810 = n809 ^ x304 ;
  assign n814 = n813 ^ n810 ;
  assign n818 = n817 ^ n814 ;
  assign n822 = n821 ^ n818 ;
  assign n826 = n825 ^ n822 ;
  assign n40091 = n37767 ^ n826 ;
  assign n33874 = n31356 ^ n818 ;
  assign n1613 = n1594 ^ n810 ;
  assign n1614 = n1613 ^ n1610 ;
  assign n935 = n865 ^ x304 ;
  assign n936 = n935 ^ x496 ;
  assign n937 = n936 ^ x240 ;
  assign n1615 = n1614 ^ n937 ;
  assign n33875 = n33874 ^ n1615 ;
  assign n934 = n867 ^ n817 ;
  assign n938 = n937 ^ n934 ;
  assign n939 = n938 ^ x495 ;
  assign n33876 = n33875 ^ n939 ;
  assign n40092 = n40091 ^ n33876 ;
  assign n941 = n871 ^ x303 ;
  assign n942 = n941 ^ x495 ;
  assign n943 = n942 ^ x239 ;
  assign n933 = n872 ^ n825 ;
  assign n940 = n939 ^ n933 ;
  assign n944 = n943 ^ n940 ;
  assign n40093 = n40092 ^ n944 ;
  assign n50096 = n48028 ^ n40093 ;
  assign n44448 = n42483 ^ n33876 ;
  assign n38564 = n36322 ^ n1615 ;
  assign n2985 = n2978 ^ n1610 ;
  assign n686 = n646 ^ x242 ;
  assign n687 = n686 ^ x434 ;
  assign n688 = n687 ^ x178 ;
  assign n685 = n648 ^ x497 ;
  assign n689 = n688 ^ n685 ;
  assign n690 = n689 ^ x433 ;
  assign n684 = n683 ^ n653 ;
  assign n691 = n690 ^ n684 ;
  assign n695 = n694 ^ n691 ;
  assign n2986 = n2985 ^ n695 ;
  assign n1642 = n1623 ^ x496 ;
  assign n1643 = n1642 ^ n694 ;
  assign n1644 = n1643 ^ x432 ;
  assign n2987 = n2986 ^ n1644 ;
  assign n38565 = n38564 ^ n2987 ;
  assign n1641 = n1625 ^ n937 ;
  assign n1645 = n1644 ^ n1641 ;
  assign n771 = n725 ^ x240 ;
  assign n772 = n771 ^ x432 ;
  assign n773 = n772 ^ x176 ;
  assign n1646 = n1645 ^ n773 ;
  assign n38566 = n38565 ^ n1646 ;
  assign n44449 = n44448 ^ n38566 ;
  assign n1640 = n1627 ^ n939 ;
  assign n1647 = n1646 ^ n1640 ;
  assign n774 = n728 ^ x495 ;
  assign n775 = n774 ^ n773 ;
  assign n776 = n775 ^ x431 ;
  assign n1648 = n1647 ^ n776 ;
  assign n44450 = n44449 ^ n1648 ;
  assign n50097 = n50096 ^ n44450 ;
  assign n1650 = n1631 ^ n943 ;
  assign n1651 = n1650 ^ n776 ;
  assign n1108 = n1013 ^ x239 ;
  assign n1109 = n1108 ^ x431 ;
  assign n1110 = n1109 ^ x175 ;
  assign n1652 = n1651 ^ n1110 ;
  assign n1639 = n1632 ^ n944 ;
  assign n1649 = n1648 ^ n1639 ;
  assign n1653 = n1652 ^ n1649 ;
  assign n50098 = n50097 ^ n1653 ;
  assign n2138 = x508 ^ x156 ;
  assign n2139 = n2138 ^ x348 ;
  assign n2140 = n2139 ^ x92 ;
  assign n2207 = n2140 ^ x251 ;
  assign n2208 = n2207 ^ x443 ;
  assign n2209 = n2208 ^ x187 ;
  assign n2284 = n2209 ^ x346 ;
  assign n1455 = x443 ^ x91 ;
  assign n1456 = n1455 ^ x283 ;
  assign n1457 = n1456 ^ x27 ;
  assign n2285 = n2284 ^ n1457 ;
  assign n2286 = n2285 ^ x282 ;
  assign n2366 = n2286 ^ x441 ;
  assign n1458 = n1457 ^ x186 ;
  assign n1459 = n1458 ^ x378 ;
  assign n1460 = n1459 ^ x122 ;
  assign n2367 = n2366 ^ n1460 ;
  assign n2368 = n2367 ^ x377 ;
  assign n564 = x441 ^ x89 ;
  assign n565 = n564 ^ x281 ;
  assign n566 = n565 ^ x25 ;
  assign n21783 = n2368 ^ n566 ;
  assign n1461 = n1460 ^ x281 ;
  assign n1462 = n1461 ^ x473 ;
  assign n1463 = n1462 ^ x217 ;
  assign n21784 = n21783 ^ n1463 ;
  assign n21785 = n21784 ^ x472 ;
  assign n567 = n566 ^ x184 ;
  assign n568 = n567 ^ x376 ;
  assign n569 = n568 ^ x120 ;
  assign n23882 = n21785 ^ n569 ;
  assign n1464 = n1463 ^ x376 ;
  assign n1465 = n1464 ^ n1451 ;
  assign n1466 = n1465 ^ x312 ;
  assign n23883 = n23882 ^ n1466 ;
  assign n23884 = n23883 ^ n13649 ;
  assign n570 = n569 ^ x279 ;
  assign n571 = n570 ^ x471 ;
  assign n572 = n571 ^ x215 ;
  assign n25825 = n23884 ^ n572 ;
  assign n1467 = n1466 ^ x471 ;
  assign n1468 = n1467 ^ n1454 ;
  assign n1469 = n1468 ^ x407 ;
  assign n25826 = n25825 ^ n1469 ;
  assign n25827 = n25826 ^ n15593 ;
  assign n573 = n572 ^ x374 ;
  assign n558 = x471 ^ x119 ;
  assign n559 = n558 ^ x311 ;
  assign n560 = n559 ^ x55 ;
  assign n574 = n573 ^ n560 ;
  assign n575 = n574 ^ x310 ;
  assign n27797 = n25827 ^ n575 ;
  assign n1470 = n1469 ^ n560 ;
  assign n1474 = n1473 ^ n1470 ;
  assign n1475 = n1474 ^ x502 ;
  assign n27798 = n27797 ^ n1475 ;
  assign n27799 = n27798 ^ n17480 ;
  assign n576 = n575 ^ x469 ;
  assign n561 = n560 ^ x214 ;
  assign n562 = n561 ^ x406 ;
  assign n563 = n562 ^ x150 ;
  assign n577 = n576 ^ n563 ;
  assign n578 = n577 ^ x405 ;
  assign n29773 = n27799 ^ n578 ;
  assign n1476 = n1475 ^ n563 ;
  assign n1483 = n1482 ^ n1476 ;
  assign n1487 = n1486 ^ n1483 ;
  assign n29774 = n29773 ^ n1487 ;
  assign n29775 = n29774 ^ n19482 ;
  assign n602 = n563 ^ x309 ;
  assign n603 = n602 ^ x501 ;
  assign n604 = n603 ^ x245 ;
  assign n601 = n578 ^ n525 ;
  assign n605 = n604 ^ n601 ;
  assign n606 = n605 ^ x500 ;
  assign n32001 = n29775 ^ n606 ;
  assign n1488 = n1487 ^ n604 ;
  assign n1495 = n1494 ^ n1488 ;
  assign n1499 = n1498 ^ n1495 ;
  assign n32002 = n32001 ^ n1499 ;
  assign n32003 = n32002 ^ n21152 ;
  assign n614 = n604 ^ x404 ;
  assign n615 = n614 ^ n613 ;
  assign n616 = n615 ^ x340 ;
  assign n610 = n606 ^ n531 ;
  assign n617 = n616 ^ n610 ;
  assign n618 = n617 ^ n555 ;
  assign n34556 = n32003 ^ n618 ;
  assign n1500 = n1499 ^ n616 ;
  assign n1513 = n1512 ^ n1500 ;
  assign n1517 = n1516 ^ n1513 ;
  assign n34557 = n34556 ^ n1517 ;
  assign n34558 = n34557 ^ n23153 ;
  assign n623 = n616 ^ x499 ;
  assign n627 = n626 ^ n623 ;
  assign n628 = n627 ^ x435 ;
  assign n622 = n618 ^ n540 ;
  assign n629 = n628 ^ n622 ;
  assign n633 = n632 ^ n629 ;
  assign n37081 = n34558 ^ n633 ;
  assign n1518 = n1517 ^ n628 ;
  assign n1531 = n1530 ^ n1518 ;
  assign n1535 = n1534 ^ n1531 ;
  assign n37082 = n37081 ^ n1535 ;
  assign n37083 = n37082 ^ n24973 ;
  assign n656 = n646 ^ n628 ;
  assign n663 = n662 ^ n656 ;
  assign n667 = n666 ^ n663 ;
  assign n655 = n648 ^ n633 ;
  assign n668 = n667 ^ n655 ;
  assign n672 = n671 ^ n668 ;
  assign n39227 = n37083 ^ n672 ;
  assign n1536 = n1535 ^ n667 ;
  assign n1549 = n1548 ^ n1536 ;
  assign n1553 = n1552 ^ n1549 ;
  assign n39228 = n39227 ^ n1553 ;
  assign n39229 = n39228 ^ n27188 ;
  assign n698 = n688 ^ n667 ;
  assign n705 = n704 ^ n698 ;
  assign n709 = n708 ^ n705 ;
  assign n697 = n690 ^ n672 ;
  assign n710 = n709 ^ n697 ;
  assign n714 = n713 ^ n710 ;
  assign n41655 = n39229 ^ n714 ;
  assign n1560 = n1559 ^ n1553 ;
  assign n1573 = n1572 ^ n1560 ;
  assign n1574 = n1573 ^ n709 ;
  assign n41656 = n41655 ^ n1574 ;
  assign n41657 = n41656 ^ n29403 ;
  assign n731 = n688 ^ x337 ;
  assign n732 = n731 ^ n678 ;
  assign n733 = n732 ^ x273 ;
  assign n746 = n733 ^ n709 ;
  assign n753 = n752 ^ n746 ;
  assign n757 = n756 ^ n753 ;
  assign n730 = n725 ^ n690 ;
  assign n734 = n733 ^ n730 ;
  assign n738 = n737 ^ n734 ;
  assign n745 = n738 ^ n714 ;
  assign n758 = n757 ^ n745 ;
  assign n762 = n761 ^ n758 ;
  assign n43766 = n41657 ^ n762 ;
  assign n1575 = n1574 ^ n757 ;
  assign n1591 = n1590 ^ n1575 ;
  assign n1595 = n1594 ^ n1591 ;
  assign n43767 = n43766 ^ n1595 ;
  assign n43768 = n43767 ^ n31356 ;
  assign n779 = n733 ^ x432 ;
  assign n780 = n779 ^ n720 ;
  assign n781 = n780 ^ x368 ;
  assign n794 = n781 ^ n757 ;
  assign n807 = n806 ^ n794 ;
  assign n811 = n810 ^ n807 ;
  assign n778 = n773 ^ n738 ;
  assign n782 = n781 ^ n778 ;
  assign n786 = n785 ^ n782 ;
  assign n793 = n786 ^ n762 ;
  assign n812 = n811 ^ n793 ;
  assign n819 = n818 ^ n812 ;
  assign n45758 = n43768 ^ n819 ;
  assign n1596 = n1595 ^ n811 ;
  assign n1612 = n1611 ^ n1596 ;
  assign n1616 = n1615 ^ n1612 ;
  assign n45759 = n45758 ^ n1616 ;
  assign n45760 = n45759 ^ n33876 ;
  assign n881 = n817 ^ x207 ;
  assign n882 = n881 ^ x399 ;
  assign n883 = n882 ^ x143 ;
  assign n849 = n785 ^ x271 ;
  assign n850 = n849 ^ x463 ;
  assign n851 = n850 ^ x207 ;
  assign n879 = n851 ^ n818 ;
  assign n874 = n810 ^ x463 ;
  assign n875 = n874 ^ n871 ;
  assign n876 = n875 ^ x399 ;
  assign n880 = n879 ^ n876 ;
  assign n884 = n883 ^ n880 ;
  assign n831 = x432 ^ x80 ;
  assign n832 = n831 ^ x272 ;
  assign n833 = n832 ^ x16 ;
  assign n845 = n833 ^ n781 ;
  assign n846 = n845 ^ n768 ;
  assign n847 = n846 ^ x463 ;
  assign n860 = n847 ^ n811 ;
  assign n873 = n872 ^ n860 ;
  assign n877 = n876 ^ n873 ;
  assign n834 = n773 ^ x335 ;
  assign n835 = n834 ^ n833 ;
  assign n836 = n835 ^ x271 ;
  assign n844 = n836 ^ n786 ;
  assign n848 = n847 ^ n844 ;
  assign n852 = n851 ^ n848 ;
  assign n859 = n852 ^ n819 ;
  assign n878 = n877 ^ n859 ;
  assign n885 = n884 ^ n878 ;
  assign n48021 = n45760 ^ n885 ;
  assign n1634 = n1615 ^ n876 ;
  assign n1635 = n1634 ^ n1631 ;
  assign n1010 = n937 ^ x399 ;
  assign n1014 = n1013 ^ n1010 ;
  assign n1015 = n1014 ^ x335 ;
  assign n1636 = n1635 ^ n1015 ;
  assign n1617 = n1616 ^ n877 ;
  assign n1633 = n1632 ^ n1617 ;
  assign n1637 = n1636 ^ n1633 ;
  assign n48022 = n48021 ^ n1637 ;
  assign n36315 = n1636 ^ n884 ;
  assign n36316 = n36315 ^ n33876 ;
  assign n1009 = n939 ^ n883 ;
  assign n1016 = n1015 ^ n1009 ;
  assign n837 = x495 ^ x143 ;
  assign n838 = n837 ^ x335 ;
  assign n839 = n838 ^ x79 ;
  assign n1017 = n1016 ^ n839 ;
  assign n36317 = n36316 ^ n1017 ;
  assign n48023 = n48022 ^ n36317 ;
  assign n953 = n883 ^ x302 ;
  assign n954 = n953 ^ x494 ;
  assign n955 = n954 ^ x238 ;
  assign n899 = x463 ^ x111 ;
  assign n900 = n899 ^ x303 ;
  assign n901 = n900 ^ x47 ;
  assign n898 = n851 ^ x366 ;
  assign n902 = n901 ^ n898 ;
  assign n903 = n902 ^ x302 ;
  assign n951 = n903 ^ n884 ;
  assign n946 = n901 ^ n876 ;
  assign n947 = n946 ^ n943 ;
  assign n948 = n947 ^ x494 ;
  assign n952 = n951 ^ n948 ;
  assign n956 = n955 ^ n952 ;
  assign n910 = n833 ^ x175 ;
  assign n911 = n910 ^ x367 ;
  assign n912 = n911 ^ x111 ;
  assign n917 = n912 ^ n847 ;
  assign n918 = n917 ^ n825 ;
  assign n919 = n918 ^ n901 ;
  assign n932 = n919 ^ n877 ;
  assign n945 = n944 ^ n932 ;
  assign n949 = n948 ^ n945 ;
  assign n913 = n836 ^ x430 ;
  assign n914 = n913 ^ n912 ;
  assign n915 = n914 ^ x366 ;
  assign n916 = n915 ^ n852 ;
  assign n920 = n919 ^ n916 ;
  assign n921 = n920 ^ n903 ;
  assign n931 = n921 ^ n885 ;
  assign n950 = n949 ^ n931 ;
  assign n957 = n956 ^ n950 ;
  assign n50090 = n48023 ^ n957 ;
  assign n1655 = n1636 ^ n948 ;
  assign n1656 = n1655 ^ n1652 ;
  assign n1107 = n1015 ^ x494 ;
  assign n1111 = n1110 ^ n1107 ;
  assign n1112 = n1111 ^ x430 ;
  assign n1657 = n1656 ^ n1112 ;
  assign n1638 = n1637 ^ n949 ;
  assign n1654 = n1653 ^ n1638 ;
  assign n1658 = n1657 ^ n1654 ;
  assign n50091 = n50090 ^ n1658 ;
  assign n38557 = n36317 ^ n956 ;
  assign n38558 = n38557 ^ n1657 ;
  assign n1106 = n1017 ^ n955 ;
  assign n1113 = n1112 ^ n1106 ;
  assign n923 = n839 ^ x238 ;
  assign n924 = n923 ^ x430 ;
  assign n925 = n924 ^ x174 ;
  assign n1114 = n1113 ^ n925 ;
  assign n38559 = n38558 ^ n1114 ;
  assign n50092 = n50091 ^ n38559 ;
  assign n50186 = n50098 ^ n50092 ;
  assign n2044 = x447 ^ x95 ;
  assign n2045 = n2044 ^ x287 ;
  assign n2046 = n2045 ^ x31 ;
  assign n2104 = n2046 ^ x190 ;
  assign n2105 = n2104 ^ x382 ;
  assign n2106 = n2105 ^ x126 ;
  assign n2173 = n2106 ^ x285 ;
  assign n2174 = n2173 ^ x477 ;
  assign n2175 = n2174 ^ x221 ;
  assign n2245 = n2175 ^ x380 ;
  assign n2242 = x477 ^ x125 ;
  assign n2243 = n2242 ^ x317 ;
  assign n2244 = n2243 ^ x61 ;
  assign n2246 = n2245 ^ n2244 ;
  assign n2247 = n2246 ^ x316 ;
  assign n2326 = n2247 ^ x475 ;
  assign n2323 = n2244 ^ x220 ;
  assign n2324 = n2323 ^ x412 ;
  assign n2325 = n2324 ^ x156 ;
  assign n2327 = n2326 ^ n2325 ;
  assign n2328 = n2327 ^ x411 ;
  assign n2256 = x475 ^ x123 ;
  assign n2257 = n2256 ^ x315 ;
  assign n2258 = n2257 ^ x59 ;
  assign n2407 = n2328 ^ n2258 ;
  assign n2404 = n2325 ^ x315 ;
  assign n2405 = n2404 ^ x507 ;
  assign n2406 = n2405 ^ x251 ;
  assign n2408 = n2407 ^ n2406 ;
  assign n2409 = n2408 ^ x506 ;
  assign n2337 = n2258 ^ x218 ;
  assign n2338 = n2337 ^ x410 ;
  assign n2339 = n2338 ^ x154 ;
  assign n24555 = n2409 ^ n2339 ;
  assign n19487 = n2406 ^ x410 ;
  assign n2144 = x507 ^ x155 ;
  assign n2145 = n2144 ^ x347 ;
  assign n2146 = n2145 ^ x91 ;
  assign n19488 = n19487 ^ n2146 ;
  assign n19489 = n19488 ^ x346 ;
  assign n24556 = n24555 ^ n19489 ;
  assign n579 = x506 ^ x154 ;
  assign n580 = n579 ^ x346 ;
  assign n581 = n580 ^ x90 ;
  assign n24557 = n24556 ^ n581 ;
  assign n2418 = n2339 ^ x313 ;
  assign n2419 = n2418 ^ x505 ;
  assign n2420 = n2419 ^ x249 ;
  assign n26484 = n24557 ^ n2420 ;
  assign n21172 = n19489 ^ x505 ;
  assign n2213 = n2146 ^ x250 ;
  assign n2214 = n2213 ^ x442 ;
  assign n2215 = n2214 ^ x186 ;
  assign n21173 = n21172 ^ n2215 ;
  assign n21174 = n21173 ^ x441 ;
  assign n26485 = n26484 ^ n21174 ;
  assign n582 = n581 ^ x249 ;
  assign n583 = n582 ^ x441 ;
  assign n584 = n583 ^ x185 ;
  assign n26486 = n26485 ^ n584 ;
  assign n19511 = n2420 ^ x408 ;
  assign n14258 = x505 ^ x153 ;
  assign n14259 = n14258 ^ x345 ;
  assign n14260 = n14259 ^ x89 ;
  assign n19512 = n19511 ^ n14260 ;
  assign n19513 = n19512 ^ x344 ;
  assign n28663 = n26486 ^ n19513 ;
  assign n23078 = n21174 ^ n14260 ;
  assign n2294 = n2215 ^ x345 ;
  assign n2295 = n2294 ^ n2291 ;
  assign n2296 = n2295 ^ x281 ;
  assign n23079 = n23078 ^ n2296 ;
  assign n23080 = n23079 ^ n566 ;
  assign n28664 = n28663 ^ n23080 ;
  assign n585 = n584 ^ x344 ;
  assign n586 = n585 ^ n566 ;
  assign n587 = n586 ^ x280 ;
  assign n28665 = n28664 ^ n587 ;
  assign n21163 = n19513 ^ x503 ;
  assign n16153 = n14260 ^ x248 ;
  assign n16154 = n16153 ^ x440 ;
  assign n16155 = n16154 ^ x184 ;
  assign n21164 = n21163 ^ n16155 ;
  assign n21165 = n21164 ^ x439 ;
  assign n30683 = n28665 ^ n21165 ;
  assign n24989 = n23080 ^ n16155 ;
  assign n2375 = n2296 ^ x440 ;
  assign n2376 = n2375 ^ n2372 ;
  assign n2377 = n2376 ^ x376 ;
  assign n24990 = n24989 ^ n2377 ;
  assign n24991 = n24990 ^ n569 ;
  assign n30684 = n30683 ^ n24991 ;
  assign n588 = n587 ^ x439 ;
  assign n589 = n588 ^ n569 ;
  assign n590 = n589 ^ x375 ;
  assign n30685 = n30684 ^ n590 ;
  assign n23131 = n21165 ^ n1480 ;
  assign n18025 = n16155 ^ x343 ;
  assign n2912 = x440 ^ x88 ;
  assign n2913 = n2912 ^ x280 ;
  assign n2914 = n2913 ^ x24 ;
  assign n18026 = n18025 ^ n2914 ;
  assign n18027 = n18026 ^ x279 ;
  assign n23132 = n23131 ^ n18027 ;
  assign n23133 = n23132 ^ n515 ;
  assign n33101 = n30685 ^ n23133 ;
  assign n27206 = n24991 ^ n18027 ;
  assign n21777 = n2914 ^ n2377 ;
  assign n21778 = n21777 ^ n16711 ;
  assign n21779 = n21778 ^ x471 ;
  assign n27207 = n27206 ^ n21779 ;
  assign n27208 = n27207 ^ n572 ;
  assign n33102 = n33101 ^ n27208 ;
  assign n591 = n590 ^ n515 ;
  assign n592 = n591 ^ n572 ;
  assign n593 = n592 ^ x470 ;
  assign n33103 = n33102 ^ n593 ;
  assign n24979 = n23133 ^ n1492 ;
  assign n19825 = n18027 ^ x438 ;
  assign n2918 = n2914 ^ x183 ;
  assign n2919 = n2918 ^ x375 ;
  assign n2920 = n2919 ^ x119 ;
  assign n19826 = n19825 ^ n2920 ;
  assign n19827 = n19826 ^ x374 ;
  assign n24980 = n24979 ^ n19827 ;
  assign n24981 = n24980 ^ n518 ;
  assign n35655 = n33103 ^ n24981 ;
  assign n28961 = n27208 ^ n19827 ;
  assign n23942 = n21779 ^ n2920 ;
  assign n23943 = n23942 ^ n18811 ;
  assign n23944 = n23943 ^ n560 ;
  assign n28962 = n28961 ^ n23944 ;
  assign n28963 = n28962 ^ n575 ;
  assign n35656 = n35655 ^ n28963 ;
  assign n594 = n593 ^ n518 ;
  assign n595 = n594 ^ n575 ;
  assign n596 = n595 ^ n545 ;
  assign n35657 = n35656 ^ n596 ;
  assign n27199 = n24981 ^ n1507 ;
  assign n21770 = n19827 ^ n1505 ;
  assign n2927 = n2920 ^ x278 ;
  assign n2928 = n2927 ^ x470 ;
  assign n2929 = n2928 ^ x214 ;
  assign n21771 = n21770 ^ n2929 ;
  assign n21772 = n21771 ^ x469 ;
  assign n27200 = n27199 ^ n21772 ;
  assign n27201 = n27200 ^ n521 ;
  assign n37656 = n35657 ^ n27201 ;
  assign n597 = n596 ^ n521 ;
  assign n598 = n597 ^ n578 ;
  assign n599 = n598 ^ n548 ;
  assign n37657 = n37656 ^ n599 ;
  assign n31394 = n28963 ^ n21772 ;
  assign n25821 = n23944 ^ n2929 ;
  assign n25822 = n25821 ^ n20760 ;
  assign n25823 = n25822 ^ n563 ;
  assign n31395 = n31394 ^ n25823 ;
  assign n31396 = n31395 ^ n578 ;
  assign n37658 = n37657 ^ n31396 ;
  assign n29414 = n27201 ^ n1525 ;
  assign n23875 = n21772 ^ n1523 ;
  assign n2936 = n2929 ^ x373 ;
  assign n2937 = n2936 ^ n545 ;
  assign n2938 = n2937 ^ x309 ;
  assign n23876 = n23875 ^ n2938 ;
  assign n23877 = n23876 ^ n525 ;
  assign n29415 = n29414 ^ n23877 ;
  assign n29416 = n29415 ^ n527 ;
  assign n40115 = n37658 ^ n29416 ;
  assign n33915 = n31396 ^ n23877 ;
  assign n27792 = n25823 ^ n2938 ;
  assign n27793 = n27792 ^ n22776 ;
  assign n27794 = n27793 ^ n604 ;
  assign n33916 = n33915 ^ n27794 ;
  assign n33917 = n33916 ^ n606 ;
  assign n40116 = n40115 ^ n33917 ;
  assign n600 = n599 ^ n527 ;
  assign n607 = n606 ^ n600 ;
  assign n608 = n607 ^ n551 ;
  assign n40117 = n40116 ^ n608 ;
  assign n31388 = n29416 ^ n1543 ;
  assign n2945 = n2938 ^ x468 ;
  assign n2946 = n2945 ^ n548 ;
  assign n2947 = n2946 ^ x404 ;
  assign n25812 = n2947 ^ n1541 ;
  assign n25813 = n25812 ^ n23877 ;
  assign n25814 = n25813 ^ n531 ;
  assign n31389 = n31388 ^ n25814 ;
  assign n31390 = n31389 ^ n533 ;
  assign n42497 = n40117 ^ n31390 ;
  assign n36333 = n33917 ^ n25814 ;
  assign n29769 = n27794 ^ n2947 ;
  assign n29770 = n29769 ^ n24537 ;
  assign n29771 = n29770 ^ n616 ;
  assign n36334 = n36333 ^ n29771 ;
  assign n36335 = n36334 ^ n618 ;
  assign n42498 = n42497 ^ n36335 ;
  assign n609 = n608 ^ n533 ;
  assign n619 = n618 ^ n609 ;
  assign n620 = n619 ^ n557 ;
  assign n42499 = n42498 ^ n620 ;
  assign n33907 = n31390 ^ n1570 ;
  assign n27784 = n25814 ^ n1567 ;
  assign n2954 = n2947 ^ n1565 ;
  assign n2955 = n2954 ^ n551 ;
  assign n2956 = n2955 ^ x499 ;
  assign n27785 = n27784 ^ n2956 ;
  assign n27786 = n27785 ^ n540 ;
  assign n33908 = n33907 ^ n27786 ;
  assign n33909 = n33908 ^ n542 ;
  assign n44326 = n42499 ^ n33909 ;
  assign n38576 = n36335 ^ n27786 ;
  assign n31996 = n29771 ^ n2956 ;
  assign n31997 = n31996 ^ n26525 ;
  assign n31998 = n31997 ^ n628 ;
  assign n38577 = n38576 ^ n31998 ;
  assign n38578 = n38577 ^ n633 ;
  assign n44327 = n44326 ^ n38578 ;
  assign n621 = n620 ^ n542 ;
  assign n634 = n633 ^ n621 ;
  assign n638 = n637 ^ n634 ;
  assign n44328 = n44327 ^ n638 ;
  assign n36325 = n33909 ^ n1585 ;
  assign n29761 = n27786 ^ n1583 ;
  assign n2963 = n2956 ^ n1581 ;
  assign n2964 = n2963 ^ n557 ;
  assign n2965 = n2964 ^ n646 ;
  assign n29762 = n29761 ^ n2965 ;
  assign n29763 = n29762 ^ n648 ;
  assign n36326 = n36325 ^ n29763 ;
  assign n36327 = n36326 ^ n653 ;
  assign n46371 = n44328 ^ n36327 ;
  assign n40867 = n38578 ^ n29763 ;
  assign n34551 = n31998 ^ n2965 ;
  assign n34552 = n34551 ^ n28622 ;
  assign n34553 = n34552 ^ n667 ;
  assign n40868 = n40867 ^ n34553 ;
  assign n40869 = n40868 ^ n672 ;
  assign n46372 = n46371 ^ n40869 ;
  assign n654 = n653 ^ n638 ;
  assign n673 = n672 ^ n654 ;
  assign n680 = n679 ^ n673 ;
  assign n46373 = n46372 ^ n680 ;
  assign n38569 = n36327 ^ n1606 ;
  assign n38570 = n38569 ^ n695 ;
  assign n31989 = n29763 ^ n1604 ;
  assign n2972 = n2965 ^ n1602 ;
  assign n2973 = n2972 ^ n637 ;
  assign n2974 = n2973 ^ n688 ;
  assign n31990 = n31989 ^ n2974 ;
  assign n31991 = n31990 ^ n690 ;
  assign n38571 = n38570 ^ n31991 ;
  assign n48730 = n46373 ^ n38571 ;
  assign n42888 = n40869 ^ n31991 ;
  assign n37076 = n34553 ^ n2974 ;
  assign n37077 = n37076 ^ n30664 ;
  assign n37078 = n37077 ^ n709 ;
  assign n42889 = n42888 ^ n37078 ;
  assign n42890 = n42889 ^ n714 ;
  assign n48731 = n48730 ^ n42890 ;
  assign n696 = n695 ^ n680 ;
  assign n715 = n714 ^ n696 ;
  assign n722 = n721 ^ n715 ;
  assign n48732 = n48731 ^ n722 ;
  assign n1357 = x427 ^ x267 ;
  assign n1358 = n1357 ^ x75 ;
  assign n1359 = n1358 ^ x11 ;
  assign n2794 = n1359 ^ x170 ;
  assign n2795 = n2794 ^ x362 ;
  assign n2796 = n2795 ^ x106 ;
  assign n1026 = x494 ^ x142 ;
  assign n1027 = n1026 ^ x334 ;
  assign n1028 = n1027 ^ x78 ;
  assign n1100 = n1028 ^ x237 ;
  assign n1101 = n1100 ^ x429 ;
  assign n1102 = n1101 ^ x173 ;
  assign n1209 = n1102 ^ x332 ;
  assign n1201 = x429 ^ x77 ;
  assign n1202 = n1201 ^ x269 ;
  assign n1203 = n1202 ^ x13 ;
  assign n1210 = n1209 ^ n1203 ;
  assign n1211 = n1210 ^ x268 ;
  assign n1311 = n1211 ^ x427 ;
  assign n1303 = n1203 ^ x172 ;
  assign n1304 = n1303 ^ x364 ;
  assign n1305 = n1304 ^ x108 ;
  assign n1312 = n1311 ^ n1305 ;
  assign n1313 = n1312 ^ x363 ;
  assign n1425 = n1359 ^ n1313 ;
  assign n1407 = n1305 ^ x267 ;
  assign n1408 = n1407 ^ x459 ;
  assign n1409 = n1408 ^ x203 ;
  assign n1426 = n1425 ^ n1409 ;
  assign n1427 = n1426 ^ x458 ;
  assign n2835 = n2796 ^ n1427 ;
  assign n2832 = n1409 ^ x362 ;
  assign n1236 = x459 ^ x107 ;
  assign n1237 = n1236 ^ x299 ;
  assign n1238 = n1237 ^ x43 ;
  assign n2833 = n2832 ^ n1238 ;
  assign n2834 = n2833 ^ x298 ;
  assign n2836 = n2835 ^ n2834 ;
  assign n2499 = x458 ^ x106 ;
  assign n2500 = n2499 ^ x298 ;
  assign n2501 = n2500 ^ x42 ;
  assign n2837 = n2836 ^ n2501 ;
  assign n2808 = n2796 ^ x265 ;
  assign n2809 = n2808 ^ x457 ;
  assign n2810 = n2809 ^ x201 ;
  assign n2880 = n2837 ^ n2810 ;
  assign n2877 = n2834 ^ x457 ;
  assign n1374 = n1238 ^ x202 ;
  assign n1375 = n1374 ^ x394 ;
  assign n1376 = n1375 ^ x138 ;
  assign n2878 = n2877 ^ n1376 ;
  assign n2879 = n2878 ^ x393 ;
  assign n2881 = n2880 ^ n2879 ;
  assign n2502 = n2501 ^ x201 ;
  assign n2503 = n2502 ^ x393 ;
  assign n2504 = n2503 ^ x137 ;
  assign n2882 = n2881 ^ n2504 ;
  assign n2854 = n2810 ^ x360 ;
  assign n2846 = x457 ^ x297 ;
  assign n2847 = n2846 ^ x105 ;
  assign n2848 = n2847 ^ x41 ;
  assign n2855 = n2854 ^ n2848 ;
  assign n2856 = n2855 ^ x296 ;
  assign n27865 = n2882 ^ n2856 ;
  assign n22746 = n2879 ^ n2848 ;
  assign n3201 = n1376 ^ x297 ;
  assign n3202 = n3201 ^ x489 ;
  assign n3203 = n3202 ^ x233 ;
  assign n22747 = n22746 ^ n3203 ;
  assign n22748 = n22747 ^ x488 ;
  assign n27866 = n27865 ^ n22748 ;
  assign n2505 = n2504 ^ x296 ;
  assign n2506 = n2505 ^ x488 ;
  assign n2507 = n2506 ^ x232 ;
  assign n27867 = n27866 ^ n2507 ;
  assign n2899 = n2856 ^ x455 ;
  assign n2891 = n2848 ^ x200 ;
  assign n2892 = n2891 ^ x392 ;
  assign n2893 = n2892 ^ x136 ;
  assign n2900 = n2899 ^ n2893 ;
  assign n2901 = n2900 ^ x391 ;
  assign n30204 = n27867 ^ n2901 ;
  assign n24510 = n22748 ^ n2893 ;
  assign n3204 = n3203 ^ x392 ;
  assign n2616 = x489 ^ x137 ;
  assign n2617 = n2616 ^ x329 ;
  assign n2618 = n2617 ^ x73 ;
  assign n3205 = n3204 ^ n2618 ;
  assign n3206 = n3205 ^ x328 ;
  assign n24511 = n24510 ^ n3206 ;
  assign n2476 = x328 ^ x136 ;
  assign n2477 = n2476 ^ x488 ;
  assign n2478 = n2477 ^ x72 ;
  assign n24512 = n24511 ^ n2478 ;
  assign n30205 = n30204 ^ n24512 ;
  assign n2508 = n2507 ^ x391 ;
  assign n2509 = n2508 ^ n2478 ;
  assign n2510 = n2509 ^ x327 ;
  assign n30206 = n30205 ^ n2510 ;
  assign n1827 = x455 ^ x39 ;
  assign n1828 = n1827 ^ x295 ;
  assign n1829 = n1828 ^ x103 ;
  assign n3099 = n2901 ^ n1829 ;
  assign n3090 = n2893 ^ x295 ;
  assign n3091 = n3090 ^ x487 ;
  assign n3092 = n3091 ^ x231 ;
  assign n3100 = n3099 ^ n3092 ;
  assign n3101 = n3100 ^ x486 ;
  assign n32516 = n30206 ^ n3101 ;
  assign n26441 = n24512 ^ n3092 ;
  assign n3207 = n3206 ^ x487 ;
  assign n2619 = n2618 ^ x232 ;
  assign n2620 = n2619 ^ x424 ;
  assign n2621 = n2620 ^ x168 ;
  assign n3208 = n3207 ^ n2621 ;
  assign n3209 = n3208 ^ x423 ;
  assign n26442 = n26441 ^ n3209 ;
  assign n2475 = x423 ^ x231 ;
  assign n2479 = n2478 ^ n2475 ;
  assign n2480 = n2479 ^ x167 ;
  assign n26443 = n26442 ^ n2480 ;
  assign n32517 = n32516 ^ n26443 ;
  assign n2511 = n2510 ^ x486 ;
  assign n2512 = n2511 ^ n2480 ;
  assign n2513 = n2512 ^ x422 ;
  assign n32518 = n32517 ^ n2513 ;
  assign n2460 = x486 ^ x134 ;
  assign n2461 = n2460 ^ x326 ;
  assign n2462 = n2461 ^ x70 ;
  assign n2514 = n2513 ^ n2462 ;
  assign n2482 = x263 ^ x71 ;
  assign n2483 = n2482 ^ x423 ;
  assign n2484 = n2483 ^ x7 ;
  assign n2481 = n2480 ^ x326 ;
  assign n2485 = n2484 ^ n2481 ;
  assign n2486 = n2485 ^ x262 ;
  assign n2515 = n2514 ^ n2486 ;
  assign n2442 = x422 ^ x70 ;
  assign n2443 = n2442 ^ x262 ;
  assign n2444 = n2443 ^ x6 ;
  assign n2516 = n2515 ^ n2444 ;
  assign n35113 = n32518 ^ n2516 ;
  assign n3094 = x487 ^ x135 ;
  assign n3095 = n3094 ^ x327 ;
  assign n3096 = n3095 ^ x71 ;
  assign n3093 = n3092 ^ x390 ;
  assign n3097 = n3096 ^ n3093 ;
  assign n3098 = n3097 ^ x326 ;
  assign n28587 = n26443 ^ n3098 ;
  assign n3210 = n3209 ^ n3096 ;
  assign n2622 = n2621 ^ x327 ;
  assign n2555 = x424 ^ x72 ;
  assign n2556 = n2555 ^ x264 ;
  assign n2557 = n2556 ^ x8 ;
  assign n2623 = n2622 ^ n2557 ;
  assign n2624 = n2623 ^ x263 ;
  assign n3211 = n3210 ^ n2624 ;
  assign n3212 = n3211 ^ n2484 ;
  assign n28588 = n28587 ^ n3212 ;
  assign n28589 = n28588 ^ n2486 ;
  assign n35114 = n35113 ^ n28589 ;
  assign n1830 = n1829 ^ x198 ;
  assign n1831 = n1830 ^ x390 ;
  assign n1832 = n1831 ^ x134 ;
  assign n3102 = n3101 ^ n1832 ;
  assign n3103 = n3102 ^ n3098 ;
  assign n3104 = n3103 ^ n2462 ;
  assign n35115 = n35114 ^ n3104 ;
  assign n1833 = n1832 ^ x293 ;
  assign n1834 = n1833 ^ x485 ;
  assign n1835 = n1834 ^ x229 ;
  assign n3136 = n3104 ^ n1835 ;
  assign n3131 = n3096 ^ x230 ;
  assign n3132 = n3131 ^ x422 ;
  assign n3133 = n3132 ^ x166 ;
  assign n3130 = n3098 ^ x485 ;
  assign n3134 = n3133 ^ n3130 ;
  assign n3135 = n3134 ^ x421 ;
  assign n3137 = n3136 ^ n3135 ;
  assign n2463 = n2462 ^ x229 ;
  assign n2464 = n2463 ^ x421 ;
  assign n2465 = n2464 ^ x165 ;
  assign n3138 = n3137 ^ n2465 ;
  assign n37385 = n35115 ^ n3138 ;
  assign n30855 = n28589 ^ n3135 ;
  assign n3213 = n3212 ^ n3133 ;
  assign n2625 = n2624 ^ x422 ;
  assign n2567 = n2557 ^ x167 ;
  assign n2568 = n2567 ^ x359 ;
  assign n2569 = n2568 ^ x103 ;
  assign n2626 = n2625 ^ n2569 ;
  assign n2627 = n2626 ^ x358 ;
  assign n3214 = n3213 ^ n2627 ;
  assign n2488 = n2484 ^ x166 ;
  assign n2489 = n2488 ^ x358 ;
  assign n2490 = n2489 ^ x102 ;
  assign n3215 = n3214 ^ n2490 ;
  assign n30856 = n30855 ^ n3215 ;
  assign n2487 = n2486 ^ x421 ;
  assign n2491 = n2490 ^ n2487 ;
  assign n2492 = n2491 ^ x357 ;
  assign n30857 = n30856 ^ n2492 ;
  assign n37386 = n37385 ^ n30857 ;
  assign n2517 = n2516 ^ n2465 ;
  assign n2518 = n2517 ^ n2492 ;
  assign n2445 = n2444 ^ x165 ;
  assign n2446 = n2445 ^ x357 ;
  assign n2447 = n2446 ^ x101 ;
  assign n2519 = n2518 ^ n2447 ;
  assign n37387 = n37386 ^ n2519 ;
  assign n1836 = n1835 ^ x388 ;
  assign n1812 = x485 ^ x133 ;
  assign n1813 = n1812 ^ x325 ;
  assign n1814 = n1813 ^ x69 ;
  assign n1837 = n1836 ^ n1814 ;
  assign n1838 = n1837 ^ x324 ;
  assign n3151 = n3138 ^ n1838 ;
  assign n3146 = n3133 ^ x325 ;
  assign n3147 = n3146 ^ n2444 ;
  assign n3148 = n3147 ^ x261 ;
  assign n3145 = n3135 ^ n1814 ;
  assign n3149 = n3148 ^ n3145 ;
  assign n2457 = x421 ^ x69 ;
  assign n2458 = n2457 ^ x261 ;
  assign n2459 = n2458 ^ x5 ;
  assign n3150 = n3149 ^ n2459 ;
  assign n3152 = n3151 ^ n3150 ;
  assign n2466 = n2465 ^ x324 ;
  assign n2467 = n2466 ^ n2459 ;
  assign n2468 = n2467 ^ x260 ;
  assign n3153 = n3152 ^ n2468 ;
  assign n39658 = n37387 ^ n3153 ;
  assign n2520 = n2519 ^ n2468 ;
  assign n2494 = n2490 ^ x261 ;
  assign n2495 = n2494 ^ x453 ;
  assign n2496 = n2495 ^ x197 ;
  assign n2493 = n2492 ^ n2459 ;
  assign n2497 = n2496 ^ n2493 ;
  assign n2498 = n2497 ^ x452 ;
  assign n2521 = n2520 ^ n2498 ;
  assign n2448 = n2447 ^ x260 ;
  assign n2449 = n2448 ^ x452 ;
  assign n2450 = n2449 ^ x196 ;
  assign n2522 = n2521 ^ n2450 ;
  assign n39659 = n39658 ^ n2522 ;
  assign n33308 = n30857 ^ n3150 ;
  assign n3216 = n3215 ^ n3148 ;
  assign n2628 = n2627 ^ n2444 ;
  assign n2579 = n2569 ^ x262 ;
  assign n2580 = n2579 ^ x454 ;
  assign n2581 = n2580 ^ x198 ;
  assign n2629 = n2628 ^ n2581 ;
  assign n2630 = n2629 ^ x453 ;
  assign n3217 = n3216 ^ n2630 ;
  assign n3218 = n3217 ^ n2496 ;
  assign n33309 = n33308 ^ n3218 ;
  assign n33310 = n33309 ^ n2498 ;
  assign n39660 = n39659 ^ n33310 ;
  assign n1839 = n1838 ^ x483 ;
  assign n1815 = n1814 ^ x228 ;
  assign n1816 = n1815 ^ x420 ;
  assign n1817 = n1816 ^ x164 ;
  assign n1840 = n1839 ^ n1817 ;
  assign n1841 = n1840 ^ x419 ;
  assign n3169 = n3153 ^ n1841 ;
  assign n3164 = n3148 ^ x420 ;
  assign n3165 = n3164 ^ n2447 ;
  assign n3166 = n3165 ^ x356 ;
  assign n3163 = n3150 ^ n1817 ;
  assign n3167 = n3166 ^ n3163 ;
  assign n2470 = n2459 ^ x164 ;
  assign n2471 = n2470 ^ x356 ;
  assign n2472 = n2471 ^ x100 ;
  assign n3168 = n3167 ^ n2472 ;
  assign n3170 = n3169 ^ n3168 ;
  assign n2469 = n2468 ^ x419 ;
  assign n2473 = n2472 ^ n2469 ;
  assign n2474 = n2473 ^ x355 ;
  assign n3171 = n3170 ^ n2474 ;
  assign n41836 = n39660 ^ n3171 ;
  assign n35934 = n33310 ^ n3168 ;
  assign n3219 = n3218 ^ n3166 ;
  assign n2631 = n2630 ^ n2447 ;
  assign n2594 = n2581 ^ x357 ;
  assign n2584 = x454 ^ x102 ;
  assign n2585 = n2584 ^ x38 ;
  assign n2586 = n2585 ^ x294 ;
  assign n2595 = n2594 ^ n2586 ;
  assign n2596 = n2595 ^ x293 ;
  assign n2632 = n2631 ^ n2596 ;
  assign n2526 = x293 ^ x101 ;
  assign n2527 = n2526 ^ x453 ;
  assign n2528 = n2527 ^ x37 ;
  assign n2633 = n2632 ^ n2528 ;
  assign n3220 = n3219 ^ n2633 ;
  assign n2525 = n2496 ^ x356 ;
  assign n2529 = n2528 ^ n2525 ;
  assign n2530 = n2529 ^ x292 ;
  assign n3221 = n3220 ^ n2530 ;
  assign n35935 = n35934 ^ n3221 ;
  assign n2524 = n2498 ^ n2472 ;
  assign n2531 = n2530 ^ n2524 ;
  assign n2452 = x452 ^ x36 ;
  assign n2453 = n2452 ^ x100 ;
  assign n2454 = n2453 ^ x292 ;
  assign n2532 = n2531 ^ n2454 ;
  assign n35936 = n35935 ^ n2532 ;
  assign n41837 = n41836 ^ n35936 ;
  assign n2523 = n2522 ^ n2474 ;
  assign n2533 = n2532 ^ n2523 ;
  assign n2451 = n2450 ^ x355 ;
  assign n2455 = n2454 ^ n2451 ;
  assign n2456 = n2455 ^ x291 ;
  assign n2534 = n2533 ^ n2456 ;
  assign n41838 = n41837 ^ n2534 ;
  assign n1776 = x483 ^ x131 ;
  assign n1777 = n1776 ^ x323 ;
  assign n1778 = n1777 ^ x67 ;
  assign n1842 = n1841 ^ n1778 ;
  assign n1818 = n1817 ^ x323 ;
  assign n1803 = x420 ^ x68 ;
  assign n1804 = n1803 ^ x260 ;
  assign n1805 = n1804 ^ x4 ;
  assign n1819 = n1818 ^ n1805 ;
  assign n1820 = n1819 ^ x259 ;
  assign n1843 = n1842 ^ n1820 ;
  assign n1794 = x419 ^ x67 ;
  assign n1795 = n1794 ^ x259 ;
  assign n1796 = n1795 ^ x3 ;
  assign n1844 = n1843 ^ n1796 ;
  assign n3191 = n3171 ^ n1844 ;
  assign n3186 = n3166 ^ n1805 ;
  assign n3187 = n3186 ^ n2450 ;
  assign n3188 = n3187 ^ x451 ;
  assign n3185 = n3168 ^ n1820 ;
  assign n3189 = n3188 ^ n3185 ;
  assign n2692 = n2472 ^ x259 ;
  assign n2693 = n2692 ^ x451 ;
  assign n2694 = n2693 ^ x195 ;
  assign n3190 = n3189 ^ n2694 ;
  assign n3192 = n3191 ^ n3190 ;
  assign n2691 = n2474 ^ n1796 ;
  assign n2695 = n2694 ^ n2691 ;
  assign n2696 = n2695 ^ x450 ;
  assign n3193 = n3192 ^ n2696 ;
  assign n43854 = n41838 ^ n3193 ;
  assign n38199 = n35936 ^ n3190 ;
  assign n2699 = n2530 ^ x451 ;
  assign n2613 = n2528 ^ x196 ;
  assign n2614 = n2613 ^ x388 ;
  assign n2615 = n2614 ^ x132 ;
  assign n2700 = n2699 ^ n2615 ;
  assign n2701 = n2700 ^ x387 ;
  assign n2698 = n2694 ^ n2532 ;
  assign n2702 = n2701 ^ n2698 ;
  assign n2686 = n2454 ^ x195 ;
  assign n2687 = n2686 ^ x387 ;
  assign n2688 = n2687 ^ x131 ;
  assign n2703 = n2702 ^ n2688 ;
  assign n38200 = n38199 ^ n2703 ;
  assign n3222 = n3221 ^ n3188 ;
  assign n2634 = n2633 ^ n2450 ;
  assign n2609 = n2596 ^ x452 ;
  assign n2599 = n2586 ^ x197 ;
  assign n2600 = n2599 ^ x389 ;
  assign n2601 = n2600 ^ x133 ;
  assign n2610 = n2609 ^ n2601 ;
  assign n2611 = n2610 ^ x388 ;
  assign n2635 = n2634 ^ n2611 ;
  assign n2636 = n2635 ^ n2615 ;
  assign n3223 = n3222 ^ n2636 ;
  assign n3224 = n3223 ^ n2701 ;
  assign n38201 = n38200 ^ n3224 ;
  assign n43855 = n43854 ^ n38201 ;
  assign n2697 = n2696 ^ n2534 ;
  assign n2704 = n2703 ^ n2697 ;
  assign n2685 = n2456 ^ x450 ;
  assign n2689 = n2688 ^ n2685 ;
  assign n2690 = n2689 ^ x386 ;
  assign n2705 = n2704 ^ n2690 ;
  assign n43856 = n43855 ^ n2705 ;
  assign n1779 = n1778 ^ x226 ;
  assign n1780 = n1779 ^ x418 ;
  assign n1781 = n1780 ^ x162 ;
  assign n1845 = n1844 ^ n1781 ;
  assign n1821 = n1820 ^ x418 ;
  assign n1806 = n1805 ^ x163 ;
  assign n1807 = n1806 ^ x355 ;
  assign n1808 = n1807 ^ x99 ;
  assign n1822 = n1821 ^ n1808 ;
  assign n1823 = n1822 ^ x354 ;
  assign n1846 = n1845 ^ n1823 ;
  assign n1797 = n1796 ^ x162 ;
  assign n1798 = n1797 ^ x354 ;
  assign n1799 = n1798 ^ x98 ;
  assign n1847 = n1846 ^ n1799 ;
  assign n35602 = n3193 ^ n1847 ;
  assign n3231 = n3190 ^ n1823 ;
  assign n3195 = n3188 ^ n1808 ;
  assign n3196 = n3195 ^ n2456 ;
  assign n2740 = x451 ^ x99 ;
  assign n2741 = n2740 ^ x291 ;
  assign n2742 = n2741 ^ x35 ;
  assign n3197 = n3196 ^ n2742 ;
  assign n3232 = n3231 ^ n3197 ;
  assign n2739 = n2694 ^ x354 ;
  assign n2743 = n2742 ^ n2739 ;
  assign n2744 = n2743 ^ x290 ;
  assign n3233 = n3232 ^ n2744 ;
  assign n35603 = n35602 ^ n3233 ;
  assign n2751 = n2696 ^ n1799 ;
  assign n2752 = n2751 ^ n2744 ;
  assign n1854 = x450 ^ x98 ;
  assign n1855 = n1854 ^ x290 ;
  assign n1856 = n1855 ^ x34 ;
  assign n2753 = n2752 ^ n1856 ;
  assign n35604 = n35603 ^ n2753 ;
  assign n45846 = n43856 ^ n35604 ;
  assign n40170 = n38201 ^ n3233 ;
  assign n3225 = n3224 ^ n3197 ;
  assign n2681 = n2636 ^ n2456 ;
  assign n2673 = n2611 ^ n2454 ;
  assign n2663 = n2601 ^ x292 ;
  assign n2664 = n2663 ^ x484 ;
  assign n2665 = n2664 ^ x228 ;
  assign n2674 = n2673 ^ n2665 ;
  assign n2675 = n2674 ^ x483 ;
  assign n2682 = n2681 ^ n2675 ;
  assign n2678 = n2615 ^ x291 ;
  assign n2679 = n2678 ^ x483 ;
  assign n2680 = n2679 ^ x227 ;
  assign n2683 = n2682 ^ n2680 ;
  assign n3226 = n3225 ^ n2683 ;
  assign n2746 = n2742 ^ n2701 ;
  assign n2747 = n2746 ^ n2680 ;
  assign n2748 = n2747 ^ x482 ;
  assign n3227 = n3226 ^ n2748 ;
  assign n40171 = n40170 ^ n3227 ;
  assign n2745 = n2744 ^ n2703 ;
  assign n2749 = n2748 ^ n2745 ;
  assign n2734 = n2688 ^ x290 ;
  assign n2735 = n2734 ^ x482 ;
  assign n2736 = n2735 ^ x226 ;
  assign n2750 = n2749 ^ n2736 ;
  assign n40172 = n40171 ^ n2750 ;
  assign n45847 = n45846 ^ n40172 ;
  assign n2754 = n2753 ^ n2750 ;
  assign n2755 = n2754 ^ n2705 ;
  assign n2733 = n2690 ^ n1856 ;
  assign n2737 = n2736 ^ n2733 ;
  assign n2738 = n2737 ^ x481 ;
  assign n2756 = n2755 ^ n2738 ;
  assign n45848 = n45847 ^ n2756 ;
  assign n1783 = x418 ^ x66 ;
  assign n1784 = n1783 ^ x258 ;
  assign n1785 = n1784 ^ x2 ;
  assign n1782 = n1781 ^ x321 ;
  assign n1786 = n1785 ^ n1782 ;
  assign n1787 = n1786 ^ x257 ;
  assign n1848 = n1847 ^ n1787 ;
  assign n1824 = n1823 ^ n1785 ;
  assign n1809 = n1808 ^ x258 ;
  assign n1810 = n1809 ^ x450 ;
  assign n1811 = n1810 ^ x194 ;
  assign n1825 = n1824 ^ n1811 ;
  assign n1826 = n1825 ^ x449 ;
  assign n1849 = n1848 ^ n1826 ;
  assign n1800 = n1799 ^ x257 ;
  assign n1801 = n1800 ^ x449 ;
  assign n1802 = n1801 ^ x193 ;
  assign n1850 = n1849 ^ n1802 ;
  assign n37702 = n35604 ^ n1850 ;
  assign n2996 = n2742 ^ x194 ;
  assign n2997 = n2996 ^ x386 ;
  assign n2998 = n2997 ^ x130 ;
  assign n2995 = n2744 ^ x449 ;
  assign n2999 = n2998 ^ n2995 ;
  assign n3000 = n2999 ^ x385 ;
  assign n2994 = n2753 ^ n1802 ;
  assign n3001 = n3000 ^ n2994 ;
  assign n1881 = n1856 ^ x193 ;
  assign n1882 = n1881 ^ x385 ;
  assign n1883 = n1882 ^ x129 ;
  assign n3002 = n3001 ^ n1883 ;
  assign n37703 = n37702 ^ n3002 ;
  assign n3234 = n3233 ^ n1826 ;
  assign n3198 = n3197 ^ n1811 ;
  assign n3199 = n3198 ^ n2690 ;
  assign n3200 = n3199 ^ n2998 ;
  assign n3235 = n3234 ^ n3200 ;
  assign n3236 = n3235 ^ n3000 ;
  assign n37704 = n37703 ^ n3236 ;
  assign n47653 = n45848 ^ n37704 ;
  assign n41974 = n40172 ^ n3236 ;
  assign n3228 = n3227 ^ n3200 ;
  assign n2728 = n2680 ^ x386 ;
  assign n2729 = n2728 ^ n1778 ;
  assign n2730 = n2729 ^ x322 ;
  assign n2726 = n2690 ^ n2683 ;
  assign n2721 = n2688 ^ n2675 ;
  assign n2709 = x484 ^ x132 ;
  assign n2710 = n2709 ^ x324 ;
  assign n2711 = n2710 ^ x68 ;
  assign n2708 = n2665 ^ x387 ;
  assign n2712 = n2711 ^ n2708 ;
  assign n2713 = n2712 ^ x323 ;
  assign n2722 = n2721 ^ n2713 ;
  assign n2723 = n2722 ^ n1778 ;
  assign n2727 = n2726 ^ n2723 ;
  assign n2731 = n2730 ^ n2727 ;
  assign n3229 = n3228 ^ n2731 ;
  assign n3007 = x482 ^ x130 ;
  assign n3008 = n3007 ^ x322 ;
  assign n3009 = n3008 ^ x66 ;
  assign n3005 = n2998 ^ n2748 ;
  assign n3006 = n3005 ^ n2730 ;
  assign n3010 = n3009 ^ n3006 ;
  assign n3230 = n3229 ^ n3010 ;
  assign n41975 = n41974 ^ n3230 ;
  assign n3012 = n2736 ^ x385 ;
  assign n3013 = n3012 ^ n3009 ;
  assign n3014 = n3013 ^ x321 ;
  assign n3004 = n3000 ^ n2750 ;
  assign n3011 = n3010 ^ n3004 ;
  assign n3015 = n3014 ^ n3011 ;
  assign n41976 = n41975 ^ n3015 ;
  assign n47654 = n47653 ^ n41976 ;
  assign n3019 = x481 ^ x129 ;
  assign n3020 = n3019 ^ x321 ;
  assign n3021 = n3020 ^ x65 ;
  assign n3017 = n2738 ^ n1883 ;
  assign n3018 = n3017 ^ n3014 ;
  assign n3022 = n3021 ^ n3018 ;
  assign n3003 = n3002 ^ n2756 ;
  assign n3016 = n3015 ^ n3003 ;
  assign n3023 = n3022 ^ n3016 ;
  assign n47655 = n47654 ^ n3023 ;
  assign n972 = x430 ^ x78 ;
  assign n973 = n972 ^ x270 ;
  assign n974 = n973 ^ x14 ;
  assign n1059 = n974 ^ x173 ;
  assign n1060 = n1059 ^ x365 ;
  assign n1061 = n1060 ^ x109 ;
  assign n1146 = n1061 ^ x268 ;
  assign n1147 = n1146 ^ x460 ;
  assign n1148 = n1147 ^ x204 ;
  assign n1248 = n1148 ^ x363 ;
  assign n1242 = x460 ^ x108 ;
  assign n1243 = n1242 ^ x300 ;
  assign n1244 = n1243 ^ x44 ;
  assign n1249 = n1248 ^ n1244 ;
  assign n1250 = n1249 ^ x299 ;
  assign n1347 = n1250 ^ x458 ;
  assign n1341 = n1244 ^ x203 ;
  assign n1342 = n1341 ^ x395 ;
  assign n1343 = n1342 ^ x139 ;
  assign n1348 = n1347 ^ n1343 ;
  assign n1349 = n1348 ^ x394 ;
  assign n2637 = n2501 ^ n1349 ;
  assign n2535 = n1343 ^ x298 ;
  assign n2536 = n2535 ^ x490 ;
  assign n2537 = n2536 ^ x234 ;
  assign n2638 = n2637 ^ n2537 ;
  assign n2639 = n2638 ^ x489 ;
  assign n975 = n974 ^ n915 ;
  assign n969 = n912 ^ x270 ;
  assign n970 = n969 ^ x462 ;
  assign n971 = n970 ^ x206 ;
  assign n976 = n975 ^ n971 ;
  assign n977 = n976 ^ x461 ;
  assign n1062 = n1061 ^ n977 ;
  assign n1056 = n971 ^ x365 ;
  assign n905 = x462 ^ x110 ;
  assign n906 = n905 ^ x302 ;
  assign n907 = n906 ^ x46 ;
  assign n1057 = n1056 ^ n907 ;
  assign n1058 = n1057 ^ x301 ;
  assign n1063 = n1062 ^ n1058 ;
  assign n1051 = x461 ^ x109 ;
  assign n1052 = n1051 ^ x301 ;
  assign n1053 = n1052 ^ x45 ;
  assign n1064 = n1063 ^ n1053 ;
  assign n1149 = n1148 ^ n1064 ;
  assign n1143 = n1058 ^ x460 ;
  assign n1000 = n907 ^ x205 ;
  assign n1001 = n1000 ^ x397 ;
  assign n1002 = n1001 ^ x141 ;
  assign n1144 = n1143 ^ n1002 ;
  assign n1145 = n1144 ^ x396 ;
  assign n1150 = n1149 ^ n1145 ;
  assign n1138 = n1053 ^ x204 ;
  assign n1139 = n1138 ^ x396 ;
  assign n1140 = n1139 ^ x140 ;
  assign n1151 = n1150 ^ n1140 ;
  assign n1251 = n1250 ^ n1151 ;
  assign n1245 = n1244 ^ n1145 ;
  assign n1087 = x492 ^ x300 ;
  assign n1088 = n1087 ^ n1002 ;
  assign n1089 = n1088 ^ x236 ;
  assign n1246 = n1245 ^ n1089 ;
  assign n1247 = n1246 ^ x491 ;
  assign n1252 = n1251 ^ n1247 ;
  assign n1233 = n1140 ^ x299 ;
  assign n1234 = n1233 ^ x491 ;
  assign n1235 = n1234 ^ x235 ;
  assign n1253 = n1252 ^ n1235 ;
  assign n1350 = n1349 ^ n1253 ;
  assign n1344 = n1343 ^ n1247 ;
  assign n1180 = n1089 ^ x395 ;
  assign n1172 = x492 ^ x140 ;
  assign n1173 = n1172 ^ x332 ;
  assign n1174 = n1173 ^ x76 ;
  assign n1181 = n1180 ^ n1174 ;
  assign n1182 = n1181 ^ x331 ;
  assign n1345 = n1344 ^ n1182 ;
  assign n1336 = x491 ^ x139 ;
  assign n1337 = n1336 ^ x331 ;
  assign n1338 = n1337 ^ x75 ;
  assign n1346 = n1345 ^ n1338 ;
  assign n1351 = n1350 ^ n1346 ;
  assign n1335 = n1235 ^ x394 ;
  assign n1339 = n1338 ^ n1335 ;
  assign n1340 = n1339 ^ x330 ;
  assign n1352 = n1351 ^ n1340 ;
  assign n32531 = n2639 ^ n1352 ;
  assign n2786 = n1338 ^ x234 ;
  assign n2787 = n2786 ^ x426 ;
  assign n2788 = n2787 ^ x170 ;
  assign n2784 = n2537 ^ n1346 ;
  assign n1282 = n1182 ^ x490 ;
  assign n1274 = n1174 ^ x235 ;
  assign n1275 = n1274 ^ x427 ;
  assign n1276 = n1275 ^ x171 ;
  assign n1283 = n1282 ^ n1276 ;
  assign n1284 = n1283 ^ x426 ;
  assign n2785 = n2784 ^ n1284 ;
  assign n2789 = n2788 ^ n2785 ;
  assign n32532 = n32531 ^ n2789 ;
  assign n21514 = n1340 ^ x489 ;
  assign n21515 = n21514 ^ n2788 ;
  assign n21516 = n21515 ^ x425 ;
  assign n32533 = n32532 ^ n21516 ;
  assign n1366 = n1276 ^ x330 ;
  assign n1367 = n1366 ^ n1359 ;
  assign n1368 = n1367 ^ x266 ;
  assign n993 = n903 ^ x461 ;
  assign n988 = n901 ^ x206 ;
  assign n989 = n988 ^ x398 ;
  assign n990 = n989 ^ x142 ;
  assign n994 = n993 ^ n990 ;
  assign n995 = n994 ^ x397 ;
  assign n1080 = n1053 ^ n995 ;
  assign n1075 = n990 ^ x301 ;
  assign n1076 = n1075 ^ x493 ;
  assign n1077 = n1076 ^ x237 ;
  assign n1081 = n1080 ^ n1077 ;
  assign n1082 = n1081 ^ x492 ;
  assign n1170 = n1140 ^ n1082 ;
  assign n1165 = n1077 ^ x396 ;
  assign n1044 = x493 ^ x141 ;
  assign n1045 = n1044 ^ x333 ;
  assign n1046 = n1045 ^ x77 ;
  assign n1166 = n1165 ^ n1046 ;
  assign n1167 = n1166 ^ x332 ;
  assign n1171 = n1170 ^ n1167 ;
  assign n1175 = n1174 ^ n1171 ;
  assign n1272 = n1235 ^ n1175 ;
  assign n1267 = n1167 ^ x491 ;
  assign n1131 = n1046 ^ x236 ;
  assign n1132 = n1131 ^ x428 ;
  assign n1133 = n1132 ^ x172 ;
  assign n1268 = n1267 ^ n1133 ;
  assign n1269 = n1268 ^ x427 ;
  assign n1273 = n1272 ^ n1269 ;
  assign n1277 = n1276 ^ n1273 ;
  assign n1364 = n1340 ^ n1277 ;
  assign n1355 = n1338 ^ n1269 ;
  assign n1227 = n1133 ^ x331 ;
  assign n1152 = x428 ^ x76 ;
  assign n1153 = n1152 ^ x268 ;
  assign n1154 = n1153 ^ x12 ;
  assign n1228 = n1227 ^ n1154 ;
  assign n1229 = n1228 ^ x267 ;
  assign n1356 = n1355 ^ n1229 ;
  assign n1360 = n1359 ^ n1356 ;
  assign n1365 = n1364 ^ n1360 ;
  assign n1369 = n1368 ^ n1365 ;
  assign n986 = n971 ^ n919 ;
  assign n889 = n825 ^ x462 ;
  assign n890 = n889 ^ n883 ;
  assign n891 = n890 ^ x398 ;
  assign n987 = n986 ^ n891 ;
  assign n991 = n990 ^ n987 ;
  assign n1073 = n1058 ^ n991 ;
  assign n961 = n955 ^ n891 ;
  assign n962 = n961 ^ n907 ;
  assign n963 = n962 ^ x493 ;
  assign n1074 = n1073 ^ n963 ;
  assign n1078 = n1077 ^ n1074 ;
  assign n1163 = n1145 ^ n1078 ;
  assign n1042 = n1002 ^ n963 ;
  assign n1034 = n955 ^ x397 ;
  assign n1035 = n1034 ^ n1028 ;
  assign n1036 = n1035 ^ x333 ;
  assign n1043 = n1042 ^ n1036 ;
  assign n1047 = n1046 ^ n1043 ;
  assign n1164 = n1163 ^ n1047 ;
  assign n1168 = n1167 ^ n1164 ;
  assign n1265 = n1247 ^ n1168 ;
  assign n1129 = n1089 ^ n1047 ;
  assign n1121 = n1036 ^ x492 ;
  assign n1122 = n1121 ^ n1102 ;
  assign n1123 = n1122 ^ x428 ;
  assign n1130 = n1129 ^ n1123 ;
  assign n1134 = n1133 ^ n1130 ;
  assign n1266 = n1265 ^ n1134 ;
  assign n1270 = n1269 ^ n1266 ;
  assign n1225 = n1182 ^ n1134 ;
  assign n1217 = n1174 ^ n1123 ;
  assign n1218 = n1217 ^ n1211 ;
  assign n1219 = n1218 ^ n1154 ;
  assign n1226 = n1225 ^ n1219 ;
  assign n1230 = n1229 ^ n1226 ;
  assign n1354 = n1270 ^ n1230 ;
  assign n1361 = n1360 ^ n1354 ;
  assign n1362 = n1361 ^ n1346 ;
  assign n985 = n977 ^ n921 ;
  assign n992 = n991 ^ n985 ;
  assign n996 = n995 ^ n992 ;
  assign n1072 = n1064 ^ n996 ;
  assign n1079 = n1078 ^ n1072 ;
  assign n1083 = n1082 ^ n1079 ;
  assign n1162 = n1151 ^ n1083 ;
  assign n1169 = n1168 ^ n1162 ;
  assign n1176 = n1175 ^ n1169 ;
  assign n1264 = n1253 ^ n1176 ;
  assign n1271 = n1270 ^ n1264 ;
  assign n1278 = n1277 ^ n1271 ;
  assign n1353 = n1352 ^ n1278 ;
  assign n1363 = n1362 ^ n1353 ;
  assign n1370 = n1369 ^ n1363 ;
  assign n43369 = n32533 ^ n1370 ;
  assign n2792 = n2788 ^ n1360 ;
  assign n1329 = n1229 ^ x426 ;
  assign n1254 = n1154 ^ x171 ;
  assign n1255 = n1254 ^ x363 ;
  assign n1256 = n1255 ^ x107 ;
  assign n1330 = n1329 ^ n1256 ;
  assign n1331 = n1330 ^ x362 ;
  assign n2793 = n2792 ^ n1331 ;
  assign n2797 = n2796 ^ n2793 ;
  assign n2790 = n2789 ^ n1362 ;
  assign n1327 = n1284 ^ n1230 ;
  assign n1319 = n1276 ^ n1219 ;
  assign n1320 = n1319 ^ n1313 ;
  assign n1321 = n1320 ^ n1256 ;
  assign n1328 = n1327 ^ n1321 ;
  assign n1332 = n1331 ^ n1328 ;
  assign n2791 = n2790 ^ n1332 ;
  assign n2798 = n2797 ^ n2791 ;
  assign n43370 = n43369 ^ n2798 ;
  assign n30641 = n21516 ^ n1369 ;
  assign n30642 = n30641 ^ n2797 ;
  assign n2814 = n1368 ^ x425 ;
  assign n2815 = n2814 ^ n2796 ;
  assign n2816 = n2815 ^ x361 ;
  assign n30643 = n30642 ^ n2816 ;
  assign n43371 = n43370 ^ n30643 ;
  assign n2640 = n2639 ^ n2504 ;
  assign n2538 = n2537 ^ x393 ;
  assign n1371 = x490 ^ x138 ;
  assign n1372 = n1371 ^ x330 ;
  assign n1373 = n1372 ^ x74 ;
  assign n2539 = n2538 ^ n1373 ;
  assign n2540 = n2539 ^ x329 ;
  assign n2641 = n2640 ^ n2540 ;
  assign n2642 = n2641 ^ n2618 ;
  assign n35055 = n32533 ^ n2642 ;
  assign n2801 = n2788 ^ x329 ;
  assign n1393 = x426 ^ x74 ;
  assign n1394 = n1393 ^ x266 ;
  assign n1395 = n1394 ^ x10 ;
  assign n2802 = n2801 ^ n1395 ;
  assign n2803 = n2802 ^ x265 ;
  assign n2799 = n2789 ^ n2540 ;
  assign n1391 = n1373 ^ n1284 ;
  assign n1392 = n1391 ^ n1368 ;
  assign n1396 = n1395 ^ n1392 ;
  assign n2800 = n2799 ^ n1396 ;
  assign n2804 = n2803 ^ n2800 ;
  assign n35056 = n35055 ^ n2804 ;
  assign n23470 = n21516 ^ n2618 ;
  assign n23471 = n23470 ^ n2803 ;
  assign n2549 = x425 ^ x73 ;
  assign n2550 = n2549 ^ x265 ;
  assign n2551 = n2550 ^ x9 ;
  assign n23472 = n23471 ^ n2551 ;
  assign n35057 = n35056 ^ n23472 ;
  assign n45292 = n43371 ^ n35057 ;
  assign n2806 = n2803 ^ n2797 ;
  assign n1443 = n1395 ^ n1331 ;
  assign n1380 = n1256 ^ x266 ;
  assign n1381 = n1380 ^ x458 ;
  assign n1382 = n1381 ^ x202 ;
  assign n1444 = n1443 ^ n1382 ;
  assign n1445 = n1444 ^ x457 ;
  assign n2807 = n2806 ^ n1445 ;
  assign n2811 = n2810 ^ n2807 ;
  assign n2805 = n2804 ^ n2798 ;
  assign n2812 = n2811 ^ n2805 ;
  assign n1441 = n1396 ^ n1332 ;
  assign n1433 = n1368 ^ n1321 ;
  assign n1434 = n1433 ^ n1427 ;
  assign n1435 = n1434 ^ n1382 ;
  assign n1442 = n1441 ^ n1435 ;
  assign n1446 = n1445 ^ n1442 ;
  assign n2813 = n2812 ^ n1446 ;
  assign n45293 = n45292 ^ n2813 ;
  assign n32971 = n30643 ^ n23472 ;
  assign n32972 = n32971 ^ n2811 ;
  assign n2859 = n2816 ^ n2551 ;
  assign n2860 = n2859 ^ n2810 ;
  assign n2861 = n2860 ^ x456 ;
  assign n32973 = n32972 ^ n2861 ;
  assign n45294 = n45293 ^ n32973 ;
  assign n2643 = n2642 ^ n2507 ;
  assign n2542 = n1373 ^ x233 ;
  assign n2543 = n2542 ^ x425 ;
  assign n2544 = n2543 ^ x169 ;
  assign n2541 = n2540 ^ x488 ;
  assign n2545 = n2544 ^ n2541 ;
  assign n2546 = n2545 ^ x424 ;
  assign n2644 = n2643 ^ n2546 ;
  assign n2645 = n2644 ^ n2621 ;
  assign n37044 = n35057 ^ n2645 ;
  assign n2825 = n2803 ^ x424 ;
  assign n2819 = n1395 ^ x169 ;
  assign n2820 = n2819 ^ x361 ;
  assign n2821 = n2820 ^ x105 ;
  assign n2826 = n2825 ^ n2821 ;
  assign n2827 = n2826 ^ x360 ;
  assign n2823 = n2804 ^ n2546 ;
  assign n2817 = n2544 ^ n1396 ;
  assign n2818 = n2817 ^ n2816 ;
  assign n2822 = n2821 ^ n2818 ;
  assign n2824 = n2823 ^ n2822 ;
  assign n2828 = n2827 ^ n2824 ;
  assign n37045 = n37044 ^ n2828 ;
  assign n25364 = n23472 ^ n2621 ;
  assign n25365 = n25364 ^ n2827 ;
  assign n2561 = n2551 ^ x168 ;
  assign n2562 = n2561 ^ x360 ;
  assign n2563 = n2562 ^ x104 ;
  assign n25366 = n25365 ^ n2563 ;
  assign n37046 = n37045 ^ n25366 ;
  assign n47395 = n45294 ^ n37046 ;
  assign n2852 = n2827 ^ n2811 ;
  assign n2844 = n2821 ^ n1445 ;
  assign n2839 = n1382 ^ x361 ;
  assign n2840 = n2839 ^ n2501 ;
  assign n2841 = n2840 ^ x297 ;
  assign n2845 = n2844 ^ n2841 ;
  assign n2849 = n2848 ^ n2845 ;
  assign n2853 = n2852 ^ n2849 ;
  assign n2857 = n2856 ^ n2853 ;
  assign n2831 = n2816 ^ n1435 ;
  assign n2838 = n2837 ^ n2831 ;
  assign n2842 = n2841 ^ n2838 ;
  assign n2830 = n2822 ^ n1446 ;
  assign n2843 = n2842 ^ n2830 ;
  assign n2850 = n2849 ^ n2843 ;
  assign n2829 = n2828 ^ n2813 ;
  assign n2851 = n2850 ^ n2829 ;
  assign n2858 = n2857 ^ n2851 ;
  assign n47396 = n47395 ^ n2858 ;
  assign n34059 = n32973 ^ n25366 ;
  assign n34060 = n34059 ^ n2857 ;
  assign n3107 = x456 ^ x104 ;
  assign n3108 = n3107 ^ x296 ;
  assign n3109 = n3108 ^ x40 ;
  assign n3105 = n2861 ^ n2563 ;
  assign n3106 = n3105 ^ n2856 ;
  assign n3110 = n3109 ^ n3106 ;
  assign n34061 = n34060 ^ n3110 ;
  assign n47397 = n47396 ^ n34061 ;
  assign n1865 = n1802 ^ x352 ;
  assign n1860 = x449 ^ x97 ;
  assign n1861 = n1860 ^ x289 ;
  assign n1862 = n1861 ^ x33 ;
  assign n1866 = n1865 ^ n1862 ;
  assign n1867 = n1866 ^ x288 ;
  assign n1853 = n1811 ^ x353 ;
  assign n1857 = n1856 ^ n1853 ;
  assign n1858 = n1857 ^ x289 ;
  assign n1789 = n1785 ^ x161 ;
  assign n1790 = n1789 ^ x353 ;
  assign n1791 = n1790 ^ x97 ;
  assign n1852 = n1826 ^ n1791 ;
  assign n1859 = n1858 ^ n1852 ;
  assign n1863 = n1862 ^ n1859 ;
  assign n1788 = n1787 ^ x416 ;
  assign n1792 = n1791 ^ n1788 ;
  assign n1793 = n1792 ^ x352 ;
  assign n1851 = n1850 ^ n1793 ;
  assign n1864 = n1863 ^ n1851 ;
  assign n1868 = n1867 ^ n1864 ;
  assign n40163 = n37704 ^ n1868 ;
  assign n3238 = n3200 ^ n1858 ;
  assign n3239 = n3238 ^ n2738 ;
  assign n3026 = n2998 ^ x289 ;
  assign n3027 = n3026 ^ x481 ;
  assign n3028 = n3027 ^ x225 ;
  assign n3240 = n3239 ^ n3028 ;
  assign n3237 = n3236 ^ n1863 ;
  assign n3241 = n3240 ^ n3237 ;
  assign n3025 = n3000 ^ n1862 ;
  assign n3029 = n3028 ^ n3025 ;
  assign n3030 = n3029 ^ x480 ;
  assign n3242 = n3241 ^ n3030 ;
  assign n40164 = n40163 ^ n3242 ;
  assign n3024 = n3002 ^ n1867 ;
  assign n3031 = n3030 ^ n3024 ;
  assign n1914 = n1883 ^ x288 ;
  assign n1915 = n1914 ^ x480 ;
  assign n1916 = n1915 ^ x224 ;
  assign n3032 = n3031 ^ n1916 ;
  assign n40165 = n40164 ^ n3032 ;
  assign n2779 = n2730 ^ x481 ;
  assign n2780 = n2779 ^ n1781 ;
  assign n2781 = n2780 ^ x417 ;
  assign n2777 = n2738 ^ n2731 ;
  assign n2761 = n2711 ^ x227 ;
  assign n2762 = n2761 ^ x419 ;
  assign n2763 = n2762 ^ x163 ;
  assign n2760 = n2713 ^ x482 ;
  assign n2764 = n2763 ^ n2760 ;
  assign n2765 = n2764 ^ x418 ;
  assign n2759 = n2736 ^ n2723 ;
  assign n2766 = n2765 ^ n2759 ;
  assign n2767 = n2766 ^ n1781 ;
  assign n2778 = n2777 ^ n2767 ;
  assign n2782 = n2781 ^ n2778 ;
  assign n1966 = x510 ^ x158 ;
  assign n1967 = n1966 ^ x350 ;
  assign n1968 = n1967 ^ x94 ;
  assign n2011 = n1968 ^ x253 ;
  assign n2012 = n2011 ^ x445 ;
  assign n2013 = n2012 ^ x189 ;
  assign n2068 = n2013 ^ x348 ;
  assign n2060 = x445 ^ x93 ;
  assign n2061 = n2060 ^ x285 ;
  assign n2062 = n2061 ^ x29 ;
  assign n2069 = n2068 ^ n2062 ;
  assign n2070 = n2069 ^ x284 ;
  assign n2128 = n2070 ^ x443 ;
  assign n2120 = n2062 ^ x188 ;
  assign n2121 = n2120 ^ x380 ;
  assign n2122 = n2121 ^ x124 ;
  assign n2129 = n2128 ^ n2122 ;
  assign n2130 = n2129 ^ x379 ;
  assign n2197 = n2130 ^ n1457 ;
  assign n2189 = n2122 ^ x283 ;
  assign n2190 = n2189 ^ x475 ;
  assign n2191 = n2190 ^ x219 ;
  assign n2198 = n2197 ^ n2191 ;
  assign n2199 = n2198 ^ x474 ;
  assign n2275 = n2199 ^ n1460 ;
  assign n2264 = n2191 ^ x378 ;
  assign n2265 = n2264 ^ n2258 ;
  assign n2266 = n2265 ^ x314 ;
  assign n2276 = n2275 ^ n2266 ;
  assign n2277 = n2276 ^ n2274 ;
  assign n2354 = n2277 ^ n1463 ;
  assign n2345 = n2266 ^ x473 ;
  assign n2346 = n2345 ^ n2339 ;
  assign n2347 = n2346 ^ x409 ;
  assign n2355 = n2354 ^ n2347 ;
  assign n2356 = n2355 ^ n2353 ;
  assign n1954 = x511 ^ x159 ;
  assign n1955 = n1954 ^ x351 ;
  assign n1956 = n1955 ^ x95 ;
  assign n1999 = n1956 ^ x254 ;
  assign n2000 = n1999 ^ x446 ;
  assign n2001 = n2000 ^ x190 ;
  assign n2053 = n2001 ^ x349 ;
  assign n2040 = x446 ^ x94 ;
  assign n2041 = n2040 ^ x286 ;
  assign n2042 = n2041 ^ x30 ;
  assign n2054 = n2053 ^ n2042 ;
  assign n2055 = n2054 ^ x285 ;
  assign n2113 = n2055 ^ x444 ;
  assign n2100 = n2042 ^ x189 ;
  assign n2101 = n2100 ^ x381 ;
  assign n2102 = n2101 ^ x125 ;
  assign n2114 = n2113 ^ n2102 ;
  assign n2115 = n2114 ^ x380 ;
  assign n2182 = n2154 ^ n2115 ;
  assign n2169 = n2102 ^ x284 ;
  assign n2170 = n2169 ^ x476 ;
  assign n2171 = n2170 ^ x220 ;
  assign n2183 = n2182 ^ n2171 ;
  assign n2184 = n2183 ^ x475 ;
  assign n2254 = n2223 ^ n2184 ;
  assign n2238 = n2171 ^ x379 ;
  assign n2073 = x476 ^ x124 ;
  assign n2074 = n2073 ^ x316 ;
  assign n2075 = n2074 ^ x60 ;
  assign n2239 = n2238 ^ n2075 ;
  assign n2240 = n2239 ^ x315 ;
  assign n2255 = n2254 ^ n2240 ;
  assign n2259 = n2258 ^ n2255 ;
  assign n2335 = n2304 ^ n2259 ;
  assign n2319 = n2240 ^ x474 ;
  assign n2133 = n2075 ^ x155 ;
  assign n2134 = n2133 ^ x411 ;
  assign n2135 = n2134 ^ x219 ;
  assign n2320 = n2319 ^ n2135 ;
  assign n2321 = n2320 ^ x410 ;
  assign n2336 = n2335 ^ n2321 ;
  assign n2340 = n2339 ^ n2336 ;
  assign n25882 = n2356 ^ n2340 ;
  assign n1019 = n943 ^ x398 ;
  assign n1020 = n1019 ^ n839 ;
  assign n1021 = n1020 ^ x334 ;
  assign n19559 = n1036 ^ n1021 ;
  assign n3244 = ~x30 & ~x31 ;
  assign n3245 = x29 & ~n3244 ;
  assign n3246 = x28 & n3245 ;
  assign n3247 = ~x27 & ~n3246 ;
  assign n3248 = ~x26 & n3247 ;
  assign n3249 = x25 & ~n3248 ;
  assign n3250 = ~x24 & ~n3249 ;
  assign n3251 = x23 & ~n3250 ;
  assign n3252 = x22 & n3251 ;
  assign n3253 = x21 & n3252 ;
  assign n3254 = ~x20 & ~n3253 ;
  assign n3255 = ~x19 & n3254 ;
  assign n3256 = x18 & ~n3255 ;
  assign n3257 = x17 & n3256 ;
  assign n3316 = n3257 ^ x16 ;
  assign n3260 = n3255 ^ x18 ;
  assign n3261 = n3254 ^ x19 ;
  assign n3262 = n3253 ^ x20 ;
  assign n3263 = n3248 ^ x25 ;
  assign n3264 = n3247 ^ x26 ;
  assign n3265 = n3246 ^ x27 ;
  assign n3266 = n3245 ^ x28 ;
  assign n3243 = x31 ^ x30 ;
  assign n3258 = ~x16 & ~n3257 ;
  assign n3267 = x15 & ~n3258 ;
  assign n3268 = x14 & n3267 ;
  assign n3269 = ~x13 & ~n3268 ;
  assign n3270 = x12 & ~n3269 ;
  assign n3271 = ~x11 & ~n3270 ;
  assign n3272 = ~x10 & n3271 ;
  assign n3273 = x9 & ~n3272 ;
  assign n3274 = ~x8 & ~n3273 ;
  assign n3275 = ~x7 & n3274 ;
  assign n3276 = ~x6 & n3275 ;
  assign n3277 = ~x5 & n3276 ;
  assign n3278 = ~x4 & n3277 ;
  assign n3279 = ~x3 & n3278 ;
  assign n3280 = x2 & ~n3279 ;
  assign n3281 = x1 & n3280 ;
  assign n3282 = n3281 ^ x0 ;
  assign n3283 = n3279 ^ x2 ;
  assign n3287 = n3280 ^ x1 ;
  assign n3292 = ~n3283 & n3287 ;
  assign n3284 = n3278 ^ x3 ;
  assign n3285 = n3283 & n3284 ;
  assign n3286 = n3285 ^ n3283 ;
  assign n3288 = n3287 ^ n3286 ;
  assign n3289 = n3288 ^ n3285 ;
  assign n3290 = ~n3288 & n3289 ;
  assign n3291 = n3290 ^ n3289 ;
  assign n3293 = n3292 ^ n3291 ;
  assign n3294 = n3282 & n3293 ;
  assign n3295 = x31 & n3294 ;
  assign n3296 = n3243 & n3295 ;
  assign n3297 = n3244 ^ x29 ;
  assign n3298 = n3296 & n3297 ;
  assign n3299 = n3266 & ~n3298 ;
  assign n3300 = n3265 & ~n3299 ;
  assign n3301 = ~n3264 & n3300 ;
  assign n3302 = n3263 & n3301 ;
  assign n3303 = n3249 ^ x24 ;
  assign n3304 = n3302 & n3303 ;
  assign n3305 = n3250 ^ x23 ;
  assign n3306 = n3304 & n3305 ;
  assign n3307 = n3251 ^ x22 ;
  assign n3308 = n3306 & ~n3307 ;
  assign n3309 = n3252 ^ x21 ;
  assign n3310 = n3308 & ~n3309 ;
  assign n3311 = n3262 & n3310 ;
  assign n3312 = ~n3261 & n3311 ;
  assign n3313 = ~n3260 & ~n3312 ;
  assign n3314 = n3256 ^ x17 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3350 = n3316 ^ n3315 ;
  assign n3319 = n3312 ^ n3260 ;
  assign n3320 = n3311 ^ n3261 ;
  assign n3321 = n3310 ^ n3262 ;
  assign n3322 = n3301 ^ n3263 ;
  assign n3323 = n3300 ^ n3264 ;
  assign n3324 = n3299 ^ n3265 ;
  assign n3325 = n3298 ^ n3266 ;
  assign n3326 = n3297 ^ n3296 ;
  assign n3327 = n3295 ^ n3243 ;
  assign n3328 = n3282 & ~n3291 ;
  assign n3329 = n3294 ^ x31 ;
  assign n3330 = n3328 & n3329 ;
  assign n3331 = n3327 & n3330 ;
  assign n3332 = ~n3326 & ~n3331 ;
  assign n3333 = ~n3325 & n3332 ;
  assign n3334 = n3324 & n3333 ;
  assign n3335 = ~n3323 & ~n3334 ;
  assign n3336 = ~n3322 & ~n3335 ;
  assign n3337 = n3303 ^ n3302 ;
  assign n3338 = ~n3336 & n3337 ;
  assign n3339 = n3305 ^ n3304 ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = n3307 ^ n3306 ;
  assign n3342 = ~n3340 & ~n3341 ;
  assign n3343 = n3309 ^ n3308 ;
  assign n3344 = ~n3342 & n3343 ;
  assign n3345 = ~n3321 & n3344 ;
  assign n3346 = ~n3320 & ~n3345 ;
  assign n3347 = n3319 & ~n3346 ;
  assign n3348 = n3314 ^ n3313 ;
  assign n3349 = n3347 & ~n3348 ;
  assign n3388 = n3350 ^ n3349 ;
  assign n3353 = n3348 ^ n3347 ;
  assign n3354 = n3346 ^ n3319 ;
  assign n3355 = n3345 ^ n3320 ;
  assign n3356 = n3344 ^ n3321 ;
  assign n3357 = n3335 ^ n3322 ;
  assign n3358 = n3334 ^ n3323 ;
  assign n3359 = n3333 ^ n3324 ;
  assign n3360 = n3292 ^ n3282 ;
  assign n3361 = n3277 ^ x4 ;
  assign n3362 = n3290 & n3361 ;
  assign n3363 = n3362 ^ n3289 ;
  assign n3364 = ~n3360 & n3363 ;
  assign n3365 = n3329 ^ n3328 ;
  assign n3366 = ~n3364 & ~n3365 ;
  assign n3367 = n3330 ^ n3327 ;
  assign n3368 = n3366 & ~n3367 ;
  assign n3369 = n3331 ^ n3326 ;
  assign n3370 = ~n3368 & ~n3369 ;
  assign n3371 = n3332 ^ n3325 ;
  assign n3372 = n3370 & n3371 ;
  assign n3373 = n3359 & ~n3372 ;
  assign n3374 = ~n3358 & n3373 ;
  assign n3375 = ~n3357 & ~n3374 ;
  assign n3376 = n3337 ^ n3336 ;
  assign n3377 = n3375 & ~n3376 ;
  assign n3378 = n3339 ^ n3338 ;
  assign n3379 = n3377 & ~n3378 ;
  assign n3380 = n3341 ^ n3340 ;
  assign n3381 = n3379 & n3380 ;
  assign n3382 = n3343 ^ n3342 ;
  assign n3383 = ~n3381 & ~n3382 ;
  assign n3384 = ~n3356 & n3383 ;
  assign n3385 = n3355 & ~n3384 ;
  assign n3386 = ~n3354 & ~n3385 ;
  assign n3387 = ~n3353 & n3386 ;
  assign n3391 = n3388 ^ n3387 ;
  assign n3392 = n3391 ^ x43 ;
  assign n3394 = n3382 ^ n3381 ;
  assign n3395 = n3394 ^ x48 ;
  assign n3397 = n3371 ^ n3370 ;
  assign n3398 = n3397 ^ x55 ;
  assign n3400 = n3365 ^ n3364 ;
  assign n3401 = n3400 ^ x58 ;
  assign n3402 = n3363 ^ n3360 ;
  assign n3403 = n3402 ^ x59 ;
  assign n3406 = n3284 & n3361 ;
  assign n3407 = n3406 ^ n3283 ;
  assign n3408 = n3407 ^ x61 ;
  assign n3409 = x63 & ~n3361 ;
  assign n3410 = n3409 ^ x62 ;
  assign n3411 = n3361 ^ n3284 ;
  assign n3412 = n3411 ^ n3409 ;
  assign n3413 = n3410 & ~n3412 ;
  assign n3414 = n3413 ^ x62 ;
  assign n3415 = n3414 ^ n3407 ;
  assign n3416 = n3408 & ~n3415 ;
  assign n3417 = n3416 ^ x61 ;
  assign n3404 = n3285 & ~n3361 ;
  assign n3405 = n3404 ^ n3288 ;
  assign n3418 = n3417 ^ n3405 ;
  assign n3717 = n3405 ^ x60 ;
  assign n3422 = ~n3418 & n3717 ;
  assign n3419 = n3402 ^ x60 ;
  assign n3423 = n3422 ^ n3419 ;
  assign n3424 = n3403 & ~n3423 ;
  assign n3425 = n3424 ^ x59 ;
  assign n3426 = n3425 ^ n3400 ;
  assign n3427 = n3401 & ~n3426 ;
  assign n3428 = n3427 ^ x58 ;
  assign n3399 = n3367 ^ n3366 ;
  assign n3429 = n3428 ^ n3399 ;
  assign n3430 = n3369 ^ n3368 ;
  assign n3431 = n3430 ^ x57 ;
  assign n3432 = n3431 ^ n3399 ;
  assign n3433 = n3432 ^ n3430 ;
  assign n3434 = n3429 & ~n3433 ;
  assign n3435 = n3434 ^ n3431 ;
  assign n3437 = n3397 ^ x56 ;
  assign n3436 = n3430 ^ n3397 ;
  assign n3438 = n3437 ^ n3436 ;
  assign n3439 = n3435 & ~n3438 ;
  assign n3440 = n3439 ^ n3437 ;
  assign n3441 = ~n3398 & n3440 ;
  assign n3442 = n3441 ^ x55 ;
  assign n3396 = n3372 ^ n3359 ;
  assign n3443 = n3442 ^ n3396 ;
  assign n3444 = n3373 ^ n3358 ;
  assign n3445 = n3444 ^ x54 ;
  assign n3446 = n3445 ^ n3396 ;
  assign n3447 = n3446 ^ n3444 ;
  assign n3448 = n3443 & ~n3447 ;
  assign n3449 = n3448 ^ n3445 ;
  assign n3450 = n3374 ^ n3357 ;
  assign n3452 = n3450 ^ x53 ;
  assign n3451 = n3450 ^ n3444 ;
  assign n3453 = n3452 ^ n3451 ;
  assign n3454 = n3449 & ~n3453 ;
  assign n3455 = n3454 ^ n3452 ;
  assign n3456 = n3376 ^ n3375 ;
  assign n3458 = n3456 ^ x52 ;
  assign n3457 = n3456 ^ n3450 ;
  assign n3459 = n3458 ^ n3457 ;
  assign n3460 = n3455 & ~n3459 ;
  assign n3461 = n3460 ^ n3458 ;
  assign n3462 = n3378 ^ n3377 ;
  assign n3464 = n3462 ^ x51 ;
  assign n3463 = n3462 ^ n3456 ;
  assign n3465 = n3464 ^ n3463 ;
  assign n3466 = ~n3461 & n3465 ;
  assign n3467 = n3466 ^ n3464 ;
  assign n3468 = n3380 ^ n3379 ;
  assign n3470 = n3468 ^ x50 ;
  assign n3469 = n3468 ^ n3462 ;
  assign n3471 = n3470 ^ n3469 ;
  assign n3472 = ~n3467 & n3471 ;
  assign n3473 = n3472 ^ n3470 ;
  assign n3475 = n3394 ^ x49 ;
  assign n3474 = n3468 ^ n3394 ;
  assign n3476 = n3475 ^ n3474 ;
  assign n3477 = n3473 & ~n3476 ;
  assign n3478 = n3477 ^ n3475 ;
  assign n3479 = n3395 & ~n3478 ;
  assign n3480 = n3479 ^ x48 ;
  assign n3393 = n3383 ^ n3356 ;
  assign n3481 = n3480 ^ n3393 ;
  assign n3695 = n3393 ^ x47 ;
  assign n3486 = n3481 & ~n3695 ;
  assign n3482 = n3384 ^ n3355 ;
  assign n3483 = n3482 ^ x47 ;
  assign n3487 = n3486 ^ n3483 ;
  assign n3488 = n3385 ^ n3354 ;
  assign n3490 = n3488 ^ x46 ;
  assign n3489 = n3488 ^ n3482 ;
  assign n3491 = n3490 ^ n3489 ;
  assign n3492 = ~n3487 & n3491 ;
  assign n3493 = n3492 ^ n3490 ;
  assign n3494 = n3386 ^ n3353 ;
  assign n3496 = n3494 ^ x45 ;
  assign n3495 = n3494 ^ n3488 ;
  assign n3497 = n3496 ^ n3495 ;
  assign n3498 = ~n3493 & n3497 ;
  assign n3499 = n3498 ^ n3496 ;
  assign n3501 = n3391 ^ x44 ;
  assign n3500 = n3494 ^ n3391 ;
  assign n3502 = n3501 ^ n3500 ;
  assign n3503 = n3499 & ~n3502 ;
  assign n3504 = n3503 ^ n3501 ;
  assign n3505 = n3392 & ~n3504 ;
  assign n3506 = n3505 ^ x43 ;
  assign n3389 = n3387 & n3388 ;
  assign n3351 = ~n3349 & n3350 ;
  assign n3317 = n3315 & n3316 ;
  assign n3259 = n3258 ^ x15 ;
  assign n3318 = n3317 ^ n3259 ;
  assign n3352 = n3351 ^ n3318 ;
  assign n3390 = n3389 ^ n3352 ;
  assign n3507 = n3506 ^ n3390 ;
  assign n3513 = ~n3352 & n3389 ;
  assign n3511 = n3318 & n3351 ;
  assign n3509 = n3259 & n3317 ;
  assign n3508 = n3267 ^ x14 ;
  assign n3510 = n3509 ^ n3508 ;
  assign n3512 = n3511 ^ n3510 ;
  assign n3514 = n3513 ^ n3512 ;
  assign n3515 = n3514 ^ x42 ;
  assign n3516 = n3515 ^ n3390 ;
  assign n3517 = n3516 ^ n3514 ;
  assign n3518 = n3507 & ~n3517 ;
  assign n3519 = n3518 ^ n3515 ;
  assign n3525 = ~n3512 & n3513 ;
  assign n3523 = n3510 & ~n3511 ;
  assign n3521 = ~n3508 & n3509 ;
  assign n3520 = n3268 ^ x13 ;
  assign n3522 = n3521 ^ n3520 ;
  assign n3524 = n3523 ^ n3522 ;
  assign n3526 = n3525 ^ n3524 ;
  assign n3528 = n3526 ^ x41 ;
  assign n3527 = n3526 ^ n3514 ;
  assign n3529 = n3528 ^ n3527 ;
  assign n3530 = n3519 & ~n3529 ;
  assign n3531 = n3530 ^ n3528 ;
  assign n3537 = n3524 & ~n3525 ;
  assign n3535 = ~n3522 & n3523 ;
  assign n3533 = n3520 & n3521 ;
  assign n3532 = n3269 ^ x12 ;
  assign n3534 = n3533 ^ n3532 ;
  assign n3536 = n3535 ^ n3534 ;
  assign n3538 = n3537 ^ n3536 ;
  assign n3540 = n3538 ^ x40 ;
  assign n3539 = n3538 ^ n3526 ;
  assign n3541 = n3540 ^ n3539 ;
  assign n3542 = ~n3531 & n3541 ;
  assign n3543 = n3542 ^ n3540 ;
  assign n3549 = ~n3536 & ~n3537 ;
  assign n3547 = ~n3534 & n3535 ;
  assign n3545 = n3532 & n3533 ;
  assign n3544 = n3270 ^ x11 ;
  assign n3546 = n3545 ^ n3544 ;
  assign n3548 = n3547 ^ n3546 ;
  assign n3550 = n3549 ^ n3548 ;
  assign n3552 = n3550 ^ x39 ;
  assign n3551 = n3550 ^ n3538 ;
  assign n3553 = n3552 ^ n3551 ;
  assign n3554 = ~n3543 & n3553 ;
  assign n3555 = n3554 ^ n3552 ;
  assign n3561 = n3548 & ~n3549 ;
  assign n3559 = ~n3546 & n3547 ;
  assign n3557 = n3544 & n3545 ;
  assign n3556 = n3271 ^ x10 ;
  assign n3558 = n3557 ^ n3556 ;
  assign n3560 = n3559 ^ n3558 ;
  assign n3562 = n3561 ^ n3560 ;
  assign n3564 = n3562 ^ x38 ;
  assign n3563 = n3562 ^ n3550 ;
  assign n3565 = n3564 ^ n3563 ;
  assign n3566 = ~n3555 & n3565 ;
  assign n3567 = n3566 ^ n3564 ;
  assign n3573 = ~n3560 & ~n3561 ;
  assign n3571 = ~n3558 & n3559 ;
  assign n3569 = n3556 & ~n3557 ;
  assign n3568 = n3272 ^ x9 ;
  assign n3570 = n3569 ^ n3568 ;
  assign n3572 = n3571 ^ n3570 ;
  assign n3574 = n3573 ^ n3572 ;
  assign n3576 = n3574 ^ x37 ;
  assign n3575 = n3574 ^ n3562 ;
  assign n3577 = n3576 ^ n3575 ;
  assign n3578 = ~n3567 & n3577 ;
  assign n3579 = n3578 ^ n3576 ;
  assign n3610 = n3579 ^ x36 ;
  assign n4078 = n3610 ^ x95 ;
  assign n3714 = n3414 ^ x61 ;
  assign n3715 = n3714 ^ n3407 ;
  assign n4541 = n3715 ^ n3297 ;
  assign n4542 = n4078 & ~n4541 ;
  assign n4543 = n4542 ^ n3297 ;
  assign n3676 = n3411 ^ n3410 ;
  assign n3666 = n3361 ^ x63 ;
  assign n3667 = n3666 ^ n3264 ;
  assign n3633 = n3276 ^ x5 ;
  assign n3634 = n3633 ^ x32 ;
  assign n3617 = n3275 ^ x6 ;
  assign n3581 = n3568 & ~n3569 ;
  assign n3580 = n3273 ^ x8 ;
  assign n3582 = n3581 ^ n3580 ;
  assign n3583 = n3570 & n3571 ;
  assign n3595 = n3582 & ~n3583 ;
  assign n3594 = n3274 ^ x7 ;
  assign n3596 = n3595 ^ n3594 ;
  assign n3597 = n3580 & n3581 ;
  assign n3598 = n3597 ^ n3596 ;
  assign n3614 = n3598 ^ n3594 ;
  assign n3615 = n3596 & ~n3614 ;
  assign n3584 = n3583 ^ n3582 ;
  assign n3585 = ~n3572 & ~n3573 ;
  assign n3599 = ~n3584 & n3585 ;
  assign n3613 = ~n3598 & ~n3599 ;
  assign n3616 = n3615 ^ n3613 ;
  assign n3618 = n3617 ^ n3616 ;
  assign n3586 = n3585 ^ n3584 ;
  assign n3588 = n3586 ^ x36 ;
  assign n3587 = n3586 ^ n3574 ;
  assign n3589 = n3588 ^ n3587 ;
  assign n3590 = n3579 & ~n3589 ;
  assign n3591 = n3590 ^ n3588 ;
  assign n3600 = n3599 ^ n3598 ;
  assign n3602 = n3600 ^ x35 ;
  assign n3601 = n3600 ^ n3586 ;
  assign n3603 = n3602 ^ n3601 ;
  assign n3604 = ~n3591 & n3603 ;
  assign n3605 = n3604 ^ n3602 ;
  assign n3620 = n3618 ^ x34 ;
  assign n3619 = n3618 ^ n3600 ;
  assign n3621 = n3620 ^ n3619 ;
  assign n3622 = ~n3605 & n3621 ;
  assign n3623 = n3622 ^ n3620 ;
  assign n3631 = n3623 ^ n3617 ;
  assign n3632 = ~n3618 & ~n3631 ;
  assign n3635 = n3634 ^ n3632 ;
  assign n3630 = x33 & ~n3623 ;
  assign n3636 = n3635 ^ n3630 ;
  assign n3624 = n3623 ^ x33 ;
  assign n3592 = n3591 ^ x35 ;
  assign n3593 = n3243 & n3592 ;
  assign n3606 = n3605 ^ x34 ;
  assign n3625 = n3593 & n3606 ;
  assign n3637 = ~n3624 & n3625 ;
  assign n3665 = ~n3636 & n3637 ;
  assign n3677 = n3666 ^ n3665 ;
  assign n3678 = n3667 & n3677 ;
  assign n3679 = n3678 ^ n3264 ;
  assign n3713 = ~n3676 & n3679 ;
  assign n3716 = n3713 & ~n3715 ;
  assign n3718 = n3717 ^ n3417 ;
  assign n3719 = ~n3716 & n3718 ;
  assign n3712 = n3423 ^ x59 ;
  assign n3720 = n3719 ^ n3712 ;
  assign n3721 = n3719 ^ n3307 ;
  assign n3722 = ~n3720 & ~n3721 ;
  assign n3723 = n3722 ^ n3307 ;
  assign n3710 = n3425 ^ x58 ;
  assign n3711 = n3710 ^ n3400 ;
  assign n3752 = n3723 ^ n3711 ;
  assign n3668 = n3667 ^ n3665 ;
  assign n3638 = n3637 ^ n3636 ;
  assign n3626 = n3625 ^ n3624 ;
  assign n3607 = n3606 ^ n3593 ;
  assign n3608 = n3592 ^ n3243 ;
  assign n3627 = ~n3607 & ~n3608 ;
  assign n3639 = n3626 & n3627 ;
  assign n3669 = n3638 & n3639 ;
  assign n3675 = ~n3668 & n3669 ;
  assign n3680 = n3679 ^ n3676 ;
  assign n3753 = n3675 & ~n3680 ;
  assign n3754 = n3715 ^ n3713 ;
  assign n3755 = n3753 & ~n3754 ;
  assign n3756 = n3718 ^ n3716 ;
  assign n3757 = ~n3755 & ~n3756 ;
  assign n3758 = n3712 ^ n3307 ;
  assign n3759 = n3758 ^ n3719 ;
  assign n3760 = n3757 & ~n3759 ;
  assign n3761 = n3752 & ~n3760 ;
  assign n3724 = n3711 & ~n3723 ;
  assign n3708 = n3428 ^ x57 ;
  assign n3709 = n3708 ^ n3399 ;
  assign n3762 = n3724 ^ n3709 ;
  assign n3763 = n3761 & ~n3762 ;
  assign n3725 = n3709 & ~n3724 ;
  assign n3707 = n3435 ^ x56 ;
  assign n3764 = n3725 ^ n3707 ;
  assign n3765 = n3763 & ~n3764 ;
  assign n3726 = ~n3707 & ~n3725 ;
  assign n3689 = n3440 ^ x55 ;
  assign n3706 = n3689 ^ n3260 ;
  assign n3751 = n3726 ^ n3706 ;
  assign n3795 = n3765 ^ n3751 ;
  assign n3796 = n3760 ^ n3752 ;
  assign n3670 = n3669 ^ n3668 ;
  assign n3609 = n3608 ^ n3607 ;
  assign n3611 = ~n3608 & ~n3610 ;
  assign n3612 = ~n3609 & n3611 ;
  assign n3628 = n3627 ^ n3626 ;
  assign n3629 = ~n3612 & n3628 ;
  assign n3640 = n3639 ^ n3638 ;
  assign n3671 = n3629 & n3640 ;
  assign n3674 = n3670 & ~n3671 ;
  assign n3681 = n3680 ^ n3675 ;
  assign n3797 = n3674 & n3681 ;
  assign n3798 = n3754 ^ n3753 ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = n3756 ^ n3755 ;
  assign n3801 = n3799 & ~n3800 ;
  assign n3802 = n3759 ^ n3757 ;
  assign n3803 = ~n3801 & ~n3802 ;
  assign n3804 = n3796 & n3803 ;
  assign n3805 = n3762 ^ n3761 ;
  assign n3806 = ~n3804 & ~n3805 ;
  assign n3807 = n3764 ^ n3763 ;
  assign n3808 = n3806 & ~n3807 ;
  assign n3809 = ~n3795 & n3808 ;
  assign n3727 = n3726 ^ n3689 ;
  assign n3728 = ~n3706 & n3727 ;
  assign n3729 = n3728 ^ n3260 ;
  assign n3704 = n3442 ^ x54 ;
  assign n3705 = n3704 ^ n3396 ;
  assign n3767 = n3729 ^ n3705 ;
  assign n3766 = ~n3751 & ~n3765 ;
  assign n3810 = n3767 ^ n3766 ;
  assign n3811 = n3809 & n3810 ;
  assign n3768 = ~n3766 & ~n3767 ;
  assign n3730 = n3705 & ~n3729 ;
  assign n3703 = n3449 ^ x53 ;
  assign n3750 = n3730 ^ n3703 ;
  assign n3794 = n3768 ^ n3750 ;
  assign n3834 = n3811 ^ n3794 ;
  assign n3835 = n3834 ^ x80 ;
  assign n3672 = n3671 ^ n3670 ;
  assign n3641 = n3640 ^ n3629 ;
  assign n3642 = n3641 ^ x91 ;
  assign n3644 = n3610 ^ n3608 ;
  assign n3643 = x95 & n3610 ;
  assign n3645 = n3644 ^ n3643 ;
  assign n4073 = n3643 ^ x94 ;
  assign n3650 = ~n3645 & n4073 ;
  assign n3646 = n3611 ^ n3609 ;
  assign n3647 = n3646 ^ x94 ;
  assign n3651 = n3650 ^ n3647 ;
  assign n3652 = n3628 ^ n3612 ;
  assign n3654 = n3652 ^ x93 ;
  assign n3653 = n3652 ^ n3646 ;
  assign n3655 = n3654 ^ n3653 ;
  assign n3656 = n3651 & ~n3655 ;
  assign n3657 = n3656 ^ n3654 ;
  assign n3659 = n3641 ^ x92 ;
  assign n3658 = n3652 ^ n3641 ;
  assign n3660 = n3659 ^ n3658 ;
  assign n3661 = ~n3657 & n3660 ;
  assign n3662 = n3661 ^ n3659 ;
  assign n3663 = ~n3642 & n3662 ;
  assign n3664 = n3663 ^ x91 ;
  assign n3673 = n3672 ^ n3664 ;
  assign n3988 = n3664 ^ x90 ;
  assign n3686 = n3673 & n3988 ;
  assign n3682 = n3681 ^ n3674 ;
  assign n3683 = n3682 ^ x90 ;
  assign n3687 = n3686 ^ n3683 ;
  assign n3836 = n3798 ^ n3797 ;
  assign n3838 = n3836 ^ x89 ;
  assign n3837 = n3836 ^ n3682 ;
  assign n3839 = n3838 ^ n3837 ;
  assign n3840 = ~n3687 & n3839 ;
  assign n3841 = n3840 ^ n3838 ;
  assign n3842 = n3800 ^ n3799 ;
  assign n3844 = n3842 ^ x88 ;
  assign n3843 = n3842 ^ n3836 ;
  assign n3845 = n3844 ^ n3843 ;
  assign n3846 = n3841 & ~n3845 ;
  assign n3847 = n3846 ^ n3844 ;
  assign n3848 = n3802 ^ n3801 ;
  assign n3850 = n3848 ^ x87 ;
  assign n3849 = n3848 ^ n3842 ;
  assign n3851 = n3850 ^ n3849 ;
  assign n3852 = ~n3847 & n3851 ;
  assign n3853 = n3852 ^ n3850 ;
  assign n3854 = n3803 ^ n3796 ;
  assign n3856 = n3854 ^ x86 ;
  assign n3855 = n3854 ^ n3848 ;
  assign n3857 = n3856 ^ n3855 ;
  assign n3858 = ~n3853 & n3857 ;
  assign n3859 = n3858 ^ n3856 ;
  assign n3860 = n3805 ^ n3804 ;
  assign n3862 = n3860 ^ x85 ;
  assign n3861 = n3860 ^ n3854 ;
  assign n3863 = n3862 ^ n3861 ;
  assign n3864 = ~n3859 & n3863 ;
  assign n3865 = n3864 ^ n3862 ;
  assign n3866 = n3807 ^ n3806 ;
  assign n3868 = n3866 ^ x84 ;
  assign n3867 = n3866 ^ n3860 ;
  assign n3869 = n3868 ^ n3867 ;
  assign n3870 = n3865 & ~n3869 ;
  assign n3871 = n3870 ^ n3868 ;
  assign n3872 = n3808 ^ n3795 ;
  assign n3874 = n3872 ^ x83 ;
  assign n3873 = n3872 ^ n3866 ;
  assign n3875 = n3874 ^ n3873 ;
  assign n3876 = ~n3871 & n3875 ;
  assign n3877 = n3876 ^ n3874 ;
  assign n3878 = n3810 ^ n3809 ;
  assign n3880 = n3878 ^ x82 ;
  assign n3879 = n3878 ^ n3872 ;
  assign n3881 = n3880 ^ n3879 ;
  assign n3882 = ~n3877 & n3881 ;
  assign n3883 = n3882 ^ n3880 ;
  assign n3885 = n3834 ^ x81 ;
  assign n3884 = n3878 ^ n3834 ;
  assign n3886 = n3885 ^ n3884 ;
  assign n3887 = n3883 & ~n3886 ;
  assign n3888 = n3887 ^ n3885 ;
  assign n3889 = ~n3835 & n3888 ;
  assign n3890 = n3889 ^ x80 ;
  assign n3812 = n3794 & ~n3811 ;
  assign n3769 = ~n3750 & n3768 ;
  assign n3731 = ~n3703 & ~n3730 ;
  assign n3702 = n3455 ^ x52 ;
  assign n3749 = n3731 ^ n3702 ;
  assign n3793 = n3769 ^ n3749 ;
  assign n3833 = n3812 ^ n3793 ;
  assign n3891 = n3890 ^ n3833 ;
  assign n4030 = n3833 ^ x79 ;
  assign n3896 = n3891 & ~n4030 ;
  assign n3813 = ~n3793 & n3812 ;
  assign n3701 = n3461 ^ x51 ;
  assign n3771 = n3701 ^ n3508 ;
  assign n3732 = n3702 & ~n3731 ;
  assign n3772 = n3771 ^ n3732 ;
  assign n3770 = n3749 & ~n3769 ;
  assign n3792 = n3772 ^ n3770 ;
  assign n3892 = n3813 ^ n3792 ;
  assign n3893 = n3892 ^ x79 ;
  assign n3897 = n3896 ^ n3893 ;
  assign n3773 = ~n3770 & ~n3772 ;
  assign n3733 = n3732 ^ n3701 ;
  assign n3734 = n3732 ^ n3508 ;
  assign n3735 = n3733 & n3734 ;
  assign n3736 = n3735 ^ n3508 ;
  assign n3700 = n3467 ^ x50 ;
  assign n3748 = n3736 ^ n3700 ;
  assign n3815 = n3773 ^ n3748 ;
  assign n3814 = n3792 & ~n3813 ;
  assign n3898 = n3815 ^ n3814 ;
  assign n3900 = n3898 ^ x78 ;
  assign n3899 = n3898 ^ n3892 ;
  assign n3901 = n3900 ^ n3899 ;
  assign n3902 = ~n3897 & n3901 ;
  assign n3903 = n3902 ^ n3900 ;
  assign n4024 = n3903 ^ x77 ;
  assign n3971 = n3531 ^ x40 ;
  assign n4023 = ~n3617 & n3971 ;
  assign n4025 = n4024 ^ n4023 ;
  assign n4027 = n3897 ^ x78 ;
  assign n4194 = n4027 ^ n4023 ;
  assign n3952 = n3519 ^ x41 ;
  assign n4026 = ~n3594 & ~n3952 ;
  assign n4028 = n4027 ^ n4026 ;
  assign n4031 = n4030 ^ n3890 ;
  assign n3941 = n3506 ^ x42 ;
  assign n3942 = n3941 ^ n3390 ;
  assign n4029 = ~n3580 & ~n3942 ;
  assign n4032 = n4031 ^ n4029 ;
  assign n4034 = n3888 ^ x80 ;
  assign n3787 = n3504 ^ x43 ;
  assign n4033 = n3568 & n3787 ;
  assign n4035 = n4034 ^ n4033 ;
  assign n4037 = n3883 ^ x81 ;
  assign n4185 = n4037 ^ n4033 ;
  assign n3693 = n3499 ^ x44 ;
  assign n4036 = n3556 & ~n3693 ;
  assign n4038 = n4037 ^ n4036 ;
  assign n4040 = n3877 ^ x82 ;
  assign n3694 = n3493 ^ x45 ;
  assign n4039 = ~n3544 & n3694 ;
  assign n4041 = n4040 ^ n4039 ;
  assign n4043 = n3871 ^ x83 ;
  assign n3743 = n3487 ^ x46 ;
  assign n4042 = ~n3532 & n3743 ;
  assign n4044 = n4043 ^ n4042 ;
  assign n4046 = n3865 ^ x84 ;
  assign n3696 = n3695 ^ n3480 ;
  assign n4045 = n3520 & ~n3696 ;
  assign n4047 = n4046 ^ n4045 ;
  assign n4049 = n3859 ^ x85 ;
  assign n3698 = n3478 ^ x48 ;
  assign n4048 = n3508 & n3698 ;
  assign n4050 = n4049 ^ n4048 ;
  assign n4052 = n3853 ^ x86 ;
  assign n3699 = n3473 ^ x49 ;
  assign n4051 = n3259 & ~n3699 ;
  assign n4053 = n4052 ^ n4051 ;
  assign n4055 = n3847 ^ x87 ;
  assign n4054 = ~n3316 & n3700 ;
  assign n4056 = n4055 ^ n4054 ;
  assign n4058 = n3841 ^ x88 ;
  assign n4057 = n3314 & n3701 ;
  assign n4059 = n4058 ^ n4057 ;
  assign n4060 = n3260 & ~n3702 ;
  assign n3688 = n3687 ^ x89 ;
  assign n4061 = n4060 ^ n3688 ;
  assign n4062 = n3261 & ~n3703 ;
  assign n3989 = n3988 ^ n3672 ;
  assign n4063 = n4062 ^ n3989 ;
  assign n4065 = ~n3262 & ~n3705 ;
  assign n4064 = n3662 ^ x91 ;
  assign n4066 = n4065 ^ n4064 ;
  assign n4068 = n3657 ^ x92 ;
  assign n4067 = n3309 & ~n3689 ;
  assign n4069 = n4068 ^ n4067 ;
  assign n4071 = n3651 ^ x93 ;
  assign n4070 = ~n3307 & ~n3707 ;
  assign n4072 = n4071 ^ n4070 ;
  assign n4075 = n3305 & ~n3709 ;
  assign n4074 = n4073 ^ n3644 ;
  assign n4076 = n4075 ^ n4074 ;
  assign n4077 = ~n3303 & n3711 ;
  assign n4079 = n4078 ^ n4077 ;
  assign n3697 = n3696 ^ n3556 ;
  assign n3737 = n3700 & ~n3736 ;
  assign n3738 = ~n3699 & n3737 ;
  assign n3739 = ~n3698 & ~n3738 ;
  assign n3740 = n3739 ^ n3696 ;
  assign n3741 = n3697 & ~n3740 ;
  assign n3742 = n3741 ^ n3556 ;
  assign n3744 = n3742 & ~n3743 ;
  assign n3745 = ~n3694 & n3744 ;
  assign n3785 = n3693 & n3745 ;
  assign n3786 = n3785 ^ n3617 ;
  assign n3938 = n3787 ^ n3785 ;
  assign n3939 = n3786 & n3938 ;
  assign n3940 = n3939 ^ n3617 ;
  assign n3953 = ~n3940 & ~n3942 ;
  assign n3972 = n3952 & ~n3953 ;
  assign n4084 = ~n3971 & n3972 ;
  assign n4019 = n3543 ^ x39 ;
  assign n4085 = n4084 ^ n4019 ;
  assign n4015 = n3555 ^ x38 ;
  assign n4086 = n4015 ^ n3283 ;
  assign n4087 = n4086 ^ n4084 ;
  assign n4088 = n4087 ^ n4015 ;
  assign n4089 = n4085 & ~n4088 ;
  assign n4090 = n4089 ^ n4086 ;
  assign n3973 = n3972 ^ n3971 ;
  assign n3954 = n3953 ^ n3952 ;
  assign n3746 = n3745 ^ n3693 ;
  assign n3747 = n3739 ^ n3697 ;
  assign n3774 = ~n3748 & ~n3773 ;
  assign n3775 = n3737 ^ n3699 ;
  assign n3776 = ~n3774 & n3775 ;
  assign n3777 = n3738 ^ n3698 ;
  assign n3778 = n3776 & n3777 ;
  assign n3779 = n3747 & n3778 ;
  assign n3780 = n3743 ^ n3742 ;
  assign n3781 = ~n3779 & n3780 ;
  assign n3782 = n3744 ^ n3694 ;
  assign n3783 = ~n3781 & ~n3782 ;
  assign n3784 = ~n3746 & ~n3783 ;
  assign n3788 = n3787 ^ n3786 ;
  assign n3937 = n3784 & n3788 ;
  assign n3943 = n3942 ^ n3940 ;
  assign n3955 = n3937 & n3943 ;
  assign n3974 = ~n3954 & ~n3955 ;
  assign n4082 = ~n3973 & n3974 ;
  assign n4091 = n4019 ^ n3283 ;
  assign n4092 = n4091 ^ n4084 ;
  assign n4115 = ~n4082 & ~n4092 ;
  assign n4119 = ~n4090 & n4115 ;
  assign n3975 = n3974 ^ n3973 ;
  assign n3956 = n3955 ^ n3954 ;
  assign n3944 = n3943 ^ n3937 ;
  assign n3789 = n3788 ^ n3784 ;
  assign n3790 = n3782 ^ n3781 ;
  assign n3791 = n3778 ^ n3747 ;
  assign n3816 = ~n3814 & n3815 ;
  assign n3817 = n3775 ^ n3774 ;
  assign n3818 = n3816 & n3817 ;
  assign n3819 = n3777 ^ n3776 ;
  assign n3820 = n3818 & ~n3819 ;
  assign n3821 = ~n3791 & n3820 ;
  assign n3822 = n3780 ^ n3779 ;
  assign n3823 = n3821 & ~n3822 ;
  assign n3824 = n3790 & ~n3823 ;
  assign n3825 = n3783 ^ n3746 ;
  assign n3826 = ~n3824 & n3825 ;
  assign n3945 = ~n3789 & ~n3826 ;
  assign n3957 = n3944 & ~n3945 ;
  assign n3976 = n3956 & ~n3957 ;
  assign n4081 = ~n3975 & n3976 ;
  assign n4083 = n4082 ^ n4081 ;
  assign n4093 = n4092 ^ n4090 ;
  assign n4094 = n4093 ^ n4081 ;
  assign n4095 = n4094 ^ n4090 ;
  assign n4096 = ~n4083 & n4095 ;
  assign n4097 = n4096 ^ n4093 ;
  assign n4116 = n4115 ^ n4015 ;
  assign n4117 = ~n4097 & ~n4116 ;
  assign n4113 = x65 ^ x64 ;
  assign n4010 = n3567 ^ x37 ;
  assign n4114 = n4113 ^ n4010 ;
  assign n4118 = n4117 ^ n4114 ;
  assign n4120 = n4119 ^ n4118 ;
  assign n4098 = n4097 ^ x65 ;
  assign n3977 = n3976 ^ n3975 ;
  assign n3828 = n3825 ^ n3824 ;
  assign n3829 = n3828 ^ x71 ;
  assign n3911 = n3819 ^ n3818 ;
  assign n3831 = n3817 ^ n3816 ;
  assign n3832 = n3831 ^ x76 ;
  assign n3905 = n3831 ^ x77 ;
  assign n3904 = n3898 ^ n3831 ;
  assign n3906 = n3905 ^ n3904 ;
  assign n3907 = n3903 & ~n3906 ;
  assign n3908 = n3907 ^ n3905 ;
  assign n3909 = n3832 & ~n3908 ;
  assign n3910 = n3909 ^ x76 ;
  assign n3912 = n3911 ^ n3910 ;
  assign n3913 = n3911 ^ x75 ;
  assign n3914 = n3912 & ~n3913 ;
  assign n3915 = n3914 ^ x75 ;
  assign n3830 = n3820 ^ n3791 ;
  assign n3916 = n3915 ^ n3830 ;
  assign n4012 = n3830 ^ x74 ;
  assign n3921 = n3916 & ~n4012 ;
  assign n3917 = n3822 ^ n3821 ;
  assign n3918 = n3917 ^ x74 ;
  assign n3922 = n3921 ^ n3918 ;
  assign n3923 = n3823 ^ n3790 ;
  assign n3925 = n3923 ^ x73 ;
  assign n3924 = n3923 ^ n3917 ;
  assign n3926 = n3925 ^ n3924 ;
  assign n3927 = n3922 & ~n3926 ;
  assign n3928 = n3927 ^ n3925 ;
  assign n3930 = n3828 ^ x72 ;
  assign n3929 = n3923 ^ n3828 ;
  assign n3931 = n3930 ^ n3929 ;
  assign n3932 = ~n3928 & n3931 ;
  assign n3933 = n3932 ^ n3930 ;
  assign n3934 = ~n3829 & n3933 ;
  assign n3935 = n3934 ^ x71 ;
  assign n3827 = n3826 ^ n3789 ;
  assign n3936 = n3935 ^ n3827 ;
  assign n3998 = n3827 ^ x70 ;
  assign n3950 = n3936 & ~n3998 ;
  assign n3946 = n3945 ^ n3944 ;
  assign n3947 = n3946 ^ x70 ;
  assign n3951 = n3950 ^ n3947 ;
  assign n3958 = n3957 ^ n3956 ;
  assign n3960 = n3958 ^ x69 ;
  assign n3959 = n3958 ^ n3946 ;
  assign n3961 = n3960 ^ n3959 ;
  assign n3962 = n3951 & ~n3961 ;
  assign n3963 = n3962 ^ n3960 ;
  assign n3967 = n3958 ^ x68 ;
  assign n3968 = ~n3963 & n3967 ;
  assign n3969 = n3968 ^ x68 ;
  assign n4099 = n3977 ^ n3969 ;
  assign n4100 = n4092 ^ n4082 ;
  assign n4101 = n4100 ^ n4081 ;
  assign n4102 = n4101 ^ x67 ;
  assign n4103 = n4102 ^ n3977 ;
  assign n4104 = n4103 ^ n4101 ;
  assign n4105 = ~n4099 & n4104 ;
  assign n4106 = n4105 ^ n4102 ;
  assign n4108 = n4097 ^ x66 ;
  assign n4107 = n4101 ^ n4097 ;
  assign n4109 = n4108 ^ n4107 ;
  assign n4110 = n4106 & ~n4109 ;
  assign n4111 = n4110 ^ n4108 ;
  assign n4112 = ~n4098 & n4111 ;
  assign n4121 = n4120 ^ n4112 ;
  assign n4080 = ~n3263 & n3712 ;
  assign n4122 = n4121 ^ n4080 ;
  assign n4124 = n4111 ^ x65 ;
  assign n4123 = n3264 & n3718 ;
  assign n4125 = n4124 ^ n4123 ;
  assign n4127 = n4106 ^ x66 ;
  assign n4126 = ~n3265 & n3715 ;
  assign n4128 = n4127 ^ n4126 ;
  assign n3964 = n3963 ^ x68 ;
  assign n3965 = ~n3297 & ~n3666 ;
  assign n3980 = n3964 & n3965 ;
  assign n3979 = n3266 & n3676 ;
  assign n3981 = n3980 ^ n3979 ;
  assign n3970 = n3969 ^ x67 ;
  assign n3978 = n3977 ^ n3970 ;
  assign n4129 = n3980 ^ n3978 ;
  assign n4130 = n3981 & n4129 ;
  assign n4131 = n4130 ^ n3980 ;
  assign n4132 = n4131 ^ n4126 ;
  assign n4133 = ~n4128 & ~n4132 ;
  assign n4134 = n4133 ^ n4127 ;
  assign n4135 = n4134 ^ n4123 ;
  assign n4136 = ~n4125 & n4135 ;
  assign n4137 = n4136 ^ n4124 ;
  assign n4138 = n4137 ^ n4080 ;
  assign n4139 = ~n4122 & n4138 ;
  assign n4140 = n4139 ^ n4121 ;
  assign n4141 = n4140 ^ n4077 ;
  assign n4142 = n4079 & n4141 ;
  assign n4143 = n4142 ^ n4078 ;
  assign n4144 = n4143 ^ n4074 ;
  assign n4145 = ~n4076 & ~n4144 ;
  assign n4146 = n4145 ^ n4075 ;
  assign n4147 = n4146 ^ n4070 ;
  assign n4148 = n4072 & ~n4147 ;
  assign n4149 = n4148 ^ n4071 ;
  assign n4150 = n4149 ^ n4067 ;
  assign n4151 = n4069 & n4150 ;
  assign n4152 = n4151 ^ n4068 ;
  assign n4153 = n4152 ^ n4064 ;
  assign n4154 = ~n4066 & n4153 ;
  assign n4155 = n4154 ^ n4065 ;
  assign n4156 = n4155 ^ n4062 ;
  assign n4157 = ~n4063 & ~n4156 ;
  assign n4158 = n4157 ^ n3989 ;
  assign n4159 = n4158 ^ n3688 ;
  assign n4160 = ~n4061 & n4159 ;
  assign n4161 = n4160 ^ n4060 ;
  assign n4162 = n4161 ^ n4057 ;
  assign n4163 = ~n4059 & n4162 ;
  assign n4164 = n4163 ^ n4058 ;
  assign n4165 = n4164 ^ n4054 ;
  assign n4166 = n4056 & n4165 ;
  assign n4167 = n4166 ^ n4055 ;
  assign n4168 = n4167 ^ n4051 ;
  assign n4169 = ~n4053 & n4168 ;
  assign n4170 = n4169 ^ n4052 ;
  assign n4171 = n4170 ^ n4048 ;
  assign n4172 = n4050 & ~n4171 ;
  assign n4173 = n4172 ^ n4049 ;
  assign n4174 = n4173 ^ n4045 ;
  assign n4175 = n4047 & n4174 ;
  assign n4176 = n4175 ^ n4046 ;
  assign n4177 = n4176 ^ n4042 ;
  assign n4178 = n4044 & n4177 ;
  assign n4179 = n4178 ^ n4043 ;
  assign n4180 = n4179 ^ n4039 ;
  assign n4181 = n4041 & ~n4180 ;
  assign n4182 = n4181 ^ n4040 ;
  assign n4183 = n4182 ^ n4037 ;
  assign n4184 = ~n4038 & ~n4183 ;
  assign n4186 = n4185 ^ n4184 ;
  assign n4187 = n4035 & ~n4186 ;
  assign n4188 = n4187 ^ n4034 ;
  assign n4189 = n4188 ^ n4031 ;
  assign n4190 = ~n4032 & n4189 ;
  assign n4191 = n4190 ^ n4031 ;
  assign n4192 = n4191 ^ n4027 ;
  assign n4193 = ~n4028 & ~n4192 ;
  assign n4195 = n4194 ^ n4193 ;
  assign n4196 = n4025 & n4195 ;
  assign n4197 = n4196 ^ n4024 ;
  assign n4021 = n3908 ^ x76 ;
  assign n4020 = ~n3633 & n4019 ;
  assign n4022 = n4021 ^ n4020 ;
  assign n4222 = n4197 ^ n4022 ;
  assign n4223 = n4195 ^ n4024 ;
  assign n4224 = n4191 ^ n4028 ;
  assign n4225 = n4188 ^ n4032 ;
  assign n4226 = n4186 ^ n4034 ;
  assign n4227 = n4182 ^ n4038 ;
  assign n4228 = n4179 ^ n4041 ;
  assign n4229 = n4176 ^ n4044 ;
  assign n4230 = n4173 ^ n4047 ;
  assign n4231 = n4158 ^ n4061 ;
  assign n4232 = n4155 ^ n4063 ;
  assign n4233 = n4140 ^ n4079 ;
  assign n4234 = n4137 ^ n4122 ;
  assign n4235 = n4134 ^ n4125 ;
  assign n3982 = n3981 ^ n3978 ;
  assign n4236 = n4131 ^ n4128 ;
  assign n4237 = n3982 & ~n4236 ;
  assign n4238 = n4235 & n4237 ;
  assign n4239 = n4234 & n4238 ;
  assign n4240 = n4233 & ~n4239 ;
  assign n4241 = n4143 ^ n4076 ;
  assign n4242 = n4240 & n4241 ;
  assign n4243 = n4146 ^ n4072 ;
  assign n4244 = n4242 & n4243 ;
  assign n4245 = n4149 ^ n4069 ;
  assign n4246 = ~n4244 & ~n4245 ;
  assign n4247 = n4152 ^ n4066 ;
  assign n4248 = ~n4246 & n4247 ;
  assign n4249 = ~n4232 & ~n4248 ;
  assign n4250 = ~n4231 & ~n4249 ;
  assign n4251 = n4161 ^ n4059 ;
  assign n4252 = ~n4250 & n4251 ;
  assign n4253 = n4164 ^ n4056 ;
  assign n4254 = ~n4252 & n4253 ;
  assign n4255 = n4167 ^ n4053 ;
  assign n4256 = n4254 & n4255 ;
  assign n4257 = n4170 ^ n4050 ;
  assign n4258 = ~n4256 & n4257 ;
  assign n4259 = ~n4230 & ~n4258 ;
  assign n4260 = n4229 & n4259 ;
  assign n4261 = n4228 & ~n4260 ;
  assign n4262 = ~n4227 & n4261 ;
  assign n4263 = n4226 & ~n4262 ;
  assign n4264 = ~n4225 & n4263 ;
  assign n4265 = ~n4224 & n4264 ;
  assign n4266 = ~n4223 & n4265 ;
  assign n4267 = ~n4222 & n4266 ;
  assign n4198 = n4197 ^ n4021 ;
  assign n4199 = ~n4022 & ~n4198 ;
  assign n4200 = n4199 ^ n4021 ;
  assign n4017 = n3913 ^ n3910 ;
  assign n4016 = n3361 & n4015 ;
  assign n4018 = n4017 ^ n4016 ;
  assign n4221 = n4200 ^ n4018 ;
  assign n4331 = n4267 ^ n4221 ;
  assign n4284 = n4259 ^ n4229 ;
  assign n4285 = n4258 ^ n4230 ;
  assign n4286 = n4249 ^ n4231 ;
  assign n4287 = n4248 ^ n4232 ;
  assign n4288 = n4243 ^ n4242 ;
  assign n3966 = n3965 ^ n3964 ;
  assign n4289 = n3966 & ~n3982 ;
  assign n4290 = n4236 ^ n3982 ;
  assign n4291 = n4289 & ~n4290 ;
  assign n4292 = n4237 ^ n4235 ;
  assign n4293 = ~n4291 & ~n4292 ;
  assign n4294 = n4238 ^ n4234 ;
  assign n4295 = n4293 & ~n4294 ;
  assign n4296 = n4239 ^ n4233 ;
  assign n4297 = ~n4295 & n4296 ;
  assign n4298 = n4241 ^ n4240 ;
  assign n4299 = n4297 & ~n4298 ;
  assign n4300 = n4288 & ~n4299 ;
  assign n4301 = n4245 ^ n4244 ;
  assign n4302 = n4300 & ~n4301 ;
  assign n4303 = n4247 ^ n4246 ;
  assign n4304 = ~n4302 & n4303 ;
  assign n4305 = n4287 & n4304 ;
  assign n4306 = n4286 & ~n4305 ;
  assign n4307 = n4251 ^ n4250 ;
  assign n4308 = n4306 & n4307 ;
  assign n4309 = n4253 ^ n4252 ;
  assign n4310 = n4308 & ~n4309 ;
  assign n4311 = n4255 ^ n4254 ;
  assign n4312 = n4310 & n4311 ;
  assign n4313 = n4257 ^ n4256 ;
  assign n4314 = ~n4312 & ~n4313 ;
  assign n4315 = ~n4285 & n4314 ;
  assign n4316 = n4284 & ~n4315 ;
  assign n4317 = n4260 ^ n4228 ;
  assign n4318 = ~n4316 & ~n4317 ;
  assign n4319 = n4261 ^ n4227 ;
  assign n4320 = n4318 & ~n4319 ;
  assign n4321 = n4262 ^ n4226 ;
  assign n4322 = n4320 & n4321 ;
  assign n4323 = n4263 ^ n4225 ;
  assign n4324 = n4322 & n4323 ;
  assign n4325 = n4264 ^ n4224 ;
  assign n4326 = n4324 & n4325 ;
  assign n4327 = n4265 ^ n4223 ;
  assign n4328 = ~n4326 & ~n4327 ;
  assign n4329 = n4266 ^ n4222 ;
  assign n4330 = ~n4328 & n4329 ;
  assign n4349 = n4331 ^ n4330 ;
  assign n4350 = n4349 ^ x102 ;
  assign n4351 = n4329 ^ n4328 ;
  assign n4352 = n4351 ^ x103 ;
  assign n4353 = n4327 ^ n4326 ;
  assign n4354 = n4353 ^ x104 ;
  assign n4377 = n4323 ^ n4322 ;
  assign n4378 = n4377 ^ x106 ;
  assign n4379 = n4321 ^ n4320 ;
  assign n4382 = n4379 ^ x107 ;
  assign n4380 = ~x107 & ~n4379 ;
  assign n4381 = n4380 ^ n4377 ;
  assign n4383 = n4382 ^ n4381 ;
  assign n4384 = n4378 & n4383 ;
  assign n4385 = n4384 ^ x106 ;
  assign n4376 = n4325 ^ n4324 ;
  assign n4386 = n4385 ^ n4376 ;
  assign n4355 = n4319 ^ n4318 ;
  assign n4356 = n4355 ^ x108 ;
  assign n4359 = n4355 ^ x109 ;
  assign n4357 = n4317 ^ n4316 ;
  assign n4358 = n4357 ^ n4355 ;
  assign n4360 = n4359 ^ n4358 ;
  assign n4361 = n4315 ^ n4284 ;
  assign n4362 = n4361 ^ x110 ;
  assign n4363 = n4314 ^ n4285 ;
  assign n4366 = n4363 ^ x111 ;
  assign n4364 = ~x111 & n4363 ;
  assign n4365 = n4364 ^ n4361 ;
  assign n4367 = n4366 ^ n4365 ;
  assign n4368 = n4362 & ~n4367 ;
  assign n4369 = n4368 ^ x110 ;
  assign n4370 = n4369 ^ n4355 ;
  assign n4371 = n4370 ^ n4359 ;
  assign n4372 = n4360 & n4371 ;
  assign n4373 = n4372 ^ n4359 ;
  assign n4374 = ~n4356 & n4373 ;
  assign n4375 = n4374 ^ x108 ;
  assign n4387 = n4386 ^ n4375 ;
  assign n4388 = n4387 ^ n4386 ;
  assign n4389 = ~x106 & ~n4377 ;
  assign n4390 = ~n4380 & n4389 ;
  assign n4391 = n4390 ^ n4380 ;
  assign n4392 = ~n4385 & ~n4391 ;
  assign n4395 = n4388 & n4392 ;
  assign n4396 = n4395 ^ n4386 ;
  assign n4398 = n4353 ^ x105 ;
  assign n4397 = n4376 ^ n4353 ;
  assign n4399 = n4398 ^ n4397 ;
  assign n4400 = ~n4396 & n4399 ;
  assign n4401 = n4400 ^ n4398 ;
  assign n4402 = ~n4354 & n4401 ;
  assign n4403 = n4402 ^ x104 ;
  assign n4404 = n4313 ^ n4312 ;
  assign n4405 = n4404 ^ x112 ;
  assign n4406 = n4311 ^ n4310 ;
  assign n4407 = n4406 ^ x113 ;
  assign n4408 = n4309 ^ n4308 ;
  assign n4409 = n4408 ^ x114 ;
  assign n4410 = n4307 ^ n4306 ;
  assign n4411 = n4410 ^ x115 ;
  assign n4412 = n4305 ^ n4286 ;
  assign n4413 = n4412 ^ x116 ;
  assign n4416 = n4303 ^ n4302 ;
  assign n4417 = n4416 ^ x118 ;
  assign n4456 = n4416 ^ x119 ;
  assign n4452 = n4301 ^ n4300 ;
  assign n4419 = n4298 ^ n4297 ;
  assign n4420 = n4419 ^ x121 ;
  assign n4421 = n4296 ^ n4295 ;
  assign n4422 = n4421 ^ x122 ;
  assign n4423 = n4294 ^ n4293 ;
  assign n4424 = n4423 ^ x123 ;
  assign n4425 = n4291 ^ n4237 ;
  assign n4426 = n4425 ^ n4235 ;
  assign n4427 = n4426 ^ x124 ;
  assign n3984 = x127 & ~n3966 ;
  assign n3985 = n3984 ^ x126 ;
  assign n3983 = n3982 ^ n3966 ;
  assign n4428 = n3984 ^ n3983 ;
  assign n4429 = n3985 & n4428 ;
  assign n4430 = n4429 ^ x126 ;
  assign n4431 = n4430 ^ x125 ;
  assign n4432 = n4290 ^ n4289 ;
  assign n4433 = n4432 ^ n4430 ;
  assign n4434 = n4431 & n4433 ;
  assign n4435 = n4434 ^ x125 ;
  assign n4436 = n4435 ^ n4426 ;
  assign n4437 = ~n4427 & n4436 ;
  assign n4438 = n4437 ^ x124 ;
  assign n4439 = n4438 ^ n4423 ;
  assign n4440 = n4424 & ~n4439 ;
  assign n4441 = n4440 ^ x123 ;
  assign n4442 = n4441 ^ n4421 ;
  assign n4443 = ~n4422 & n4442 ;
  assign n4444 = n4443 ^ x122 ;
  assign n4445 = n4444 ^ n4419 ;
  assign n4446 = ~n4420 & n4445 ;
  assign n4447 = n4446 ^ x121 ;
  assign n4418 = n4299 ^ n4288 ;
  assign n4448 = n4447 ^ n4418 ;
  assign n4449 = n4447 ^ x120 ;
  assign n4450 = ~n4448 & n4449 ;
  assign n4451 = n4450 ^ x120 ;
  assign n4453 = n4452 ^ n4451 ;
  assign n4454 = n4452 ^ x119 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4457 = n4456 ^ n4455 ;
  assign n4458 = ~n4417 & n4457 ;
  assign n4459 = n4458 ^ x118 ;
  assign n4415 = n4304 ^ n4287 ;
  assign n4460 = n4459 ^ n4415 ;
  assign n4744 = n4415 ^ x117 ;
  assign n4465 = ~n4460 & n4744 ;
  assign n4414 = n4412 ^ x117 ;
  assign n4466 = n4465 ^ n4414 ;
  assign n4467 = n4413 & ~n4466 ;
  assign n4468 = n4467 ^ x116 ;
  assign n4469 = n4468 ^ n4410 ;
  assign n4470 = ~n4411 & n4469 ;
  assign n4471 = n4470 ^ x115 ;
  assign n4472 = n4471 ^ n4408 ;
  assign n4473 = n4409 & ~n4472 ;
  assign n4474 = n4473 ^ x114 ;
  assign n4475 = n4474 ^ n4406 ;
  assign n4476 = ~n4407 & n4475 ;
  assign n4477 = n4476 ^ x113 ;
  assign n4478 = n4477 ^ n4404 ;
  assign n4479 = n4405 & ~n4478 ;
  assign n4480 = n4479 ^ x112 ;
  assign n4481 = ~x110 & ~n4361 ;
  assign n4482 = ~n4364 & n4481 ;
  assign n4483 = n4482 ^ n4364 ;
  assign n4484 = n4483 ^ n4355 ;
  assign n4485 = ~x109 & ~n4357 ;
  assign n4486 = ~n4483 & n4485 ;
  assign n4487 = n4486 ^ n4483 ;
  assign n4488 = ~x108 & ~n4487 ;
  assign n4489 = n4484 & n4488 ;
  assign n4490 = n4489 ^ n4487 ;
  assign n4491 = ~n4354 & ~n4490 ;
  assign n4492 = ~n4391 & n4491 ;
  assign n4493 = n4480 & n4492 ;
  assign n4494 = ~n4403 & n4493 ;
  assign n4497 = n4494 ^ n4403 ;
  assign n4495 = ~x105 & ~n4376 ;
  assign n4496 = n4494 & n4495 ;
  assign n4498 = n4497 ^ n4496 ;
  assign n4499 = n4498 ^ n4351 ;
  assign n4500 = ~n4352 & n4499 ;
  assign n4501 = n4500 ^ x103 ;
  assign n4502 = n4501 ^ n4349 ;
  assign n4503 = n4350 & ~n4502 ;
  assign n4504 = n4503 ^ x102 ;
  assign n4201 = n4200 ^ n4016 ;
  assign n4202 = ~n4018 & ~n4201 ;
  assign n4203 = n4202 ^ n4017 ;
  assign n4013 = n4012 ^ n3915 ;
  assign n4011 = n3284 & n4010 ;
  assign n4014 = n4013 ^ n4011 ;
  assign n4269 = n4203 ^ n4014 ;
  assign n4268 = n4221 & n4267 ;
  assign n4333 = n4269 ^ n4268 ;
  assign n4332 = ~n4330 & n4331 ;
  assign n4348 = n4333 ^ n4332 ;
  assign n4505 = n4504 ^ n4348 ;
  assign n4334 = ~n4332 & ~n4333 ;
  assign n4270 = ~n4268 & n4269 ;
  assign n4204 = n4203 ^ n4011 ;
  assign n4205 = ~n4014 & n4204 ;
  assign n4206 = n4205 ^ n4013 ;
  assign n4008 = n3922 ^ x73 ;
  assign n4007 = n3283 & ~n3610 ;
  assign n4009 = n4008 ^ n4007 ;
  assign n4220 = n4206 ^ n4009 ;
  assign n4283 = n4270 ^ n4220 ;
  assign n4346 = n4334 ^ n4283 ;
  assign n4506 = n4346 ^ x101 ;
  assign n4507 = n4506 ^ n4346 ;
  assign n4508 = n4507 ^ n4348 ;
  assign n4509 = ~n4505 & n4508 ;
  assign n4510 = n4509 ^ n4506 ;
  assign n4540 = n4510 ^ x100 ;
  assign n4581 = n4543 ^ n4540 ;
  assign n4639 = x159 & ~n4581 ;
  assign n4207 = n4206 ^ n4007 ;
  assign n4208 = n4009 & ~n4207 ;
  assign n4209 = n4208 ^ n4008 ;
  assign n4005 = n3928 ^ x72 ;
  assign n4004 = ~n3287 & n3592 ;
  assign n4006 = n4005 ^ n4004 ;
  assign n4272 = n4209 ^ n4006 ;
  assign n4271 = n4220 & ~n4270 ;
  assign n4336 = n4272 ^ n4271 ;
  assign n4335 = ~n4283 & ~n4334 ;
  assign n4514 = n4336 ^ n4335 ;
  assign n4347 = n4346 ^ x100 ;
  assign n4511 = ~n4347 & n4510 ;
  assign n4512 = n4511 ^ x100 ;
  assign n4513 = n4512 ^ x99 ;
  assign n4550 = n4514 ^ n4513 ;
  assign n4544 = ~n4540 & ~n4543 ;
  assign n4545 = n4544 ^ n3266 ;
  assign n4546 = n4545 ^ n3718 ;
  assign n4547 = n4546 ^ n4544 ;
  assign n4548 = n4074 & n4547 ;
  assign n4549 = n4548 ^ n4545 ;
  assign n4580 = n4550 ^ n4549 ;
  assign n4638 = n4581 ^ n4580 ;
  assign n4640 = n4639 ^ n4638 ;
  assign n4641 = n4639 ^ x158 ;
  assign n4642 = ~n4640 & n4641 ;
  assign n4643 = n4642 ^ x158 ;
  assign n4536 = n3712 ^ n3265 ;
  assign n4537 = ~n4071 & ~n4536 ;
  assign n4538 = n4537 ^ n3265 ;
  assign n4553 = n4544 ^ n4538 ;
  assign n4551 = n4550 ^ n4544 ;
  assign n4552 = n4549 & n4551 ;
  assign n4554 = n4553 ^ n4552 ;
  assign n4210 = n4209 ^ n4004 ;
  assign n4211 = ~n4006 & ~n4210 ;
  assign n4212 = n4211 ^ n4005 ;
  assign n4002 = n3933 ^ x71 ;
  assign n4001 = ~n3282 & n3606 ;
  assign n4003 = n4002 ^ n4001 ;
  assign n4274 = n4212 ^ n4003 ;
  assign n4273 = n4271 & ~n4272 ;
  assign n4338 = n4274 ^ n4273 ;
  assign n4337 = n4335 & ~n4336 ;
  assign n4345 = n4338 ^ n4337 ;
  assign n4534 = n4345 ^ x98 ;
  assign n4515 = n4514 ^ n4512 ;
  assign n4516 = n4513 & ~n4515 ;
  assign n4517 = n4516 ^ x99 ;
  assign n4535 = n4534 ^ n4517 ;
  assign n4583 = n4554 ^ n4535 ;
  assign n4582 = n4580 & n4581 ;
  assign n4637 = n4583 ^ n4582 ;
  assign n4644 = n4643 ^ n4637 ;
  assign n4645 = n4643 ^ x157 ;
  assign n4646 = n4644 & n4645 ;
  assign n4647 = n4646 ^ x157 ;
  assign n4584 = n4582 & ~n4583 ;
  assign n4539 = n4538 ^ n4535 ;
  assign n4555 = ~n4539 & ~n4554 ;
  assign n4556 = n4555 ^ n4538 ;
  assign n4518 = n4517 ^ n4345 ;
  assign n4519 = n4517 ^ x98 ;
  assign n4520 = ~n4518 & n4519 ;
  assign n4521 = n4520 ^ x98 ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4213 = n4212 ^ n4001 ;
  assign n4214 = ~n4003 & ~n4213 ;
  assign n4215 = n4214 ^ n4002 ;
  assign n3999 = n3998 ^ n3935 ;
  assign n3997 = x31 & ~n3624 ;
  assign n4000 = n3999 ^ n3997 ;
  assign n4281 = n4215 ^ n4000 ;
  assign n4275 = n4273 & n4274 ;
  assign n4282 = n4281 ^ n4275 ;
  assign n4343 = n4339 ^ n4282 ;
  assign n4344 = n4343 ^ x97 ;
  assign n4532 = n4521 ^ n4344 ;
  assign n4529 = n3711 ^ n3264 ;
  assign n4530 = n4068 & n4529 ;
  assign n4531 = n4530 ^ n3264 ;
  assign n4533 = n4532 ^ n4531 ;
  assign n4579 = n4556 ^ n4533 ;
  assign n4635 = n4584 ^ n4579 ;
  assign n4636 = n4635 ^ x156 ;
  assign n5323 = n4647 ^ n4636 ;
  assign n4706 = n4454 ^ n4451 ;
  assign n5290 = n4049 ^ n3703 ;
  assign n5291 = n4706 & ~n5290 ;
  assign n5292 = n5291 ^ n3703 ;
  assign n5395 = n5323 ^ n5292 ;
  assign n5312 = n4637 ^ x157 ;
  assign n5313 = n5312 ^ n4643 ;
  assign n4683 = n4444 ^ n4420 ;
  assign n5304 = n4055 ^ n3689 ;
  assign n5305 = ~n4683 & ~n5304 ;
  assign n5306 = n5305 ^ n3689 ;
  assign n4673 = n4441 ^ n4422 ;
  assign n5296 = n4058 ^ n3707 ;
  assign n5297 = ~n4673 & n5296 ;
  assign n5298 = n5297 ^ n3707 ;
  assign n4609 = n4438 ^ n4424 ;
  assign n4218 = n3951 ^ x69 ;
  assign n4944 = n4480 & ~n4490 ;
  assign n4945 = ~n4375 & n4944 ;
  assign n4946 = n4945 ^ n4375 ;
  assign n4956 = n4946 ^ n4382 ;
  assign n4953 = n3610 ^ n3361 ;
  assign n4954 = ~n3999 & ~n4953 ;
  assign n4955 = n4954 ^ n3361 ;
  assign n4957 = n4956 ^ n4955 ;
  assign n4929 = ~n4369 & n4480 ;
  assign n4930 = ~n4483 & n4929 ;
  assign n4931 = n4930 ^ n4369 ;
  assign n4928 = n4357 ^ x109 ;
  assign n4932 = n4931 ^ n4928 ;
  assign n4933 = n4932 ^ n3617 ;
  assign n4934 = n4933 ^ n4015 ;
  assign n4935 = n4934 ^ n4932 ;
  assign n4936 = n4005 & n4935 ;
  assign n4937 = n4936 ^ n4933 ;
  assign n4885 = n4480 ^ n4366 ;
  assign n4886 = n4885 ^ n3580 ;
  assign n4887 = n4886 ^ n3971 ;
  assign n4888 = n4887 ^ n4885 ;
  assign n4889 = ~n4013 & ~n4888 ;
  assign n4890 = n4889 ^ n4886 ;
  assign n4877 = n4477 ^ n4405 ;
  assign n4874 = n3952 ^ n3568 ;
  assign n4875 = ~n4017 & n4874 ;
  assign n4876 = n4875 ^ n3568 ;
  assign n4878 = n4877 ^ n4876 ;
  assign n4862 = n4474 ^ n4407 ;
  assign n4859 = n3942 ^ n3556 ;
  assign n4860 = n4021 & ~n4859 ;
  assign n4861 = n4860 ^ n3556 ;
  assign n4863 = n4862 ^ n4861 ;
  assign n4851 = n4471 ^ n4409 ;
  assign n4848 = n3787 ^ n3544 ;
  assign n4849 = ~n4024 & ~n4848 ;
  assign n4850 = n4849 ^ n3544 ;
  assign n4852 = n4851 ^ n4850 ;
  assign n4828 = n4468 ^ x115 ;
  assign n4829 = n4828 ^ n4410 ;
  assign n4825 = n3693 ^ n3532 ;
  assign n4826 = n4027 & n4825 ;
  assign n4827 = n4826 ^ n3532 ;
  assign n4830 = n4829 ^ n4827 ;
  assign n4813 = n3694 ^ n3520 ;
  assign n4814 = ~n4031 & ~n4813 ;
  assign n4815 = n4814 ^ n3520 ;
  assign n4745 = n4744 ^ n4459 ;
  assign n4746 = n4745 ^ n3508 ;
  assign n4747 = n4746 ^ n3743 ;
  assign n4748 = n4747 ^ n4745 ;
  assign n4749 = ~n4034 & n4748 ;
  assign n4750 = n4749 ^ n4746 ;
  assign n4726 = n3696 ^ n3259 ;
  assign n4727 = ~n4037 & n4726 ;
  assign n4728 = n4727 ^ n3259 ;
  assign n4723 = x119 ^ x118 ;
  assign n4724 = n4723 ^ n4416 ;
  assign n4725 = n4724 ^ n4455 ;
  assign n4729 = n4728 ^ n4725 ;
  assign n4703 = n3698 ^ n3316 ;
  assign n4704 = n4040 & ~n4703 ;
  assign n4705 = n4704 ^ n3316 ;
  assign n4707 = n4706 ^ n4705 ;
  assign n4711 = n4418 ^ x120 ;
  assign n4712 = n4711 ^ n4447 ;
  assign n4708 = n3699 ^ n3314 ;
  assign n4709 = n4043 & ~n4708 ;
  assign n4710 = n4709 ^ n3314 ;
  assign n4713 = n4712 ^ n4710 ;
  assign n4684 = n4683 ^ n4673 ;
  assign n4670 = n3701 ^ n3261 ;
  assign n4671 = n4049 & n4670 ;
  assign n4672 = n4671 ^ n3261 ;
  assign n4674 = n4673 ^ n4672 ;
  assign n4598 = n4435 ^ x124 ;
  assign n4599 = n4598 ^ n4426 ;
  assign n4610 = n4609 ^ n4599 ;
  assign n4595 = n3703 ^ n3309 ;
  assign n4596 = n4055 & ~n4595 ;
  assign n4597 = n4596 ^ n3309 ;
  assign n4600 = n4599 ^ n4597 ;
  assign n4570 = n3705 ^ n3307 ;
  assign n4571 = ~n4058 & ~n4570 ;
  assign n4572 = n4571 ^ n3307 ;
  assign n4569 = n4432 ^ n4431 ;
  assign n4573 = n4572 ^ n4569 ;
  assign n3986 = n3985 ^ n3983 ;
  assign n3690 = n3689 ^ n3305 ;
  assign n3691 = n3688 & n3690 ;
  assign n3692 = n3691 ^ n3305 ;
  assign n3987 = n3986 ^ n3692 ;
  assign n3990 = n3966 ^ x127 ;
  assign n3991 = n3990 ^ n3303 ;
  assign n3992 = n3991 ^ n3707 ;
  assign n3993 = n3992 ^ n3990 ;
  assign n3994 = ~n3989 & n3993 ;
  assign n3995 = n3994 ^ n3991 ;
  assign n4525 = n3709 ^ n3263 ;
  assign n4526 = ~n4064 & n4525 ;
  assign n4527 = n4526 ^ n3263 ;
  assign n4522 = n4521 ^ n4343 ;
  assign n4523 = n4344 & ~n4522 ;
  assign n4340 = n4339 ^ n4275 ;
  assign n4341 = n4282 & ~n4340 ;
  assign n4276 = n4275 ^ x96 ;
  assign n4219 = n4218 ^ n3999 ;
  assign n4277 = n4276 ^ n4219 ;
  assign n4278 = n4277 ^ x97 ;
  assign n4216 = n4215 ^ n3999 ;
  assign n4217 = n4000 & n4216 ;
  assign n4279 = n4278 ^ n4217 ;
  assign n3996 = ~n3243 & ~n3636 ;
  assign n4280 = n4279 ^ n3996 ;
  assign n4342 = n4341 ^ n4280 ;
  assign n4524 = n4523 ^ n4342 ;
  assign n4528 = n4527 ^ n4524 ;
  assign n4557 = n4556 ^ n4531 ;
  assign n4558 = n4533 & n4557 ;
  assign n4559 = n4558 ^ n4532 ;
  assign n4560 = n4559 ^ n4524 ;
  assign n4561 = ~n4528 & ~n4560 ;
  assign n4562 = n4561 ^ n4527 ;
  assign n4563 = n4562 ^ n3990 ;
  assign n4564 = n3995 & n4563 ;
  assign n4565 = n4564 ^ n3990 ;
  assign n4566 = n4565 ^ n3692 ;
  assign n4567 = n3987 & ~n4566 ;
  assign n4568 = n4567 ^ n3986 ;
  assign n4592 = n4569 ^ n4568 ;
  assign n4593 = ~n4573 & ~n4592 ;
  assign n4594 = n4593 ^ n4572 ;
  assign n4607 = n4597 ^ n4594 ;
  assign n4608 = ~n4600 & ~n4607 ;
  assign n4611 = n4610 ^ n4608 ;
  assign n4612 = n3702 ^ n3262 ;
  assign n4613 = ~n4052 & n4612 ;
  assign n4614 = n4613 ^ n3702 ;
  assign n4667 = n4614 ^ n4609 ;
  assign n4668 = ~n4611 & ~n4667 ;
  assign n4669 = n4668 ^ n4609 ;
  assign n4681 = n4672 ^ n4669 ;
  assign n4682 = ~n4674 & ~n4681 ;
  assign n4685 = n4684 ^ n4682 ;
  assign n4686 = n3700 ^ n3260 ;
  assign n4687 = ~n4046 & ~n4686 ;
  assign n4688 = n4687 ^ n3260 ;
  assign n4714 = n4688 ^ n4683 ;
  assign n4715 = n4685 & n4714 ;
  assign n4716 = n4715 ^ n4683 ;
  assign n4717 = n4716 ^ n4710 ;
  assign n4718 = n4713 & n4717 ;
  assign n4719 = n4718 ^ n4712 ;
  assign n4720 = n4719 ^ n4705 ;
  assign n4721 = ~n4707 & n4720 ;
  assign n4722 = n4721 ^ n4706 ;
  assign n4751 = n4725 ^ n4722 ;
  assign n4752 = n4729 & n4751 ;
  assign n4753 = n4752 ^ n4728 ;
  assign n4810 = n4753 ^ n4745 ;
  assign n4811 = n4750 & ~n4810 ;
  assign n4812 = n4811 ^ n4745 ;
  assign n4816 = n4815 ^ n4812 ;
  assign n4817 = n4413 ^ x117 ;
  assign n4821 = n4817 ^ n4465 ;
  assign n4822 = n4821 ^ n4812 ;
  assign n4823 = ~n4816 & ~n4822 ;
  assign n4824 = n4823 ^ n4815 ;
  assign n4845 = n4827 ^ n4824 ;
  assign n4846 = n4830 & ~n4845 ;
  assign n4847 = n4846 ^ n4829 ;
  assign n4856 = n4850 ^ n4847 ;
  assign n4857 = ~n4852 & ~n4856 ;
  assign n4858 = n4857 ^ n4851 ;
  assign n4879 = n4861 ^ n4858 ;
  assign n4880 = ~n4863 & ~n4879 ;
  assign n4881 = n4880 ^ n4862 ;
  assign n4882 = n4881 ^ n4876 ;
  assign n4883 = ~n4878 & ~n4882 ;
  assign n4884 = n4883 ^ n4877 ;
  assign n4904 = n4885 ^ n4884 ;
  assign n4905 = n4890 & ~n4904 ;
  assign n4900 = n4480 ^ n4363 ;
  assign n4901 = ~n4366 & n4900 ;
  assign n4898 = x111 ^ x110 ;
  assign n4899 = n4898 ^ n4361 ;
  assign n4902 = n4901 ^ n4899 ;
  assign n4903 = n4902 ^ n4885 ;
  assign n4906 = n4905 ^ n4903 ;
  assign n4907 = n4019 ^ n3594 ;
  assign n4908 = ~n4008 & n4907 ;
  assign n4909 = n4908 ^ n3594 ;
  assign n4925 = n4909 ^ n4902 ;
  assign n4926 = ~n4906 & n4925 ;
  assign n4927 = n4926 ^ n4902 ;
  assign n4962 = n4932 ^ n4927 ;
  assign n4963 = n4937 & n4962 ;
  assign n4958 = n4010 ^ n3633 ;
  assign n4959 = ~n4002 & n4958 ;
  assign n4960 = n4959 ^ n3633 ;
  assign n4961 = n4960 ^ n4932 ;
  assign n4964 = n4963 ^ n4961 ;
  assign n4967 = n4931 ^ n4357 ;
  assign n4968 = n4356 ^ x109 ;
  assign n4969 = n4968 ^ n4356 ;
  assign n4970 = n4969 ^ n4931 ;
  assign n4971 = ~n4967 & n4970 ;
  assign n4972 = n4971 ^ n4968 ;
  assign n4973 = n4972 ^ n4960 ;
  assign n4974 = n4964 & ~n4973 ;
  assign n4965 = n4960 ^ n4956 ;
  assign n4975 = n4974 ^ n4965 ;
  assign n4976 = n4957 & n4975 ;
  assign n4977 = n4976 ^ n4956 ;
  assign n4978 = n4977 ^ n3284 ;
  assign n4979 = n4978 ^ n3592 ;
  assign n4980 = n4979 ^ n4977 ;
  assign n4981 = ~n4218 & n4980 ;
  assign n4982 = n4981 ^ n4978 ;
  assign n5066 = n4376 ^ x105 ;
  assign n5064 = n4392 & n4946 ;
  assign n5065 = n5064 ^ n4385 ;
  assign n5067 = n5066 ^ n5065 ;
  assign n5068 = n5067 ^ n4977 ;
  assign n5069 = n5068 ^ n5067 ;
  assign n4947 = n4946 ^ n4379 ;
  assign n4948 = n4378 ^ x107 ;
  assign n4949 = n4948 ^ n4378 ;
  assign n4950 = n4949 ^ n4946 ;
  assign n4951 = ~n4947 & n4950 ;
  assign n4952 = n4951 ^ n4948 ;
  assign n5070 = n5069 ^ n4952 ;
  assign n5071 = n4982 & n5070 ;
  assign n5072 = n5071 ^ n5068 ;
  assign n5096 = n5065 ^ n4376 ;
  assign n5097 = n4354 ^ x105 ;
  assign n5098 = n5097 ^ n4354 ;
  assign n5099 = n5098 ^ n5065 ;
  assign n5100 = ~n5096 & n5099 ;
  assign n5101 = n5100 ^ n5097 ;
  assign n5102 = n5101 ^ n5067 ;
  assign n5073 = n3606 ^ n3283 ;
  assign n5074 = n3964 & ~n5073 ;
  assign n5075 = n5074 ^ n3283 ;
  assign n5103 = n5102 ^ n5075 ;
  assign n5104 = n5103 ^ n5101 ;
  assign n5105 = n5072 & ~n5104 ;
  assign n5106 = n5105 ^ n5102 ;
  assign n5107 = n3624 ^ n3287 ;
  assign n5108 = n3978 & ~n5107 ;
  assign n5109 = n5108 ^ n3287 ;
  assign n5136 = n5109 ^ n5101 ;
  assign n5137 = n5106 & ~n5136 ;
  assign n5138 = n5137 ^ n5109 ;
  assign n5129 = n4498 ^ x103 ;
  assign n5130 = n5129 ^ n4351 ;
  assign n5131 = n5130 ^ n3282 ;
  assign n5132 = n5131 ^ n3636 ;
  assign n5133 = n5132 ^ n5130 ;
  assign n5134 = ~n4127 & n5133 ;
  assign n5135 = n5134 ^ n5131 ;
  assign n5139 = n5138 ^ n5135 ;
  assign n5076 = n5075 ^ n5072 ;
  assign n4983 = n4982 ^ n4952 ;
  assign n4984 = n4975 ^ n4955 ;
  assign n4985 = n4972 ^ n4964 ;
  assign n4891 = n4890 ^ n4884 ;
  assign n4892 = n4881 ^ n4878 ;
  assign n4897 = n4891 & n4892 ;
  assign n4910 = n4909 ^ n4906 ;
  assign n4924 = ~n4897 & n4910 ;
  assign n4938 = n4937 ^ n4927 ;
  assign n4986 = n4924 & ~n4938 ;
  assign n4987 = n4985 & n4986 ;
  assign n4988 = n4984 & ~n4987 ;
  assign n5077 = n4983 & n4988 ;
  assign n5095 = n5076 & ~n5077 ;
  assign n5110 = n5109 ^ n5106 ;
  assign n5140 = n5095 & n5110 ;
  assign n5174 = n5139 & ~n5140 ;
  assign n5170 = n3666 ^ x31 ;
  assign n5171 = ~n4124 & n5170 ;
  assign n5172 = n5171 ^ x31 ;
  assign n5164 = n4501 ^ n4350 ;
  assign n5166 = n5164 ^ n5130 ;
  assign n5165 = n5164 ^ n5138 ;
  assign n5167 = n5166 ^ n5165 ;
  assign n5168 = n5135 & ~n5167 ;
  assign n5169 = n5168 ^ n5166 ;
  assign n5173 = n5172 ^ n5169 ;
  assign n5175 = n5174 ^ n5173 ;
  assign n5141 = n5140 ^ n5139 ;
  assign n5078 = n5077 ^ n5076 ;
  assign n4989 = n4988 ^ n4983 ;
  assign n4990 = n4987 ^ n4984 ;
  assign n4991 = n4986 ^ n4985 ;
  assign n4893 = n4892 ^ n4891 ;
  assign n4853 = n4852 ^ n4847 ;
  assign n4831 = n4830 ^ n4824 ;
  assign n4832 = n4821 ^ n4816 ;
  assign n4754 = n4753 ^ n4750 ;
  assign n4730 = n4729 ^ n4722 ;
  assign n4731 = n4719 ^ n4707 ;
  assign n4732 = n4716 ^ n4713 ;
  assign n4689 = n4688 ^ n4685 ;
  assign n4675 = n4674 ^ n4669 ;
  assign n4615 = n4614 ^ n4611 ;
  assign n4574 = n4573 ^ n4568 ;
  assign n4575 = n4565 ^ n3987 ;
  assign n4576 = n4575 ^ n4574 ;
  assign n4577 = n4574 & ~n4576 ;
  assign n4591 = n4577 ^ n4575 ;
  assign n4601 = n4600 ^ n4594 ;
  assign n4616 = ~n4591 & ~n4601 ;
  assign n4676 = n4615 & n4616 ;
  assign n4690 = ~n4675 & n4676 ;
  assign n4733 = n4689 & ~n4690 ;
  assign n4734 = ~n4732 & ~n4733 ;
  assign n4735 = ~n4731 & n4734 ;
  assign n4743 = ~n4730 & ~n4735 ;
  assign n4755 = n4754 ^ n4743 ;
  assign n4736 = n4735 ^ n4730 ;
  assign n4737 = n4734 ^ n4731 ;
  assign n4738 = n4733 ^ n4732 ;
  assign n4691 = n4690 ^ n4689 ;
  assign n4677 = n4676 ^ n4675 ;
  assign n4617 = n4616 ^ n4615 ;
  assign n4578 = n4559 ^ n4528 ;
  assign n4585 = n4579 & ~n4584 ;
  assign n4586 = n4578 & n4585 ;
  assign n4587 = n4562 ^ n3995 ;
  assign n4588 = ~n4586 & ~n4587 ;
  assign n4589 = n4577 & n4588 ;
  assign n4590 = n4589 ^ n4576 ;
  assign n4602 = n4601 ^ n4591 ;
  assign n4618 = ~n4590 & ~n4602 ;
  assign n4678 = n4617 & ~n4618 ;
  assign n4692 = ~n4677 & n4678 ;
  assign n4739 = ~n4691 & ~n4692 ;
  assign n4740 = ~n4738 & n4739 ;
  assign n4741 = n4737 & n4740 ;
  assign n4742 = n4736 & n4741 ;
  assign n4833 = n4743 ^ n4742 ;
  assign n4834 = n4755 & n4833 ;
  assign n4835 = n4834 ^ n4743 ;
  assign n4836 = n4832 & n4835 ;
  assign n4854 = n4831 & n4836 ;
  assign n4855 = n4853 & ~n4854 ;
  assign n4864 = n4863 ^ n4858 ;
  assign n4894 = n4855 & ~n4864 ;
  assign n4895 = ~n4892 & n4894 ;
  assign n4896 = n4893 & n4895 ;
  assign n4911 = n4910 ^ n4897 ;
  assign n4923 = n4896 & n4911 ;
  assign n4939 = n4938 ^ n4924 ;
  assign n4992 = ~n4923 & ~n4939 ;
  assign n4993 = ~n4991 & ~n4992 ;
  assign n4994 = n4990 & ~n4993 ;
  assign n5079 = n4989 & ~n4994 ;
  assign n5094 = ~n5078 & ~n5079 ;
  assign n5111 = n5110 ^ n5095 ;
  assign n5142 = n5094 & n5111 ;
  assign n5163 = ~n5141 & ~n5142 ;
  assign n5203 = n5174 ^ n5163 ;
  assign n5204 = n5175 & n5203 ;
  assign n5196 = n4348 ^ x101 ;
  assign n5197 = n5196 ^ n4504 ;
  assign n5195 = n5172 ^ n3243 ;
  assign n5198 = n5197 ^ n5195 ;
  assign n5194 = n5174 ^ x128 ;
  assign n5199 = n5198 ^ n5194 ;
  assign n5200 = n5199 ^ x129 ;
  assign n5192 = n3676 ^ n3243 ;
  assign n5193 = ~n4121 & ~n5192 ;
  assign n5201 = n5200 ^ n5193 ;
  assign n5190 = n5172 ^ n5164 ;
  assign n5191 = n5169 & ~n5190 ;
  assign n5202 = n5201 ^ n5191 ;
  assign n5205 = n5204 ^ n5202 ;
  assign n5143 = n5142 ^ n5141 ;
  assign n5144 = n5143 ^ x130 ;
  assign n5112 = n5111 ^ n5094 ;
  assign n5113 = n5112 ^ x131 ;
  assign n5080 = n5079 ^ n5078 ;
  assign n5081 = n5080 ^ x132 ;
  assign n4756 = n4755 ^ n4742 ;
  assign n4757 = n4756 ^ x144 ;
  assign n4774 = n4741 ^ n4736 ;
  assign n4767 = n4739 ^ n4738 ;
  assign n4768 = x147 & n4767 ;
  assign n4769 = n4768 ^ x146 ;
  assign n4770 = n4740 ^ n4737 ;
  assign n4771 = n4770 ^ n4768 ;
  assign n4772 = n4769 & n4771 ;
  assign n4773 = n4772 ^ x146 ;
  assign n4775 = n4774 ^ n4773 ;
  assign n4693 = n4692 ^ n4691 ;
  assign n4694 = n4693 ^ x148 ;
  assign n4759 = n4693 ^ x149 ;
  assign n4679 = n4678 ^ n4677 ;
  assign n4758 = n4693 ^ n4679 ;
  assign n4760 = n4759 ^ n4758 ;
  assign n4603 = n4602 ^ n4590 ;
  assign n4605 = x151 & ~n4603 ;
  assign n4623 = n4605 ^ x150 ;
  assign n4619 = n4618 ^ n4617 ;
  assign n4624 = n4619 ^ n4605 ;
  assign n4625 = n4623 & n4624 ;
  assign n4626 = n4625 ^ x150 ;
  assign n4761 = n4693 ^ n4626 ;
  assign n4762 = n4761 ^ n4759 ;
  assign n4763 = ~n4760 & n4762 ;
  assign n4764 = n4763 ^ n4759 ;
  assign n4765 = ~n4694 & n4764 ;
  assign n4766 = n4765 ^ x148 ;
  assign n4776 = n4775 ^ n4766 ;
  assign n4777 = n4776 ^ n4775 ;
  assign n4778 = n4767 ^ x147 ;
  assign n4779 = n4778 ^ n4768 ;
  assign n4780 = ~x146 & n4770 ;
  assign n4781 = n4779 & n4780 ;
  assign n4782 = n4781 ^ n4779 ;
  assign n4783 = ~n4773 & n4782 ;
  assign n4786 = n4777 & n4783 ;
  assign n4787 = n4786 ^ n4775 ;
  assign n4789 = n4756 ^ x145 ;
  assign n4788 = n4774 ^ n4756 ;
  assign n4790 = n4789 ^ n4788 ;
  assign n4791 = n4787 & ~n4790 ;
  assign n4792 = n4791 ^ n4789 ;
  assign n4793 = ~n4757 & n4792 ;
  assign n4794 = n4793 ^ x144 ;
  assign n4627 = n4575 & n4588 ;
  assign n4628 = n4627 ^ n4576 ;
  assign n4629 = n4628 ^ x152 ;
  assign n4630 = n4588 ^ n4575 ;
  assign n4631 = n4630 ^ x153 ;
  assign n4632 = n4587 ^ n4586 ;
  assign n4633 = n4632 ^ x154 ;
  assign n4648 = n4647 ^ n4635 ;
  assign n4649 = n4636 & ~n4648 ;
  assign n4650 = n4649 ^ x156 ;
  assign n4634 = n4585 ^ n4578 ;
  assign n4651 = n4650 ^ n4634 ;
  assign n4652 = n4650 ^ x155 ;
  assign n4653 = n4651 & n4652 ;
  assign n4654 = n4653 ^ x155 ;
  assign n4655 = n4654 ^ n4632 ;
  assign n4656 = n4633 & ~n4655 ;
  assign n4657 = n4656 ^ x154 ;
  assign n4658 = n4657 ^ n4630 ;
  assign n4659 = n4631 & ~n4658 ;
  assign n4660 = n4659 ^ x153 ;
  assign n4661 = n4660 ^ n4628 ;
  assign n4662 = ~n4629 & n4661 ;
  assign n4663 = n4662 ^ x152 ;
  assign n4604 = n4603 ^ x151 ;
  assign n4606 = n4605 ^ n4604 ;
  assign n4620 = ~x150 & n4619 ;
  assign n4621 = ~n4606 & n4620 ;
  assign n4622 = n4621 ^ n4606 ;
  assign n4795 = n4694 ^ n4622 ;
  assign n4796 = ~x149 & n4679 ;
  assign n4797 = ~n4622 & n4796 ;
  assign n4798 = n4797 ^ n4622 ;
  assign n4799 = n4693 & ~n4798 ;
  assign n4800 = n4795 & n4799 ;
  assign n4801 = n4800 ^ n4798 ;
  assign n4802 = ~n4757 & ~n4801 ;
  assign n4803 = n4782 & n4802 ;
  assign n4804 = n4663 & n4803 ;
  assign n4805 = ~n4794 & n4804 ;
  assign n4808 = n4805 ^ n4794 ;
  assign n4806 = ~x145 & n4774 ;
  assign n4807 = n4805 & n4806 ;
  assign n4809 = n4808 ^ n4807 ;
  assign n4837 = n4836 ^ n4831 ;
  assign n4838 = n4832 ^ n4743 ;
  assign n4839 = n4838 ^ n4834 ;
  assign n4840 = ~x143 & n4839 ;
  assign n4841 = ~x142 & ~n4840 ;
  assign n4842 = n4837 & n4841 ;
  assign n4843 = n4842 ^ n4840 ;
  assign n4844 = n4843 ^ x140 ;
  assign n4865 = n4864 ^ n4855 ;
  assign n4866 = n4854 ^ n4853 ;
  assign n4867 = ~x141 & n4866 ;
  assign n4868 = ~n4843 & n4867 ;
  assign n4869 = n4868 ^ n4843 ;
  assign n4870 = n4865 & ~n4869 ;
  assign n4871 = ~n4844 & n4870 ;
  assign n4872 = n4871 ^ n4869 ;
  assign n4873 = n4809 & ~n4872 ;
  assign n4912 = n4911 ^ n4896 ;
  assign n4913 = n4895 ^ n4893 ;
  assign n4914 = n4894 ^ n4892 ;
  assign n4915 = ~x139 & n4914 ;
  assign n4916 = ~x138 & ~n4915 ;
  assign n4917 = ~n4913 & n4916 ;
  assign n4918 = n4917 ^ n4915 ;
  assign n4919 = ~n4872 & ~n4918 ;
  assign n4920 = ~x137 & n4919 ;
  assign n4921 = ~n4912 & n4920 ;
  assign n4922 = n4921 ^ n4919 ;
  assign n4940 = n4939 ^ n4923 ;
  assign n4941 = ~x136 & n4940 ;
  assign n4942 = n4922 & n4941 ;
  assign n4943 = n4942 ^ n4922 ;
  assign n4995 = n4994 ^ n4989 ;
  assign n4996 = n4995 ^ x133 ;
  assign n4997 = n4943 & ~n4996 ;
  assign n4998 = n4992 ^ n4991 ;
  assign n5000 = n4998 ^ x135 ;
  assign n4999 = x135 & n4998 ;
  assign n5001 = n5000 ^ n4999 ;
  assign n5002 = n4993 ^ n4990 ;
  assign n5003 = ~x134 & ~n5002 ;
  assign n5004 = n5001 & n5003 ;
  assign n5005 = n5004 ^ n5001 ;
  assign n5006 = n4997 & n5005 ;
  assign n5007 = n4873 & n5006 ;
  assign n5049 = n5002 ^ n4999 ;
  assign n5050 = n5002 ^ x134 ;
  assign n5051 = ~n5049 & n5050 ;
  assign n5052 = n5051 ^ x134 ;
  assign n5053 = n5052 ^ n4995 ;
  assign n5008 = n4940 ^ x136 ;
  assign n5045 = n4940 ^ x137 ;
  assign n5009 = n4912 ^ x137 ;
  assign n5010 = n4913 ^ x138 ;
  assign n5012 = n4914 ^ x139 ;
  assign n5011 = n4915 ^ n4913 ;
  assign n5013 = n5012 ^ n5011 ;
  assign n5014 = n5010 & ~n5013 ;
  assign n5015 = n5014 ^ x138 ;
  assign n5019 = n4865 ^ x140 ;
  assign n5021 = n4837 ^ x142 ;
  assign n5023 = n4840 ^ n4837 ;
  assign n5022 = n4839 ^ x143 ;
  assign n5024 = n5023 ^ n5022 ;
  assign n5025 = ~n5021 & n5024 ;
  assign n5026 = n5025 ^ x142 ;
  assign n5020 = n4866 ^ n4865 ;
  assign n5027 = n5026 ^ n5020 ;
  assign n5028 = n5027 ^ x141 ;
  assign n5029 = n5028 ^ n5020 ;
  assign n5030 = n5026 ^ n4865 ;
  assign n5031 = n5030 ^ n5020 ;
  assign n5032 = ~n5029 & ~n5031 ;
  assign n5033 = n5032 ^ n5020 ;
  assign n5034 = ~n5019 & ~n5033 ;
  assign n5035 = n5034 ^ x140 ;
  assign n5016 = n5015 ^ n4912 ;
  assign n5038 = n5016 ^ n4918 ;
  assign n5039 = n5038 ^ n5016 ;
  assign n5040 = n5035 & ~n5039 ;
  assign n5041 = ~n5015 & n5040 ;
  assign n5042 = n5041 ^ n5015 ;
  assign n5017 = n5016 ^ n5015 ;
  assign n5043 = n5042 ^ n5017 ;
  assign n5044 = n5009 & ~n5043 ;
  assign n5046 = n5045 ^ n5044 ;
  assign n5047 = ~n5008 & n5046 ;
  assign n5048 = n5047 ^ x136 ;
  assign n5054 = n5053 ^ n5048 ;
  assign n5055 = n5054 ^ n5053 ;
  assign n5056 = n5005 & ~n5052 ;
  assign n5059 = n5055 & n5056 ;
  assign n5060 = n5059 ^ n5053 ;
  assign n5061 = ~n4996 & n5060 ;
  assign n5062 = n5061 ^ x133 ;
  assign n5063 = ~n5007 & ~n5062 ;
  assign n5091 = n5080 ^ n5063 ;
  assign n5092 = ~n5081 & ~n5091 ;
  assign n5093 = n5092 ^ x132 ;
  assign n5126 = n5112 ^ n5093 ;
  assign n5127 = ~n5113 & n5126 ;
  assign n5128 = n5127 ^ x131 ;
  assign n5178 = n5143 ^ n5128 ;
  assign n5179 = n5144 & ~n5178 ;
  assign n5180 = n5179 ^ x130 ;
  assign n5176 = n5175 ^ n5163 ;
  assign n5187 = n5180 ^ n5176 ;
  assign n5188 = n5180 ^ x129 ;
  assign n5189 = ~n5187 & n5188 ;
  assign n5206 = n5205 ^ n5189 ;
  assign n5207 = n5206 ^ n3709 ;
  assign n5208 = n5207 ^ n3688 ;
  assign n5209 = n5208 ^ n5206 ;
  assign n5210 = n4609 & ~n5209 ;
  assign n5211 = n5210 ^ n5207 ;
  assign n5177 = n5176 ^ x129 ;
  assign n5181 = n5180 ^ n5177 ;
  assign n5160 = n3989 ^ n3711 ;
  assign n5161 = ~n4599 & ~n5160 ;
  assign n5162 = n5161 ^ n3711 ;
  assign n5182 = n5181 ^ n5162 ;
  assign n5145 = n5144 ^ n5128 ;
  assign n5123 = n4064 ^ n3712 ;
  assign n5124 = ~n4569 & ~n5123 ;
  assign n5125 = n5124 ^ n3712 ;
  assign n5146 = n5145 ^ n5125 ;
  assign n4700 = n4071 ^ n3715 ;
  assign n4701 = ~n3990 & ~n4700 ;
  assign n4702 = n4701 ^ n3715 ;
  assign n5082 = n5081 ^ n5063 ;
  assign n5085 = n4702 & n5082 ;
  assign n5086 = n5085 ^ n3718 ;
  assign n5087 = n5086 ^ n4068 ;
  assign n5088 = n5087 ^ n5085 ;
  assign n5089 = ~n3986 & n5088 ;
  assign n5090 = n5089 ^ n5086 ;
  assign n5114 = n5113 ^ n5093 ;
  assign n5120 = n5114 ^ n5085 ;
  assign n5121 = n5090 & ~n5120 ;
  assign n5122 = n5121 ^ n5085 ;
  assign n5157 = n5125 ^ n5122 ;
  assign n5158 = n5146 & ~n5157 ;
  assign n5159 = n5158 ^ n5145 ;
  assign n5212 = n5162 ^ n5159 ;
  assign n5213 = n5182 & ~n5212 ;
  assign n5214 = n5213 ^ n5181 ;
  assign n5293 = n5214 ^ n5206 ;
  assign n5294 = ~n5211 & ~n5293 ;
  assign n5295 = n5294 ^ n5214 ;
  assign n5299 = n5298 ^ n5295 ;
  assign n5300 = n4581 ^ x159 ;
  assign n5301 = n5300 ^ n5298 ;
  assign n5302 = n5299 & n5301 ;
  assign n5303 = n5302 ^ n5300 ;
  assign n5307 = n5306 ^ n5303 ;
  assign n5308 = n4641 ^ n4638 ;
  assign n5309 = n5308 ^ n5306 ;
  assign n5310 = ~n5307 & ~n5309 ;
  assign n5311 = n5310 ^ n5308 ;
  assign n5314 = n5313 ^ n5311 ;
  assign n5315 = n5313 ^ n3705 ;
  assign n5316 = n5315 ^ n4052 ;
  assign n5317 = n5316 ^ n5313 ;
  assign n5318 = n4712 & ~n5317 ;
  assign n5319 = n5318 ^ n5315 ;
  assign n5320 = ~n5314 & n5319 ;
  assign n5321 = n5320 ^ n5313 ;
  assign n5396 = n5395 ^ n5321 ;
  assign n5398 = n5396 ^ n3309 ;
  assign n5386 = n5309 ^ n5303 ;
  assign n5378 = n5301 ^ n5295 ;
  assign n5379 = n5378 ^ n3303 ;
  assign n5215 = n5214 ^ n5211 ;
  assign n5216 = n5215 ^ n3263 ;
  assign n5183 = n5182 ^ n5159 ;
  assign n5184 = n5183 ^ n3264 ;
  assign n5147 = n5146 ^ n5122 ;
  assign n5148 = n5147 ^ n3265 ;
  assign n5083 = n5082 ^ n4702 ;
  assign n5116 = ~n3297 & n5083 ;
  assign n5117 = n5116 ^ n3266 ;
  assign n5115 = n5114 ^ n5090 ;
  assign n5149 = n5116 ^ n5115 ;
  assign n5150 = n5117 & n5149 ;
  assign n5151 = n5150 ^ n3266 ;
  assign n5154 = n5151 ^ n5147 ;
  assign n5155 = ~n5148 & ~n5154 ;
  assign n5156 = n5155 ^ n3265 ;
  assign n5217 = n5183 ^ n5156 ;
  assign n5218 = n5184 & n5217 ;
  assign n5219 = n5218 ^ n3264 ;
  assign n5380 = n5219 ^ n5215 ;
  assign n5381 = ~n5216 & ~n5380 ;
  assign n5382 = n5381 ^ n3263 ;
  assign n5383 = n5382 ^ n5378 ;
  assign n5384 = ~n5379 & n5383 ;
  assign n5385 = n5384 ^ n3303 ;
  assign n5387 = n5386 ^ n5385 ;
  assign n5388 = n5386 ^ n3305 ;
  assign n5389 = n5387 & ~n5388 ;
  assign n5390 = n5389 ^ n3305 ;
  assign n5377 = n5319 ^ n5311 ;
  assign n5391 = n5390 ^ n5377 ;
  assign n5392 = n5390 ^ n3307 ;
  assign n5393 = n5391 & ~n5392 ;
  assign n5394 = n5393 ^ n3307 ;
  assign n5552 = n5398 ^ n5394 ;
  assign n5542 = n5377 ^ n3307 ;
  assign n5543 = n5542 ^ n5390 ;
  assign n5544 = n5382 ^ n5379 ;
  assign n5084 = n5083 ^ n3297 ;
  assign n5118 = n5117 ^ n5115 ;
  assign n5119 = ~n5084 & ~n5118 ;
  assign n5152 = n5151 ^ n5148 ;
  assign n5153 = n5119 & ~n5152 ;
  assign n5185 = n5184 ^ n5156 ;
  assign n5186 = ~n5153 & n5185 ;
  assign n5220 = n5219 ^ n5216 ;
  assign n5545 = n5186 & n5220 ;
  assign n5546 = n5544 & ~n5545 ;
  assign n5547 = n5388 ^ n5385 ;
  assign n5548 = n5547 ^ n5546 ;
  assign n5549 = n5546 & ~n5548 ;
  assign n5550 = n5549 ^ n5543 ;
  assign n5551 = n5543 & n5550 ;
  assign n5603 = n5552 ^ n5551 ;
  assign n5605 = x183 & n5603 ;
  assign n5604 = n5603 ^ x183 ;
  assign n5606 = n5605 ^ n5604 ;
  assign n5553 = n5551 & ~n5552 ;
  assign n5322 = n5321 ^ n5292 ;
  assign n5324 = n5323 ^ n5321 ;
  assign n5325 = ~n5322 & ~n5324 ;
  assign n5326 = n5325 ^ n5323 ;
  assign n5287 = n4634 ^ x155 ;
  assign n5288 = n5287 ^ n4650 ;
  assign n5284 = n4046 ^ n3702 ;
  assign n5285 = ~n4725 & n5284 ;
  assign n5286 = n5285 ^ n3702 ;
  assign n5289 = n5288 ^ n5286 ;
  assign n5376 = n5326 ^ n5289 ;
  assign n5540 = n5376 ^ n3262 ;
  assign n5397 = n5396 ^ n5394 ;
  assign n5399 = ~n5397 & n5398 ;
  assign n5400 = n5399 ^ n3309 ;
  assign n5541 = n5540 ^ n5400 ;
  assign n5607 = n5553 ^ n5541 ;
  assign n5608 = ~x182 & ~n5607 ;
  assign n5609 = n5606 & n5608 ;
  assign n5610 = n5609 ^ n5606 ;
  assign n5581 = n5550 ^ x184 ;
  assign n5582 = n5548 ^ x185 ;
  assign n5583 = n5545 ^ n5544 ;
  assign n5584 = n5583 ^ x186 ;
  assign n5223 = n5185 ^ n5153 ;
  assign n5224 = n5223 ^ x188 ;
  assign n5225 = x191 & n5084 ;
  assign n5226 = n5225 ^ x190 ;
  assign n5227 = n5118 ^ n5084 ;
  assign n5228 = n5227 ^ n5225 ;
  assign n5229 = n5226 & ~n5228 ;
  assign n5230 = n5229 ^ x190 ;
  assign n5231 = n5230 ^ x189 ;
  assign n5232 = n5152 ^ n5119 ;
  assign n5233 = n5232 ^ n5230 ;
  assign n5234 = n5231 & n5233 ;
  assign n5235 = n5234 ^ x189 ;
  assign n5236 = n5235 ^ n5223 ;
  assign n5237 = n5224 & ~n5236 ;
  assign n5238 = n5237 ^ x188 ;
  assign n5221 = n5220 ^ n5186 ;
  assign n5586 = n5238 ^ n5221 ;
  assign n5589 = n5583 ^ n5221 ;
  assign n5585 = n5583 ^ x187 ;
  assign n5590 = n5589 ^ n5585 ;
  assign n5591 = n5586 & ~n5590 ;
  assign n5592 = n5591 ^ n5585 ;
  assign n5593 = ~n5584 & n5592 ;
  assign n5594 = n5593 ^ x186 ;
  assign n5595 = n5594 ^ n5548 ;
  assign n5596 = n5582 & ~n5595 ;
  assign n5597 = n5596 ^ x185 ;
  assign n5598 = n5597 ^ n5550 ;
  assign n5599 = n5581 & ~n5598 ;
  assign n5600 = n5599 ^ x184 ;
  assign n5616 = n5607 ^ n5605 ;
  assign n5617 = n5607 ^ x182 ;
  assign n5618 = ~n5616 & n5617 ;
  assign n5619 = n5618 ^ x182 ;
  assign n5705 = n5600 & ~n5619 ;
  assign n5706 = n5610 & n5705 ;
  assign n5707 = n5706 ^ n5619 ;
  assign n5554 = ~n5541 & ~n5553 ;
  assign n5401 = n5400 ^ n5376 ;
  assign n5402 = n5400 ^ n3262 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = n5403 ^ n3262 ;
  assign n5327 = n5326 ^ n5286 ;
  assign n5328 = n5289 & n5327 ;
  assign n5329 = n5328 ^ n5288 ;
  assign n5280 = n4043 ^ n3701 ;
  assign n5281 = n4745 & n5280 ;
  assign n5282 = n5281 ^ n3701 ;
  assign n5279 = n4654 ^ n4633 ;
  assign n5283 = n5282 ^ n5279 ;
  assign n5374 = n5329 ^ n5283 ;
  assign n5375 = n5374 ^ n3261 ;
  assign n5539 = n5404 ^ n5375 ;
  assign n5601 = n5554 ^ n5539 ;
  assign n5602 = n5601 ^ x181 ;
  assign n6181 = n5707 ^ n5602 ;
  assign n6171 = x183 ^ x182 ;
  assign n6172 = n6171 ^ n5607 ;
  assign n6168 = n5603 ^ n5600 ;
  assign n6169 = n5600 ^ x183 ;
  assign n6170 = ~n6168 & n6169 ;
  assign n6173 = n6172 ^ n6170 ;
  assign n6182 = n6181 ^ n6173 ;
  assign n5718 = n5604 ^ n5600 ;
  assign n6174 = n6173 ^ n5718 ;
  assign n5439 = x147 ^ x146 ;
  assign n5440 = n5439 ^ n4770 ;
  assign n5247 = n4663 & ~n4801 ;
  assign n5248 = ~n4766 & n5247 ;
  assign n5249 = n5248 ^ n4766 ;
  assign n5437 = n5249 ^ n4767 ;
  assign n5438 = n4778 & ~n5437 ;
  assign n5441 = n5440 ^ n5438 ;
  assign n5719 = n5718 ^ n4034 ;
  assign n5720 = n5719 ^ n4877 ;
  assign n5721 = n5720 ^ n5718 ;
  assign n5722 = ~n5441 & ~n5721 ;
  assign n5723 = n5722 ^ n5719 ;
  assign n5727 = n5597 ^ n5581 ;
  assign n5250 = n5249 ^ n4778 ;
  assign n5724 = n4862 ^ n4037 ;
  assign n5725 = n5250 & n5724 ;
  assign n5726 = n5725 ^ n4037 ;
  assign n5728 = n5727 ^ n5726 ;
  assign n5732 = n5594 ^ n5582 ;
  assign n4664 = ~n4626 & n4663 ;
  assign n4665 = ~n4622 & n4664 ;
  assign n4666 = n4665 ^ n4626 ;
  assign n4680 = n4679 ^ n4666 ;
  assign n4695 = n4694 ^ x149 ;
  assign n4696 = n4695 ^ n4694 ;
  assign n4697 = n4696 ^ n4666 ;
  assign n4698 = n4680 & n4697 ;
  assign n4699 = n4698 ^ n4695 ;
  assign n5729 = n4851 ^ n4040 ;
  assign n5730 = ~n4699 & n5729 ;
  assign n5731 = n5730 ^ n4040 ;
  assign n5733 = n5732 ^ n5731 ;
  assign n5345 = n4679 ^ x149 ;
  assign n5346 = n5345 ^ n4666 ;
  assign n5739 = n4829 ^ n4043 ;
  assign n5740 = ~n5346 & ~n5739 ;
  assign n5741 = n5740 ^ n4043 ;
  assign n5734 = n5584 ^ x187 ;
  assign n5735 = n5734 ^ n5584 ;
  assign n5736 = n5735 ^ n5221 ;
  assign n5737 = n5586 & ~n5736 ;
  assign n5738 = n5737 ^ n5734 ;
  assign n5742 = n5741 ^ n5738 ;
  assign n5258 = n4663 ^ n4603 ;
  assign n5259 = ~n4604 & n5258 ;
  assign n5256 = x151 ^ x150 ;
  assign n5257 = n5256 ^ n4619 ;
  assign n5260 = n5259 ^ n5257 ;
  assign n5743 = n4821 ^ n4046 ;
  assign n5744 = ~n5260 & ~n5743 ;
  assign n5745 = n5744 ^ n4046 ;
  assign n5222 = n5221 ^ x187 ;
  assign n5239 = n5238 ^ n5222 ;
  assign n5746 = n5745 ^ n5239 ;
  assign n5750 = n5235 ^ n5224 ;
  assign n5268 = n4663 ^ n4604 ;
  assign n5747 = n4745 ^ n4049 ;
  assign n5748 = ~n5268 & n5747 ;
  assign n5749 = n5748 ^ n4049 ;
  assign n5751 = n5750 ^ n5749 ;
  assign n5270 = n4660 ^ n4629 ;
  assign n5754 = n4725 ^ n4052 ;
  assign n5755 = ~n5270 & ~n5754 ;
  assign n5756 = n5755 ^ n4052 ;
  assign n5752 = n5232 ^ x189 ;
  assign n5753 = n5752 ^ n5230 ;
  assign n5757 = n5756 ^ n5753 ;
  assign n6139 = n5227 ^ n5226 ;
  assign n6130 = n5084 ^ x191 ;
  assign n5686 = n4809 & n4943 ;
  assign n5687 = ~n5048 & n5686 ;
  assign n5688 = n5687 ^ n5048 ;
  assign n5773 = n5688 ^ n5000 ;
  assign n5770 = n4121 ^ n3636 ;
  assign n5771 = n4535 & n5770 ;
  assign n5772 = n5771 ^ n3636 ;
  assign n5774 = n5773 ^ n5772 ;
  assign n5785 = n4124 ^ n3624 ;
  assign n5786 = n4550 & n5785 ;
  assign n5787 = n5786 ^ n3624 ;
  assign n5775 = ~n4873 & ~n5035 ;
  assign n5776 = ~n5015 & ~n5775 ;
  assign n5777 = ~n4918 & n5776 ;
  assign n5778 = n5777 ^ n5015 ;
  assign n5779 = n5778 ^ n4912 ;
  assign n5780 = n5008 ^ x137 ;
  assign n5781 = n5780 ^ n5008 ;
  assign n5782 = n5781 ^ n5778 ;
  assign n5783 = ~n5779 & n5782 ;
  assign n5784 = n5783 ^ n5780 ;
  assign n5788 = n5787 ^ n5784 ;
  assign n5795 = n4866 ^ x141 ;
  assign n5792 = n4809 & ~n5026 ;
  assign n5793 = ~n4843 & n5792 ;
  assign n5794 = n5793 ^ n5026 ;
  assign n5796 = n5795 ^ n5794 ;
  assign n5789 = n4015 ^ n3999 ;
  assign n5790 = ~n5101 & ~n5789 ;
  assign n5791 = n5790 ^ n4015 ;
  assign n5797 = n5796 ^ n5791 ;
  assign n5672 = n4005 ^ n3971 ;
  assign n5673 = n4952 & n5672 ;
  assign n5674 = n5673 ^ n3971 ;
  assign n5461 = n4783 & n5249 ;
  assign n5462 = n5461 ^ n4773 ;
  assign n5520 = n5462 ^ n4774 ;
  assign n5521 = n4757 ^ x145 ;
  assign n5522 = n5521 ^ n4757 ;
  assign n5523 = n5522 ^ n5462 ;
  assign n5524 = n5520 & n5523 ;
  assign n5525 = n5524 ^ n5521 ;
  assign n5526 = n4008 ^ n3952 ;
  assign n5527 = n4956 & n5526 ;
  assign n5528 = n5527 ^ n3952 ;
  assign n5667 = ~n5525 & ~n5528 ;
  assign n5803 = n5674 ^ n5667 ;
  assign n5671 = n5022 ^ n4809 ;
  assign n5804 = n5671 ^ n5667 ;
  assign n5805 = n5803 & n5804 ;
  assign n5806 = n5805 ^ n5674 ;
  assign n5798 = n4019 ^ n4002 ;
  assign n5799 = n5067 & ~n5798 ;
  assign n5800 = n5799 ^ n4019 ;
  assign n5801 = n5800 ^ n5796 ;
  assign n5697 = n4839 ^ n4809 ;
  assign n5698 = n5021 ^ x143 ;
  assign n5699 = n5698 ^ n4839 ;
  assign n5700 = n5699 ^ n5021 ;
  assign n5701 = n5697 & ~n5700 ;
  assign n5702 = n5701 ^ n5698 ;
  assign n5802 = n5801 ^ n5702 ;
  assign n5807 = n5806 ^ n5802 ;
  assign n5808 = n5807 ^ n5801 ;
  assign n5809 = n5791 ^ n5702 ;
  assign n5810 = n5809 ^ n5801 ;
  assign n5811 = n5808 & ~n5810 ;
  assign n5812 = n5811 ^ n5801 ;
  assign n5813 = ~n5797 & ~n5812 ;
  assign n5814 = n5813 ^ n5796 ;
  assign n5529 = n5528 ^ n5525 ;
  assign n5668 = n5667 ^ n5529 ;
  assign n5815 = n5671 & ~n5674 ;
  assign n5816 = n5668 & ~n5815 ;
  assign n5817 = ~n5791 & n5796 ;
  assign n5818 = n5816 & n5817 ;
  assign n5819 = n5818 ^ n5816 ;
  assign n5820 = ~n5800 & n5819 ;
  assign n5821 = n5702 & n5820 ;
  assign n5822 = n5821 ^ n5819 ;
  assign n5261 = n4031 ^ n3696 ;
  assign n5262 = ~n4862 & n5261 ;
  assign n5263 = n5262 ^ n3696 ;
  assign n5264 = n5263 ^ n5260 ;
  assign n5265 = n4034 ^ n3698 ;
  assign n5266 = n4851 & ~n5265 ;
  assign n5267 = n5266 ^ n3698 ;
  assign n5269 = n5268 ^ n5267 ;
  assign n5271 = n4037 ^ n3699 ;
  assign n5272 = ~n4829 & n5271 ;
  assign n5273 = n5272 ^ n3699 ;
  assign n5274 = n5273 ^ n5270 ;
  assign n5275 = n4040 ^ n3700 ;
  assign n5276 = n4821 & n5275 ;
  assign n5277 = n5276 ^ n3700 ;
  assign n5240 = n4657 ^ n4631 ;
  assign n5278 = n5277 ^ n5240 ;
  assign n5330 = n5329 ^ n5282 ;
  assign n5331 = ~n5283 & ~n5330 ;
  assign n5332 = n5331 ^ n5329 ;
  assign n5333 = n5332 ^ n5277 ;
  assign n5334 = n5278 & n5333 ;
  assign n5335 = n5334 ^ n5240 ;
  assign n5336 = n5335 ^ n5270 ;
  assign n5337 = n5274 & n5336 ;
  assign n5338 = n5337 ^ n5273 ;
  assign n5339 = n5338 ^ n5267 ;
  assign n5340 = ~n5269 & n5339 ;
  assign n5341 = n5340 ^ n5268 ;
  assign n5342 = n5341 ^ n5260 ;
  assign n5343 = n5264 & ~n5342 ;
  assign n5344 = n5343 ^ n5263 ;
  assign n5347 = n5346 ^ n5344 ;
  assign n5348 = n5346 ^ n3743 ;
  assign n5349 = n5348 ^ n4027 ;
  assign n5350 = n5349 ^ n5346 ;
  assign n5351 = n4877 & n5350 ;
  assign n5352 = n5351 ^ n5348 ;
  assign n5353 = n5347 & ~n5352 ;
  assign n5354 = n5353 ^ n5346 ;
  assign n5823 = n5814 ^ n5354 ;
  assign n5824 = n5823 ^ n5822 ;
  assign n5460 = n4774 ^ x145 ;
  assign n5463 = n5462 ^ n5460 ;
  assign n5457 = n4013 ^ n3942 ;
  assign n5458 = ~n4972 & n5457 ;
  assign n5459 = n5458 ^ n3942 ;
  assign n5464 = n5463 ^ n5459 ;
  assign n5434 = n4017 ^ n3787 ;
  assign n5435 = n4932 & ~n5434 ;
  assign n5436 = n5435 ^ n3787 ;
  assign n5499 = n5459 ^ n5436 ;
  assign n5500 = n5499 ^ n5441 ;
  assign n5244 = n4021 ^ n3693 ;
  assign n5245 = n4902 & ~n5244 ;
  assign n5246 = n5245 ^ n3693 ;
  assign n5251 = n5250 ^ n5246 ;
  assign n5252 = n4024 ^ n3694 ;
  assign n5253 = ~n4885 & ~n5252 ;
  assign n5254 = n5253 ^ n3694 ;
  assign n5255 = ~n4699 & n5254 ;
  assign n5427 = n5255 ^ n5250 ;
  assign n5428 = n5251 & n5427 ;
  assign n5429 = n5428 ^ n5255 ;
  assign n5501 = n5500 ^ n5429 ;
  assign n5502 = n5501 ^ n5499 ;
  assign n5503 = n5459 ^ n5441 ;
  assign n5504 = n5503 ^ n5499 ;
  assign n5505 = n5502 & ~n5504 ;
  assign n5506 = n5505 ^ n5499 ;
  assign n5507 = n5464 & n5506 ;
  assign n5508 = n5507 ^ n5463 ;
  assign n5825 = n5508 ^ n5354 ;
  assign n5826 = n5825 ^ n5822 ;
  assign n5355 = n5254 ^ n4699 ;
  assign n5356 = n5355 ^ n5255 ;
  assign n5430 = n5246 & ~n5250 ;
  assign n5509 = ~n5356 & ~n5430 ;
  assign n5510 = n5459 & n5509 ;
  assign n5511 = n5463 & n5510 ;
  assign n5512 = n5511 ^ n5509 ;
  assign n5513 = n5441 & n5512 ;
  assign n5514 = n5511 ^ n5436 ;
  assign n5515 = n5513 & ~n5514 ;
  assign n5516 = n5515 ^ n5512 ;
  assign n5827 = n5516 ^ n5508 ;
  assign n5828 = n5827 ^ n5814 ;
  assign n5829 = ~n5826 & n5828 ;
  assign n5830 = ~n5824 & n5829 ;
  assign n5831 = n5830 ^ n5508 ;
  assign n5832 = n5831 ^ n5814 ;
  assign n5833 = n5822 & n5832 ;
  assign n5834 = n5814 & n5833 ;
  assign n5835 = n5834 ^ n5814 ;
  assign n5836 = n4218 ^ n4010 ;
  assign n5837 = ~n5130 & ~n5836 ;
  assign n5838 = n5837 ^ n4010 ;
  assign n5839 = n5794 ^ n4866 ;
  assign n5840 = n5019 ^ x141 ;
  assign n5841 = n5840 ^ n5019 ;
  assign n5842 = n5841 ^ n5794 ;
  assign n5843 = n5839 & n5842 ;
  assign n5844 = n5843 ^ n5840 ;
  assign n5845 = ~n5838 & n5844 ;
  assign n5846 = ~n5835 & ~n5845 ;
  assign n5853 = n3978 ^ n3592 ;
  assign n5854 = n5197 & n5853 ;
  assign n5855 = n5854 ^ n3592 ;
  assign n5847 = n5775 ^ n4914 ;
  assign n5848 = n5010 ^ x139 ;
  assign n5849 = n5848 ^ n5010 ;
  assign n5850 = n5849 ^ n5775 ;
  assign n5851 = ~n5847 & ~n5850 ;
  assign n5852 = n5851 ^ n5848 ;
  assign n5856 = n5855 ^ n5852 ;
  assign n5857 = n3964 ^ n3610 ;
  assign n5858 = n5164 & ~n5857 ;
  assign n5859 = n5858 ^ n3610 ;
  assign n5860 = n5775 ^ n5012 ;
  assign n5861 = n5859 & ~n5860 ;
  assign n5865 = n5778 ^ n5009 ;
  assign n5862 = n4127 ^ n3606 ;
  assign n5863 = ~n4540 & ~n5862 ;
  assign n5864 = n5863 ^ n3606 ;
  assign n5866 = n5865 ^ n5864 ;
  assign n5867 = ~n5861 & n5866 ;
  assign n5868 = ~n5845 & n5867 ;
  assign n5869 = n5856 & n5868 ;
  assign n5870 = n5846 & n5869 ;
  assign n5877 = n5865 ^ n5855 ;
  assign n5871 = n5860 ^ n5859 ;
  assign n5872 = n5844 ^ n5838 ;
  assign n5873 = n5872 ^ n5845 ;
  assign n5874 = n5873 ^ n5860 ;
  assign n5875 = ~n5871 & ~n5874 ;
  assign n5876 = n5875 ^ n5859 ;
  assign n5878 = n5877 ^ n5876 ;
  assign n5879 = n5878 ^ n5852 ;
  assign n5880 = n5879 ^ n5877 ;
  assign n5881 = n5876 ^ n5864 ;
  assign n5882 = n5881 ^ n5877 ;
  assign n5883 = n5880 & n5882 ;
  assign n5884 = n5883 ^ n5877 ;
  assign n5885 = n5866 & n5884 ;
  assign n5886 = n5885 ^ n5865 ;
  assign n5887 = ~n5870 & ~n5886 ;
  assign n5888 = n5887 ^ n5787 ;
  assign n5889 = ~n5788 & n5888 ;
  assign n5890 = n5889 ^ n5887 ;
  assign n5891 = n5890 ^ n5772 ;
  assign n5892 = ~n5774 & ~n5891 ;
  assign n5893 = n5892 ^ n5773 ;
  assign n5766 = n4078 ^ n3666 ;
  assign n5767 = n4532 & ~n5766 ;
  assign n5768 = n5767 ^ n3666 ;
  assign n5763 = x135 ^ x134 ;
  assign n5764 = n5763 ^ n5002 ;
  assign n5761 = n5688 ^ n4998 ;
  assign n5762 = n5000 & ~n5761 ;
  assign n5765 = n5764 ^ n5762 ;
  assign n5769 = n5768 ^ n5765 ;
  assign n6034 = n5893 ^ n5769 ;
  assign n6086 = n6034 ^ x31 ;
  assign n5992 = n5890 ^ n5774 ;
  assign n5993 = n5992 ^ n3282 ;
  assign n5906 = n5872 ^ n5835 ;
  assign n5907 = ~n3633 & ~n5906 ;
  assign n5517 = ~n5354 & n5516 ;
  assign n5518 = n5508 & n5517 ;
  assign n5519 = n5518 ^ n5508 ;
  assign n5669 = ~n5519 & n5668 ;
  assign n5909 = n5669 & ~n5815 ;
  assign n5910 = ~n5806 & n5909 ;
  assign n5911 = n5910 ^ n5806 ;
  assign n5912 = n5911 ^ n5702 ;
  assign n5913 = n5911 ^ n5800 ;
  assign n5914 = n5912 & n5913 ;
  assign n5908 = n5800 ^ n5797 ;
  assign n5915 = n5914 ^ n5908 ;
  assign n5916 = n5915 ^ n3617 ;
  assign n5920 = n5915 ^ n3594 ;
  assign n5917 = n5800 ^ n5702 ;
  assign n5918 = n5917 ^ n5911 ;
  assign n5919 = n5918 ^ n5915 ;
  assign n5921 = n5920 ^ n5919 ;
  assign n5530 = n5529 ^ n5519 ;
  assign n5678 = ~n3568 & ~n5530 ;
  assign n5675 = n5674 ^ n5671 ;
  assign n5670 = ~n5667 & ~n5669 ;
  assign n5676 = n5675 ^ n5670 ;
  assign n5922 = n5678 ^ n5676 ;
  assign n5923 = n5678 ^ n3580 ;
  assign n5924 = ~n5922 & ~n5923 ;
  assign n5925 = n5924 ^ n3580 ;
  assign n5926 = n5925 ^ n5915 ;
  assign n5927 = n5926 ^ n5920 ;
  assign n5928 = ~n5921 & ~n5927 ;
  assign n5929 = n5928 ^ n5920 ;
  assign n5930 = ~n5916 & n5929 ;
  assign n5931 = n5930 ^ n3617 ;
  assign n5531 = n5530 ^ n3568 ;
  assign n5679 = n5678 ^ n5531 ;
  assign n5932 = n3580 & ~n5676 ;
  assign n5933 = n5679 & ~n5932 ;
  assign n5934 = ~n3617 & n5915 ;
  assign n5935 = n5933 & n5934 ;
  assign n5936 = n5935 ^ n5933 ;
  assign n5937 = ~n3594 & n5918 ;
  assign n5938 = n5936 & n5937 ;
  assign n5939 = n5938 ^ n5936 ;
  assign n5365 = n5352 ^ n5344 ;
  assign n5366 = n5365 ^ n3508 ;
  assign n5367 = n5341 ^ n5264 ;
  assign n5368 = n5367 ^ n3259 ;
  assign n5369 = n5338 ^ n5269 ;
  assign n5370 = n5369 ^ n3316 ;
  assign n5371 = n5335 ^ n5274 ;
  assign n5372 = n5371 ^ n3314 ;
  assign n5405 = n5404 ^ n5374 ;
  assign n5406 = ~n5375 & ~n5405 ;
  assign n5407 = n5406 ^ n3261 ;
  assign n5373 = n5332 ^ n5278 ;
  assign n5408 = n5407 ^ n5373 ;
  assign n5409 = n5407 ^ n3260 ;
  assign n5410 = n5408 & ~n5409 ;
  assign n5411 = n5410 ^ n3260 ;
  assign n5412 = n5411 ^ n5371 ;
  assign n5413 = n5372 & n5412 ;
  assign n5414 = n5413 ^ n3314 ;
  assign n5415 = n5414 ^ n5369 ;
  assign n5416 = ~n5370 & ~n5415 ;
  assign n5417 = n5416 ^ n3316 ;
  assign n5418 = n5417 ^ n5367 ;
  assign n5419 = n5368 & ~n5418 ;
  assign n5420 = n5419 ^ n3259 ;
  assign n5421 = n5420 ^ n5365 ;
  assign n5422 = n5366 & n5421 ;
  assign n5423 = n5422 ^ n3508 ;
  assign n5940 = n5931 ^ n5423 ;
  assign n5941 = n5940 ^ n5939 ;
  assign n5357 = ~n5354 & ~n5356 ;
  assign n5431 = n5357 & ~n5430 ;
  assign n5432 = ~n5429 & n5431 ;
  assign n5433 = n5432 ^ n5429 ;
  assign n5456 = n5436 ^ n5433 ;
  assign n5465 = n5464 ^ n5441 ;
  assign n5466 = n5465 ^ n5464 ;
  assign n5467 = n5466 ^ n5433 ;
  assign n5468 = ~n5456 & ~n5467 ;
  assign n5469 = n5468 ^ n5465 ;
  assign n5486 = n5469 ^ n3556 ;
  assign n5488 = n5469 ^ n3544 ;
  assign n5361 = n5355 ^ n5354 ;
  assign n5362 = ~n3520 & n5361 ;
  assign n5446 = n5362 ^ n3532 ;
  assign n5358 = ~n5255 & ~n5357 ;
  assign n5359 = n5358 ^ n5251 ;
  assign n5447 = n5362 ^ n5359 ;
  assign n5448 = ~n5446 & ~n5447 ;
  assign n5449 = n5448 ^ n3532 ;
  assign n5487 = n5469 ^ n5449 ;
  assign n5489 = n5488 ^ n5487 ;
  assign n5442 = n5441 ^ n5436 ;
  assign n5443 = n5442 ^ n5433 ;
  assign n5490 = n5469 ^ n5443 ;
  assign n5491 = n5490 ^ n5488 ;
  assign n5492 = n5489 & n5491 ;
  assign n5493 = n5492 ^ n5488 ;
  assign n5494 = ~n5486 & ~n5493 ;
  assign n5495 = n5494 ^ n3556 ;
  assign n5942 = n5495 ^ n5423 ;
  assign n5943 = n5942 ^ n5939 ;
  assign n5363 = n5361 ^ n3520 ;
  assign n5364 = n5363 ^ n5362 ;
  assign n5445 = n3532 & ~n5359 ;
  assign n5478 = ~n5364 & ~n5445 ;
  assign n5479 = ~n3556 & n5478 ;
  assign n5480 = n5469 & n5479 ;
  assign n5481 = n5480 ^ n5478 ;
  assign n5482 = n5443 & n5481 ;
  assign n5483 = n5480 ^ n3544 ;
  assign n5484 = n5482 & n5483 ;
  assign n5485 = n5484 ^ n5481 ;
  assign n5944 = n5495 ^ n5485 ;
  assign n5945 = n5944 ^ n5931 ;
  assign n5946 = ~n5943 & n5945 ;
  assign n5947 = ~n5941 & n5946 ;
  assign n5948 = n5947 ^ n5495 ;
  assign n5949 = n5948 ^ n5931 ;
  assign n5950 = n5939 & n5949 ;
  assign n5951 = ~n5931 & n5950 ;
  assign n5952 = n5951 ^ n5931 ;
  assign n5953 = ~n5907 & n5952 ;
  assign n5954 = n5846 & ~n5861 ;
  assign n5955 = n5876 & n5954 ;
  assign n5956 = n5955 ^ n5876 ;
  assign n5957 = n5956 ^ n5856 ;
  assign n5958 = n5957 ^ n3284 ;
  assign n5959 = ~n5846 & ~n5873 ;
  assign n5960 = n5959 ^ n5871 ;
  assign n5961 = ~n3361 & ~n5960 ;
  assign n5964 = n5956 ^ n5852 ;
  assign n5965 = ~n5856 & ~n5964 ;
  assign n5962 = n5956 ^ n5866 ;
  assign n5966 = n5965 ^ n5962 ;
  assign n5967 = n5966 ^ n3283 ;
  assign n5968 = ~n5907 & n5967 ;
  assign n5969 = ~n5961 & n5968 ;
  assign n5970 = ~n5958 & n5969 ;
  assign n5971 = n5953 & n5970 ;
  assign n5979 = n5966 ^ n5957 ;
  assign n5972 = n5906 ^ n3633 ;
  assign n5973 = n5972 ^ n5907 ;
  assign n5974 = n5973 ^ n5960 ;
  assign n5975 = n5973 ^ n3361 ;
  assign n5976 = n5974 & ~n5975 ;
  assign n5977 = n5976 ^ n3361 ;
  assign n5978 = n5977 ^ n5966 ;
  assign n5980 = n5979 ^ n5978 ;
  assign n5981 = n5966 ^ n3284 ;
  assign n5982 = n5981 ^ n5979 ;
  assign n5983 = ~n5980 & ~n5982 ;
  assign n5984 = n5983 ^ n5979 ;
  assign n5985 = n5967 & ~n5984 ;
  assign n5986 = n5985 ^ n3283 ;
  assign n5987 = ~n5971 & n5986 ;
  assign n5905 = n5887 ^ n5788 ;
  assign n5988 = n5987 ^ n5905 ;
  assign n5989 = n5987 ^ n3287 ;
  assign n5990 = ~n5988 & ~n5989 ;
  assign n5991 = n5990 ^ n3287 ;
  assign n6036 = n5992 ^ n5991 ;
  assign n6037 = ~n5993 & ~n6036 ;
  assign n6038 = n6037 ^ n3282 ;
  assign n6087 = n6086 ^ n6038 ;
  assign n5994 = n5993 ^ n5991 ;
  assign n5995 = n5953 & ~n5961 ;
  assign n5996 = ~n5977 & n5995 ;
  assign n5997 = n5996 ^ n5977 ;
  assign n5998 = n5997 ^ n5958 ;
  assign n6000 = n5960 ^ n3361 ;
  assign n5999 = ~n5953 & n5973 ;
  assign n6001 = n6000 ^ n5999 ;
  assign n6002 = n5972 ^ n5952 ;
  assign n5496 = n5485 & ~n5495 ;
  assign n5497 = n5423 & n5496 ;
  assign n5498 = n5497 ^ n5495 ;
  assign n5532 = n5531 ^ n5498 ;
  assign n5424 = ~n5364 & n5423 ;
  assign n5425 = ~n5362 & ~n5424 ;
  assign n5360 = n5359 ^ n3532 ;
  assign n5426 = n5425 ^ n5360 ;
  assign n5534 = n5420 ^ n5366 ;
  assign n5535 = n5417 ^ n5368 ;
  assign n5536 = n5414 ^ n5370 ;
  assign n5537 = n5373 ^ n3260 ;
  assign n5538 = n5537 ^ n5407 ;
  assign n5555 = n5539 & n5554 ;
  assign n5556 = n5555 ^ n5538 ;
  assign n5557 = ~n5538 & ~n5556 ;
  assign n5558 = n5411 ^ n5372 ;
  assign n5559 = n5557 & n5558 ;
  assign n5560 = n5536 & n5559 ;
  assign n5561 = n5535 & n5560 ;
  assign n5562 = n5561 ^ n5534 ;
  assign n5563 = ~n5534 & ~n5562 ;
  assign n5450 = ~n5445 & n5449 ;
  assign n5451 = n5424 & n5450 ;
  assign n5452 = n5451 ^ n5449 ;
  assign n5455 = n5452 ^ n5443 ;
  assign n5470 = n3556 ^ n3544 ;
  assign n5471 = n5470 ^ n5469 ;
  assign n5472 = n5471 ^ n3556 ;
  assign n5473 = n5472 ^ n5452 ;
  assign n5474 = n5473 ^ n5469 ;
  assign n5475 = ~n5455 & n5474 ;
  assign n5476 = n5475 ^ n5471 ;
  assign n5444 = n5443 ^ n3544 ;
  assign n5453 = n5452 ^ n5444 ;
  assign n5564 = n5423 ^ n5363 ;
  assign n5565 = ~n5453 & ~n5564 ;
  assign n5566 = n5476 & n5565 ;
  assign n5567 = n5563 & n5566 ;
  assign n5568 = ~n5426 & n5567 ;
  assign n5454 = n5426 & ~n5453 ;
  assign n5477 = n5454 & n5476 ;
  assign n5665 = n5568 ^ n5477 ;
  assign n5666 = n5532 & n5665 ;
  assign n5680 = n5498 & n5679 ;
  assign n5681 = ~n5678 & ~n5680 ;
  assign n5677 = n5676 ^ n3580 ;
  assign n5682 = n5681 ^ n5677 ;
  assign n6003 = n5666 & n5682 ;
  assign n6007 = n5918 ^ n3594 ;
  assign n6004 = n5925 & ~n5932 ;
  assign n6005 = n5680 & n6004 ;
  assign n6006 = n6005 ^ n5925 ;
  assign n6008 = n6007 ^ n6006 ;
  assign n6009 = n6008 ^ n6003 ;
  assign n6010 = n6003 & ~n6009 ;
  assign n6011 = n6006 ^ n5918 ;
  assign n6015 = n6006 ^ n3594 ;
  assign n6016 = ~n6011 & ~n6015 ;
  assign n6012 = n3617 ^ n3594 ;
  assign n6013 = n6012 ^ n5915 ;
  assign n6017 = n6016 ^ n6013 ;
  assign n6018 = ~n6010 & n6017 ;
  assign n6019 = n6002 & ~n6018 ;
  assign n6020 = n6001 & ~n6019 ;
  assign n6021 = ~n5998 & ~n6020 ;
  assign n6022 = n5997 ^ n5957 ;
  assign n6023 = n5967 ^ n3284 ;
  assign n6024 = n6023 ^ n5957 ;
  assign n6025 = n6024 ^ n5967 ;
  assign n6026 = n6022 & ~n6025 ;
  assign n6027 = n6026 ^ n6023 ;
  assign n6028 = ~n6021 & ~n6027 ;
  assign n6029 = n5905 ^ n3287 ;
  assign n6030 = n6029 ^ n5987 ;
  assign n6031 = n6028 & ~n6030 ;
  assign n6032 = n6031 ^ n5994 ;
  assign n6033 = ~n5994 & ~n6032 ;
  assign n6088 = n6087 ^ n6033 ;
  assign n6045 = n6032 ^ x162 ;
  assign n6046 = n6030 ^ n6028 ;
  assign n6047 = n6046 ^ x163 ;
  assign n6075 = n6027 ^ n6021 ;
  assign n6048 = n6020 ^ n5998 ;
  assign n6049 = n6048 ^ x165 ;
  assign n6050 = n6019 ^ n6001 ;
  assign n6051 = n6050 ^ x166 ;
  assign n6052 = n6018 ^ n6002 ;
  assign n6053 = n6052 ^ x167 ;
  assign n6054 = n6017 ^ n6010 ;
  assign n6055 = n6054 ^ x168 ;
  assign n6056 = n6009 ^ x169 ;
  assign n5683 = n5682 ^ n5666 ;
  assign n5684 = n5683 ^ x170 ;
  assign n5533 = n5532 ^ n5477 ;
  assign n5569 = n5568 ^ n5533 ;
  assign n5570 = n5569 ^ x171 ;
  assign n5571 = n5563 & ~n5564 ;
  assign n5572 = ~n5426 & ~n5571 ;
  assign n5573 = n5572 ^ n5453 ;
  assign n5574 = n5573 ^ x173 ;
  assign n5575 = n5571 ^ n5426 ;
  assign n5576 = n5575 ^ x174 ;
  assign n5577 = n5564 ^ n5563 ;
  assign n5578 = n5577 ^ x175 ;
  assign n5579 = n5560 ^ n5535 ;
  assign n5580 = n5579 ^ x177 ;
  assign n5635 = n5559 ^ n5536 ;
  assign n5630 = n5558 ^ n5557 ;
  assign n5611 = n5602 & n5610 ;
  assign n5612 = n5556 ^ x180 ;
  assign n5613 = n5611 & ~n5612 ;
  assign n5614 = n5600 & n5613 ;
  assign n5615 = n5601 ^ n5556 ;
  assign n5620 = n5619 ^ n5615 ;
  assign n5621 = n5620 ^ x181 ;
  assign n5622 = n5621 ^ n5615 ;
  assign n5623 = n5619 ^ n5556 ;
  assign n5624 = n5623 ^ n5615 ;
  assign n5625 = ~n5622 & n5624 ;
  assign n5626 = n5625 ^ n5615 ;
  assign n5627 = ~n5612 & n5626 ;
  assign n5628 = n5627 ^ x180 ;
  assign n5629 = ~n5614 & ~n5628 ;
  assign n5631 = n5630 ^ n5629 ;
  assign n5632 = n5630 ^ x179 ;
  assign n5633 = ~n5631 & ~n5632 ;
  assign n5634 = n5633 ^ x179 ;
  assign n5636 = n5635 ^ n5634 ;
  assign n5637 = n5635 ^ x178 ;
  assign n5638 = n5636 & ~n5637 ;
  assign n5639 = n5638 ^ x178 ;
  assign n5640 = n5639 ^ n5579 ;
  assign n5641 = ~n5580 & n5640 ;
  assign n5642 = n5641 ^ x177 ;
  assign n5643 = n5642 ^ n5562 ;
  assign n5644 = n5562 ^ x176 ;
  assign n5645 = ~n5643 & n5644 ;
  assign n5646 = n5645 ^ x176 ;
  assign n5647 = n5646 ^ n5577 ;
  assign n5648 = ~n5578 & n5647 ;
  assign n5649 = n5648 ^ x175 ;
  assign n5650 = n5649 ^ n5575 ;
  assign n5651 = ~n5576 & n5650 ;
  assign n5652 = n5651 ^ x174 ;
  assign n5653 = n5652 ^ n5573 ;
  assign n5654 = n5574 & ~n5653 ;
  assign n5655 = n5654 ^ x173 ;
  assign n5656 = n5655 ^ x172 ;
  assign n5657 = ~n5453 & ~n5572 ;
  assign n5658 = n5657 ^ n5476 ;
  assign n5659 = n5658 ^ n5655 ;
  assign n5660 = n5656 & ~n5659 ;
  assign n5661 = n5660 ^ x172 ;
  assign n5662 = n5661 ^ n5569 ;
  assign n5663 = n5570 & ~n5662 ;
  assign n5664 = n5663 ^ x171 ;
  assign n6057 = n5683 ^ n5664 ;
  assign n6058 = n5684 & ~n6057 ;
  assign n6059 = n6058 ^ x170 ;
  assign n6060 = n6059 ^ n6009 ;
  assign n6061 = n6056 & ~n6060 ;
  assign n6062 = n6061 ^ x169 ;
  assign n6063 = n6062 ^ n6054 ;
  assign n6064 = n6055 & ~n6063 ;
  assign n6065 = n6064 ^ x168 ;
  assign n6066 = n6065 ^ n6052 ;
  assign n6067 = ~n6053 & n6066 ;
  assign n6068 = n6067 ^ x167 ;
  assign n6069 = n6068 ^ n6050 ;
  assign n6070 = n6051 & ~n6069 ;
  assign n6071 = n6070 ^ x166 ;
  assign n6072 = n6071 ^ n6048 ;
  assign n6073 = n6049 & ~n6072 ;
  assign n6074 = n6073 ^ x165 ;
  assign n6076 = n6075 ^ n6074 ;
  assign n6077 = n6075 ^ x164 ;
  assign n6078 = n6076 & ~n6077 ;
  assign n6079 = n6078 ^ x164 ;
  assign n6080 = n6079 ^ n6046 ;
  assign n6081 = n6047 & ~n6080 ;
  assign n6082 = n6081 ^ x163 ;
  assign n6083 = n6082 ^ n6032 ;
  assign n6084 = n6045 & ~n6083 ;
  assign n6085 = n6084 ^ x162 ;
  assign n6089 = n6088 ^ n6085 ;
  assign n6090 = n6088 ^ x161 ;
  assign n6091 = ~n6089 & n6090 ;
  assign n6035 = n6034 ^ n6033 ;
  assign n6042 = n6038 ^ n6034 ;
  assign n6043 = n6035 & ~n6042 ;
  assign n6039 = n6038 ^ n6035 ;
  assign n6040 = ~x31 & ~n6039 ;
  assign n5901 = n4074 ^ n3676 ;
  assign n5902 = n4524 & n5901 ;
  assign n5899 = x161 ^ x160 ;
  assign n5690 = n5052 ^ n4996 ;
  assign n5689 = n5056 & n5688 ;
  assign n5691 = n5690 ^ n5689 ;
  assign n5896 = n5691 ^ n3676 ;
  assign n5897 = n5896 ^ n3243 ;
  assign n5898 = n5897 ^ n5768 ;
  assign n5900 = n5899 ^ n5898 ;
  assign n5903 = n5902 ^ n5900 ;
  assign n5894 = n5893 ^ n5765 ;
  assign n5895 = ~n5769 & ~n5894 ;
  assign n5904 = n5903 ^ n5895 ;
  assign n6041 = n6040 ^ n5904 ;
  assign n6044 = n6043 ^ n6041 ;
  assign n6092 = n6091 ^ n6044 ;
  assign n5758 = n4683 ^ n3688 ;
  assign n5759 = ~n5288 & ~n5758 ;
  assign n5760 = n5759 ^ n3688 ;
  assign n6093 = n6092 ^ n5760 ;
  assign n6097 = n6085 ^ x161 ;
  assign n6098 = n6097 ^ n6088 ;
  assign n6094 = n4673 ^ n3989 ;
  assign n6095 = n5323 & n6094 ;
  assign n6096 = n6095 ^ n3989 ;
  assign n6099 = n6098 ^ n6096 ;
  assign n6102 = n4569 ^ n4071 ;
  assign n6103 = ~n5300 & n6102 ;
  assign n6104 = n6103 ^ n4071 ;
  assign n6105 = n6074 ^ x164 ;
  assign n6106 = n6105 ^ n6075 ;
  assign n6107 = ~n6104 & ~n6106 ;
  assign n6101 = n6079 ^ n6047 ;
  assign n6108 = n6107 ^ n6101 ;
  assign n6109 = n6107 ^ n4068 ;
  assign n6110 = n6109 ^ n4599 ;
  assign n6111 = n6110 ^ n6107 ;
  assign n6112 = n5308 & ~n6111 ;
  assign n6113 = n6112 ^ n6109 ;
  assign n6114 = n6108 & n6113 ;
  assign n6115 = n6114 ^ n6107 ;
  assign n6100 = n6082 ^ n6045 ;
  assign n6116 = n6115 ^ n6100 ;
  assign n6117 = n6100 ^ n4064 ;
  assign n6118 = n6117 ^ n4609 ;
  assign n6119 = n6118 ^ n6100 ;
  assign n6120 = ~n5313 & ~n6119 ;
  assign n6121 = n6120 ^ n6117 ;
  assign n6122 = n6116 & n6121 ;
  assign n6123 = n6122 ^ n6115 ;
  assign n6124 = n6123 ^ n6096 ;
  assign n6125 = ~n6099 & n6124 ;
  assign n6126 = n6125 ^ n6098 ;
  assign n6127 = n6126 ^ n5760 ;
  assign n6128 = n6093 & ~n6127 ;
  assign n6129 = n6128 ^ n6092 ;
  assign n6131 = n6130 ^ n6129 ;
  assign n6132 = n6130 ^ n4058 ;
  assign n6133 = n6132 ^ n4712 ;
  assign n6134 = n6133 ^ n6130 ;
  assign n6135 = n5279 & ~n6134 ;
  assign n6136 = n6135 ^ n6132 ;
  assign n6137 = n6131 & ~n6136 ;
  assign n6138 = n6137 ^ n6130 ;
  assign n6140 = n6139 ^ n6138 ;
  assign n6141 = n6139 ^ n4055 ;
  assign n6142 = n6141 ^ n4706 ;
  assign n6143 = n6142 ^ n6139 ;
  assign n6144 = n5240 & n6143 ;
  assign n6145 = n6144 ^ n6141 ;
  assign n6146 = n6140 & n6145 ;
  assign n6147 = n6146 ^ n6139 ;
  assign n6148 = n6147 ^ n5753 ;
  assign n6149 = ~n5757 & n6148 ;
  assign n6150 = n6149 ^ n5756 ;
  assign n6151 = n6150 ^ n5749 ;
  assign n6152 = n5751 & ~n6151 ;
  assign n6153 = n6152 ^ n5750 ;
  assign n6154 = n6153 ^ n5239 ;
  assign n6155 = n5746 & n6154 ;
  assign n6156 = n6155 ^ n5745 ;
  assign n6157 = n6156 ^ n5738 ;
  assign n6158 = ~n5742 & ~n6157 ;
  assign n6159 = n6158 ^ n5741 ;
  assign n6160 = n6159 ^ n5731 ;
  assign n6161 = n5733 & ~n6160 ;
  assign n6162 = n6161 ^ n5732 ;
  assign n6163 = n6162 ^ n5726 ;
  assign n6164 = ~n5728 & n6163 ;
  assign n6165 = n6164 ^ n5727 ;
  assign n6166 = n6165 ^ n5718 ;
  assign n6167 = ~n5723 & n6166 ;
  assign n6175 = n6174 ^ n6167 ;
  assign n6176 = n4885 ^ n4031 ;
  assign n6177 = ~n5463 & n6176 ;
  assign n6178 = n6177 ^ n4031 ;
  assign n6179 = n6178 ^ n6173 ;
  assign n6180 = n6175 & ~n6179 ;
  assign n6183 = n6182 ^ n6180 ;
  assign n5708 = n5707 ^ n5601 ;
  assign n5709 = n5612 ^ x181 ;
  assign n5710 = n5709 ^ n5612 ;
  assign n5711 = n5710 ^ n5707 ;
  assign n5712 = ~n5708 & n5711 ;
  assign n5713 = n5712 ^ n5709 ;
  assign n6187 = n6181 ^ n5713 ;
  assign n6184 = n4902 ^ n4027 ;
  assign n6185 = ~n5525 & n6184 ;
  assign n6186 = n6185 ^ n4027 ;
  assign n6188 = n6187 ^ n6186 ;
  assign n6189 = n6188 ^ n5713 ;
  assign n6190 = n6183 & n6189 ;
  assign n6191 = n6190 ^ n6187 ;
  assign n5714 = n4932 ^ n4024 ;
  assign n5715 = ~n5671 & ~n5714 ;
  assign n5716 = n5715 ^ n4024 ;
  assign n6293 = n6191 ^ n5716 ;
  assign n6294 = n6293 ^ n3694 ;
  assign n6367 = n6186 ^ n6183 ;
  assign n6295 = n6178 ^ n6175 ;
  assign n6296 = n6295 ^ n3696 ;
  assign n6355 = n6162 ^ n5728 ;
  assign n6298 = n6159 ^ n5733 ;
  assign n6299 = n6298 ^ n3700 ;
  assign n6347 = n6156 ^ n5742 ;
  assign n6300 = n6153 ^ n5746 ;
  assign n6301 = n6300 ^ n3702 ;
  assign n6339 = n6150 ^ n5751 ;
  assign n6302 = n6147 ^ n5757 ;
  assign n6303 = n6302 ^ n3705 ;
  assign n6304 = n6145 ^ n6138 ;
  assign n6305 = n6304 ^ n3689 ;
  assign n6328 = n6136 ^ n6129 ;
  assign n6306 = n6126 ^ n6093 ;
  assign n6307 = n6306 ^ n3709 ;
  assign n6320 = n6123 ^ n6099 ;
  assign n6310 = n6106 ^ n6104 ;
  assign n6311 = n3715 & n6310 ;
  assign n6309 = n6113 ^ n6101 ;
  assign n6312 = n6311 ^ n6309 ;
  assign n6313 = n6311 ^ n3718 ;
  assign n6314 = ~n6312 & n6313 ;
  assign n6315 = n6314 ^ n3718 ;
  assign n6308 = n6121 ^ n6115 ;
  assign n6316 = n6315 ^ n6308 ;
  assign n6317 = n6315 ^ n3712 ;
  assign n6318 = n6316 & n6317 ;
  assign n6319 = n6318 ^ n3712 ;
  assign n6321 = n6320 ^ n6319 ;
  assign n6322 = n6320 ^ n3711 ;
  assign n6323 = n6321 & ~n6322 ;
  assign n6324 = n6323 ^ n3711 ;
  assign n6325 = n6324 ^ n6306 ;
  assign n6326 = ~n6307 & ~n6325 ;
  assign n6327 = n6326 ^ n3709 ;
  assign n6329 = n6328 ^ n6327 ;
  assign n6330 = n6328 ^ n3707 ;
  assign n6331 = ~n6329 & n6330 ;
  assign n6332 = n6331 ^ n3707 ;
  assign n6333 = n6332 ^ n6304 ;
  assign n6334 = ~n6305 & n6333 ;
  assign n6335 = n6334 ^ n3689 ;
  assign n6336 = n6335 ^ n6302 ;
  assign n6337 = n6303 & ~n6336 ;
  assign n6338 = n6337 ^ n3705 ;
  assign n6340 = n6339 ^ n6338 ;
  assign n6341 = n6339 ^ n3703 ;
  assign n6342 = n6340 & ~n6341 ;
  assign n6343 = n6342 ^ n3703 ;
  assign n6344 = n6343 ^ n6300 ;
  assign n6345 = ~n6301 & n6344 ;
  assign n6346 = n6345 ^ n3702 ;
  assign n6348 = n6347 ^ n6346 ;
  assign n6349 = n6347 ^ n3701 ;
  assign n6350 = n6348 & n6349 ;
  assign n6351 = n6350 ^ n3701 ;
  assign n6352 = n6351 ^ n6298 ;
  assign n6353 = n6299 & ~n6352 ;
  assign n6354 = n6353 ^ n3700 ;
  assign n6356 = n6355 ^ n6354 ;
  assign n6357 = n6355 ^ n3699 ;
  assign n6358 = n6356 & n6357 ;
  assign n6359 = n6358 ^ n3699 ;
  assign n6297 = n6165 ^ n5723 ;
  assign n6360 = n6359 ^ n6297 ;
  assign n6361 = n6359 ^ n3698 ;
  assign n6362 = ~n6360 & ~n6361 ;
  assign n6363 = n6362 ^ n3698 ;
  assign n6364 = n6363 ^ n6295 ;
  assign n6365 = n6296 & n6364 ;
  assign n6366 = n6365 ^ n3696 ;
  assign n6368 = n6367 ^ n6366 ;
  assign n6369 = n6367 ^ n3743 ;
  assign n6370 = n6368 & n6369 ;
  assign n6371 = n6370 ^ n3743 ;
  assign n6372 = n6371 ^ n6293 ;
  assign n6373 = n6294 & ~n6372 ;
  assign n6374 = n6373 ^ n3694 ;
  assign n6375 = n6374 ^ n3693 ;
  assign n6196 = n5629 ^ x179 ;
  assign n6197 = n6196 ^ n5630 ;
  assign n5696 = n4972 ^ n4021 ;
  assign n5703 = ~n5696 & ~n5702 ;
  assign n5704 = n5703 ^ n4021 ;
  assign n6376 = n6197 ^ n5704 ;
  assign n5717 = n5716 ^ n5713 ;
  assign n6192 = n5717 & n6191 ;
  assign n6193 = n6192 ^ n5716 ;
  assign n6377 = n6376 ^ n6193 ;
  assign n6378 = n6377 ^ n6374 ;
  assign n6379 = ~n6375 & n6378 ;
  assign n6380 = n6379 ^ n3693 ;
  assign n6381 = n6380 ^ n3787 ;
  assign n6204 = n4956 ^ n4017 ;
  assign n6205 = ~n5796 & ~n6204 ;
  assign n6206 = n6205 ^ n4017 ;
  assign n6194 = n6193 ^ n5704 ;
  assign n6201 = n6194 & n6376 ;
  assign n6195 = n5637 ^ n5634 ;
  assign n6198 = n6197 ^ n6195 ;
  assign n6202 = n6201 ^ n6198 ;
  assign n6382 = n6206 ^ n6202 ;
  assign n6383 = n6382 ^ n6380 ;
  assign n6384 = ~n6381 & n6383 ;
  assign n6385 = n6384 ^ n3787 ;
  assign n6212 = n4952 ^ n4013 ;
  assign n6213 = ~n5844 & ~n6212 ;
  assign n6214 = n6213 ^ n4013 ;
  assign n6203 = n5639 ^ n5580 ;
  assign n6208 = n6203 ^ n6195 ;
  assign n6207 = n6206 ^ n6203 ;
  assign n6209 = n6208 ^ n6207 ;
  assign n6210 = ~n6202 & n6209 ;
  assign n6211 = n6210 ^ n6208 ;
  assign n6292 = n6214 ^ n6211 ;
  assign n6386 = n6385 ^ n6292 ;
  assign n6387 = n6385 ^ n3942 ;
  assign n6388 = n6386 & ~n6387 ;
  assign n6389 = n6388 ^ n3942 ;
  assign n6221 = n5067 ^ n4008 ;
  assign n6222 = n5860 & ~n6221 ;
  assign n6223 = n6222 ^ n4008 ;
  assign n6215 = n5644 ^ n5642 ;
  assign n6217 = n6215 ^ n6203 ;
  assign n6216 = n6215 ^ n6214 ;
  assign n6218 = n6217 ^ n6216 ;
  assign n6219 = n6211 & n6218 ;
  assign n6220 = n6219 ^ n6217 ;
  assign n6291 = n6223 ^ n6220 ;
  assign n6390 = n6389 ^ n6291 ;
  assign n6391 = n6389 ^ n3952 ;
  assign n6392 = n6390 & n6391 ;
  assign n6393 = n6392 ^ n3952 ;
  assign n6231 = n5101 ^ n4005 ;
  assign n6232 = n5852 & ~n6231 ;
  assign n6233 = n6232 ^ n4005 ;
  assign n6224 = n5646 ^ n5578 ;
  assign n6226 = n6224 ^ n6215 ;
  assign n6225 = n6224 ^ n6223 ;
  assign n6227 = n6226 ^ n6225 ;
  assign n6228 = ~n6220 & ~n6227 ;
  assign n6229 = n6228 ^ n6226 ;
  assign n6290 = n6233 ^ n6229 ;
  assign n6394 = n6393 ^ n6290 ;
  assign n6395 = n6393 ^ n3971 ;
  assign n6396 = ~n6394 & ~n6395 ;
  assign n6397 = n6396 ^ n3971 ;
  assign n6242 = n5130 ^ n4002 ;
  assign n6243 = n5865 & n6242 ;
  assign n6244 = n6243 ^ n4002 ;
  assign n6230 = n5649 ^ n5576 ;
  assign n6235 = n6230 ^ n6224 ;
  assign n6234 = n6233 ^ n6230 ;
  assign n6236 = n6235 ^ n6234 ;
  assign n6237 = ~n6229 & ~n6236 ;
  assign n6238 = n6237 ^ n6235 ;
  assign n6289 = n6244 ^ n6238 ;
  assign n6398 = n6397 ^ n6289 ;
  assign n6399 = n6397 ^ n4019 ;
  assign n6400 = n6398 & n6399 ;
  assign n6401 = n6400 ^ n4019 ;
  assign n6403 = n6401 ^ n4015 ;
  assign n6250 = n5164 ^ n3999 ;
  assign n6251 = ~n5784 & ~n6250 ;
  assign n6252 = n6251 ^ n3999 ;
  assign n6239 = n5652 ^ n5574 ;
  assign n6240 = n6239 ^ n6230 ;
  assign n6241 = n6240 ^ n6239 ;
  assign n6245 = n6244 ^ n6241 ;
  assign n6246 = n6238 & n6245 ;
  assign n6247 = n6246 ^ n6240 ;
  assign n6288 = n6252 ^ n6247 ;
  assign n6489 = n6403 ^ n6288 ;
  assign n6436 = n6395 ^ n6290 ;
  assign n6437 = n6387 ^ n6292 ;
  assign n6438 = n6366 ^ n3743 ;
  assign n6439 = n6438 ^ n6367 ;
  assign n6440 = n6363 ^ n6296 ;
  assign n6441 = n6332 ^ n6305 ;
  assign n6442 = n6308 ^ n3712 ;
  assign n6443 = n6442 ^ n6315 ;
  assign n6444 = n6310 ^ n3715 ;
  assign n6445 = n6313 ^ n6309 ;
  assign n6446 = n6444 & n6445 ;
  assign n6447 = ~n6443 & n6446 ;
  assign n6448 = n6319 ^ n3711 ;
  assign n6449 = n6448 ^ n6320 ;
  assign n6450 = ~n6447 & n6449 ;
  assign n6451 = n6324 ^ n6307 ;
  assign n6452 = n6450 & n6451 ;
  assign n6453 = n6327 ^ n3707 ;
  assign n6454 = n6453 ^ n6328 ;
  assign n6455 = ~n6452 & ~n6454 ;
  assign n6456 = n6441 & n6455 ;
  assign n6457 = n6335 ^ n3705 ;
  assign n6458 = n6457 ^ n6302 ;
  assign n6459 = ~n6456 & n6458 ;
  assign n6460 = n6341 ^ n6338 ;
  assign n6461 = n6459 & ~n6460 ;
  assign n6462 = n6343 ^ n3702 ;
  assign n6463 = n6462 ^ n6300 ;
  assign n6464 = ~n6461 & n6463 ;
  assign n6465 = n6349 ^ n6346 ;
  assign n6466 = n6464 & ~n6465 ;
  assign n6467 = n6351 ^ n3700 ;
  assign n6468 = n6467 ^ n6298 ;
  assign n6469 = ~n6466 & ~n6468 ;
  assign n6470 = n6357 ^ n6354 ;
  assign n6471 = n6469 & ~n6470 ;
  assign n6472 = n6361 ^ n6297 ;
  assign n6473 = n6471 & ~n6472 ;
  assign n6474 = ~n6440 & n6473 ;
  assign n6475 = ~n6439 & ~n6474 ;
  assign n6476 = n6371 ^ n3694 ;
  assign n6477 = n6476 ^ n6293 ;
  assign n6478 = n6475 & n6477 ;
  assign n6479 = n6377 ^ n6375 ;
  assign n6480 = ~n6478 & ~n6479 ;
  assign n6481 = n6382 ^ n6381 ;
  assign n6482 = ~n6480 & ~n6481 ;
  assign n6483 = n6437 & n6482 ;
  assign n6484 = n6391 ^ n6291 ;
  assign n6485 = n6483 & n6484 ;
  assign n6486 = n6436 & n6485 ;
  assign n6487 = n6399 ^ n6289 ;
  assign n6488 = n6486 & ~n6487 ;
  assign n6505 = n6489 ^ n6488 ;
  assign n6506 = n6505 ^ x200 ;
  assign n6507 = n6487 ^ n6486 ;
  assign n6508 = n6507 ^ x201 ;
  assign n6607 = n6484 ^ n6483 ;
  assign n6510 = n6482 ^ n6437 ;
  assign n6511 = n6510 ^ x204 ;
  assign n6512 = n6481 ^ n6480 ;
  assign n6513 = n6512 ^ x205 ;
  assign n6514 = n6479 ^ n6478 ;
  assign n6515 = n6514 ^ x206 ;
  assign n6516 = n6477 ^ n6475 ;
  assign n6517 = n6516 ^ x207 ;
  assign n6585 = n6473 ^ n6440 ;
  assign n6519 = n6470 ^ n6469 ;
  assign n6520 = n6519 ^ x211 ;
  assign n6521 = n6468 ^ n6466 ;
  assign n6522 = n6521 ^ x212 ;
  assign n6523 = n6465 ^ n6464 ;
  assign n6524 = n6523 ^ x213 ;
  assign n6525 = n6463 ^ n6461 ;
  assign n6526 = n6525 ^ x214 ;
  assign n6527 = n6460 ^ n6459 ;
  assign n6528 = n6527 ^ x215 ;
  assign n6529 = n6458 ^ n6456 ;
  assign n6530 = n6529 ^ x216 ;
  assign n6549 = n6451 ^ n6450 ;
  assign n6533 = n6449 ^ n6447 ;
  assign n6534 = n6533 ^ x220 ;
  assign n6535 = n6446 ^ n6443 ;
  assign n6536 = n6535 ^ x221 ;
  assign n6537 = x223 & ~n6444 ;
  assign n6538 = n6537 ^ x222 ;
  assign n6539 = n6445 ^ n6444 ;
  assign n6540 = n6539 ^ n6537 ;
  assign n6541 = n6538 & ~n6540 ;
  assign n6542 = n6541 ^ x222 ;
  assign n6543 = n6542 ^ n6535 ;
  assign n6544 = ~n6536 & n6543 ;
  assign n6545 = n6544 ^ x221 ;
  assign n6546 = n6545 ^ n6533 ;
  assign n6547 = n6534 & ~n6546 ;
  assign n6548 = n6547 ^ x220 ;
  assign n6550 = n6549 ^ n6548 ;
  assign n6551 = n6549 ^ x219 ;
  assign n6552 = n6550 & ~n6551 ;
  assign n6553 = n6552 ^ x219 ;
  assign n6532 = n6454 ^ n6452 ;
  assign n6554 = n6553 ^ n6532 ;
  assign n6555 = n6553 ^ x218 ;
  assign n6556 = ~n6554 & n6555 ;
  assign n6557 = n6556 ^ x218 ;
  assign n6531 = n6455 ^ n6441 ;
  assign n6558 = n6557 ^ n6531 ;
  assign n6559 = n6557 ^ x217 ;
  assign n6560 = ~n6558 & n6559 ;
  assign n6561 = n6560 ^ x217 ;
  assign n6562 = n6561 ^ n6529 ;
  assign n6563 = n6530 & ~n6562 ;
  assign n6564 = n6563 ^ x216 ;
  assign n6565 = n6564 ^ n6527 ;
  assign n6566 = n6528 & ~n6565 ;
  assign n6567 = n6566 ^ x215 ;
  assign n6568 = n6567 ^ n6525 ;
  assign n6569 = ~n6526 & n6568 ;
  assign n6570 = n6569 ^ x214 ;
  assign n6571 = n6570 ^ n6523 ;
  assign n6572 = ~n6524 & n6571 ;
  assign n6573 = n6572 ^ x213 ;
  assign n6574 = n6573 ^ n6521 ;
  assign n6575 = ~n6522 & n6574 ;
  assign n6576 = n6575 ^ x212 ;
  assign n6577 = n6576 ^ n6519 ;
  assign n6578 = n6520 & ~n6577 ;
  assign n6579 = n6578 ^ x211 ;
  assign n6580 = n6579 ^ x210 ;
  assign n6581 = n6472 ^ n6471 ;
  assign n6582 = n6581 ^ n6579 ;
  assign n6583 = n6580 & ~n6582 ;
  assign n6584 = n6583 ^ x210 ;
  assign n6586 = n6585 ^ n6584 ;
  assign n6587 = n6585 ^ x209 ;
  assign n6588 = ~n6586 & n6587 ;
  assign n6589 = n6588 ^ x209 ;
  assign n6518 = n6474 ^ n6439 ;
  assign n6590 = n6589 ^ n6518 ;
  assign n6591 = n6516 ^ x208 ;
  assign n6592 = n6591 ^ n6516 ;
  assign n6593 = n6592 ^ n6518 ;
  assign n6594 = ~n6590 & n6593 ;
  assign n6595 = n6594 ^ n6591 ;
  assign n6596 = n6517 & ~n6595 ;
  assign n6597 = n6596 ^ x207 ;
  assign n6598 = n6597 ^ n6514 ;
  assign n6599 = ~n6515 & n6598 ;
  assign n6600 = n6599 ^ x206 ;
  assign n6601 = n6600 ^ n6512 ;
  assign n6602 = n6513 & ~n6601 ;
  assign n6603 = n6602 ^ x205 ;
  assign n6604 = n6603 ^ n6510 ;
  assign n6605 = n6511 & ~n6604 ;
  assign n6606 = n6605 ^ x204 ;
  assign n6608 = n6607 ^ n6606 ;
  assign n6609 = n6607 ^ x203 ;
  assign n6610 = ~n6608 & n6609 ;
  assign n6611 = n6610 ^ x203 ;
  assign n6509 = n6485 ^ n6436 ;
  assign n6612 = n6611 ^ n6509 ;
  assign n6613 = n6611 ^ x202 ;
  assign n6614 = ~n6612 & n6613 ;
  assign n6615 = n6614 ^ x202 ;
  assign n6616 = n6615 ^ n6507 ;
  assign n6617 = ~n6508 & n6616 ;
  assign n6618 = n6617 ^ x201 ;
  assign n6619 = n6618 ^ n6505 ;
  assign n6620 = ~n6506 & n6619 ;
  assign n6621 = n6620 ^ x200 ;
  assign n7335 = n6621 ^ x199 ;
  assign n6402 = n6401 ^ n6288 ;
  assign n6404 = ~n6402 & n6403 ;
  assign n6405 = n6404 ^ n4015 ;
  assign n6407 = n6405 ^ n4010 ;
  assign n6258 = n5197 ^ n4218 ;
  assign n6259 = n5773 & ~n6258 ;
  assign n6260 = n6259 ^ n4218 ;
  assign n6248 = n5658 ^ x172 ;
  assign n6249 = n6248 ^ n5655 ;
  assign n6254 = n6249 ^ n6239 ;
  assign n6253 = n6252 ^ n6249 ;
  assign n6255 = n6254 ^ n6253 ;
  assign n6256 = ~n6247 & ~n6255 ;
  assign n6257 = n6256 ^ n6254 ;
  assign n6287 = n6260 ^ n6257 ;
  assign n6491 = n6407 ^ n6287 ;
  assign n6490 = ~n6488 & ~n6489 ;
  assign n6503 = n6491 ^ n6490 ;
  assign n7336 = n7335 ^ n6503 ;
  assign n6905 = n6576 ^ n6520 ;
  assign n6994 = n6905 ^ n4972 ;
  assign n6992 = n5844 ^ n4972 ;
  assign n6993 = ~n6230 & n6992 ;
  assign n6995 = n6994 ^ n6993 ;
  assign n6906 = n6573 ^ x212 ;
  assign n6907 = n6906 ^ n6521 ;
  assign n6908 = n6907 ^ n4932 ;
  assign n6909 = n6908 ^ n5796 ;
  assign n6910 = n6909 ^ n6907 ;
  assign n6911 = ~n6224 & ~n6910 ;
  assign n6912 = n6911 ^ n6908 ;
  assign n6914 = n5702 ^ n4902 ;
  assign n6915 = n6215 & ~n6914 ;
  assign n6916 = n6915 ^ n4902 ;
  assign n6913 = n6570 ^ n6524 ;
  assign n6917 = n6916 ^ n6913 ;
  assign n6920 = n5441 ^ n4851 ;
  assign n6921 = ~n5713 & ~n6920 ;
  assign n6922 = n6921 ^ n4851 ;
  assign n6918 = n6531 ^ x217 ;
  assign n6919 = n6918 ^ n6557 ;
  assign n6923 = n6922 ^ n6919 ;
  assign n6929 = n6551 ^ n6548 ;
  assign n6926 = n4821 ^ n4699 ;
  assign n6927 = n6173 & ~n6926 ;
  assign n6928 = n6927 ^ n4821 ;
  assign n6930 = n6929 ^ n6928 ;
  assign n6934 = n6545 ^ x220 ;
  assign n6935 = n6934 ^ n6533 ;
  assign n6842 = n5260 ^ n4725 ;
  assign n6843 = ~n5727 & n6842 ;
  assign n6844 = n6843 ^ n5260 ;
  assign n6841 = n6542 ^ n6536 ;
  assign n6845 = n6844 ^ n6841 ;
  assign n6823 = n6539 ^ n6538 ;
  assign n6820 = n5268 ^ n4706 ;
  assign n6821 = n5732 & ~n6820 ;
  assign n6822 = n6821 ^ n4706 ;
  assign n6824 = n6823 ^ n6822 ;
  assign n6744 = n6444 ^ x223 ;
  assign n6746 = n6744 ^ n4712 ;
  assign n6745 = n6744 ^ n5270 ;
  assign n6747 = n6746 ^ n6745 ;
  assign n6748 = ~n5738 & ~n6747 ;
  assign n6749 = n6748 ^ n6746 ;
  assign n6430 = n6062 ^ x168 ;
  assign n6431 = n6430 ^ n6054 ;
  assign n6277 = n6059 ^ x169 ;
  assign n6278 = n6277 ^ n6009 ;
  assign n6279 = n6278 ^ n4127 ;
  assign n6280 = n6279 ^ n4535 ;
  assign n6281 = n6280 ^ n6278 ;
  assign n6282 = n5082 & ~n6281 ;
  assign n6283 = n6282 ^ n6279 ;
  assign n6422 = n4532 ^ n4124 ;
  assign n6423 = ~n5114 & ~n6422 ;
  assign n6424 = n6423 ^ n4124 ;
  assign n6425 = n6424 ^ n6278 ;
  assign n6426 = n6425 ^ n6424 ;
  assign n5692 = n4550 ^ n3978 ;
  assign n5693 = ~n5691 & n5692 ;
  assign n5694 = n5693 ^ n3978 ;
  assign n5685 = n5684 ^ n5664 ;
  assign n5695 = n5694 ^ n5685 ;
  assign n6261 = n4540 ^ n3964 ;
  assign n6262 = n5765 & ~n6261 ;
  assign n6263 = n6262 ^ n3964 ;
  assign n6273 = n6263 ^ n5694 ;
  assign n6265 = n6263 ^ n6249 ;
  assign n6264 = n6263 ^ n6260 ;
  assign n6266 = n6265 ^ n6264 ;
  assign n6267 = n6257 & ~n6266 ;
  assign n6268 = n6267 ^ n6265 ;
  assign n6269 = n5661 ^ x171 ;
  assign n6270 = n6269 ^ n5569 ;
  assign n6271 = n6270 ^ n6263 ;
  assign n6272 = n6268 & n6271 ;
  assign n6274 = n6273 ^ n6272 ;
  assign n6275 = n5695 & n6274 ;
  assign n6276 = n6275 ^ n5694 ;
  assign n6427 = n6426 ^ n6276 ;
  assign n6428 = ~n6283 & n6427 ;
  assign n6429 = n6428 ^ n6425 ;
  assign n6432 = n6431 ^ n6429 ;
  assign n6406 = n6405 ^ n6287 ;
  assign n6408 = n6406 & n6407 ;
  assign n6409 = n6408 ^ n4010 ;
  assign n6286 = n6270 ^ n6268 ;
  assign n6410 = n6409 ^ n6286 ;
  assign n6411 = n6409 ^ n3610 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = n6412 ^ n3610 ;
  assign n6285 = n6274 ^ n5685 ;
  assign n6414 = n6413 ^ n6285 ;
  assign n6415 = n6413 ^ n3592 ;
  assign n6416 = n6414 & ~n6415 ;
  assign n6417 = n6416 ^ n3592 ;
  assign n6284 = n6283 ^ n6276 ;
  assign n6418 = n6417 ^ n6284 ;
  assign n6419 = n6417 ^ n3606 ;
  assign n6420 = n6418 & n6419 ;
  assign n6421 = n6420 ^ n3606 ;
  assign n6640 = n6432 ^ n6421 ;
  assign n6643 = n6421 ^ n3624 ;
  assign n6644 = n6640 & ~n6643 ;
  assign n6641 = n3636 ^ n3624 ;
  assign n6645 = n6644 ^ n6641 ;
  assign n6670 = n4078 ^ n3990 ;
  assign n6671 = n5181 & ~n6670 ;
  assign n6672 = n6671 ^ n4078 ;
  assign n6646 = n6065 ^ n6053 ;
  assign n6648 = n6646 ^ n6431 ;
  assign n6647 = n6646 ^ n6424 ;
  assign n6649 = n6648 ^ n6647 ;
  assign n6650 = ~n6429 & ~n6649 ;
  assign n6651 = n6650 ^ n6647 ;
  assign n6663 = n6068 ^ x166 ;
  assign n6664 = n6663 ^ n6050 ;
  assign n6666 = n6664 ^ n6646 ;
  assign n6652 = n4524 ^ n4121 ;
  assign n6653 = n5145 & ~n6652 ;
  assign n6654 = n6653 ^ n4121 ;
  assign n6665 = n6664 ^ n6654 ;
  assign n6667 = n6666 ^ n6665 ;
  assign n6668 = n6651 & n6667 ;
  assign n6669 = n6668 ^ n6666 ;
  assign n6673 = n6672 ^ n6669 ;
  assign n6675 = n6673 ^ n3636 ;
  assign n6655 = n6654 ^ n6651 ;
  assign n6674 = n6673 ^ n6655 ;
  assign n6676 = n6675 ^ n6674 ;
  assign n6677 = n6645 & n6676 ;
  assign n6678 = n6677 ^ n6675 ;
  assign n6656 = n6655 ^ n6645 ;
  assign n6433 = n6432 ^ n3624 ;
  assign n6434 = n6433 ^ n6421 ;
  assign n6435 = n6419 ^ n6284 ;
  assign n6492 = ~n6490 & ~n6491 ;
  assign n6493 = n6411 ^ n6286 ;
  assign n6494 = ~n6492 & n6493 ;
  assign n6495 = n6415 ^ n6285 ;
  assign n6496 = ~n6494 & ~n6495 ;
  assign n6497 = n6435 & ~n6496 ;
  assign n6657 = ~n6434 & n6497 ;
  assign n6680 = ~n6656 & ~n6657 ;
  assign n6700 = n6680 ^ n6673 ;
  assign n6703 = ~n6678 & n6700 ;
  assign n6699 = n6678 ^ n6673 ;
  assign n6701 = n6700 ^ n6699 ;
  assign n6702 = ~n3666 & n6701 ;
  assign n6704 = n6703 ^ n6702 ;
  assign n6695 = n6672 ^ n6664 ;
  assign n6696 = n6669 & n6695 ;
  assign n6692 = n4074 ^ n3986 ;
  assign n6693 = ~n5206 & ~n6692 ;
  assign n6688 = n6672 ^ n3676 ;
  assign n6686 = n6071 ^ n6049 ;
  assign n6687 = n6686 ^ n4074 ;
  assign n6689 = n6688 ^ n6687 ;
  assign n6690 = n6689 ^ n3666 ;
  assign n6685 = x193 ^ x192 ;
  assign n6691 = n6690 ^ n6685 ;
  assign n6694 = n6693 ^ n6691 ;
  assign n6697 = n6696 ^ n6694 ;
  assign n6679 = n6678 ^ n3666 ;
  assign n6681 = n6680 ^ n6679 ;
  assign n6658 = n6657 ^ n6656 ;
  assign n6499 = n6495 ^ n6494 ;
  assign n6500 = n6499 ^ x197 ;
  assign n6501 = n6493 ^ n6492 ;
  assign n6502 = n6501 ^ x198 ;
  assign n6504 = n6503 ^ x199 ;
  assign n6622 = n6621 ^ n6503 ;
  assign n6623 = n6504 & ~n6622 ;
  assign n6624 = n6623 ^ x199 ;
  assign n6625 = n6624 ^ n6501 ;
  assign n6626 = n6502 & ~n6625 ;
  assign n6627 = n6626 ^ x198 ;
  assign n6628 = n6627 ^ n6499 ;
  assign n6629 = n6500 & ~n6628 ;
  assign n6630 = n6629 ^ x197 ;
  assign n6631 = n6630 ^ x196 ;
  assign n6632 = n6496 ^ n6435 ;
  assign n6633 = n6632 ^ n6630 ;
  assign n6634 = n6631 & ~n6633 ;
  assign n6635 = n6634 ^ x196 ;
  assign n6498 = n6497 ^ n6434 ;
  assign n6636 = n6635 ^ n6498 ;
  assign n6637 = n6635 ^ x195 ;
  assign n6638 = ~n6636 & n6637 ;
  assign n6639 = n6638 ^ x195 ;
  assign n6659 = n6658 ^ n6639 ;
  assign n6660 = n6658 ^ x194 ;
  assign n6661 = ~n6659 & n6660 ;
  assign n6662 = n6661 ^ x194 ;
  assign n6682 = n6681 ^ n6662 ;
  assign n6683 = n6681 ^ x193 ;
  assign n6684 = ~n6682 & n6683 ;
  assign n6698 = n6697 ^ n6684 ;
  assign n6705 = n6704 ^ n6698 ;
  assign n5241 = n5240 ^ n4683 ;
  assign n5242 = ~n5239 & ~n5241 ;
  assign n5243 = n5242 ^ n4683 ;
  assign n6706 = n6705 ^ n5243 ;
  assign n6710 = n6662 ^ x193 ;
  assign n6711 = n6710 ^ n6681 ;
  assign n6707 = n5279 ^ n4673 ;
  assign n6708 = n5750 & ~n6707 ;
  assign n6709 = n6708 ^ n4673 ;
  assign n6712 = n6711 ^ n6709 ;
  assign n6728 = n6639 ^ x194 ;
  assign n6729 = n6728 ^ n6658 ;
  assign n6715 = n6632 ^ n6631 ;
  assign n6716 = n5313 ^ n4569 ;
  assign n6717 = ~n6130 & n6716 ;
  assign n6718 = n6717 ^ n5313 ;
  assign n6719 = n6715 & ~n6718 ;
  assign n6713 = n6498 ^ x195 ;
  assign n6714 = n6713 ^ n6635 ;
  assign n6720 = n6719 ^ n6714 ;
  assign n6721 = n6719 ^ n5323 ;
  assign n6722 = n6721 ^ n4599 ;
  assign n6723 = n6722 ^ n6719 ;
  assign n6724 = ~n6139 & ~n6723 ;
  assign n6725 = n6724 ^ n6721 ;
  assign n6726 = n6720 & n6725 ;
  assign n6727 = n6726 ^ n6719 ;
  assign n6730 = n6729 ^ n6727 ;
  assign n6731 = n6729 ^ n5288 ;
  assign n6732 = n6731 ^ n4609 ;
  assign n6733 = n6732 ^ n6729 ;
  assign n6734 = n5753 & ~n6733 ;
  assign n6735 = n6734 ^ n6731 ;
  assign n6736 = n6730 & ~n6735 ;
  assign n6737 = n6736 ^ n6729 ;
  assign n6738 = n6737 ^ n6709 ;
  assign n6739 = ~n6712 & n6738 ;
  assign n6740 = n6739 ^ n6711 ;
  assign n6741 = n6740 ^ n5243 ;
  assign n6742 = ~n6706 & n6741 ;
  assign n6743 = n6742 ^ n6705 ;
  assign n6817 = n6744 ^ n6743 ;
  assign n6818 = ~n6749 & ~n6817 ;
  assign n6819 = n6818 ^ n6744 ;
  assign n6838 = n6822 ^ n6819 ;
  assign n6839 = n6824 & n6838 ;
  assign n6840 = n6839 ^ n6823 ;
  assign n6931 = n6841 ^ n6840 ;
  assign n6932 = n6845 & n6931 ;
  assign n6933 = n6932 ^ n6844 ;
  assign n6936 = n6935 ^ n6933 ;
  assign n6937 = n6935 ^ n4745 ;
  assign n6938 = n6937 ^ n5346 ;
  assign n6939 = n6938 ^ n6935 ;
  assign n6940 = n5718 & ~n6939 ;
  assign n6941 = n6940 ^ n6937 ;
  assign n6942 = ~n6936 & n6941 ;
  assign n6943 = n6942 ^ n6935 ;
  assign n6944 = n6943 ^ n6928 ;
  assign n6945 = ~n6930 & ~n6944 ;
  assign n6946 = n6945 ^ n6929 ;
  assign n6924 = n6555 ^ n6532 ;
  assign n6947 = n6946 ^ n6924 ;
  assign n6948 = n6924 ^ n4829 ;
  assign n6949 = n6948 ^ n5250 ;
  assign n6950 = n6949 ^ n6924 ;
  assign n6951 = n6181 & ~n6950 ;
  assign n6952 = n6951 ^ n6948 ;
  assign n6953 = ~n6947 & ~n6952 ;
  assign n6925 = n6924 ^ n6922 ;
  assign n6954 = n6953 ^ n6925 ;
  assign n6955 = n6923 & n6954 ;
  assign n6956 = n6955 ^ n6922 ;
  assign n6957 = n6956 ^ n4862 ;
  assign n6958 = n6957 ^ n5463 ;
  assign n6959 = n6958 ^ n6956 ;
  assign n6960 = n6197 & n6959 ;
  assign n6961 = n6960 ^ n6957 ;
  assign n6966 = n6561 ^ x216 ;
  assign n6967 = n6966 ^ n6529 ;
  assign n6962 = n5525 ^ n4877 ;
  assign n6963 = ~n6195 & ~n6962 ;
  assign n6964 = n6963 ^ n4877 ;
  assign n6968 = n6967 ^ n6964 ;
  assign n6965 = n6964 ^ n6956 ;
  assign n6969 = n6968 ^ n6965 ;
  assign n6970 = n6961 & n6969 ;
  assign n6971 = n6970 ^ n6968 ;
  assign n6972 = n5671 ^ n4885 ;
  assign n6973 = ~n6203 & n6972 ;
  assign n6974 = n6973 ^ n4885 ;
  assign n6975 = n6974 ^ n6964 ;
  assign n6853 = n6564 ^ x215 ;
  assign n6854 = n6853 ^ n6527 ;
  assign n6976 = n6975 ^ n6854 ;
  assign n6977 = n6976 ^ n6974 ;
  assign n6978 = n6971 & n6977 ;
  assign n6979 = n6978 ^ n6975 ;
  assign n6981 = n6567 ^ n6526 ;
  assign n6982 = n6981 ^ n6916 ;
  assign n6980 = n6974 ^ n6916 ;
  assign n6983 = n6982 ^ n6980 ;
  assign n6984 = n6979 & n6983 ;
  assign n6985 = n6984 ^ n6982 ;
  assign n6986 = ~n6917 & ~n6985 ;
  assign n6987 = n6986 ^ n6916 ;
  assign n6988 = n6987 ^ n6907 ;
  assign n6989 = ~n6912 & ~n6988 ;
  assign n6990 = n6989 ^ n6907 ;
  assign n7028 = n6995 ^ n6990 ;
  assign n7029 = n7028 ^ n4021 ;
  assign n7069 = n6985 ^ n6913 ;
  assign n7064 = n6981 ^ n6979 ;
  assign n7031 = n6954 ^ n6919 ;
  assign n7032 = n7031 ^ n4040 ;
  assign n7033 = n6952 ^ n6946 ;
  assign n7034 = n7033 ^ n4043 ;
  assign n7036 = n6941 ^ n6933 ;
  assign n7037 = n7036 ^ n4049 ;
  assign n6846 = n6845 ^ n6840 ;
  assign n6847 = n6846 ^ n4052 ;
  assign n6825 = n6824 ^ n6819 ;
  assign n6752 = n6737 ^ n6712 ;
  assign n6753 = n6752 ^ n3989 ;
  assign n6761 = n6735 ^ n6727 ;
  assign n6756 = n6725 ^ n6714 ;
  assign n6754 = n6718 ^ n6715 ;
  assign n6755 = ~n4071 & ~n6754 ;
  assign n6757 = n6756 ^ n6755 ;
  assign n6758 = n6756 ^ n4068 ;
  assign n6759 = ~n6757 & n6758 ;
  assign n6760 = n6759 ^ n4068 ;
  assign n6762 = n6761 ^ n6760 ;
  assign n6763 = n6761 ^ n4064 ;
  assign n6764 = n6762 & n6763 ;
  assign n6765 = n6764 ^ n4064 ;
  assign n6766 = n6765 ^ n6752 ;
  assign n6767 = n6753 & ~n6766 ;
  assign n6768 = n6767 ^ n3989 ;
  assign n6769 = n6768 ^ n3688 ;
  assign n6770 = n6740 ^ n6706 ;
  assign n6771 = n6770 ^ n6768 ;
  assign n6772 = ~n6769 & ~n6771 ;
  assign n6773 = n6772 ^ n3688 ;
  assign n6750 = n6749 ^ n6743 ;
  assign n6812 = n6773 ^ n6750 ;
  assign n6813 = n6773 ^ n4058 ;
  assign n6814 = n6812 & ~n6813 ;
  assign n6815 = n6814 ^ n4058 ;
  assign n6834 = n6825 ^ n6815 ;
  assign n6835 = n6825 ^ n4055 ;
  assign n6836 = ~n6834 & ~n6835 ;
  assign n6837 = n6836 ^ n4055 ;
  assign n7038 = n6846 ^ n6837 ;
  assign n7039 = n6847 & ~n7038 ;
  assign n7040 = n7039 ^ n4052 ;
  assign n7041 = n7040 ^ n7036 ;
  assign n7042 = ~n7037 & n7041 ;
  assign n7043 = n7042 ^ n4049 ;
  assign n7035 = n6943 ^ n6930 ;
  assign n7044 = n7043 ^ n7035 ;
  assign n7045 = n7043 ^ n4046 ;
  assign n7046 = n7044 & ~n7045 ;
  assign n7047 = n7046 ^ n4046 ;
  assign n7048 = n7047 ^ n7033 ;
  assign n7049 = n7034 & n7048 ;
  assign n7050 = n7049 ^ n4043 ;
  assign n7051 = n7050 ^ n7031 ;
  assign n7052 = n7032 & ~n7051 ;
  assign n7053 = n7052 ^ n4040 ;
  assign n7054 = n7053 ^ n4037 ;
  assign n7055 = n6967 ^ n6961 ;
  assign n7056 = n7055 ^ n7053 ;
  assign n7057 = ~n7054 & n7056 ;
  assign n7058 = n7057 ^ n4037 ;
  assign n7059 = n7058 ^ n4034 ;
  assign n7060 = n6971 ^ n6854 ;
  assign n7061 = n7060 ^ n7058 ;
  assign n7062 = n7059 & n7061 ;
  assign n7063 = n7062 ^ n4034 ;
  assign n7065 = n7064 ^ n7063 ;
  assign n7066 = n7064 ^ n4031 ;
  assign n7067 = n7065 & ~n7066 ;
  assign n7068 = n7067 ^ n4031 ;
  assign n7070 = n7069 ^ n7068 ;
  assign n7071 = n7069 ^ n4027 ;
  assign n7072 = n7070 & n7071 ;
  assign n7073 = n7072 ^ n4027 ;
  assign n7030 = n6987 ^ n6912 ;
  assign n7074 = n7073 ^ n7030 ;
  assign n7075 = n7073 ^ n4024 ;
  assign n7076 = n7074 & ~n7075 ;
  assign n7077 = n7076 ^ n4024 ;
  assign n7078 = n7077 ^ n7028 ;
  assign n7079 = n7029 & n7078 ;
  assign n7080 = n7079 ^ n4021 ;
  assign n7151 = n7080 ^ n4017 ;
  assign n6991 = n6990 ^ n6905 ;
  assign n6996 = ~n6991 & n6995 ;
  assign n6997 = n6996 ^ n6990 ;
  assign n6901 = n5860 ^ n4956 ;
  assign n6902 = n6239 & n6901 ;
  assign n6903 = n6902 ^ n4956 ;
  assign n6900 = n6581 ^ n6580 ;
  assign n6904 = n6903 ^ n6900 ;
  assign n7081 = n6997 ^ n6904 ;
  assign n7152 = n7151 ^ n7081 ;
  assign n7124 = n7030 ^ n4024 ;
  assign n7125 = n7124 ^ n7073 ;
  assign n7126 = n7063 ^ n4031 ;
  assign n7127 = n7126 ^ n7064 ;
  assign n6848 = n6847 ^ n6837 ;
  assign n6816 = n6815 ^ n4055 ;
  assign n6826 = n6825 ^ n6816 ;
  assign n6751 = n6750 ^ n4058 ;
  assign n6774 = n6773 ^ n6751 ;
  assign n6775 = n6754 ^ n4071 ;
  assign n6776 = n6755 ^ n4068 ;
  assign n6777 = n6776 ^ n6756 ;
  assign n6778 = n6775 & n6777 ;
  assign n6779 = n6760 ^ n4064 ;
  assign n6780 = n6779 ^ n6761 ;
  assign n6781 = n6778 & n6780 ;
  assign n6782 = n6765 ^ n6753 ;
  assign n6783 = ~n6781 & n6782 ;
  assign n6784 = n6770 ^ n6769 ;
  assign n6785 = n6783 & ~n6784 ;
  assign n6827 = n6774 & ~n6785 ;
  assign n6849 = n6826 & n6827 ;
  assign n7128 = ~n6848 & ~n6849 ;
  assign n7129 = n7040 ^ n4049 ;
  assign n7130 = n7129 ^ n7036 ;
  assign n7131 = n7128 & n7130 ;
  assign n7132 = n7035 ^ n4046 ;
  assign n7133 = n7132 ^ n7043 ;
  assign n7134 = ~n7131 & n7133 ;
  assign n7135 = n7047 ^ n4043 ;
  assign n7136 = n7135 ^ n7033 ;
  assign n7137 = n7134 & ~n7136 ;
  assign n7138 = n7050 ^ n7032 ;
  assign n7139 = ~n7137 & ~n7138 ;
  assign n7140 = n7055 ^ n7054 ;
  assign n7141 = n7139 & ~n7140 ;
  assign n7142 = n7060 ^ n7059 ;
  assign n7143 = n7141 & ~n7142 ;
  assign n7144 = ~n7127 & n7143 ;
  assign n7145 = n7068 ^ n4027 ;
  assign n7146 = n7145 ^ n7069 ;
  assign n7147 = ~n7144 & ~n7146 ;
  assign n7148 = n7125 & n7147 ;
  assign n7149 = n7077 ^ n7029 ;
  assign n7150 = ~n7148 & n7149 ;
  assign n7202 = n7152 ^ n7150 ;
  assign n7203 = n7202 ^ x237 ;
  assign n7204 = n7149 ^ n7148 ;
  assign n7205 = n7204 ^ x238 ;
  assign n7206 = n7147 ^ n7125 ;
  assign n7207 = n7206 ^ x239 ;
  assign n7209 = n7143 ^ n7127 ;
  assign n7210 = n7209 ^ x241 ;
  assign n7211 = n7142 ^ n7141 ;
  assign n7212 = n7211 ^ x242 ;
  assign n7236 = n7140 ^ n7139 ;
  assign n7213 = n7136 ^ n7134 ;
  assign n7214 = n7213 ^ x245 ;
  assign n7215 = n7133 ^ n7131 ;
  assign n7216 = n7215 ^ x246 ;
  assign n7217 = n7130 ^ n7128 ;
  assign n7218 = n7217 ^ x247 ;
  assign n6828 = n6827 ^ n6826 ;
  assign n6786 = n6785 ^ n6774 ;
  assign n6787 = n6786 ^ x250 ;
  assign n6804 = n6784 ^ n6783 ;
  assign n6788 = n6782 ^ n6781 ;
  assign n6789 = n6788 ^ x252 ;
  assign n6796 = n6780 ^ n6778 ;
  assign n6790 = x255 & ~n6775 ;
  assign n6791 = n6790 ^ x254 ;
  assign n6792 = n6777 ^ n6775 ;
  assign n6793 = n6792 ^ n6790 ;
  assign n6794 = n6791 & ~n6793 ;
  assign n6795 = n6794 ^ x254 ;
  assign n6797 = n6796 ^ n6795 ;
  assign n6798 = n6796 ^ x253 ;
  assign n6799 = ~n6797 & n6798 ;
  assign n6800 = n6799 ^ x253 ;
  assign n6801 = n6800 ^ n6788 ;
  assign n6802 = n6789 & ~n6801 ;
  assign n6803 = n6802 ^ x252 ;
  assign n6805 = n6804 ^ n6803 ;
  assign n6806 = n6804 ^ x251 ;
  assign n6807 = ~n6805 & n6806 ;
  assign n6808 = n6807 ^ x251 ;
  assign n6809 = n6808 ^ n6786 ;
  assign n6810 = ~n6787 & n6809 ;
  assign n6811 = n6810 ^ x250 ;
  assign n6829 = n6828 ^ n6811 ;
  assign n6830 = n6828 ^ x249 ;
  assign n6831 = ~n6829 & n6830 ;
  assign n6832 = n6831 ^ x249 ;
  assign n6833 = n6832 ^ x248 ;
  assign n6850 = n6849 ^ n6848 ;
  assign n7219 = n6850 ^ n6832 ;
  assign n7220 = n6833 & n7219 ;
  assign n7221 = n7220 ^ x248 ;
  assign n7222 = n7221 ^ n7217 ;
  assign n7223 = ~n7218 & n7222 ;
  assign n7224 = n7223 ^ x247 ;
  assign n7225 = n7224 ^ n7215 ;
  assign n7226 = ~n7216 & n7225 ;
  assign n7227 = n7226 ^ x246 ;
  assign n7228 = n7227 ^ n7213 ;
  assign n7229 = ~n7214 & n7228 ;
  assign n7230 = n7229 ^ x245 ;
  assign n7231 = n7230 ^ x244 ;
  assign n7232 = n7138 ^ n7137 ;
  assign n7233 = n7232 ^ n7230 ;
  assign n7234 = n7231 & n7233 ;
  assign n7235 = n7234 ^ x244 ;
  assign n7237 = n7236 ^ n7235 ;
  assign n7238 = n7236 ^ x243 ;
  assign n7239 = ~n7237 & n7238 ;
  assign n7240 = n7239 ^ x243 ;
  assign n7241 = n7240 ^ n7211 ;
  assign n7242 = n7212 & ~n7241 ;
  assign n7243 = n7242 ^ x242 ;
  assign n7244 = n7243 ^ n7209 ;
  assign n7245 = n7210 & ~n7244 ;
  assign n7246 = n7245 ^ x241 ;
  assign n7208 = n7146 ^ n7144 ;
  assign n7247 = n7246 ^ n7208 ;
  assign n7248 = n7206 ^ x240 ;
  assign n7249 = n7248 ^ n7208 ;
  assign n7250 = n7249 ^ n7206 ;
  assign n7251 = ~n7247 & n7250 ;
  assign n7252 = n7251 ^ n7248 ;
  assign n7253 = n7207 & ~n7252 ;
  assign n7254 = n7253 ^ x239 ;
  assign n7255 = n7254 ^ n7204 ;
  assign n7256 = n7205 & ~n7255 ;
  assign n7257 = n7256 ^ x238 ;
  assign n7258 = n7257 ^ n7202 ;
  assign n7259 = ~n7203 & n7258 ;
  assign n7260 = n7259 ^ x237 ;
  assign n7337 = n7260 ^ x236 ;
  assign n7082 = n7081 ^ n7080 ;
  assign n7083 = n7081 ^ n4017 ;
  assign n7084 = n7082 & n7083 ;
  assign n7085 = n7084 ^ n4017 ;
  assign n6998 = n6997 ^ n6900 ;
  assign n6999 = n6904 & n6998 ;
  assign n7000 = n6999 ^ n6903 ;
  assign n6898 = n6587 ^ n6584 ;
  assign n6895 = n5852 ^ n4952 ;
  assign n6896 = n6249 & n6895 ;
  assign n6897 = n6896 ^ n4952 ;
  assign n6899 = n6898 ^ n6897 ;
  assign n7026 = n7000 ^ n6899 ;
  assign n7027 = n7026 ^ n4013 ;
  assign n7154 = n7085 ^ n7027 ;
  assign n7153 = ~n7150 & n7152 ;
  assign n7200 = n7154 ^ n7153 ;
  assign n7338 = n7337 ^ n7200 ;
  assign n7339 = n7338 ^ n5691 ;
  assign n7340 = n7339 ^ n6686 ;
  assign n7341 = n7340 ^ n7338 ;
  assign n7342 = n7336 & ~n7341 ;
  assign n7343 = n7342 ^ n7339 ;
  assign n7420 = n6624 ^ x198 ;
  assign n7421 = n7420 ^ n6501 ;
  assign n7723 = n6106 ^ n5082 ;
  assign n7724 = n7421 & ~n7723 ;
  assign n7725 = n7724 ^ n5082 ;
  assign n7305 = n6618 ^ x200 ;
  assign n7306 = n7305 ^ n6505 ;
  assign n7182 = n6615 ^ n6508 ;
  assign n7346 = n6646 ^ n5773 ;
  assign n7347 = ~n7182 & ~n7346 ;
  assign n7348 = n7347 ^ n5773 ;
  assign n7344 = n7254 ^ x238 ;
  assign n7345 = n7344 ^ n7204 ;
  assign n7349 = n7348 ^ n7345 ;
  assign n6861 = n6609 ^ n6606 ;
  assign n7350 = n7246 ^ x240 ;
  assign n7351 = n7350 ^ n7208 ;
  assign n7353 = n7351 ^ n5865 ;
  assign n7352 = n7351 ^ n6278 ;
  assign n7354 = n7353 ^ n7352 ;
  assign n7355 = n6861 & n7354 ;
  assign n7356 = n7355 ^ n7353 ;
  assign n7363 = n7243 ^ n7210 ;
  assign n6867 = n6603 ^ x204 ;
  assign n6868 = n6867 ^ n6510 ;
  assign n7360 = n5852 ^ n5685 ;
  assign n7361 = ~n6868 & n7360 ;
  assign n7362 = n7361 ^ n5685 ;
  assign n7364 = n7363 ^ n7362 ;
  assign n7568 = n7240 ^ x242 ;
  assign n7569 = n7568 ^ n7211 ;
  assign n7559 = n7238 ^ n7235 ;
  assign n7368 = n7232 ^ n7231 ;
  assign n6887 = n6595 ^ x207 ;
  assign n7365 = n6239 ^ n5796 ;
  assign n7366 = n6887 & ~n7365 ;
  assign n7367 = n7366 ^ n5796 ;
  assign n7369 = n7368 ^ n7367 ;
  assign n7547 = n7227 ^ n7214 ;
  assign n7327 = n6808 ^ x250 ;
  assign n7328 = n7327 ^ n6786 ;
  assign n7371 = n7328 ^ n6197 ;
  assign n7372 = n7371 ^ n5250 ;
  assign n7373 = n7372 ^ n7328 ;
  assign n7374 = n6913 & n7373 ;
  assign n7375 = n7374 ^ n7371 ;
  assign n7376 = n6800 ^ x252 ;
  assign n7377 = n7376 ^ n6788 ;
  assign n7378 = n7377 ^ n5346 ;
  assign n7379 = n7378 ^ n6181 ;
  assign n7380 = n7379 ^ n7377 ;
  assign n7381 = n6854 & ~n7380 ;
  assign n7382 = n7381 ^ n7378 ;
  assign n7387 = n6173 ^ n5260 ;
  assign n7388 = n6967 & ~n7387 ;
  assign n7389 = n7388 ^ n5260 ;
  assign n7386 = n6798 ^ n6795 ;
  assign n7390 = n7389 ^ n7386 ;
  assign n7334 = n6792 ^ n6791 ;
  assign n7391 = n7334 ^ n5268 ;
  assign n7392 = n7391 ^ n5718 ;
  assign n7393 = n7392 ^ n7334 ;
  assign n7394 = n6919 & ~n7393 ;
  assign n7395 = n7394 ^ n7391 ;
  assign n7401 = n6775 ^ x255 ;
  assign n7398 = n5727 ^ n5270 ;
  assign n7399 = n6924 & ~n7398 ;
  assign n7400 = n7399 ^ n5270 ;
  assign n7402 = n7401 ^ n7400 ;
  assign n7465 = n5732 ^ n5240 ;
  assign n7466 = ~n6929 & n7465 ;
  assign n7467 = n7466 ^ n5240 ;
  assign n7458 = n5308 ^ n3986 ;
  assign n7459 = n6092 & ~n7458 ;
  assign n7453 = n6627 ^ n6500 ;
  assign n7454 = n7453 ^ n6692 ;
  assign n7427 = n5300 ^ n3990 ;
  assign n7428 = n6098 & n7427 ;
  assign n7429 = n7428 ^ n3990 ;
  assign n7455 = n7454 ^ n7429 ;
  assign n7456 = n7455 ^ n4078 ;
  assign n7452 = x225 ^ x224 ;
  assign n7457 = n7456 ^ n7452 ;
  assign n7460 = n7459 ^ n7457 ;
  assign n6862 = n6861 ^ n4540 ;
  assign n6863 = n6862 ^ n5082 ;
  assign n6864 = n6863 ^ n6861 ;
  assign n6865 = n6664 & ~n6864 ;
  assign n6866 = n6865 ^ n6862 ;
  assign n7113 = n5114 ^ n4550 ;
  assign n7114 = n6686 & ~n7113 ;
  assign n7115 = n7114 ^ n4550 ;
  assign n7117 = n7115 ^ n6861 ;
  assign n6869 = n5691 ^ n5197 ;
  assign n6870 = ~n6646 & ~n6869 ;
  assign n6871 = n6870 ^ n5197 ;
  assign n6872 = n6871 ^ n6868 ;
  assign n6874 = n5765 ^ n5164 ;
  assign n6875 = n6431 & n6874 ;
  assign n6876 = n6875 ^ n5164 ;
  assign n6873 = n6600 ^ n6513 ;
  assign n6877 = n6876 ^ n6873 ;
  assign n6880 = n5773 ^ n5130 ;
  assign n6881 = n6278 & ~n6880 ;
  assign n6882 = n6881 ^ n5130 ;
  assign n6878 = n6597 ^ x206 ;
  assign n6879 = n6878 ^ n6514 ;
  assign n6883 = n6882 ^ n6879 ;
  assign n6884 = n5784 ^ n5101 ;
  assign n6885 = n5685 & n6884 ;
  assign n6886 = n6885 ^ n5101 ;
  assign n6888 = n6887 ^ n6886 ;
  assign n6891 = n5865 ^ n5067 ;
  assign n6892 = n6270 & n6891 ;
  assign n6893 = n6892 ^ n5067 ;
  assign n6889 = n6589 ^ x208 ;
  assign n6890 = n6889 ^ n6518 ;
  assign n6894 = n6893 ^ n6890 ;
  assign n7001 = n7000 ^ n6897 ;
  assign n7002 = n6899 & ~n7001 ;
  assign n7003 = n7002 ^ n6898 ;
  assign n7004 = n7003 ^ n6890 ;
  assign n7005 = n6894 & ~n7004 ;
  assign n7006 = n7005 ^ n6893 ;
  assign n7007 = n7006 ^ n6886 ;
  assign n7008 = ~n6888 & n7007 ;
  assign n7009 = n7008 ^ n6887 ;
  assign n7010 = n7009 ^ n6879 ;
  assign n7011 = n6883 & n7010 ;
  assign n7012 = n7011 ^ n6882 ;
  assign n7013 = n7012 ^ n6873 ;
  assign n7014 = n6877 & n7013 ;
  assign n7015 = n7014 ^ n6876 ;
  assign n7016 = n7015 ^ n6868 ;
  assign n7017 = n6872 & ~n7016 ;
  assign n7018 = n7017 ^ n6871 ;
  assign n7116 = n7115 ^ n7018 ;
  assign n7118 = n7117 ^ n7116 ;
  assign n7119 = ~n6866 & n7118 ;
  assign n7120 = n7119 ^ n7117 ;
  assign n7174 = n5145 ^ n4535 ;
  assign n7175 = ~n6106 & n7174 ;
  assign n7176 = n7175 ^ n4535 ;
  assign n7178 = n7176 ^ n7115 ;
  assign n7121 = n6613 ^ n6509 ;
  assign n7177 = n7176 ^ n7121 ;
  assign n7179 = n7178 ^ n7177 ;
  assign n7180 = n7120 & n7179 ;
  assign n7181 = n7180 ^ n7178 ;
  assign n7297 = n5181 ^ n4532 ;
  assign n7298 = n6101 & n7297 ;
  assign n7299 = n7298 ^ n4532 ;
  assign n7301 = n7299 ^ n7176 ;
  assign n7300 = n7299 ^ n7182 ;
  assign n7302 = n7301 ^ n7300 ;
  assign n7303 = n7181 & ~n7302 ;
  assign n7304 = n7303 ^ n7301 ;
  assign n7404 = n7336 ^ n7299 ;
  assign n7403 = n7336 ^ n7306 ;
  assign n7405 = n7404 ^ n7403 ;
  assign n7406 = n7304 & ~n7405 ;
  assign n7407 = n7406 ^ n7404 ;
  assign n7423 = n7421 ^ n7336 ;
  assign n7408 = n5206 ^ n4524 ;
  assign n7409 = n6100 & ~n7408 ;
  assign n7410 = n7409 ^ n4524 ;
  assign n7422 = n7421 ^ n7410 ;
  assign n7424 = n7423 ^ n7422 ;
  assign n7425 = ~n7407 & n7424 ;
  assign n7426 = n7425 ^ n7422 ;
  assign n7450 = n7429 ^ n7421 ;
  assign n7451 = ~n7426 & ~n7450 ;
  assign n7461 = n7460 ^ n7451 ;
  assign n7019 = n7018 ^ n6866 ;
  assign n7020 = n7019 ^ n3964 ;
  assign n7022 = n7012 ^ n6877 ;
  assign n7023 = n7022 ^ n3999 ;
  assign n7024 = n7006 ^ n6888 ;
  assign n7025 = n7024 ^ n4005 ;
  assign n7086 = n7085 ^ n7026 ;
  assign n7087 = ~n7027 & n7086 ;
  assign n7088 = n7087 ^ n4013 ;
  assign n7089 = n7088 ^ n4008 ;
  assign n7090 = n7003 ^ n6894 ;
  assign n7091 = n7090 ^ n7088 ;
  assign n7092 = n7089 & n7091 ;
  assign n7093 = n7092 ^ n4008 ;
  assign n7094 = n7093 ^ n7024 ;
  assign n7095 = ~n7025 & ~n7094 ;
  assign n7096 = n7095 ^ n4005 ;
  assign n7097 = n7096 ^ n4002 ;
  assign n7098 = n7009 ^ n6883 ;
  assign n7099 = n7098 ^ n7096 ;
  assign n7100 = ~n7097 & ~n7099 ;
  assign n7101 = n7100 ^ n4002 ;
  assign n7102 = n7101 ^ n7022 ;
  assign n7103 = n7023 & ~n7102 ;
  assign n7104 = n7103 ^ n3999 ;
  assign n7021 = n7015 ^ n6872 ;
  assign n7105 = n7104 ^ n7021 ;
  assign n7106 = n7104 ^ n4218 ;
  assign n7107 = n7105 & n7106 ;
  assign n7108 = n7107 ^ n4218 ;
  assign n7109 = n7108 ^ n7019 ;
  assign n7110 = ~n7020 & ~n7109 ;
  assign n7111 = n7110 ^ n3964 ;
  assign n7112 = n7111 ^ n3978 ;
  assign n7122 = n7121 ^ n7120 ;
  assign n7170 = n7122 ^ n7111 ;
  assign n7171 = n7112 & ~n7170 ;
  assign n7172 = n7171 ^ n3978 ;
  assign n7173 = n7172 ^ n4127 ;
  assign n7183 = n7182 ^ n7181 ;
  assign n7293 = n7183 ^ n7172 ;
  assign n7294 = ~n7173 & n7293 ;
  assign n7295 = n7294 ^ n4127 ;
  assign n7296 = n7295 ^ n4124 ;
  assign n7307 = n7306 ^ n7304 ;
  assign n7412 = n7307 ^ n7295 ;
  assign n7413 = n7296 & ~n7412 ;
  assign n7414 = n7413 ^ n4124 ;
  assign n7416 = n7414 ^ n4121 ;
  assign n7411 = n7410 ^ n7407 ;
  assign n7433 = n7416 ^ n7411 ;
  assign n7308 = n7307 ^ n7296 ;
  assign n7123 = n7122 ^ n7112 ;
  assign n7155 = n7153 & n7154 ;
  assign n7156 = n7090 ^ n7089 ;
  assign n7157 = n7155 & n7156 ;
  assign n7158 = n7093 ^ n7025 ;
  assign n7159 = n7157 & n7158 ;
  assign n7160 = n7098 ^ n7097 ;
  assign n7161 = n7159 & ~n7160 ;
  assign n7162 = n7101 ^ n7023 ;
  assign n7163 = ~n7161 & n7162 ;
  assign n7164 = n7021 ^ n4218 ;
  assign n7165 = n7164 ^ n7104 ;
  assign n7166 = ~n7163 & n7165 ;
  assign n7167 = n7108 ^ n7020 ;
  assign n7168 = ~n7166 & ~n7167 ;
  assign n7169 = n7123 & ~n7168 ;
  assign n7184 = n7183 ^ n7173 ;
  assign n7309 = ~n7169 & ~n7184 ;
  assign n7434 = n7308 & n7309 ;
  assign n7443 = n7433 & ~n7434 ;
  assign n7430 = n7429 ^ n7426 ;
  assign n7415 = n7414 ^ n7411 ;
  assign n7417 = n7415 & n7416 ;
  assign n7418 = n7417 ^ n4121 ;
  assign n7419 = n7418 ^ n4078 ;
  assign n7444 = n7430 ^ n7419 ;
  assign n7449 = ~n7443 & ~n7444 ;
  assign n7462 = n7461 ^ n7449 ;
  assign n7445 = n7444 ^ n7443 ;
  assign n7310 = n7309 ^ n7308 ;
  assign n7311 = n7310 ^ x227 ;
  assign n7186 = n7168 ^ n7123 ;
  assign n7187 = n7186 ^ x229 ;
  assign n7188 = n7167 ^ n7166 ;
  assign n7189 = n7188 ^ x230 ;
  assign n7190 = n7165 ^ n7163 ;
  assign n7191 = n7190 ^ x231 ;
  assign n7192 = n7162 ^ n7161 ;
  assign n7193 = n7192 ^ x232 ;
  assign n7194 = n7160 ^ n7159 ;
  assign n7195 = n7194 ^ x233 ;
  assign n7196 = n7158 ^ n7157 ;
  assign n7197 = n7196 ^ x234 ;
  assign n7198 = n7156 ^ n7155 ;
  assign n7199 = n7198 ^ x235 ;
  assign n7201 = n7200 ^ x236 ;
  assign n7261 = n7260 ^ n7200 ;
  assign n7262 = n7201 & ~n7261 ;
  assign n7263 = n7262 ^ x236 ;
  assign n7264 = n7263 ^ n7198 ;
  assign n7265 = n7199 & ~n7264 ;
  assign n7266 = n7265 ^ x235 ;
  assign n7267 = n7266 ^ n7196 ;
  assign n7268 = n7197 & ~n7267 ;
  assign n7269 = n7268 ^ x234 ;
  assign n7270 = n7269 ^ n7194 ;
  assign n7271 = ~n7195 & n7270 ;
  assign n7272 = n7271 ^ x233 ;
  assign n7273 = n7272 ^ n7192 ;
  assign n7274 = n7193 & ~n7273 ;
  assign n7275 = n7274 ^ x232 ;
  assign n7276 = n7275 ^ n7190 ;
  assign n7277 = ~n7191 & n7276 ;
  assign n7278 = n7277 ^ x231 ;
  assign n7279 = n7278 ^ n7188 ;
  assign n7280 = ~n7189 & n7279 ;
  assign n7281 = n7280 ^ x230 ;
  assign n7282 = n7281 ^ n7186 ;
  assign n7283 = ~n7187 & n7282 ;
  assign n7284 = n7283 ^ x229 ;
  assign n7285 = n7284 ^ x228 ;
  assign n7185 = n7184 ^ n7169 ;
  assign n7312 = n7284 ^ n7185 ;
  assign n7313 = n7285 & n7312 ;
  assign n7314 = n7313 ^ x228 ;
  assign n7436 = n7314 ^ n7310 ;
  assign n7437 = ~n7311 & n7436 ;
  assign n7438 = n7437 ^ x227 ;
  assign n7435 = n7434 ^ n7433 ;
  assign n7439 = n7438 ^ n7435 ;
  assign n7440 = n7438 ^ x226 ;
  assign n7441 = n7439 & n7440 ;
  assign n7442 = n7441 ^ x226 ;
  assign n7446 = n7445 ^ n7442 ;
  assign n7447 = n7445 ^ x225 ;
  assign n7448 = n7446 & ~n7447 ;
  assign n7463 = n7462 ^ n7448 ;
  assign n7431 = n7430 ^ n7418 ;
  assign n7432 = ~n7419 & ~n7431 ;
  assign n7464 = n7463 ^ n7432 ;
  assign n7468 = n7467 ^ n7464 ;
  assign n7472 = n7442 ^ x225 ;
  assign n7473 = n7472 ^ n7445 ;
  assign n7469 = n5738 ^ n5279 ;
  assign n7470 = n6935 & ~n7469 ;
  assign n7471 = n7470 ^ n5279 ;
  assign n7474 = n7473 ^ n7471 ;
  assign n7475 = n7440 ^ n7435 ;
  assign n7486 = n7475 ^ n7471 ;
  assign n7476 = n7475 ^ n5288 ;
  assign n7477 = n7476 ^ n5239 ;
  assign n7478 = n7477 ^ n7475 ;
  assign n7479 = ~n6841 & n7478 ;
  assign n7480 = n7479 ^ n7476 ;
  assign n6858 = n5753 ^ n5313 ;
  assign n6859 = ~n6744 & n6858 ;
  assign n6860 = n6859 ^ n5313 ;
  assign n7286 = n7285 ^ n7185 ;
  assign n7287 = ~n6860 & ~n7286 ;
  assign n7288 = n7287 ^ n5323 ;
  assign n7289 = n7288 ^ n5750 ;
  assign n7290 = n7289 ^ n7287 ;
  assign n7291 = n6823 & n7290 ;
  assign n7292 = n7291 ^ n7288 ;
  assign n7315 = n7314 ^ n7311 ;
  assign n7481 = n7315 ^ n7287 ;
  assign n7482 = ~n7292 & ~n7481 ;
  assign n7483 = n7482 ^ n7315 ;
  assign n7484 = n7483 ^ n7475 ;
  assign n7485 = n7480 & n7484 ;
  assign n7487 = n7486 ^ n7485 ;
  assign n7488 = ~n7474 & n7487 ;
  assign n7489 = n7488 ^ n7473 ;
  assign n7490 = n7489 ^ n7464 ;
  assign n7491 = ~n7468 & ~n7490 ;
  assign n7492 = n7491 ^ n7467 ;
  assign n7493 = n7492 ^ n7400 ;
  assign n7494 = n7402 & n7493 ;
  assign n7495 = n7494 ^ n7401 ;
  assign n7396 = n7389 ^ n7334 ;
  assign n7397 = n7396 ^ n7389 ;
  assign n7496 = n7495 ^ n7397 ;
  assign n7497 = ~n7395 & ~n7496 ;
  assign n7498 = n7497 ^ n7396 ;
  assign n7499 = ~n7390 & ~n7498 ;
  assign n7500 = n7499 ^ n7389 ;
  assign n7383 = n5713 ^ n4699 ;
  assign n7384 = n6981 & n7383 ;
  assign n7385 = n7384 ^ n5713 ;
  assign n7501 = n7500 ^ n7385 ;
  assign n7502 = n7501 ^ n7377 ;
  assign n7503 = n7502 ^ n7385 ;
  assign n7504 = n7382 & ~n7503 ;
  assign n7505 = n7504 ^ n7501 ;
  assign n7506 = n6806 ^ n6803 ;
  assign n7507 = n7506 ^ n7385 ;
  assign n7508 = ~n7505 & ~n7507 ;
  assign n7509 = n7508 ^ n7506 ;
  assign n7510 = n7509 ^ n7328 ;
  assign n7511 = ~n7375 & ~n7510 ;
  assign n7512 = n7511 ^ n7328 ;
  assign n6852 = n6830 ^ n6811 ;
  assign n7513 = n7512 ^ n6852 ;
  assign n7514 = n7512 ^ n5441 ;
  assign n7515 = n7514 ^ n6195 ;
  assign n7516 = n7515 ^ n7512 ;
  assign n7517 = ~n6907 & n7516 ;
  assign n7518 = n7517 ^ n7514 ;
  assign n7519 = ~n7513 & ~n7518 ;
  assign n7520 = n7519 ^ n6852 ;
  assign n6851 = n6850 ^ n6833 ;
  assign n7521 = n7520 ^ n6851 ;
  assign n7522 = n6851 ^ n5463 ;
  assign n7523 = n7522 ^ n6203 ;
  assign n7524 = n7523 ^ n6851 ;
  assign n7525 = n6905 & n7524 ;
  assign n7526 = n7525 ^ n7522 ;
  assign n7527 = ~n7521 & ~n7526 ;
  assign n7528 = n7527 ^ n7520 ;
  assign n7529 = n7528 ^ n6215 ;
  assign n7530 = n7529 ^ n5525 ;
  assign n7531 = n7530 ^ n7528 ;
  assign n7532 = ~n6900 & ~n7531 ;
  assign n7533 = n7532 ^ n7529 ;
  assign n7534 = n7221 ^ x247 ;
  assign n7535 = n7534 ^ n7217 ;
  assign n7536 = n7535 ^ n7528 ;
  assign n7537 = ~n7533 & ~n7536 ;
  assign n7538 = n7537 ^ n7535 ;
  assign n7370 = n7224 ^ n7216 ;
  assign n7539 = n7538 ^ n7370 ;
  assign n7540 = n7370 ^ n5671 ;
  assign n7541 = n7540 ^ n6224 ;
  assign n7542 = n7541 ^ n7370 ;
  assign n7543 = n6898 & n7542 ;
  assign n7544 = n7543 ^ n7540 ;
  assign n7545 = n7539 & ~n7544 ;
  assign n7546 = n7545 ^ n7538 ;
  assign n7548 = n7547 ^ n7546 ;
  assign n7549 = n7546 ^ n6230 ;
  assign n7550 = n7549 ^ n5702 ;
  assign n7551 = n7550 ^ n7546 ;
  assign n7552 = ~n6890 & n7551 ;
  assign n7553 = n7552 ^ n7549 ;
  assign n7554 = n7548 & ~n7553 ;
  assign n7555 = n7554 ^ n7547 ;
  assign n7556 = n7555 ^ n7367 ;
  assign n7557 = n7369 & ~n7556 ;
  assign n7558 = n7557 ^ n7368 ;
  assign n7560 = n7559 ^ n7558 ;
  assign n7561 = n7558 ^ n6249 ;
  assign n7562 = n7561 ^ n5844 ;
  assign n7563 = n7562 ^ n7558 ;
  assign n7564 = n6879 & ~n7563 ;
  assign n7565 = n7564 ^ n7561 ;
  assign n7566 = ~n7560 & n7565 ;
  assign n7567 = n7566 ^ n7559 ;
  assign n7570 = n7569 ^ n7567 ;
  assign n7571 = n7569 ^ n5860 ;
  assign n7572 = n7571 ^ n6270 ;
  assign n7573 = n7572 ^ n7569 ;
  assign n7574 = n6873 & n7573 ;
  assign n7575 = n7574 ^ n7571 ;
  assign n7576 = n7570 & n7575 ;
  assign n7577 = n7576 ^ n7569 ;
  assign n7578 = n7577 ^ n7362 ;
  assign n7579 = n7364 & ~n7578 ;
  assign n7580 = n7579 ^ n7363 ;
  assign n7357 = n7252 ^ x239 ;
  assign n7358 = n7357 ^ n7351 ;
  assign n7359 = n7358 ^ n7357 ;
  assign n7581 = n7580 ^ n7359 ;
  assign n7582 = n7356 & n7581 ;
  assign n7583 = n7582 ^ n7358 ;
  assign n7588 = n7357 ^ n7345 ;
  assign n7584 = n6431 ^ n5784 ;
  assign n7585 = ~n7121 & ~n7584 ;
  assign n7586 = n7585 ^ n6431 ;
  assign n7587 = n7586 ^ n7345 ;
  assign n7589 = n7588 ^ n7587 ;
  assign n7590 = n7583 & n7589 ;
  assign n7591 = n7590 ^ n7588 ;
  assign n7592 = n7349 & ~n7591 ;
  assign n7593 = n7592 ^ n7348 ;
  assign n7594 = n7593 ^ n5765 ;
  assign n7595 = n7594 ^ n6664 ;
  assign n7596 = n7595 ^ n7593 ;
  assign n7597 = ~n7306 & n7596 ;
  assign n7598 = n7597 ^ n7594 ;
  assign n7599 = n7257 ^ n7203 ;
  assign n7600 = n7599 ^ n7593 ;
  assign n7601 = ~n7598 & ~n7600 ;
  assign n7602 = n7601 ^ n7599 ;
  assign n7727 = n7725 ^ n7602 ;
  assign n7726 = n7725 ^ n7338 ;
  assign n7728 = n7727 ^ n7726 ;
  assign n7729 = ~n7343 & ~n7728 ;
  assign n7730 = n7729 ^ n7726 ;
  assign n7737 = n6101 ^ n5114 ;
  assign n7738 = n7453 & ~n7737 ;
  assign n7739 = n7738 ^ n5114 ;
  assign n7741 = n7739 ^ n7725 ;
  assign n7731 = n7263 ^ n7199 ;
  assign n7740 = n7739 ^ n7731 ;
  assign n7742 = n7741 ^ n7740 ;
  assign n7743 = n7730 & n7742 ;
  assign n7744 = n7743 ^ n7741 ;
  assign n7939 = n6100 ^ n5145 ;
  assign n7940 = n6715 & n7939 ;
  assign n7941 = n7940 ^ n5145 ;
  assign n7943 = n7941 ^ n7739 ;
  assign n7745 = n7266 ^ x234 ;
  assign n7746 = n7745 ^ n7196 ;
  assign n7942 = n7941 ^ n7746 ;
  assign n7944 = n7943 ^ n7942 ;
  assign n7945 = ~n7744 & ~n7944 ;
  assign n7946 = n7945 ^ n7943 ;
  assign n7979 = n6098 ^ n5181 ;
  assign n7980 = n6714 & n7979 ;
  assign n7981 = n7980 ^ n5181 ;
  assign n7947 = n7269 ^ n7195 ;
  assign n7983 = n7981 ^ n7947 ;
  assign n7982 = n7981 ^ n7941 ;
  assign n7984 = n7983 ^ n7982 ;
  assign n7985 = ~n7946 & ~n7984 ;
  assign n7986 = n7985 ^ n7982 ;
  assign n8011 = n7275 ^ n7191 ;
  assign n8013 = n8011 ^ n7981 ;
  assign n7987 = n7272 ^ x232 ;
  assign n7988 = n7987 ^ n7192 ;
  assign n8012 = n8011 ^ n7988 ;
  assign n8014 = n8013 ^ n8012 ;
  assign n8015 = n7986 & n8014 ;
  assign n8016 = n8015 ^ n8013 ;
  assign n8008 = n6092 ^ n5206 ;
  assign n8009 = ~n6729 & ~n8008 ;
  assign n8010 = n8009 ^ n6092 ;
  assign n8017 = n8016 ^ n8010 ;
  assign n7603 = n7602 ^ n7343 ;
  assign n7604 = n7603 ^ n5197 ;
  assign n7605 = n7591 ^ n7348 ;
  assign n7606 = n7605 ^ n5130 ;
  assign n7701 = n7580 ^ n7356 ;
  assign n7608 = n7565 ^ n7559 ;
  assign n7609 = n7608 ^ n4972 ;
  assign n7679 = n7553 ^ n7547 ;
  assign n7611 = n7535 ^ n7533 ;
  assign n7612 = n7611 ^ n4877 ;
  assign n7613 = n7526 ^ n7520 ;
  assign n7614 = n7613 ^ n4862 ;
  assign n7615 = n7518 ^ n6852 ;
  assign n7616 = n7615 ^ n4851 ;
  assign n7617 = n7509 ^ n7375 ;
  assign n7618 = n7617 ^ n4829 ;
  assign n7619 = n7506 ^ n7505 ;
  assign n7620 = n7619 ^ n4821 ;
  assign n7654 = n7500 ^ n7382 ;
  assign n7649 = n7498 ^ n7386 ;
  assign n7621 = n7495 ^ n7395 ;
  assign n7622 = n7621 ^ n4706 ;
  assign n7623 = n7492 ^ n7402 ;
  assign n7624 = n7623 ^ n4712 ;
  assign n7625 = n7489 ^ n7468 ;
  assign n7626 = n7625 ^ n4683 ;
  assign n7627 = n7487 ^ n7473 ;
  assign n7628 = n7627 ^ n4673 ;
  assign n7317 = n7286 ^ n6860 ;
  assign n7318 = ~n4569 & n7317 ;
  assign n7319 = n7318 ^ n4599 ;
  assign n7316 = n7315 ^ n7292 ;
  assign n7630 = n7318 ^ n7316 ;
  assign n7631 = ~n7319 & n7630 ;
  assign n7632 = n7631 ^ n4599 ;
  assign n7629 = n7483 ^ n7480 ;
  assign n7633 = n7632 ^ n7629 ;
  assign n7634 = n7632 ^ n4609 ;
  assign n7635 = ~n7633 & ~n7634 ;
  assign n7636 = n7635 ^ n4609 ;
  assign n7637 = n7636 ^ n7627 ;
  assign n7638 = ~n7628 & ~n7637 ;
  assign n7639 = n7638 ^ n4673 ;
  assign n7640 = n7639 ^ n7625 ;
  assign n7641 = ~n7626 & n7640 ;
  assign n7642 = n7641 ^ n4683 ;
  assign n7643 = n7642 ^ n7623 ;
  assign n7644 = n7624 & n7643 ;
  assign n7645 = n7644 ^ n4712 ;
  assign n7646 = n7645 ^ n7621 ;
  assign n7647 = n7622 & ~n7646 ;
  assign n7648 = n7647 ^ n4706 ;
  assign n7650 = n7649 ^ n7648 ;
  assign n7651 = n7648 ^ n4725 ;
  assign n7652 = ~n7650 & n7651 ;
  assign n7653 = n7652 ^ n7649 ;
  assign n7655 = n7654 ^ n7653 ;
  assign n7656 = n7654 ^ n4745 ;
  assign n7657 = n7655 & n7656 ;
  assign n7658 = n7657 ^ n4745 ;
  assign n7659 = n7658 ^ n7619 ;
  assign n7660 = ~n7620 & n7659 ;
  assign n7661 = n7660 ^ n7658 ;
  assign n7662 = n7661 ^ n7617 ;
  assign n7663 = n7618 & n7662 ;
  assign n7664 = n7663 ^ n4829 ;
  assign n7665 = n7664 ^ n7615 ;
  assign n7666 = n7616 & n7665 ;
  assign n7667 = n7666 ^ n4851 ;
  assign n7668 = n7667 ^ n7613 ;
  assign n7669 = ~n7614 & ~n7668 ;
  assign n7670 = n7669 ^ n4862 ;
  assign n7671 = n7670 ^ n7611 ;
  assign n7672 = ~n7612 & ~n7671 ;
  assign n7673 = n7672 ^ n4877 ;
  assign n7674 = n7673 ^ n4885 ;
  assign n7675 = n7544 ^ n7538 ;
  assign n7676 = n7675 ^ n7673 ;
  assign n7677 = ~n7674 & n7676 ;
  assign n7678 = n7677 ^ n4885 ;
  assign n7680 = n7679 ^ n7678 ;
  assign n7681 = n7679 ^ n4902 ;
  assign n7682 = ~n7680 & ~n7681 ;
  assign n7683 = n7682 ^ n4902 ;
  assign n7610 = n7555 ^ n7369 ;
  assign n7684 = n7683 ^ n7610 ;
  assign n7685 = n4972 ^ n4932 ;
  assign n7686 = n7685 ^ n7610 ;
  assign n7687 = n7686 ^ n4972 ;
  assign n7688 = n7684 & ~n7687 ;
  assign n7689 = n7688 ^ n7685 ;
  assign n7690 = n7609 & n7689 ;
  assign n7691 = n7690 ^ n7608 ;
  assign n7607 = n7575 ^ n7567 ;
  assign n7692 = n7691 ^ n7607 ;
  assign n7693 = n7691 ^ n4956 ;
  assign n7694 = n7692 & ~n7693 ;
  assign n7695 = n7694 ^ n4956 ;
  assign n7696 = n7695 ^ n4952 ;
  assign n7697 = n7577 ^ n7364 ;
  assign n7698 = n7697 ^ n7695 ;
  assign n7699 = ~n7696 & n7698 ;
  assign n7700 = n7699 ^ n7697 ;
  assign n7702 = n7701 ^ n7700 ;
  assign n7703 = n7701 ^ n5067 ;
  assign n7704 = ~n7702 & n7703 ;
  assign n7705 = n7704 ^ n5067 ;
  assign n7706 = n7705 ^ n5101 ;
  assign n7707 = n7586 ^ n7583 ;
  assign n7708 = n7707 ^ n5101 ;
  assign n7709 = n7706 & ~n7708 ;
  assign n7710 = n7709 ^ n7707 ;
  assign n7711 = n7710 ^ n7605 ;
  assign n7712 = ~n7606 & ~n7711 ;
  assign n7713 = n7712 ^ n5130 ;
  assign n7714 = n7713 ^ n5164 ;
  assign n7715 = n7599 ^ n7598 ;
  assign n7716 = n7715 ^ n7713 ;
  assign n7717 = ~n7714 & ~n7716 ;
  assign n7718 = n7717 ^ n5164 ;
  assign n7719 = n7718 ^ n7603 ;
  assign n7720 = n7604 & ~n7719 ;
  assign n7721 = n7720 ^ n5197 ;
  assign n7722 = n7721 ^ n4540 ;
  assign n7732 = n7731 ^ n7730 ;
  assign n7733 = n7732 ^ n7721 ;
  assign n7734 = ~n7722 & ~n7733 ;
  assign n7735 = n7734 ^ n4540 ;
  assign n7736 = n7735 ^ n4550 ;
  assign n7747 = n7746 ^ n7744 ;
  assign n7949 = n7747 ^ n7735 ;
  assign n7950 = ~n7736 & ~n7949 ;
  assign n7951 = n7950 ^ n4550 ;
  assign n7952 = n7951 ^ n4535 ;
  assign n7948 = n7947 ^ n7946 ;
  assign n7975 = n7951 ^ n7948 ;
  assign n7976 = n7952 & ~n7975 ;
  assign n7977 = n7976 ^ n4535 ;
  assign n7978 = n7977 ^ n4532 ;
  assign n7989 = n7988 ^ n7986 ;
  assign n8002 = n7989 ^ n7977 ;
  assign n8006 = n7978 & ~n8002 ;
  assign n8003 = n4532 ^ n4524 ;
  assign n8007 = n8006 ^ n8003 ;
  assign n8018 = n8017 ^ n8007 ;
  assign n7748 = n7747 ^ n7736 ;
  assign n7749 = n7718 ^ n7604 ;
  assign n7750 = n7715 ^ n7714 ;
  assign n7751 = n7700 ^ n5067 ;
  assign n7752 = n7751 ^ n7701 ;
  assign n7753 = n7661 ^ n4829 ;
  assign n7754 = n7753 ^ n7617 ;
  assign n7755 = n7658 ^ n7620 ;
  assign n7320 = n7319 ^ n7316 ;
  assign n7321 = n7317 ^ n4569 ;
  assign n7756 = n7320 & ~n7321 ;
  assign n7757 = n7634 ^ n7629 ;
  assign n7758 = n7756 & n7757 ;
  assign n7759 = n7636 ^ n7628 ;
  assign n7760 = ~n7758 & n7759 ;
  assign n7761 = n7639 ^ n4683 ;
  assign n7762 = n7761 ^ n7625 ;
  assign n7763 = n7760 & ~n7762 ;
  assign n7764 = n7642 ^ n7624 ;
  assign n7765 = ~n7763 & ~n7764 ;
  assign n7766 = n7645 ^ n4706 ;
  assign n7767 = n7766 ^ n7621 ;
  assign n7768 = n7765 & n7767 ;
  assign n7769 = n7649 ^ n4725 ;
  assign n7770 = n7769 ^ n7648 ;
  assign n7771 = ~n7768 & ~n7770 ;
  assign n7772 = n7653 ^ n4745 ;
  assign n7773 = n7772 ^ n7654 ;
  assign n7774 = n7771 & n7773 ;
  assign n7775 = n7755 & ~n7774 ;
  assign n7776 = n7754 & n7775 ;
  assign n7777 = n7664 ^ n7616 ;
  assign n7778 = ~n7776 & n7777 ;
  assign n7779 = n7667 ^ n4862 ;
  assign n7780 = n7779 ^ n7613 ;
  assign n7781 = n7778 & n7780 ;
  assign n7782 = n7670 ^ n7612 ;
  assign n7783 = n7781 & ~n7782 ;
  assign n7784 = n7675 ^ n7674 ;
  assign n7785 = n7783 & ~n7784 ;
  assign n7786 = n7681 ^ n7678 ;
  assign n7787 = ~n7785 & n7786 ;
  assign n7788 = n7610 ^ n4932 ;
  assign n7789 = n7788 ^ n7683 ;
  assign n7790 = n7787 & ~n7789 ;
  assign n7791 = n7689 ^ n7608 ;
  assign n7792 = ~n7790 & ~n7791 ;
  assign n7793 = n7693 ^ n7607 ;
  assign n7794 = ~n7792 & ~n7793 ;
  assign n7795 = n7697 ^ n4952 ;
  assign n7796 = n7795 ^ n7695 ;
  assign n7797 = n7794 & n7796 ;
  assign n7798 = n7752 & n7797 ;
  assign n7799 = n7708 ^ n7705 ;
  assign n7800 = n7798 & ~n7799 ;
  assign n7801 = n7710 ^ n5130 ;
  assign n7802 = n7801 ^ n7605 ;
  assign n7803 = n7800 & ~n7802 ;
  assign n7804 = ~n7750 & ~n7803 ;
  assign n7805 = n7749 & ~n7804 ;
  assign n7806 = n7732 ^ n7722 ;
  assign n7807 = ~n7805 & n7806 ;
  assign n7938 = n7748 & ~n7807 ;
  assign n7953 = n7952 ^ n7948 ;
  assign n7974 = ~n7938 & ~n7953 ;
  assign n7990 = n7989 ^ n7978 ;
  assign n8001 = n7974 & ~n7990 ;
  assign n8019 = n8018 ^ n8001 ;
  assign n8020 = n8019 ^ x258 ;
  assign n7991 = n7990 ^ n7974 ;
  assign n7954 = n7953 ^ n7938 ;
  assign n7808 = n7807 ^ n7748 ;
  assign n7809 = n7808 ^ x261 ;
  assign n7810 = n7806 ^ n7805 ;
  assign n7811 = n7810 ^ x262 ;
  assign n7926 = n7804 ^ n7749 ;
  assign n7812 = n7803 ^ n7750 ;
  assign n7813 = n7812 ^ x264 ;
  assign n7814 = n7802 ^ n7800 ;
  assign n7815 = n7814 ^ x265 ;
  assign n7816 = n7799 ^ n7798 ;
  assign n7817 = n7816 ^ x266 ;
  assign n7912 = n7797 ^ n7752 ;
  assign n7818 = n7793 ^ n7792 ;
  assign n7819 = n7818 ^ x269 ;
  assign n7820 = n7791 ^ n7790 ;
  assign n7821 = n7820 ^ x270 ;
  assign n7822 = n7789 ^ n7787 ;
  assign n7823 = n7822 ^ x271 ;
  assign n7825 = n7784 ^ n7783 ;
  assign n7826 = n7825 ^ x273 ;
  assign n7827 = n7782 ^ n7781 ;
  assign n7828 = n7827 ^ x274 ;
  assign n7829 = n7780 ^ n7778 ;
  assign n7830 = n7829 ^ x275 ;
  assign n7831 = n7777 ^ n7776 ;
  assign n7832 = n7831 ^ x276 ;
  assign n7834 = n7774 ^ n7755 ;
  assign n7835 = n7834 ^ x278 ;
  assign n7836 = n7773 ^ n7771 ;
  assign n7837 = n7836 ^ x279 ;
  assign n7838 = n7770 ^ n7768 ;
  assign n7839 = n7838 ^ x280 ;
  assign n7840 = n7767 ^ n7765 ;
  assign n7841 = n7840 ^ x281 ;
  assign n7842 = n7764 ^ n7763 ;
  assign n7843 = n7842 ^ x282 ;
  assign n7857 = n7762 ^ n7760 ;
  assign n7844 = n7759 ^ n7758 ;
  assign n7845 = n7844 ^ x284 ;
  assign n7323 = x287 & n7321 ;
  assign n7324 = n7323 ^ x286 ;
  assign n7322 = n7321 ^ n7320 ;
  assign n7847 = n7323 ^ n7322 ;
  assign n7848 = n7324 & n7847 ;
  assign n7849 = n7848 ^ x286 ;
  assign n7846 = n7757 ^ n7756 ;
  assign n7850 = n7849 ^ n7846 ;
  assign n7851 = n7849 ^ x285 ;
  assign n7852 = ~n7850 & n7851 ;
  assign n7853 = n7852 ^ x285 ;
  assign n7854 = n7853 ^ n7844 ;
  assign n7855 = n7845 & ~n7854 ;
  assign n7856 = n7855 ^ x284 ;
  assign n7858 = n7857 ^ n7856 ;
  assign n7859 = n7857 ^ x283 ;
  assign n7860 = ~n7858 & n7859 ;
  assign n7861 = n7860 ^ x283 ;
  assign n7862 = n7861 ^ n7842 ;
  assign n7863 = n7843 & ~n7862 ;
  assign n7864 = n7863 ^ x282 ;
  assign n7865 = n7864 ^ n7840 ;
  assign n7866 = n7841 & ~n7865 ;
  assign n7867 = n7866 ^ x281 ;
  assign n7868 = n7867 ^ n7838 ;
  assign n7869 = ~n7839 & n7868 ;
  assign n7870 = n7869 ^ x280 ;
  assign n7871 = n7870 ^ n7836 ;
  assign n7872 = ~n7837 & n7871 ;
  assign n7873 = n7872 ^ x279 ;
  assign n7874 = n7873 ^ n7834 ;
  assign n7875 = ~n7835 & n7874 ;
  assign n7876 = n7875 ^ x278 ;
  assign n7833 = n7775 ^ n7754 ;
  assign n7877 = n7876 ^ n7833 ;
  assign n7878 = n7876 ^ x277 ;
  assign n7879 = ~n7877 & n7878 ;
  assign n7880 = n7879 ^ x277 ;
  assign n7881 = n7880 ^ n7831 ;
  assign n7882 = n7832 & ~n7881 ;
  assign n7883 = n7882 ^ x276 ;
  assign n7884 = n7883 ^ n7829 ;
  assign n7885 = ~n7830 & n7884 ;
  assign n7886 = n7885 ^ x275 ;
  assign n7887 = n7886 ^ n7827 ;
  assign n7888 = n7828 & ~n7887 ;
  assign n7889 = n7888 ^ x274 ;
  assign n7890 = n7889 ^ n7825 ;
  assign n7891 = n7826 & ~n7890 ;
  assign n7892 = n7891 ^ x273 ;
  assign n7824 = n7786 ^ n7785 ;
  assign n7893 = n7892 ^ n7824 ;
  assign n7894 = n7822 ^ x272 ;
  assign n7895 = n7894 ^ n7822 ;
  assign n7896 = n7895 ^ n7824 ;
  assign n7897 = n7893 & ~n7896 ;
  assign n7898 = n7897 ^ n7894 ;
  assign n7899 = ~n7823 & n7898 ;
  assign n7900 = n7899 ^ x271 ;
  assign n7901 = n7900 ^ n7820 ;
  assign n7902 = ~n7821 & n7901 ;
  assign n7903 = n7902 ^ x270 ;
  assign n7904 = n7903 ^ n7818 ;
  assign n7905 = n7819 & ~n7904 ;
  assign n7906 = n7905 ^ x269 ;
  assign n7907 = n7906 ^ x268 ;
  assign n7908 = n7796 ^ n7794 ;
  assign n7909 = n7908 ^ n7906 ;
  assign n7910 = n7907 & ~n7909 ;
  assign n7911 = n7910 ^ x268 ;
  assign n7913 = n7912 ^ n7911 ;
  assign n7914 = n7912 ^ x267 ;
  assign n7915 = ~n7913 & n7914 ;
  assign n7916 = n7915 ^ x267 ;
  assign n7917 = n7916 ^ n7816 ;
  assign n7918 = ~n7817 & n7917 ;
  assign n7919 = n7918 ^ x266 ;
  assign n7920 = n7919 ^ n7814 ;
  assign n7921 = ~n7815 & n7920 ;
  assign n7922 = n7921 ^ x265 ;
  assign n7923 = n7922 ^ n7812 ;
  assign n7924 = ~n7813 & n7923 ;
  assign n7925 = n7924 ^ x264 ;
  assign n7927 = n7926 ^ n7925 ;
  assign n7928 = n7926 ^ x263 ;
  assign n7929 = n7927 & ~n7928 ;
  assign n7930 = n7929 ^ x263 ;
  assign n7931 = n7930 ^ n7810 ;
  assign n7932 = n7811 & ~n7931 ;
  assign n7933 = n7932 ^ x262 ;
  assign n7934 = n7933 ^ n7808 ;
  assign n7935 = ~n7809 & n7934 ;
  assign n7936 = n7935 ^ x261 ;
  assign n7969 = n7954 ^ n7936 ;
  assign n7970 = n7954 ^ x260 ;
  assign n7971 = n7969 & ~n7970 ;
  assign n7972 = n7971 ^ x260 ;
  assign n7997 = n7991 ^ n7972 ;
  assign n7998 = n7991 ^ x259 ;
  assign n7999 = ~n7997 & n7998 ;
  assign n8000 = n7999 ^ x259 ;
  assign n8021 = n8020 ^ n8000 ;
  assign n7937 = n7936 ^ x260 ;
  assign n7955 = n7954 ^ n7937 ;
  assign n7956 = n6841 ^ n5753 ;
  assign n7957 = n7401 & n7956 ;
  assign n7958 = n7957 ^ n6841 ;
  assign n7959 = ~n7955 & ~n7958 ;
  assign n7960 = n7959 ^ n5750 ;
  assign n7961 = n7960 ^ n6935 ;
  assign n7962 = n7961 ^ n7959 ;
  assign n7963 = n7334 & n7962 ;
  assign n7964 = n7963 ^ n7960 ;
  assign n7973 = n7972 ^ x259 ;
  assign n7992 = n7991 ^ n7973 ;
  assign n7965 = n6929 ^ n5239 ;
  assign n7966 = ~n7386 & n7965 ;
  assign n7967 = n7966 ^ n6929 ;
  assign n7968 = n7967 ^ n7959 ;
  assign n7993 = n7992 ^ n7968 ;
  assign n7994 = n7993 ^ n7967 ;
  assign n7995 = n7964 & n7994 ;
  assign n7996 = n7995 ^ n7968 ;
  assign n8120 = n8021 ^ n7996 ;
  assign n8112 = n7958 ^ n7955 ;
  assign n8113 = ~n5313 & n8112 ;
  assign n8114 = n8113 ^ n5323 ;
  assign n8115 = n7992 ^ n7964 ;
  assign n8116 = n8115 ^ n8113 ;
  assign n8117 = n8114 & ~n8116 ;
  assign n8118 = n8117 ^ n5323 ;
  assign n8119 = n8118 ^ n5288 ;
  assign n8165 = n8120 ^ n8119 ;
  assign n8162 = n8112 ^ n5313 ;
  assign n8163 = n8115 ^ n8114 ;
  assign n8164 = ~n8162 & n8163 ;
  assign n8212 = n8165 ^ n8164 ;
  assign n8206 = x319 & n8162 ;
  assign n8207 = n8206 ^ x318 ;
  assign n8208 = n8163 ^ n8162 ;
  assign n8209 = n8208 ^ n8206 ;
  assign n8210 = n8207 & n8209 ;
  assign n8211 = n8210 ^ x318 ;
  assign n8213 = n8212 ^ n8211 ;
  assign n8214 = n8212 ^ x317 ;
  assign n8215 = ~n8213 & n8214 ;
  assign n8216 = n8215 ^ x317 ;
  assign n8925 = n8216 ^ x316 ;
  assign n8051 = n8019 ^ n8000 ;
  assign n8052 = n8020 & ~n8051 ;
  assign n8053 = n8052 ^ x258 ;
  assign n8054 = n8053 ^ x257 ;
  assign n8049 = ~n8001 & ~n8018 ;
  assign n8044 = n8017 ^ n4524 ;
  assign n8045 = n8007 & ~n8044 ;
  assign n8046 = n8045 ^ n4524 ;
  assign n8047 = n8046 ^ n3990 ;
  assign n8040 = n6130 ^ n5300 ;
  assign n8041 = n6711 & ~n8040 ;
  assign n8042 = n8041 ^ n5300 ;
  assign n8033 = n7278 ^ x230 ;
  assign n8034 = n8033 ^ n7188 ;
  assign n8035 = n8034 ^ n8011 ;
  assign n8036 = n8035 ^ n8034 ;
  assign n8037 = n8036 ^ n8010 ;
  assign n8038 = ~n8016 & ~n8037 ;
  assign n8039 = n8038 ^ n8035 ;
  assign n8043 = n8042 ^ n8039 ;
  assign n8048 = n8047 ^ n8043 ;
  assign n8050 = n8049 ^ n8048 ;
  assign n8055 = n8054 ^ n8050 ;
  assign n8024 = n6924 ^ n5738 ;
  assign n8025 = ~n7377 & ~n8024 ;
  assign n8026 = n8025 ^ n6924 ;
  assign n8027 = n8026 ^ n8021 ;
  assign n8022 = n8021 ^ n7967 ;
  assign n8023 = n7996 & ~n8022 ;
  assign n8028 = n8027 ^ n8023 ;
  assign n8124 = n8055 ^ n8028 ;
  assign n8126 = n8124 ^ n5279 ;
  assign n8121 = n8120 ^ n8118 ;
  assign n8122 = ~n8119 & n8121 ;
  assign n8123 = n8122 ^ n5288 ;
  assign n8167 = n8126 ^ n8123 ;
  assign n8166 = n8164 & n8165 ;
  assign n8204 = n8167 ^ n8166 ;
  assign n8926 = n8925 ^ n8204 ;
  assign n8322 = n7870 ^ x279 ;
  assign n8323 = n8322 ^ n7836 ;
  assign n8922 = n7547 ^ n6913 ;
  assign n8923 = ~n8323 & n8922 ;
  assign n8924 = n8923 ^ n6913 ;
  assign n8927 = n8926 ^ n8924 ;
  assign n8931 = n8214 ^ n8211 ;
  assign n8305 = n7867 ^ x280 ;
  assign n8306 = n8305 ^ n7838 ;
  assign n8928 = n7370 ^ n6981 ;
  assign n8929 = ~n8306 & n8928 ;
  assign n8930 = n8929 ^ n6981 ;
  assign n8932 = n8931 ^ n8930 ;
  assign n8936 = n8208 ^ n8207 ;
  assign n8308 = n7864 ^ n7841 ;
  assign n8933 = n7535 ^ n6854 ;
  assign n8934 = n8308 & ~n8933 ;
  assign n8935 = n8934 ^ n6854 ;
  assign n8937 = n8936 ^ n8935 ;
  assign n8770 = n8162 ^ x319 ;
  assign n8184 = n7861 ^ x282 ;
  assign n8185 = n8184 ^ n7842 ;
  assign n8767 = n6967 ^ n6851 ;
  assign n8768 = n8185 & ~n8767 ;
  assign n8769 = n8768 ^ n6967 ;
  assign n8771 = n8770 ^ n8769 ;
  assign n8156 = n7859 ^ n7856 ;
  assign n8738 = n6919 ^ n6852 ;
  assign n8739 = n8156 & n8738 ;
  assign n8740 = n8739 ^ n6919 ;
  assign n8496 = n7922 ^ x264 ;
  assign n8497 = n8496 ^ n7812 ;
  assign n8245 = n7908 ^ n7907 ;
  assign n8246 = n8245 ^ n6686 ;
  assign n8247 = n8246 ^ n7453 ;
  assign n8248 = n8247 ^ n8245 ;
  assign n8249 = ~n8011 & n8248 ;
  assign n8250 = n8249 ^ n8246 ;
  assign n8257 = n7421 ^ n6664 ;
  assign n8258 = n7988 & n8257 ;
  assign n8259 = n8258 ^ n6664 ;
  assign n8256 = n7903 ^ n7819 ;
  assign n8260 = n8259 ^ n8256 ;
  assign n8263 = n7336 ^ n6646 ;
  assign n8264 = ~n7947 & ~n8263 ;
  assign n8265 = n8264 ^ n6646 ;
  assign n8261 = n7900 ^ x270 ;
  assign n8262 = n8261 ^ n7820 ;
  assign n8266 = n8265 ^ n8262 ;
  assign n8268 = n7306 ^ n6431 ;
  assign n8269 = n7746 & ~n8268 ;
  assign n8270 = n8269 ^ n6431 ;
  assign n8267 = n7898 ^ x271 ;
  assign n8271 = n8270 ^ n8267 ;
  assign n8274 = n7182 ^ n6278 ;
  assign n8275 = n7731 & ~n8274 ;
  assign n8276 = n8275 ^ n6278 ;
  assign n8272 = n7892 ^ x272 ;
  assign n8273 = n8272 ^ n7824 ;
  assign n8277 = n8276 ^ n8273 ;
  assign n8279 = n7121 ^ n5685 ;
  assign n8280 = n7338 & n8279 ;
  assign n8281 = n8280 ^ n5685 ;
  assign n8278 = n7889 ^ n7826 ;
  assign n8282 = n8281 ^ n8278 ;
  assign n8290 = n7880 ^ x276 ;
  assign n8291 = n8290 ^ n7831 ;
  assign n8287 = n6873 ^ n6239 ;
  assign n8288 = n7357 & n8287 ;
  assign n8289 = n8288 ^ n6239 ;
  assign n8292 = n8291 ^ n8289 ;
  assign n8293 = n7833 ^ x277 ;
  assign n8294 = n8293 ^ n7876 ;
  assign n8295 = n8294 ^ n6230 ;
  assign n8296 = n8295 ^ n6879 ;
  assign n8297 = n8296 ^ n8294 ;
  assign n8298 = n7351 & n8297 ;
  assign n8299 = n8298 ^ n8295 ;
  assign n8332 = n7873 ^ n7835 ;
  assign n8302 = n6898 ^ n6203 ;
  assign n8303 = n7559 & ~n8302 ;
  assign n8304 = n8303 ^ n6203 ;
  assign n8307 = n8306 ^ n8304 ;
  assign n8309 = n6900 ^ n6195 ;
  assign n8310 = ~n7368 & ~n8309 ;
  assign n8311 = n8310 ^ n6195 ;
  assign n8312 = n8311 ^ n8308 ;
  assign n8187 = n8185 ^ n6197 ;
  assign n8186 = n8185 ^ n6905 ;
  assign n8188 = n8187 ^ n8186 ;
  assign n8189 = ~n7547 & n8188 ;
  assign n8190 = n8189 ^ n8187 ;
  assign n8098 = n6913 ^ n6181 ;
  assign n8099 = ~n7535 & ~n8098 ;
  assign n8100 = n8099 ^ n6181 ;
  assign n8094 = n7846 ^ x285 ;
  assign n8095 = n8094 ^ n7849 ;
  assign n8101 = n8100 ^ n8095 ;
  assign n7325 = n7324 ^ n7322 ;
  assign n6855 = n6854 ^ n5718 ;
  assign n6856 = n6852 & n6855 ;
  assign n6857 = n6856 ^ n5718 ;
  assign n7326 = n7325 ^ n6857 ;
  assign n7332 = n7321 ^ x287 ;
  assign n8085 = n7332 ^ n7325 ;
  assign n7329 = n6967 ^ n5727 ;
  assign n7330 = ~n7328 & n7329 ;
  assign n7331 = n7330 ^ n5727 ;
  assign n7333 = n7332 ^ n7331 ;
  assign n8074 = n8042 ^ n8034 ;
  assign n8075 = ~n8039 & n8074 ;
  assign n8071 = n6139 ^ n5308 ;
  assign n8072 = n6705 & n8071 ;
  assign n8067 = n8042 ^ n7458 ;
  assign n8066 = n7281 ^ n7187 ;
  assign n8068 = n8067 ^ n8066 ;
  assign n8069 = n8068 ^ n3990 ;
  assign n8065 = x257 ^ x256 ;
  assign n8070 = n8069 ^ n8065 ;
  assign n8073 = n8072 ^ n8070 ;
  assign n8076 = n8075 ^ n8073 ;
  assign n8064 = ~n8048 & ~n8049 ;
  assign n8077 = n8076 ^ n8064 ;
  assign n8062 = n8053 ^ n8050 ;
  assign n8063 = n8054 & n8062 ;
  assign n8078 = n8077 ^ n8063 ;
  assign n8060 = n8046 ^ n8043 ;
  assign n8061 = ~n8047 & n8060 ;
  assign n8079 = n8078 ^ n8061 ;
  assign n8082 = n8079 ^ n7331 ;
  assign n8029 = n6919 ^ n5732 ;
  assign n8030 = ~n7506 & n8029 ;
  assign n8031 = n8030 ^ n6919 ;
  assign n8032 = n8031 ^ n8026 ;
  assign n8056 = n8055 ^ n8032 ;
  assign n8057 = n8056 ^ n8031 ;
  assign n8058 = n8028 & ~n8057 ;
  assign n8059 = n8058 ^ n8032 ;
  assign n8080 = n8079 ^ n8031 ;
  assign n8081 = ~n8059 & ~n8080 ;
  assign n8083 = n8082 ^ n8081 ;
  assign n8084 = n7333 & n8083 ;
  assign n8086 = n8085 ^ n8084 ;
  assign n8087 = ~n7326 & ~n8086 ;
  assign n8088 = n8087 ^ n7325 ;
  assign n8089 = n8088 ^ n6173 ;
  assign n8090 = n8089 ^ n6981 ;
  assign n8091 = n8090 ^ n8088 ;
  assign n8092 = ~n6851 & ~n8091 ;
  assign n8093 = n8092 ^ n8089 ;
  assign n8096 = n8095 ^ n8088 ;
  assign n8097 = n8093 & ~n8096 ;
  assign n8102 = n8101 ^ n8097 ;
  assign n8103 = n7853 ^ x284 ;
  assign n8104 = n8103 ^ n7844 ;
  assign n8148 = n8104 ^ n8100 ;
  assign n8149 = n8102 & n8148 ;
  assign n8150 = n8149 ^ n8100 ;
  assign n8151 = n8150 ^ n6907 ;
  assign n8152 = n8151 ^ n5713 ;
  assign n8153 = n8152 ^ n8150 ;
  assign n8154 = n7370 & n8153 ;
  assign n8155 = n8154 ^ n8151 ;
  assign n8191 = n8156 ^ n8150 ;
  assign n8192 = n8155 & n8191 ;
  assign n8193 = n8192 ^ n8156 ;
  assign n8313 = n8193 ^ n8185 ;
  assign n8314 = n8190 & n8313 ;
  assign n8315 = n8314 ^ n8185 ;
  assign n8316 = n8315 ^ n8308 ;
  assign n8317 = ~n8312 & ~n8316 ;
  assign n8318 = n8317 ^ n8311 ;
  assign n8319 = n8318 ^ n8304 ;
  assign n8320 = n8307 & ~n8319 ;
  assign n8321 = n8320 ^ n8306 ;
  assign n8324 = n8323 ^ n8321 ;
  assign n8326 = n8323 ^ n6215 ;
  assign n8325 = n8323 ^ n6890 ;
  assign n8327 = n8326 ^ n8325 ;
  assign n8328 = n7569 & n8327 ;
  assign n8329 = n8328 ^ n8326 ;
  assign n8330 = n8324 & ~n8329 ;
  assign n8331 = n8330 ^ n8323 ;
  assign n8333 = n8332 ^ n8331 ;
  assign n8334 = n8332 ^ n6224 ;
  assign n8335 = n8334 ^ n6887 ;
  assign n8336 = n8335 ^ n8332 ;
  assign n8337 = n7363 & ~n8336 ;
  assign n8338 = n8337 ^ n8334 ;
  assign n8339 = n8333 & n8338 ;
  assign n8340 = n8339 ^ n8332 ;
  assign n8341 = n8340 ^ n8294 ;
  assign n8342 = ~n8299 & ~n8341 ;
  assign n8300 = n8294 ^ n8289 ;
  assign n8343 = n8342 ^ n8300 ;
  assign n8344 = n8292 & ~n8343 ;
  assign n8345 = n8344 ^ n8291 ;
  assign n8286 = n7883 ^ n7830 ;
  assign n8346 = n8345 ^ n8286 ;
  assign n8347 = n6868 ^ n6249 ;
  assign n8348 = n7345 & n8347 ;
  assign n8349 = n8348 ^ n6249 ;
  assign n8350 = n8349 ^ n8286 ;
  assign n8351 = ~n8346 & n8350 ;
  assign n8352 = n8351 ^ n8345 ;
  assign n8283 = n6861 ^ n6270 ;
  assign n8284 = ~n7599 & n8283 ;
  assign n8285 = n8284 ^ n6270 ;
  assign n8353 = n8352 ^ n8285 ;
  assign n8354 = n7886 ^ x274 ;
  assign n8355 = n8354 ^ n7827 ;
  assign n8356 = n8355 ^ n8352 ;
  assign n8357 = ~n8353 & n8356 ;
  assign n8358 = n8357 ^ n8355 ;
  assign n8359 = n8358 ^ n8278 ;
  assign n8360 = n8282 & ~n8359 ;
  assign n8361 = n8360 ^ n8281 ;
  assign n8362 = n8361 ^ n8273 ;
  assign n8363 = ~n8277 & n8362 ;
  assign n8364 = n8363 ^ n8276 ;
  assign n8365 = n8364 ^ n8267 ;
  assign n8366 = ~n8271 & n8365 ;
  assign n8367 = n8366 ^ n8270 ;
  assign n8368 = n8367 ^ n8262 ;
  assign n8369 = n8266 & n8368 ;
  assign n8370 = n8369 ^ n8265 ;
  assign n8371 = n8370 ^ n8256 ;
  assign n8372 = n8260 & n8371 ;
  assign n8373 = n8372 ^ n8259 ;
  assign n8251 = n6715 ^ n6106 ;
  assign n8252 = ~n8034 & ~n8251 ;
  assign n8253 = n8252 ^ n6106 ;
  assign n8254 = n8253 ^ n8245 ;
  assign n8255 = n8254 ^ n8253 ;
  assign n8374 = n8373 ^ n8255 ;
  assign n8375 = n8250 & n8374 ;
  assign n8376 = n8375 ^ n8254 ;
  assign n8458 = n6714 ^ n6101 ;
  assign n8459 = ~n8066 & n8458 ;
  assign n8460 = n8459 ^ n6101 ;
  assign n8377 = n7914 ^ n7911 ;
  assign n8462 = n8460 ^ n8377 ;
  assign n8461 = n8460 ^ n8253 ;
  assign n8463 = n8462 ^ n8461 ;
  assign n8464 = ~n8376 & ~n8463 ;
  assign n8465 = n8464 ^ n8461 ;
  assign n8473 = n6729 ^ n6100 ;
  assign n8474 = ~n7286 & n8473 ;
  assign n8475 = n8474 ^ n6100 ;
  assign n8477 = n8475 ^ n8460 ;
  assign n8466 = n7916 ^ x266 ;
  assign n8467 = n8466 ^ n7816 ;
  assign n8476 = n8475 ^ n8467 ;
  assign n8478 = n8477 ^ n8476 ;
  assign n8479 = ~n8465 & ~n8478 ;
  assign n8480 = n8479 ^ n8477 ;
  assign n8488 = n6711 ^ n6098 ;
  assign n8489 = ~n7315 & n8488 ;
  assign n8490 = n8489 ^ n6098 ;
  assign n8492 = n8490 ^ n8475 ;
  assign n8481 = n7919 ^ n7815 ;
  assign n8491 = n8490 ^ n8481 ;
  assign n8493 = n8492 ^ n8491 ;
  assign n8494 = n8480 & ~n8493 ;
  assign n8495 = n8494 ^ n8492 ;
  assign n8498 = n8497 ^ n8495 ;
  assign n8482 = n8481 ^ n8480 ;
  assign n8468 = n8467 ^ n8465 ;
  assign n8378 = n8377 ^ n8376 ;
  assign n8379 = n8378 ^ n5082 ;
  assign n8380 = n8373 ^ n8250 ;
  assign n8381 = n8380 ^ n5691 ;
  assign n8383 = n8367 ^ n8266 ;
  assign n8384 = n8383 ^ n5773 ;
  assign n8386 = n8361 ^ n8277 ;
  assign n8387 = n8386 ^ n5865 ;
  assign n8433 = n8358 ^ n8282 ;
  assign n8388 = n8355 ^ n8285 ;
  assign n8389 = n8388 ^ n8352 ;
  assign n8390 = n8389 ^ n5860 ;
  assign n8392 = n8343 ^ n8291 ;
  assign n8393 = n8392 ^ n5796 ;
  assign n8418 = n8340 ^ n8299 ;
  assign n8394 = n8338 ^ n8331 ;
  assign n8395 = n8394 ^ n5671 ;
  assign n8397 = n8318 ^ n8307 ;
  assign n8398 = n8397 ^ n5463 ;
  assign n8194 = n8193 ^ n8190 ;
  assign n8400 = n8194 ^ n5250 ;
  assign n8105 = n8104 ^ n8102 ;
  assign n8106 = n8105 ^ n5346 ;
  assign n8108 = n8086 ^ n6857 ;
  assign n8109 = n8108 ^ n5268 ;
  assign n8110 = n8079 ^ n8059 ;
  assign n8111 = n8110 ^ n5240 ;
  assign n8125 = n8124 ^ n8123 ;
  assign n8127 = ~n8125 & ~n8126 ;
  assign n8128 = n8127 ^ n5279 ;
  assign n8129 = n8128 ^ n8110 ;
  assign n8130 = ~n8111 & n8129 ;
  assign n8131 = n8130 ^ n5240 ;
  assign n8132 = n8131 ^ n5270 ;
  assign n8133 = n8083 ^ n7332 ;
  assign n8134 = n8133 ^ n8131 ;
  assign n8135 = ~n8132 & n8134 ;
  assign n8136 = n8135 ^ n5270 ;
  assign n8137 = n8136 ^ n8108 ;
  assign n8138 = n8109 & ~n8137 ;
  assign n8139 = n8138 ^ n5268 ;
  assign n8107 = n8095 ^ n8093 ;
  assign n8140 = n8139 ^ n8107 ;
  assign n8141 = n8139 ^ n5260 ;
  assign n8142 = ~n8140 & n8141 ;
  assign n8143 = n8142 ^ n5260 ;
  assign n8144 = n8143 ^ n8105 ;
  assign n8145 = ~n8106 & n8144 ;
  assign n8146 = n8145 ^ n5346 ;
  assign n8147 = n8146 ^ n4699 ;
  assign n8157 = n8156 ^ n8155 ;
  assign n8180 = n8157 ^ n8146 ;
  assign n8181 = ~n8147 & n8180 ;
  assign n8182 = n8181 ^ n8157 ;
  assign n8401 = n8194 ^ n8182 ;
  assign n8402 = n8400 & n8401 ;
  assign n8403 = n8402 ^ n5250 ;
  assign n8399 = n8315 ^ n8312 ;
  assign n8404 = n8403 ^ n8399 ;
  assign n8405 = n8403 ^ n5441 ;
  assign n8406 = n8404 & ~n8405 ;
  assign n8407 = n8406 ^ n5441 ;
  assign n8408 = n8407 ^ n8397 ;
  assign n8409 = n8398 & ~n8408 ;
  assign n8410 = n8409 ^ n5463 ;
  assign n8396 = n8329 ^ n8321 ;
  assign n8411 = n8410 ^ n8396 ;
  assign n8412 = n8396 ^ n5525 ;
  assign n8413 = ~n8411 & n8412 ;
  assign n8414 = n8413 ^ n8410 ;
  assign n8415 = n8414 ^ n8394 ;
  assign n8416 = n8395 & ~n8415 ;
  assign n8417 = n8416 ^ n5671 ;
  assign n8419 = n8418 ^ n8417 ;
  assign n8420 = n8417 ^ n5702 ;
  assign n8421 = ~n8419 & ~n8420 ;
  assign n8422 = n8421 ^ n8418 ;
  assign n8423 = n8422 ^ n8392 ;
  assign n8424 = ~n8393 & ~n8423 ;
  assign n8425 = n8424 ^ n5796 ;
  assign n8391 = n8350 ^ n8345 ;
  assign n8426 = n8425 ^ n8391 ;
  assign n8427 = n8391 ^ n5844 ;
  assign n8428 = n8426 & ~n8427 ;
  assign n8429 = n8428 ^ n8425 ;
  assign n8430 = n8429 ^ n8389 ;
  assign n8431 = n8390 & n8430 ;
  assign n8432 = n8431 ^ n5860 ;
  assign n8434 = n8433 ^ n8432 ;
  assign n8435 = n8432 ^ n5852 ;
  assign n8436 = n8434 & ~n8435 ;
  assign n8437 = n8436 ^ n8433 ;
  assign n8438 = n8437 ^ n8386 ;
  assign n8439 = ~n8387 & n8438 ;
  assign n8440 = n8439 ^ n5865 ;
  assign n8385 = n8364 ^ n8271 ;
  assign n8441 = n8440 ^ n8385 ;
  assign n8442 = n8385 ^ n5784 ;
  assign n8443 = ~n8441 & ~n8442 ;
  assign n8444 = n8443 ^ n8440 ;
  assign n8445 = n8444 ^ n8383 ;
  assign n8446 = n8384 & ~n8445 ;
  assign n8447 = n8446 ^ n5773 ;
  assign n8382 = n8370 ^ n8260 ;
  assign n8448 = n8447 ^ n8382 ;
  assign n8449 = n8447 ^ n5765 ;
  assign n8450 = n8448 & n8449 ;
  assign n8451 = n8450 ^ n5765 ;
  assign n8452 = n8451 ^ n8380 ;
  assign n8453 = ~n8381 & ~n8452 ;
  assign n8454 = n8453 ^ n5691 ;
  assign n8455 = n8454 ^ n8378 ;
  assign n8456 = ~n8379 & ~n8455 ;
  assign n8457 = n8456 ^ n5082 ;
  assign n8469 = n8468 ^ n8457 ;
  assign n8470 = n8468 ^ n5114 ;
  assign n8471 = ~n8469 & ~n8470 ;
  assign n8472 = n8471 ^ n5114 ;
  assign n8483 = n8482 ^ n8472 ;
  assign n8484 = n8482 ^ n5145 ;
  assign n8485 = ~n8483 & ~n8484 ;
  assign n8486 = n8485 ^ n5145 ;
  assign n8556 = n8498 ^ n8486 ;
  assign n8557 = n8498 ^ n5181 ;
  assign n8558 = n8556 & ~n8557 ;
  assign n8559 = n8558 ^ n5181 ;
  assign n8560 = n8559 ^ n5206 ;
  assign n8552 = n6705 ^ n6092 ;
  assign n8553 = ~n7475 & n8552 ;
  assign n8554 = n8553 ^ n6092 ;
  assign n8546 = n7928 ^ n7925 ;
  assign n8548 = n8546 ^ n8490 ;
  assign n8547 = n8546 ^ n8497 ;
  assign n8549 = n8548 ^ n8547 ;
  assign n8550 = n8495 & ~n8549 ;
  assign n8551 = n8550 ^ n8548 ;
  assign n8555 = n8554 ^ n8551 ;
  assign n8561 = n8560 ^ n8555 ;
  assign n8487 = n8486 ^ n5181 ;
  assign n8499 = n8498 ^ n8487 ;
  assign n8500 = n8457 ^ n5114 ;
  assign n8501 = n8500 ^ n8468 ;
  assign n8502 = n8444 ^ n5773 ;
  assign n8503 = n8502 ^ n8383 ;
  assign n8504 = n8429 ^ n5860 ;
  assign n8505 = n8504 ^ n8389 ;
  assign n8506 = n8420 ^ n8418 ;
  assign n8507 = n8414 ^ n5671 ;
  assign n8508 = n8507 ^ n8394 ;
  assign n8158 = n8157 ^ n8147 ;
  assign n8159 = n8143 ^ n5346 ;
  assign n8160 = n8159 ^ n8105 ;
  assign n8161 = n8141 ^ n8107 ;
  assign n8168 = ~n8166 & ~n8167 ;
  assign n8169 = n8128 ^ n5240 ;
  assign n8170 = n8169 ^ n8110 ;
  assign n8171 = n8168 & n8170 ;
  assign n8172 = n8133 ^ n8132 ;
  assign n8173 = ~n8171 & n8172 ;
  assign n8174 = n8136 ^ n5268 ;
  assign n8175 = n8174 ^ n8108 ;
  assign n8176 = n8173 & ~n8175 ;
  assign n8177 = n8161 & ~n8176 ;
  assign n8178 = ~n8160 & n8177 ;
  assign n8179 = ~n8158 & ~n8178 ;
  assign n8183 = n8182 ^ n5250 ;
  assign n8195 = n8194 ^ n8183 ;
  assign n8509 = n8179 & ~n8195 ;
  assign n8510 = n8399 ^ n5441 ;
  assign n8511 = n8510 ^ n8403 ;
  assign n8512 = ~n8509 & ~n8511 ;
  assign n8513 = n8407 ^ n5463 ;
  assign n8514 = n8513 ^ n8397 ;
  assign n8515 = n8512 & n8514 ;
  assign n8516 = n8412 ^ n8410 ;
  assign n8517 = n8515 & ~n8516 ;
  assign n8518 = n8508 & n8517 ;
  assign n8519 = n8506 & ~n8518 ;
  assign n8520 = n8422 ^ n8393 ;
  assign n8521 = n8519 & ~n8520 ;
  assign n8522 = n8427 ^ n8425 ;
  assign n8523 = ~n8521 & n8522 ;
  assign n8524 = ~n8505 & ~n8523 ;
  assign n8525 = n8433 ^ n5852 ;
  assign n8526 = n8525 ^ n8432 ;
  assign n8527 = n8524 & n8526 ;
  assign n8528 = n8437 ^ n5865 ;
  assign n8529 = n8528 ^ n8386 ;
  assign n8530 = n8527 & ~n8529 ;
  assign n8531 = n8442 ^ n8440 ;
  assign n8532 = n8530 & n8531 ;
  assign n8533 = n8503 & n8532 ;
  assign n8534 = n8382 ^ n5765 ;
  assign n8535 = n8534 ^ n8447 ;
  assign n8536 = ~n8533 & n8535 ;
  assign n8537 = n8451 ^ n8381 ;
  assign n8538 = ~n8536 & ~n8537 ;
  assign n8539 = n8454 ^ n8379 ;
  assign n8540 = ~n8538 & ~n8539 ;
  assign n8541 = ~n8501 & ~n8540 ;
  assign n8542 = n8472 ^ n5145 ;
  assign n8543 = n8542 ^ n8482 ;
  assign n8544 = ~n8541 & ~n8543 ;
  assign n8545 = n8499 & n8544 ;
  assign n8580 = n8561 ^ n8545 ;
  assign n8581 = n8580 ^ x290 ;
  assign n8673 = n8544 ^ n8499 ;
  assign n8668 = n8543 ^ n8541 ;
  assign n8582 = n8540 ^ n8501 ;
  assign n8583 = n8582 ^ x293 ;
  assign n8584 = n8539 ^ n8538 ;
  assign n8585 = n8584 ^ x294 ;
  assign n8586 = n8537 ^ n8536 ;
  assign n8587 = n8586 ^ x295 ;
  assign n8588 = n8535 ^ n8533 ;
  assign n8589 = n8588 ^ x296 ;
  assign n8590 = n8532 ^ n8503 ;
  assign n8591 = n8590 ^ x297 ;
  assign n8592 = n8531 ^ n8530 ;
  assign n8593 = n8592 ^ x298 ;
  assign n8594 = n8529 ^ n8527 ;
  assign n8595 = n8594 ^ x299 ;
  assign n8642 = n8526 ^ n8524 ;
  assign n8596 = n8523 ^ n8505 ;
  assign n8597 = n8596 ^ x301 ;
  assign n8598 = n8522 ^ n8521 ;
  assign n8599 = n8598 ^ x302 ;
  assign n8600 = n8520 ^ n8519 ;
  assign n8601 = n8600 ^ x303 ;
  assign n8627 = n8518 ^ n8506 ;
  assign n8602 = n8517 ^ n8508 ;
  assign n8603 = n8602 ^ x305 ;
  assign n8604 = n8516 ^ n8515 ;
  assign n8605 = n8604 ^ x306 ;
  assign n8606 = n8514 ^ n8512 ;
  assign n8607 = n8606 ^ x307 ;
  assign n8608 = n8511 ^ n8509 ;
  assign n8609 = n8608 ^ x308 ;
  assign n8198 = n8178 ^ n8158 ;
  assign n8199 = n8198 ^ x310 ;
  assign n8200 = n8176 ^ n8161 ;
  assign n8201 = n8200 ^ x312 ;
  assign n8228 = n8175 ^ n8173 ;
  assign n8202 = n8172 ^ n8171 ;
  assign n8203 = n8202 ^ x314 ;
  assign n8220 = n8170 ^ n8168 ;
  assign n8205 = n8204 ^ x316 ;
  assign n8217 = n8216 ^ n8204 ;
  assign n8218 = ~n8205 & n8217 ;
  assign n8219 = n8218 ^ x316 ;
  assign n8221 = n8220 ^ n8219 ;
  assign n8222 = n8220 ^ x315 ;
  assign n8223 = n8221 & ~n8222 ;
  assign n8224 = n8223 ^ x315 ;
  assign n8225 = n8224 ^ n8202 ;
  assign n8226 = ~n8203 & n8225 ;
  assign n8227 = n8226 ^ x314 ;
  assign n8229 = n8228 ^ n8227 ;
  assign n8230 = n8228 ^ x313 ;
  assign n8231 = n8229 & ~n8230 ;
  assign n8232 = n8231 ^ x313 ;
  assign n8233 = n8232 ^ n8200 ;
  assign n8234 = n8201 & ~n8233 ;
  assign n8235 = n8234 ^ x312 ;
  assign n8236 = n8235 ^ x311 ;
  assign n8237 = n8177 ^ n8160 ;
  assign n8238 = n8237 ^ n8235 ;
  assign n8239 = n8236 & ~n8238 ;
  assign n8240 = n8239 ^ x311 ;
  assign n8241 = n8240 ^ n8198 ;
  assign n8242 = n8199 & ~n8241 ;
  assign n8243 = n8242 ^ x310 ;
  assign n8196 = n8195 ^ n8179 ;
  assign n8610 = n8243 ^ n8196 ;
  assign n8611 = n8608 ^ x309 ;
  assign n8612 = n8611 ^ n8608 ;
  assign n8613 = n8612 ^ n8243 ;
  assign n8614 = n8610 & n8613 ;
  assign n8615 = n8614 ^ n8611 ;
  assign n8616 = ~n8609 & n8615 ;
  assign n8617 = n8616 ^ x308 ;
  assign n8618 = n8617 ^ n8606 ;
  assign n8619 = ~n8607 & n8618 ;
  assign n8620 = n8619 ^ x307 ;
  assign n8621 = n8620 ^ n8604 ;
  assign n8622 = n8605 & ~n8621 ;
  assign n8623 = n8622 ^ x306 ;
  assign n8624 = n8623 ^ n8602 ;
  assign n8625 = ~n8603 & n8624 ;
  assign n8626 = n8625 ^ x305 ;
  assign n8628 = n8627 ^ n8626 ;
  assign n8629 = n8600 ^ x304 ;
  assign n8630 = n8629 ^ n8600 ;
  assign n8631 = n8630 ^ n8626 ;
  assign n8632 = n8628 & n8631 ;
  assign n8633 = n8632 ^ n8629 ;
  assign n8634 = ~n8601 & n8633 ;
  assign n8635 = n8634 ^ x303 ;
  assign n8636 = n8635 ^ n8598 ;
  assign n8637 = n8599 & ~n8636 ;
  assign n8638 = n8637 ^ x302 ;
  assign n8639 = n8638 ^ n8596 ;
  assign n8640 = n8597 & ~n8639 ;
  assign n8641 = n8640 ^ x301 ;
  assign n8643 = n8642 ^ n8641 ;
  assign n8644 = n8642 ^ x300 ;
  assign n8645 = ~n8643 & n8644 ;
  assign n8646 = n8645 ^ x300 ;
  assign n8647 = n8646 ^ n8594 ;
  assign n8648 = ~n8595 & n8647 ;
  assign n8649 = n8648 ^ x299 ;
  assign n8650 = n8649 ^ n8592 ;
  assign n8651 = n8593 & ~n8650 ;
  assign n8652 = n8651 ^ x298 ;
  assign n8653 = n8652 ^ n8590 ;
  assign n8654 = n8591 & ~n8653 ;
  assign n8655 = n8654 ^ x297 ;
  assign n8656 = n8655 ^ n8588 ;
  assign n8657 = n8589 & ~n8656 ;
  assign n8658 = n8657 ^ x296 ;
  assign n8659 = n8658 ^ n8586 ;
  assign n8660 = n8587 & ~n8659 ;
  assign n8661 = n8660 ^ x295 ;
  assign n8662 = n8661 ^ n8584 ;
  assign n8663 = ~n8585 & n8662 ;
  assign n8664 = n8663 ^ x294 ;
  assign n8665 = n8664 ^ n8582 ;
  assign n8666 = n8583 & ~n8665 ;
  assign n8667 = n8666 ^ x293 ;
  assign n8669 = n8668 ^ n8667 ;
  assign n8670 = n8668 ^ x292 ;
  assign n8671 = n8669 & ~n8670 ;
  assign n8672 = n8671 ^ x292 ;
  assign n8674 = n8673 ^ n8672 ;
  assign n8675 = n8580 ^ x291 ;
  assign n8676 = n8675 ^ n8580 ;
  assign n8677 = n8676 ^ n8672 ;
  assign n8678 = n8674 & n8677 ;
  assign n8679 = n8678 ^ n8675 ;
  assign n8680 = ~n8581 & n8679 ;
  assign n8681 = n8680 ^ x290 ;
  assign n8682 = n8681 ^ x289 ;
  assign n8574 = n8555 ^ n5206 ;
  assign n8575 = n8560 & n8574 ;
  assign n8576 = n8575 ^ n8555 ;
  assign n8577 = n8576 ^ n5300 ;
  assign n8570 = n6744 ^ n6130 ;
  assign n8571 = ~n7473 & ~n8570 ;
  assign n8572 = n8571 ^ n6130 ;
  assign n8563 = n7930 ^ x262 ;
  assign n8564 = n8563 ^ n7810 ;
  assign n8566 = n8564 ^ n8546 ;
  assign n8565 = n8564 ^ n8554 ;
  assign n8567 = n8566 ^ n8565 ;
  assign n8568 = ~n8551 & ~n8567 ;
  assign n8569 = n8568 ^ n8566 ;
  assign n8573 = n8572 ^ n8569 ;
  assign n8578 = n8577 ^ n8573 ;
  assign n8562 = ~n8545 & n8561 ;
  assign n8579 = n8578 ^ n8562 ;
  assign n8734 = n8681 ^ n8579 ;
  assign n8735 = n8682 & ~n8734 ;
  assign n8730 = n8572 ^ n8564 ;
  assign n8731 = n8569 & n8730 ;
  assign n8727 = n6823 ^ n6139 ;
  assign n8728 = ~n7464 & n8727 ;
  assign n8723 = n8572 ^ n8071 ;
  assign n8722 = n7933 ^ n7809 ;
  assign n8724 = n8723 ^ n8722 ;
  assign n8725 = n8724 ^ n5300 ;
  assign n8721 = x289 ^ x288 ;
  assign n8726 = n8725 ^ n8721 ;
  assign n8729 = n8728 ^ n8726 ;
  assign n8732 = n8731 ^ n8729 ;
  assign n8720 = ~n8562 & n8578 ;
  assign n8733 = n8732 ^ n8720 ;
  assign n8736 = n8735 ^ n8733 ;
  assign n8717 = n8576 ^ n8573 ;
  assign n8718 = n8573 ^ n5300 ;
  assign n8719 = ~n8717 & n8718 ;
  assign n8737 = n8736 ^ n8719 ;
  assign n8741 = n8740 ^ n8737 ;
  assign n8684 = n8679 ^ x290 ;
  assign n8685 = n8684 ^ n6929 ;
  assign n8686 = n8685 ^ n7506 ;
  assign n8687 = n8686 ^ n8684 ;
  assign n8688 = n8095 & ~n8687 ;
  assign n8689 = n8688 ^ n8685 ;
  assign n8692 = n7386 ^ n6841 ;
  assign n8693 = n7332 & ~n8692 ;
  assign n8694 = n8693 ^ n6841 ;
  assign n8695 = n8667 ^ x292 ;
  assign n8696 = n8695 ^ n8668 ;
  assign n8697 = ~n8694 & ~n8696 ;
  assign n8690 = n8673 ^ x291 ;
  assign n8691 = n8690 ^ n8672 ;
  assign n8698 = n8697 ^ n8691 ;
  assign n8699 = n8697 ^ n6935 ;
  assign n8700 = n8699 ^ n7377 ;
  assign n8701 = n8700 ^ n8697 ;
  assign n8702 = ~n7325 & n8701 ;
  assign n8703 = n8702 ^ n8699 ;
  assign n8704 = ~n8698 & n8703 ;
  assign n8705 = n8704 ^ n8697 ;
  assign n8706 = n8705 ^ n8684 ;
  assign n8707 = n8689 & ~n8706 ;
  assign n8708 = n8707 ^ n8684 ;
  assign n8683 = n8682 ^ n8579 ;
  assign n8709 = n8708 ^ n8683 ;
  assign n8710 = n8683 ^ n6924 ;
  assign n8711 = n8710 ^ n7328 ;
  assign n8712 = n8711 ^ n8683 ;
  assign n8713 = n8104 & ~n8712 ;
  assign n8714 = n8713 ^ n8710 ;
  assign n8715 = ~n8709 & ~n8714 ;
  assign n8716 = n8715 ^ n8708 ;
  assign n8764 = n8737 ^ n8716 ;
  assign n8765 = ~n8741 & ~n8764 ;
  assign n8766 = n8765 ^ n8740 ;
  assign n8938 = n8769 ^ n8766 ;
  assign n8939 = n8771 & ~n8938 ;
  assign n8940 = n8939 ^ n8770 ;
  assign n8941 = n8940 ^ n8935 ;
  assign n8942 = ~n8937 & ~n8941 ;
  assign n8943 = n8942 ^ n8936 ;
  assign n8944 = n8943 ^ n8930 ;
  assign n8945 = ~n8932 & ~n8944 ;
  assign n8946 = n8945 ^ n8931 ;
  assign n8947 = n8946 ^ n8924 ;
  assign n8948 = n8927 & n8947 ;
  assign n8949 = n8948 ^ n8926 ;
  assign n8918 = n7368 ^ n6907 ;
  assign n8919 = ~n8332 & n8918 ;
  assign n8920 = n8919 ^ n6907 ;
  assign n8835 = n8222 ^ n8219 ;
  assign n8921 = n8920 ^ n8835 ;
  assign n9081 = n8949 ^ n8921 ;
  assign n9101 = n9081 ^ n5713 ;
  assign n9082 = n8946 ^ n8927 ;
  assign n9083 = n9082 ^ n6181 ;
  assign n9085 = n8940 ^ n8937 ;
  assign n9086 = n9085 ^ n5718 ;
  assign n8772 = n8771 ^ n8766 ;
  assign n8773 = n8772 ^ n5727 ;
  assign n8742 = n8741 ^ n8716 ;
  assign n8743 = n8742 ^ n5732 ;
  assign n8745 = n8696 ^ n8694 ;
  assign n8746 = ~n5753 & n8745 ;
  assign n8747 = n8746 ^ n5750 ;
  assign n8748 = n8703 ^ n8691 ;
  assign n8749 = n8748 ^ n8746 ;
  assign n8750 = n8747 & n8749 ;
  assign n8751 = n8750 ^ n5750 ;
  assign n8752 = n8751 ^ n5239 ;
  assign n8753 = n8705 ^ n8689 ;
  assign n8754 = n8753 ^ n8751 ;
  assign n8755 = ~n8752 & ~n8754 ;
  assign n8756 = n8755 ^ n5239 ;
  assign n8744 = n8714 ^ n8708 ;
  assign n8757 = n8756 ^ n8744 ;
  assign n8758 = n8744 ^ n5738 ;
  assign n8759 = n8757 & ~n8758 ;
  assign n8760 = n8759 ^ n8756 ;
  assign n8761 = n8760 ^ n8742 ;
  assign n8762 = n8743 & n8761 ;
  assign n8763 = n8762 ^ n5732 ;
  assign n9087 = n8772 ^ n8763 ;
  assign n9088 = n8773 & ~n9087 ;
  assign n9089 = n9088 ^ n5727 ;
  assign n9090 = n9089 ^ n9085 ;
  assign n9091 = ~n9086 & n9090 ;
  assign n9092 = n9091 ^ n5718 ;
  assign n9084 = n8943 ^ n8932 ;
  assign n9093 = n9092 ^ n9084 ;
  assign n9094 = n9092 ^ n6173 ;
  assign n9095 = ~n9093 & n9094 ;
  assign n9096 = n9095 ^ n6173 ;
  assign n9097 = n9096 ^ n9082 ;
  assign n9098 = n9083 & ~n9097 ;
  assign n9099 = n9098 ^ n6181 ;
  assign n9198 = n9101 ^ n9099 ;
  assign n9190 = n9089 ^ n9086 ;
  assign n8774 = n8773 ^ n8763 ;
  assign n8775 = n8760 ^ n8743 ;
  assign n8776 = n8745 ^ n5753 ;
  assign n8777 = n8748 ^ n8747 ;
  assign n8778 = ~n8776 & ~n8777 ;
  assign n8779 = n8753 ^ n8752 ;
  assign n8780 = n8778 & ~n8779 ;
  assign n8781 = n8758 ^ n8756 ;
  assign n8782 = ~n8780 & n8781 ;
  assign n8783 = n8775 & n8782 ;
  assign n9191 = n8774 & ~n8783 ;
  assign n9192 = ~n9190 & n9191 ;
  assign n9193 = n9084 ^ n6173 ;
  assign n9194 = n9193 ^ n9092 ;
  assign n9195 = ~n9192 & ~n9194 ;
  assign n9196 = n9096 ^ n9083 ;
  assign n9197 = n9195 & ~n9196 ;
  assign n9258 = n9198 ^ n9197 ;
  assign n9259 = n9258 ^ x342 ;
  assign n9260 = n9196 ^ n9195 ;
  assign n9261 = n9260 ^ x343 ;
  assign n9262 = n9194 ^ n9192 ;
  assign n9263 = n9262 ^ x344 ;
  assign n9267 = n9191 ^ n9190 ;
  assign n8785 = n8782 ^ n8775 ;
  assign n8786 = n8785 ^ x347 ;
  assign n8787 = x351 & n8776 ;
  assign n8788 = n8787 ^ x350 ;
  assign n8789 = n8777 ^ n8776 ;
  assign n8790 = n8789 ^ n8787 ;
  assign n8791 = n8788 & ~n8790 ;
  assign n8792 = n8791 ^ x350 ;
  assign n8793 = n8792 ^ x349 ;
  assign n8794 = n8779 ^ n8778 ;
  assign n8795 = n8794 ^ n8792 ;
  assign n8796 = n8793 & n8795 ;
  assign n8797 = n8796 ^ x349 ;
  assign n8798 = n8797 ^ x348 ;
  assign n8799 = n8781 ^ n8780 ;
  assign n8800 = n8799 ^ n8797 ;
  assign n8801 = n8798 & ~n8800 ;
  assign n8802 = n8801 ^ x348 ;
  assign n8803 = n8802 ^ n8785 ;
  assign n8804 = ~n8786 & n8803 ;
  assign n8805 = n8804 ^ x347 ;
  assign n8806 = n8805 ^ x346 ;
  assign n8784 = n8783 ^ n8774 ;
  assign n9264 = n8805 ^ n8784 ;
  assign n9265 = n8806 & n9264 ;
  assign n9266 = n9265 ^ x346 ;
  assign n9268 = n9267 ^ n9266 ;
  assign n9269 = n9267 ^ x345 ;
  assign n9270 = n9268 & ~n9269 ;
  assign n9271 = n9270 ^ x345 ;
  assign n9272 = n9271 ^ n9262 ;
  assign n9273 = ~n9263 & n9272 ;
  assign n9274 = n9273 ^ x344 ;
  assign n9275 = n9274 ^ n9260 ;
  assign n9276 = n9261 & ~n9275 ;
  assign n9277 = n9276 ^ x343 ;
  assign n9278 = n9277 ^ n9258 ;
  assign n9279 = ~n9259 & n9278 ;
  assign n9280 = n9279 ^ x342 ;
  assign n9100 = n9099 ^ n9081 ;
  assign n9102 = ~n9100 & ~n9101 ;
  assign n9103 = n9102 ^ n9099 ;
  assign n8950 = n8949 ^ n8920 ;
  assign n8951 = n8921 & ~n8950 ;
  assign n8952 = n8951 ^ n8835 ;
  assign n8914 = n7559 ^ n6905 ;
  assign n8915 = n8294 & n8914 ;
  assign n8916 = n8915 ^ n6905 ;
  assign n8828 = n8224 ^ x314 ;
  assign n8829 = n8828 ^ n8202 ;
  assign n8917 = n8916 ^ n8829 ;
  assign n9079 = n8952 ^ n8917 ;
  assign n9080 = n9079 ^ n6197 ;
  assign n9200 = n9103 ^ n9080 ;
  assign n9199 = ~n9197 & n9198 ;
  assign n9256 = n9200 ^ n9199 ;
  assign n9257 = n9256 ^ x341 ;
  assign n9649 = n9280 ^ n9257 ;
  assign n8980 = n8617 ^ n8607 ;
  assign n10279 = n8980 ^ n8286 ;
  assign n10280 = n9649 & n10279 ;
  assign n10281 = n10280 ^ n8286 ;
  assign n9041 = n7464 ^ n6705 ;
  assign n9042 = n8021 & ~n9041 ;
  assign n9043 = n9042 ^ n6705 ;
  assign n8839 = n8649 ^ x298 ;
  assign n8840 = n8839 ^ n8592 ;
  assign n8841 = n8840 ^ n6714 ;
  assign n8842 = n8841 ^ n7315 ;
  assign n8843 = n8842 ^ n8840 ;
  assign n8844 = ~n8722 & ~n8843 ;
  assign n8845 = n8844 ^ n8841 ;
  assign n8854 = n8646 ^ n8595 ;
  assign n8851 = n7286 ^ n6715 ;
  assign n8852 = n8564 & ~n8851 ;
  assign n8853 = n8852 ^ n6715 ;
  assign n8855 = n8854 ^ n8853 ;
  assign n8856 = n8641 ^ x300 ;
  assign n8857 = n8856 ^ n8642 ;
  assign n8859 = n8857 ^ n7453 ;
  assign n8858 = n8857 ^ n8066 ;
  assign n8860 = n8859 ^ n8858 ;
  assign n8861 = ~n8546 & ~n8860 ;
  assign n8862 = n8861 ^ n8859 ;
  assign n9015 = n8857 ^ n8853 ;
  assign n8866 = n8638 ^ n8597 ;
  assign n8863 = n8034 ^ n7421 ;
  assign n8864 = ~n8497 & ~n8863 ;
  assign n8865 = n8864 ^ n7421 ;
  assign n8867 = n8866 ^ n8865 ;
  assign n8871 = n8635 ^ x302 ;
  assign n8872 = n8871 ^ n8598 ;
  assign n8868 = n8011 ^ n7336 ;
  assign n8869 = ~n8481 & ~n8868 ;
  assign n8870 = n8869 ^ n7336 ;
  assign n8873 = n8872 ^ n8870 ;
  assign n8877 = n8633 ^ x303 ;
  assign n8874 = n7988 ^ n7306 ;
  assign n8875 = ~n8467 & ~n8874 ;
  assign n8876 = n8875 ^ n7306 ;
  assign n8878 = n8877 ^ n8876 ;
  assign n8882 = n8626 ^ x304 ;
  assign n8883 = n8882 ^ n8627 ;
  assign n8879 = n7947 ^ n7182 ;
  assign n8880 = n8377 & n8879 ;
  assign n8881 = n8880 ^ n7182 ;
  assign n8884 = n8883 ^ n8881 ;
  assign n8888 = n8623 ^ n8603 ;
  assign n8885 = n7746 ^ n7121 ;
  assign n8886 = n8245 & n8885 ;
  assign n8887 = n8886 ^ n7121 ;
  assign n8889 = n8888 ^ n8887 ;
  assign n8989 = n8620 ^ x306 ;
  assign n8990 = n8989 ^ n8604 ;
  assign n8893 = n8615 ^ x308 ;
  assign n8890 = n7599 ^ n6873 ;
  assign n8891 = ~n8267 & ~n8890 ;
  assign n8892 = n8891 ^ n6873 ;
  assign n8894 = n8893 ^ n8892 ;
  assign n8197 = n8196 ^ x309 ;
  assign n8244 = n8243 ^ n8197 ;
  assign n8976 = n8892 ^ n8244 ;
  assign n8895 = n7345 ^ n6879 ;
  assign n8896 = ~n8273 & ~n8895 ;
  assign n8897 = n8896 ^ n6879 ;
  assign n8898 = n8897 ^ n8244 ;
  assign n8814 = n8240 ^ x310 ;
  assign n8815 = n8814 ^ n8198 ;
  assign n8899 = n8815 ^ n6887 ;
  assign n8900 = n8899 ^ n7357 ;
  assign n8901 = n8900 ^ n8815 ;
  assign n8902 = n8278 & n8901 ;
  assign n8903 = n8902 ^ n8899 ;
  assign n8971 = n8897 ^ n8815 ;
  assign n8962 = n8237 ^ n8236 ;
  assign n8904 = n7363 ^ n6898 ;
  assign n8905 = ~n8286 & n8904 ;
  assign n8906 = n8905 ^ n6898 ;
  assign n8821 = n8232 ^ x312 ;
  assign n8822 = n8821 ^ n8200 ;
  assign n8907 = n8906 ^ n8822 ;
  assign n8908 = n8230 ^ n8227 ;
  assign n8909 = n8908 ^ n6900 ;
  assign n8910 = n8909 ^ n7569 ;
  assign n8911 = n8910 ^ n8908 ;
  assign n8912 = n8291 & n8911 ;
  assign n8913 = n8912 ^ n8909 ;
  assign n8953 = n8952 ^ n8916 ;
  assign n8954 = ~n8917 & n8953 ;
  assign n8955 = n8954 ^ n8829 ;
  assign n8956 = n8955 ^ n8908 ;
  assign n8957 = ~n8913 & n8956 ;
  assign n8958 = n8957 ^ n8908 ;
  assign n8959 = n8958 ^ n8906 ;
  assign n8960 = n8907 & n8959 ;
  assign n8961 = n8960 ^ n8822 ;
  assign n8963 = n8962 ^ n8961 ;
  assign n8964 = n7351 ^ n6890 ;
  assign n8965 = ~n8355 & n8964 ;
  assign n8966 = n8965 ^ n7351 ;
  assign n8967 = n8966 ^ n8961 ;
  assign n8968 = n8963 & ~n8967 ;
  assign n8969 = n8968 ^ n8962 ;
  assign n8970 = n8969 ^ n8897 ;
  assign n8972 = n8971 ^ n8970 ;
  assign n8973 = n8903 & n8972 ;
  assign n8974 = n8973 ^ n8971 ;
  assign n8975 = n8898 & n8974 ;
  assign n8977 = n8976 ^ n8975 ;
  assign n8978 = ~n8894 & n8977 ;
  assign n8979 = n8978 ^ n8893 ;
  assign n8981 = n8980 ^ n8979 ;
  assign n8982 = n8980 ^ n6868 ;
  assign n8983 = n8982 ^ n7338 ;
  assign n8984 = n8983 ^ n8980 ;
  assign n8985 = ~n8262 & n8984 ;
  assign n8986 = n8985 ^ n8982 ;
  assign n8987 = n8981 & ~n8986 ;
  assign n8988 = n8987 ^ n8980 ;
  assign n8991 = n8990 ^ n8988 ;
  assign n8992 = n8990 ^ n6861 ;
  assign n8993 = n8992 ^ n7731 ;
  assign n8994 = n8993 ^ n8990 ;
  assign n8995 = n8256 & n8994 ;
  assign n8996 = n8995 ^ n8992 ;
  assign n8997 = ~n8991 & n8996 ;
  assign n8998 = n8997 ^ n8990 ;
  assign n8999 = n8998 ^ n8887 ;
  assign n9000 = ~n8889 & ~n8999 ;
  assign n9001 = n9000 ^ n8888 ;
  assign n9002 = n9001 ^ n8881 ;
  assign n9003 = n8884 & ~n9002 ;
  assign n9004 = n9003 ^ n8883 ;
  assign n9005 = n9004 ^ n8876 ;
  assign n9006 = n8878 & ~n9005 ;
  assign n9007 = n9006 ^ n8877 ;
  assign n9008 = n9007 ^ n8870 ;
  assign n9009 = n8873 & n9008 ;
  assign n9010 = n9009 ^ n8872 ;
  assign n9011 = n9010 ^ n8865 ;
  assign n9012 = n8867 & ~n9011 ;
  assign n9013 = n9012 ^ n8866 ;
  assign n9014 = n9013 ^ n8853 ;
  assign n9016 = n9015 ^ n9014 ;
  assign n9017 = n8862 & n9016 ;
  assign n9018 = n9017 ^ n9015 ;
  assign n9019 = ~n8855 & ~n9018 ;
  assign n9020 = n9019 ^ n8854 ;
  assign n8846 = n7475 ^ n6729 ;
  assign n8847 = ~n7955 & ~n8846 ;
  assign n8848 = n8847 ^ n6729 ;
  assign n8849 = n8848 ^ n8840 ;
  assign n8850 = n8849 ^ n8848 ;
  assign n9021 = n9020 ^ n8850 ;
  assign n9022 = n8845 & ~n9021 ;
  assign n9023 = n9022 ^ n8849 ;
  assign n9025 = n7473 ^ n6711 ;
  assign n9026 = n7992 & ~n9025 ;
  assign n9027 = n9026 ^ n6711 ;
  assign n9029 = n9027 ^ n8848 ;
  assign n9024 = n8652 ^ n8591 ;
  assign n9028 = n9027 ^ n9024 ;
  assign n9030 = n9029 ^ n9028 ;
  assign n9031 = n9023 & n9030 ;
  assign n9032 = n9031 ^ n9029 ;
  assign n9035 = n8658 ^ n8587 ;
  assign n9037 = n9035 ^ n9027 ;
  assign n9033 = n8655 ^ x296 ;
  assign n9034 = n9033 ^ n8588 ;
  assign n9036 = n9035 ^ n9034 ;
  assign n9038 = n9037 ^ n9036 ;
  assign n9039 = n9032 & n9038 ;
  assign n9040 = n9039 ^ n9037 ;
  assign n9176 = n9043 ^ n9040 ;
  assign n9058 = n9018 ^ n8854 ;
  assign n9059 = n9058 ^ n6106 ;
  assign n9154 = n9013 ^ n8862 ;
  assign n9060 = n9010 ^ n8867 ;
  assign n9061 = n9060 ^ n6664 ;
  assign n9146 = n9007 ^ n8873 ;
  assign n9062 = n9004 ^ n8878 ;
  assign n9063 = n9062 ^ n6431 ;
  assign n9064 = n9001 ^ n8884 ;
  assign n9065 = n9064 ^ n6278 ;
  assign n9066 = n8996 ^ n8988 ;
  assign n9067 = n9066 ^ n6270 ;
  assign n9069 = n8977 ^ n8893 ;
  assign n9070 = n9069 ^ n6239 ;
  assign n9120 = n8974 ^ n8244 ;
  assign n9071 = n8969 ^ n8903 ;
  assign n9072 = n9071 ^ n6224 ;
  assign n9075 = n8958 ^ n8907 ;
  assign n9076 = n9075 ^ n6203 ;
  assign n9077 = n8955 ^ n8913 ;
  assign n9078 = n9077 ^ n6195 ;
  assign n9104 = n9103 ^ n9079 ;
  assign n9105 = n9080 & ~n9104 ;
  assign n9106 = n9105 ^ n6197 ;
  assign n9107 = n9106 ^ n9077 ;
  assign n9108 = ~n9078 & ~n9107 ;
  assign n9109 = n9108 ^ n6195 ;
  assign n9110 = n9109 ^ n9075 ;
  assign n9111 = n9076 & ~n9110 ;
  assign n9112 = n9111 ^ n6203 ;
  assign n9073 = n8966 ^ n8962 ;
  assign n9074 = n9073 ^ n8961 ;
  assign n9113 = n9112 ^ n9074 ;
  assign n9114 = n9112 ^ n6215 ;
  assign n9115 = n9113 & ~n9114 ;
  assign n9116 = n9115 ^ n6215 ;
  assign n9117 = n9116 ^ n9071 ;
  assign n9118 = ~n9072 & ~n9117 ;
  assign n9119 = n9118 ^ n6224 ;
  assign n9121 = n9120 ^ n9119 ;
  assign n9122 = n9120 ^ n6230 ;
  assign n9123 = n9121 & ~n9122 ;
  assign n9124 = n9123 ^ n6230 ;
  assign n9125 = n9124 ^ n9069 ;
  assign n9126 = n9070 & n9125 ;
  assign n9127 = n9126 ^ n6239 ;
  assign n9068 = n8986 ^ n8979 ;
  assign n9128 = n9127 ^ n9068 ;
  assign n9129 = n9127 ^ n6249 ;
  assign n9130 = ~n9128 & n9129 ;
  assign n9131 = n9130 ^ n6249 ;
  assign n9132 = n9131 ^ n9066 ;
  assign n9133 = ~n9067 & n9132 ;
  assign n9134 = n9133 ^ n6270 ;
  assign n9135 = n9134 ^ n5685 ;
  assign n9136 = n8998 ^ n8889 ;
  assign n9137 = n9136 ^ n9134 ;
  assign n9138 = n9135 & n9137 ;
  assign n9139 = n9138 ^ n5685 ;
  assign n9140 = n9139 ^ n9064 ;
  assign n9141 = ~n9065 & n9140 ;
  assign n9142 = n9141 ^ n6278 ;
  assign n9143 = n9142 ^ n9062 ;
  assign n9144 = ~n9063 & n9143 ;
  assign n9145 = n9144 ^ n6431 ;
  assign n9147 = n9146 ^ n9145 ;
  assign n9148 = n9146 ^ n6646 ;
  assign n9149 = n9147 & n9148 ;
  assign n9150 = n9149 ^ n6646 ;
  assign n9151 = n9150 ^ n9060 ;
  assign n9152 = n9061 & n9151 ;
  assign n9153 = n9152 ^ n6664 ;
  assign n9155 = n9154 ^ n9153 ;
  assign n9156 = n9154 ^ n6686 ;
  assign n9157 = ~n9155 & n9156 ;
  assign n9158 = n9157 ^ n6686 ;
  assign n9159 = n9158 ^ n9058 ;
  assign n9160 = n9059 & n9159 ;
  assign n9161 = n9160 ^ n6106 ;
  assign n9162 = n9161 ^ n6101 ;
  assign n9163 = n9020 ^ n8845 ;
  assign n9164 = n9163 ^ n9161 ;
  assign n9165 = ~n9162 & ~n9164 ;
  assign n9166 = n9165 ^ n6101 ;
  assign n9057 = n9024 ^ n9023 ;
  assign n9167 = n9166 ^ n9057 ;
  assign n9168 = n9166 ^ n6100 ;
  assign n9169 = ~n9167 & n9168 ;
  assign n9170 = n9169 ^ n6100 ;
  assign n9056 = n9034 ^ n9032 ;
  assign n9171 = n9170 ^ n9056 ;
  assign n9172 = n9170 ^ n6098 ;
  assign n9173 = ~n9171 & n9172 ;
  assign n9174 = n9173 ^ n6098 ;
  assign n9175 = n9174 ^ n6092 ;
  assign n9352 = n9176 ^ n9175 ;
  assign n9182 = n9168 ^ n9057 ;
  assign n9183 = n9142 ^ n9063 ;
  assign n9184 = n9136 ^ n9135 ;
  assign n9185 = n9068 ^ n6249 ;
  assign n9186 = n9185 ^ n9127 ;
  assign n9187 = n9116 ^ n9072 ;
  assign n9188 = n9074 ^ n6215 ;
  assign n9189 = n9188 ^ n9112 ;
  assign n9201 = n9199 & n9200 ;
  assign n9202 = n9106 ^ n9078 ;
  assign n9203 = ~n9201 & n9202 ;
  assign n9204 = n9109 ^ n9076 ;
  assign n9205 = n9203 & n9204 ;
  assign n9206 = n9189 & n9205 ;
  assign n9207 = n9187 & n9206 ;
  assign n9208 = n9122 ^ n9119 ;
  assign n9209 = ~n9207 & n9208 ;
  assign n9210 = n9124 ^ n9070 ;
  assign n9211 = n9209 & ~n9210 ;
  assign n9212 = ~n9186 & ~n9211 ;
  assign n9213 = n9131 ^ n9067 ;
  assign n9214 = ~n9212 & ~n9213 ;
  assign n9215 = ~n9184 & n9214 ;
  assign n9216 = n9139 ^ n9065 ;
  assign n9217 = n9215 & ~n9216 ;
  assign n9218 = ~n9183 & n9217 ;
  assign n9219 = n9148 ^ n9145 ;
  assign n9220 = n9218 & n9219 ;
  assign n9221 = n9150 ^ n9061 ;
  assign n9222 = ~n9220 & n9221 ;
  assign n9223 = n9156 ^ n9153 ;
  assign n9224 = ~n9222 & n9223 ;
  assign n9225 = n9158 ^ n9059 ;
  assign n9226 = ~n9224 & ~n9225 ;
  assign n9227 = n9163 ^ n9162 ;
  assign n9228 = ~n9226 & n9227 ;
  assign n9229 = ~n9182 & ~n9228 ;
  assign n9230 = n9172 ^ n9056 ;
  assign n9351 = n9229 & ~n9230 ;
  assign n9353 = n9352 ^ n9351 ;
  assign n9231 = n9230 ^ n9229 ;
  assign n9232 = n9231 ^ x323 ;
  assign n9233 = n9228 ^ n9182 ;
  assign n9234 = n9233 ^ x324 ;
  assign n9339 = n9227 ^ n9226 ;
  assign n9235 = n9225 ^ n9224 ;
  assign n9236 = n9235 ^ x326 ;
  assign n9237 = n9223 ^ n9222 ;
  assign n9238 = n9237 ^ x327 ;
  assign n9239 = n9221 ^ n9220 ;
  assign n9240 = n9239 ^ x328 ;
  assign n9241 = n9219 ^ n9218 ;
  assign n9242 = n9241 ^ x329 ;
  assign n9318 = n9216 ^ n9215 ;
  assign n9313 = n9214 ^ n9184 ;
  assign n9245 = n9211 ^ n9186 ;
  assign n9246 = n9245 ^ x334 ;
  assign n9247 = n9210 ^ n9209 ;
  assign n9248 = n9247 ^ x335 ;
  assign n9297 = n9208 ^ n9207 ;
  assign n9250 = n9205 ^ n9189 ;
  assign n9251 = n9250 ^ x338 ;
  assign n9252 = n9204 ^ n9203 ;
  assign n9253 = n9252 ^ x339 ;
  assign n9254 = n9202 ^ n9201 ;
  assign n9255 = n9254 ^ x340 ;
  assign n9281 = n9280 ^ n9256 ;
  assign n9282 = n9257 & ~n9281 ;
  assign n9283 = n9282 ^ x341 ;
  assign n9284 = n9283 ^ n9254 ;
  assign n9285 = n9255 & ~n9284 ;
  assign n9286 = n9285 ^ x340 ;
  assign n9287 = n9286 ^ n9252 ;
  assign n9288 = ~n9253 & n9287 ;
  assign n9289 = n9288 ^ x339 ;
  assign n9290 = n9289 ^ n9250 ;
  assign n9291 = ~n9251 & n9290 ;
  assign n9292 = n9291 ^ x338 ;
  assign n9249 = n9206 ^ n9187 ;
  assign n9293 = n9292 ^ n9249 ;
  assign n9294 = n9292 ^ x337 ;
  assign n9295 = n9293 & n9294 ;
  assign n9296 = n9295 ^ x337 ;
  assign n9298 = n9297 ^ n9296 ;
  assign n9299 = n9247 ^ x336 ;
  assign n9300 = n9299 ^ n9247 ;
  assign n9301 = n9300 ^ n9296 ;
  assign n9302 = n9298 & n9301 ;
  assign n9303 = n9302 ^ n9299 ;
  assign n9304 = ~n9248 & n9303 ;
  assign n9305 = n9304 ^ x335 ;
  assign n9306 = n9305 ^ n9245 ;
  assign n9307 = ~n9246 & n9306 ;
  assign n9308 = n9307 ^ x334 ;
  assign n9244 = n9213 ^ n9212 ;
  assign n9309 = n9308 ^ n9244 ;
  assign n9310 = n9308 ^ x333 ;
  assign n9311 = ~n9309 & n9310 ;
  assign n9312 = n9311 ^ x333 ;
  assign n9314 = n9313 ^ n9312 ;
  assign n9315 = n9313 ^ x332 ;
  assign n9316 = n9314 & ~n9315 ;
  assign n9317 = n9316 ^ x332 ;
  assign n9319 = n9318 ^ n9317 ;
  assign n9320 = n9318 ^ x331 ;
  assign n9321 = n9319 & ~n9320 ;
  assign n9322 = n9321 ^ x331 ;
  assign n9243 = n9217 ^ n9183 ;
  assign n9323 = n9322 ^ n9243 ;
  assign n9324 = n9322 ^ x330 ;
  assign n9325 = n9323 & n9324 ;
  assign n9326 = n9325 ^ x330 ;
  assign n9327 = n9326 ^ n9241 ;
  assign n9328 = n9242 & ~n9327 ;
  assign n9329 = n9328 ^ x329 ;
  assign n9330 = n9329 ^ n9239 ;
  assign n9331 = n9240 & ~n9330 ;
  assign n9332 = n9331 ^ x328 ;
  assign n9333 = n9332 ^ n9237 ;
  assign n9334 = ~n9238 & n9333 ;
  assign n9335 = n9334 ^ x327 ;
  assign n9336 = n9335 ^ n9235 ;
  assign n9337 = ~n9236 & n9336 ;
  assign n9338 = n9337 ^ x326 ;
  assign n9340 = n9339 ^ n9338 ;
  assign n9341 = n9339 ^ x325 ;
  assign n9342 = n9340 & ~n9341 ;
  assign n9343 = n9342 ^ x325 ;
  assign n9344 = n9343 ^ n9233 ;
  assign n9345 = ~n9234 & n9344 ;
  assign n9346 = n9345 ^ x324 ;
  assign n9347 = n9346 ^ n9231 ;
  assign n9348 = n9232 & ~n9347 ;
  assign n9349 = n9348 ^ x323 ;
  assign n9350 = n9349 ^ x322 ;
  assign n9386 = n9353 ^ n9350 ;
  assign n9381 = n8185 ^ n7328 ;
  assign n9382 = ~n8926 & ~n9381 ;
  assign n9383 = n9382 ^ n7328 ;
  assign n9409 = n9386 ^ n9383 ;
  assign n9387 = n9386 ^ n7506 ;
  assign n9388 = n9387 ^ n8156 ;
  assign n9389 = n9388 ^ n9386 ;
  assign n9390 = n8931 & n9389 ;
  assign n9391 = n9390 ^ n9387 ;
  assign n9398 = n9346 ^ n9232 ;
  assign n9392 = n9343 ^ x324 ;
  assign n9393 = n9392 ^ n9233 ;
  assign n9394 = n8095 ^ n7386 ;
  assign n9395 = n8770 & n9394 ;
  assign n9396 = n9395 ^ n7386 ;
  assign n9397 = ~n9393 & n9396 ;
  assign n9399 = n9398 ^ n9397 ;
  assign n9400 = n9397 ^ n7377 ;
  assign n9401 = n9400 ^ n8104 ;
  assign n9402 = n9401 ^ n9397 ;
  assign n9403 = ~n8936 & n9402 ;
  assign n9404 = n9403 ^ n9400 ;
  assign n9405 = n9399 & ~n9404 ;
  assign n9406 = n9405 ^ n9398 ;
  assign n9407 = n9406 ^ n9386 ;
  assign n9408 = ~n9391 & ~n9407 ;
  assign n9410 = n9409 ^ n9408 ;
  assign n9360 = ~n9351 & n9352 ;
  assign n9177 = n9176 ^ n9174 ;
  assign n9178 = n9175 & ~n9177 ;
  assign n9179 = n9178 ^ n6092 ;
  assign n9358 = n9179 ^ n6130 ;
  assign n9051 = n7401 ^ n6744 ;
  assign n9052 = ~n8055 & n9051 ;
  assign n9053 = n9052 ^ n6744 ;
  assign n9044 = n8661 ^ x294 ;
  assign n9045 = n9044 ^ n8584 ;
  assign n9047 = n9045 ^ n9035 ;
  assign n9046 = n9045 ^ n9043 ;
  assign n9048 = n9047 ^ n9046 ;
  assign n9049 = n9040 & n9048 ;
  assign n9050 = n9049 ^ n9047 ;
  assign n9054 = n9053 ^ n9050 ;
  assign n9359 = n9358 ^ n9054 ;
  assign n9361 = n9360 ^ n9359 ;
  assign n9354 = n9353 ^ n9349 ;
  assign n9355 = n9350 & n9354 ;
  assign n9356 = n9355 ^ x322 ;
  assign n9357 = n9356 ^ x321 ;
  assign n9384 = n9361 ^ n9357 ;
  assign n9476 = n9410 ^ n9384 ;
  assign n9464 = n9396 ^ n9393 ;
  assign n9465 = ~n6841 & ~n9464 ;
  assign n9466 = n9465 ^ n6935 ;
  assign n9467 = n9404 ^ n9398 ;
  assign n9468 = n9467 ^ n9465 ;
  assign n9469 = n9466 & ~n9468 ;
  assign n9470 = n9469 ^ n6935 ;
  assign n9471 = n9470 ^ n6929 ;
  assign n9472 = n9406 ^ n9391 ;
  assign n9473 = n9472 ^ n9470 ;
  assign n9474 = ~n9471 & n9473 ;
  assign n9475 = n9474 ^ n6929 ;
  assign n9477 = n9476 ^ n9475 ;
  assign n9478 = n9476 ^ n6924 ;
  assign n9479 = ~n9477 & ~n9478 ;
  assign n9480 = n9479 ^ n6924 ;
  assign n9385 = n9384 ^ n9383 ;
  assign n9411 = n9385 & ~n9410 ;
  assign n9412 = n9411 ^ n9384 ;
  assign n9374 = n9053 ^ n9045 ;
  assign n9375 = n9050 & n9374 ;
  assign n9371 = n7334 ^ n6823 ;
  assign n9372 = ~n8079 & n9371 ;
  assign n9367 = n9053 ^ n8727 ;
  assign n9366 = n8664 ^ n8583 ;
  assign n9368 = n9367 ^ n9366 ;
  assign n9369 = n9368 ^ n6130 ;
  assign n9365 = x321 ^ x320 ;
  assign n9370 = n9369 ^ n9365 ;
  assign n9373 = n9372 ^ n9370 ;
  assign n9376 = n9375 ^ n9373 ;
  assign n9364 = ~n9359 & ~n9360 ;
  assign n9377 = n9376 ^ n9364 ;
  assign n9362 = n9361 ^ n9356 ;
  assign n9363 = n9357 & n9362 ;
  assign n9378 = n9377 ^ n9363 ;
  assign n9055 = n9054 ^ n6130 ;
  assign n9180 = n9179 ^ n9054 ;
  assign n9181 = n9055 & ~n9180 ;
  assign n9379 = n9378 ^ n9181 ;
  assign n8836 = n8308 ^ n6852 ;
  assign n8837 = n8835 & n8836 ;
  assign n8838 = n8837 ^ n8308 ;
  assign n9380 = n9379 ^ n8838 ;
  assign n9462 = n9412 ^ n9380 ;
  assign n9463 = n9462 ^ n6919 ;
  assign n9516 = n9480 ^ n9463 ;
  assign n9509 = n9467 ^ n9466 ;
  assign n9510 = n9464 ^ n6841 ;
  assign n9511 = n9509 & n9510 ;
  assign n9512 = n9472 ^ n9471 ;
  assign n9513 = n9511 & n9512 ;
  assign n9514 = n9478 ^ n9475 ;
  assign n9515 = ~n9513 & ~n9514 ;
  assign n9575 = n9516 ^ n9515 ;
  assign n9559 = n9514 ^ n9513 ;
  assign n9560 = n9559 ^ x380 ;
  assign n9563 = x383 & ~n9510 ;
  assign n9562 = n9510 ^ n9509 ;
  assign n9564 = n9563 ^ n9562 ;
  assign n9565 = n9563 ^ x382 ;
  assign n9566 = ~n9564 & n9565 ;
  assign n9567 = n9566 ^ x382 ;
  assign n9561 = n9512 ^ n9511 ;
  assign n9568 = n9567 ^ n9561 ;
  assign n9569 = n9567 ^ x381 ;
  assign n9570 = ~n9568 & n9569 ;
  assign n9571 = n9570 ^ x381 ;
  assign n9572 = n9571 ^ n9559 ;
  assign n9573 = ~n9560 & n9572 ;
  assign n9574 = n9573 ^ x380 ;
  assign n9576 = n9575 ^ n9574 ;
  assign n9577 = n9575 ^ x379 ;
  assign n9578 = n9576 & ~n9577 ;
  assign n9579 = n9578 ^ x379 ;
  assign n10206 = n9579 ^ x378 ;
  assign n9413 = n9412 ^ n8838 ;
  assign n9414 = n9380 & n9413 ;
  assign n9415 = n9414 ^ n9379 ;
  assign n8833 = n8776 ^ x351 ;
  assign n8830 = n8306 ^ n6851 ;
  assign n8831 = n8829 & n8830 ;
  assign n8832 = n8831 ^ n8306 ;
  assign n8834 = n8833 ^ n8832 ;
  assign n9484 = n9415 ^ n8834 ;
  assign n9486 = n9484 ^ n6967 ;
  assign n9481 = n9480 ^ n9462 ;
  assign n9482 = ~n9463 & n9481 ;
  assign n9483 = n9482 ^ n6919 ;
  assign n9518 = n9486 ^ n9483 ;
  assign n9517 = n9515 & n9516 ;
  assign n9557 = n9518 ^ n9517 ;
  assign n10207 = n10206 ^ n9557 ;
  assign n10282 = n10281 ^ n10207 ;
  assign n9678 = n9283 ^ x340 ;
  assign n9679 = n9678 ^ n9254 ;
  assign n10275 = n8990 ^ n8355 ;
  assign n10276 = n9679 & n10275 ;
  assign n10277 = n10276 ^ n8355 ;
  assign n10305 = n10277 ^ n10207 ;
  assign n9660 = n9274 ^ x343 ;
  assign n9661 = n9660 ^ n9260 ;
  assign n10283 = n9571 ^ x380 ;
  assign n10284 = n10283 ^ n9559 ;
  assign n10285 = n10284 ^ n8294 ;
  assign n10286 = n10285 ^ n8244 ;
  assign n10287 = n10286 ^ n10284 ;
  assign n10288 = n9661 & ~n10287 ;
  assign n10289 = n10288 ^ n10285 ;
  assign n8820 = n8799 ^ n8798 ;
  assign n9991 = n7401 ^ n7332 ;
  assign n9992 = n8683 & ~n9991 ;
  assign n9993 = n9992 ^ n7401 ;
  assign n9609 = n9326 ^ n9242 ;
  assign n9606 = n8021 ^ n7475 ;
  assign n9607 = ~n8696 & ~n9606 ;
  assign n9608 = n9607 ^ n7475 ;
  assign n9610 = n9609 ^ n9608 ;
  assign n9731 = n7992 ^ n7315 ;
  assign n9732 = n9366 & ~n9731 ;
  assign n9733 = n9732 ^ n7315 ;
  assign n9742 = n9733 ^ n9608 ;
  assign n9611 = n9312 ^ x332 ;
  assign n9612 = n9611 ^ n9313 ;
  assign n9613 = n9612 ^ n8066 ;
  assign n9614 = n9613 ^ n8722 ;
  assign n9615 = n9614 ^ n9612 ;
  assign n9616 = n9035 & n9615 ;
  assign n9617 = n9616 ^ n9613 ;
  assign n9626 = n9244 ^ x333 ;
  assign n9627 = n9626 ^ n9308 ;
  assign n9623 = n8564 ^ n8034 ;
  assign n9624 = n9034 & ~n9623 ;
  assign n9625 = n9624 ^ n8034 ;
  assign n9628 = n9627 ^ n9625 ;
  assign n9635 = n9303 ^ x335 ;
  assign n9632 = n8497 ^ n7988 ;
  assign n9633 = n8840 & ~n9632 ;
  assign n9634 = n9633 ^ n7988 ;
  assign n9636 = n9635 ^ n9634 ;
  assign n9637 = n9249 ^ x337 ;
  assign n9638 = n9637 ^ n9292 ;
  assign n9639 = n9638 ^ n7746 ;
  assign n9640 = n9639 ^ n8467 ;
  assign n9641 = n9640 ^ n9638 ;
  assign n9642 = n8857 & ~n9641 ;
  assign n9643 = n9642 ^ n9639 ;
  assign n9696 = n8377 ^ n7731 ;
  assign n9697 = n8866 & n9696 ;
  assign n9698 = n9697 ^ n7731 ;
  assign n9688 = n8245 ^ n7338 ;
  assign n9689 = n8872 & n9688 ;
  assign n9690 = n9689 ^ n7338 ;
  assign n9650 = n8262 ^ n7345 ;
  assign n9651 = ~n8883 & ~n9650 ;
  assign n9652 = n9651 ^ n7345 ;
  assign n9653 = n9652 ^ n9649 ;
  assign n9654 = n9277 ^ n9259 ;
  assign n9674 = n9654 ^ n9652 ;
  assign n9655 = n9654 ^ n7357 ;
  assign n9656 = n9655 ^ n8267 ;
  assign n9657 = n9656 ^ n9654 ;
  assign n9658 = ~n8888 & ~n9657 ;
  assign n9659 = n9658 ^ n9655 ;
  assign n9662 = n8273 ^ n7351 ;
  assign n9663 = n8990 & ~n9662 ;
  assign n9664 = n9663 ^ n7351 ;
  assign n9665 = n9664 ^ n9661 ;
  assign n9537 = n9271 ^ x344 ;
  assign n9538 = n9537 ^ n9262 ;
  assign n9668 = n9664 ^ n9538 ;
  assign n9539 = n9538 ^ n7363 ;
  assign n9540 = n9539 ^ n8278 ;
  assign n9541 = n9540 ^ n9538 ;
  assign n9542 = ~n8980 & n9541 ;
  assign n9543 = n9542 ^ n9539 ;
  assign n9444 = n8355 ^ n7569 ;
  assign n9445 = ~n8893 & n9444 ;
  assign n9446 = n9445 ^ n7569 ;
  assign n8807 = n8806 ^ n8784 ;
  assign n9447 = n9446 ^ n8807 ;
  assign n8809 = n8807 ^ n7559 ;
  assign n8808 = n8807 ^ n8286 ;
  assign n8810 = n8809 ^ n8808 ;
  assign n8811 = ~n8244 & ~n8810 ;
  assign n8812 = n8811 ^ n8809 ;
  assign n8816 = n8291 ^ n7368 ;
  assign n8817 = n8815 & ~n8816 ;
  assign n8818 = n8817 ^ n7368 ;
  assign n8813 = n8802 ^ n8786 ;
  assign n8819 = n8818 ^ n8813 ;
  assign n8826 = n8794 ^ n8793 ;
  assign n8823 = n8332 ^ n7370 ;
  assign n8824 = ~n8822 & n8823 ;
  assign n8825 = n8824 ^ n8332 ;
  assign n8827 = n8826 ^ n8825 ;
  assign n9419 = n8323 ^ n7535 ;
  assign n9420 = n8908 & n9419 ;
  assign n9421 = n9420 ^ n8323 ;
  assign n9416 = n9415 ^ n8832 ;
  assign n9417 = ~n8834 & n9416 ;
  assign n9418 = n9417 ^ n8833 ;
  assign n9422 = n9421 ^ n9418 ;
  assign n9423 = n8789 ^ n8788 ;
  assign n9426 = n9423 ^ n9418 ;
  assign n9427 = n9422 & n9426 ;
  assign n9424 = n9423 ^ n8825 ;
  assign n9428 = n9427 ^ n9424 ;
  assign n9429 = n8827 & n9428 ;
  assign n9430 = n9429 ^ n8826 ;
  assign n9438 = n9430 ^ n8818 ;
  assign n9431 = n9430 ^ n8820 ;
  assign n9432 = n9430 ^ n8294 ;
  assign n9433 = n9432 ^ n7547 ;
  assign n9434 = n9433 ^ n9430 ;
  assign n9435 = ~n8962 & ~n9434 ;
  assign n9436 = n9435 ^ n9432 ;
  assign n9437 = ~n9431 & ~n9436 ;
  assign n9439 = n9438 ^ n9437 ;
  assign n9440 = n8819 & n9439 ;
  assign n9441 = n9440 ^ n8818 ;
  assign n9442 = n9441 ^ n8807 ;
  assign n9443 = ~n8812 & n9442 ;
  assign n9448 = n9447 ^ n9443 ;
  assign n9449 = n9269 ^ n9266 ;
  assign n9534 = n9449 ^ n9446 ;
  assign n9535 = ~n9448 & ~n9534 ;
  assign n9536 = n9535 ^ n9446 ;
  assign n9666 = n9538 ^ n9536 ;
  assign n9667 = ~n9543 & ~n9666 ;
  assign n9669 = n9668 ^ n9667 ;
  assign n9670 = n9665 & ~n9669 ;
  assign n9671 = n9670 ^ n9664 ;
  assign n9672 = n9671 ^ n9654 ;
  assign n9673 = ~n9659 & ~n9672 ;
  assign n9675 = n9674 ^ n9673 ;
  assign n9676 = n9653 & ~n9675 ;
  assign n9677 = n9676 ^ n9652 ;
  assign n9680 = n9679 ^ n9677 ;
  assign n9681 = n9679 ^ n7599 ;
  assign n9682 = n9681 ^ n8256 ;
  assign n9683 = n9682 ^ n9679 ;
  assign n9684 = ~n8877 & ~n9683 ;
  assign n9685 = n9684 ^ n9681 ;
  assign n9686 = n9680 & ~n9685 ;
  assign n9687 = n9686 ^ n9679 ;
  assign n9691 = n9690 ^ n9687 ;
  assign n9692 = n9286 ^ n9253 ;
  assign n9693 = n9692 ^ n9687 ;
  assign n9694 = n9691 & n9693 ;
  assign n9695 = n9694 ^ n9690 ;
  assign n9699 = n9698 ^ n9695 ;
  assign n9700 = n9289 ^ x338 ;
  assign n9701 = n9700 ^ n9250 ;
  assign n9702 = n9701 ^ n9698 ;
  assign n9703 = ~n9699 & ~n9702 ;
  assign n9704 = n9703 ^ n9701 ;
  assign n9644 = n8481 ^ n7947 ;
  assign n9645 = ~n8854 & n9644 ;
  assign n9646 = n9645 ^ n7947 ;
  assign n9647 = n9646 ^ n9638 ;
  assign n9648 = n9647 ^ n9646 ;
  assign n9705 = n9704 ^ n9648 ;
  assign n9706 = ~n9643 & n9705 ;
  assign n9707 = n9706 ^ n9647 ;
  assign n9711 = n9646 ^ n9635 ;
  assign n9708 = n9296 ^ x336 ;
  assign n9709 = n9708 ^ n9297 ;
  assign n9710 = n9709 ^ n9635 ;
  assign n9712 = n9711 ^ n9710 ;
  assign n9713 = n9707 & n9712 ;
  assign n9714 = n9713 ^ n9711 ;
  assign n9715 = ~n9636 & n9714 ;
  assign n9716 = n9715 ^ n9635 ;
  assign n9629 = n9305 ^ x334 ;
  assign n9630 = n9629 ^ n9245 ;
  assign n9717 = n9716 ^ n9630 ;
  assign n9718 = n9630 ^ n8011 ;
  assign n9719 = n9718 ^ n8546 ;
  assign n9720 = n9719 ^ n9630 ;
  assign n9721 = n9024 & n9720 ;
  assign n9722 = n9721 ^ n9718 ;
  assign n9723 = n9717 & n9722 ;
  assign n9631 = n9630 ^ n9627 ;
  assign n9724 = n9723 ^ n9631 ;
  assign n9725 = ~n9628 & ~n9724 ;
  assign n9726 = n9725 ^ n9627 ;
  assign n9618 = n7955 ^ n7286 ;
  assign n9619 = ~n9045 & n9618 ;
  assign n9620 = n9619 ^ n7286 ;
  assign n9621 = n9620 ^ n9612 ;
  assign n9622 = n9621 ^ n9620 ;
  assign n9727 = n9726 ^ n9622 ;
  assign n9728 = n9617 & ~n9727 ;
  assign n9729 = n9728 ^ n9621 ;
  assign n9735 = n9733 ^ n9620 ;
  assign n9730 = n9320 ^ n9317 ;
  assign n9734 = n9733 ^ n9730 ;
  assign n9736 = n9735 ^ n9734 ;
  assign n9737 = n9729 & n9736 ;
  assign n9738 = n9737 ^ n9735 ;
  assign n9739 = n9324 ^ n9243 ;
  assign n9740 = n9739 ^ n9733 ;
  assign n9741 = n9738 & n9740 ;
  assign n9743 = n9742 ^ n9741 ;
  assign n9744 = ~n9610 & ~n9743 ;
  assign n9745 = n9744 ^ n9609 ;
  assign n9746 = n9745 ^ n7473 ;
  assign n9747 = n9746 ^ n8055 ;
  assign n9748 = n9747 ^ n9745 ;
  assign n9749 = ~n8691 & n9748 ;
  assign n9750 = n9749 ^ n9746 ;
  assign n9842 = n9332 ^ n9238 ;
  assign n9751 = n9329 ^ x328 ;
  assign n9752 = n9751 ^ n9239 ;
  assign n9844 = n9842 ^ n9752 ;
  assign n9843 = n9842 ^ n9745 ;
  assign n9845 = n9844 ^ n9843 ;
  assign n9846 = n9750 & n9845 ;
  assign n9847 = n9846 ^ n9844 ;
  assign n9984 = n9335 ^ x326 ;
  assign n9985 = n9984 ^ n9235 ;
  assign n9986 = n9985 ^ n9842 ;
  assign n9987 = n9986 ^ n9985 ;
  assign n9839 = n8079 ^ n7464 ;
  assign n9840 = ~n8684 & n9839 ;
  assign n9841 = n9840 ^ n7464 ;
  assign n9988 = n9987 ^ n9841 ;
  assign n9989 = ~n9847 & n9988 ;
  assign n9990 = n9989 ^ n9986 ;
  assign n9994 = n9993 ^ n9990 ;
  assign n9754 = n9739 ^ n9738 ;
  assign n9755 = n9754 ^ n6714 ;
  assign n9756 = n9730 ^ n9729 ;
  assign n9757 = n9756 ^ n6715 ;
  assign n9818 = n9726 ^ n9617 ;
  assign n9758 = n9724 ^ n9625 ;
  assign n9759 = n9758 ^ n7421 ;
  assign n9809 = n9722 ^ n9716 ;
  assign n9761 = n9709 ^ n9707 ;
  assign n9762 = n9761 ^ n7182 ;
  assign n9763 = n9704 ^ n9643 ;
  assign n9764 = n9763 ^ n7121 ;
  assign n9794 = n9702 ^ n9695 ;
  assign n9765 = n9692 ^ n9690 ;
  assign n9766 = n9765 ^ n9687 ;
  assign n9767 = n9766 ^ n6868 ;
  assign n9769 = n9675 ^ n9649 ;
  assign n9770 = n9769 ^ n6879 ;
  assign n9772 = n9669 ^ n9661 ;
  assign n9773 = n9772 ^ n6890 ;
  assign n9544 = n9543 ^ n9536 ;
  assign n9545 = n9544 ^ n6898 ;
  assign n9452 = n9441 ^ n8812 ;
  assign n9453 = n9452 ^ n6905 ;
  assign n9454 = n9439 ^ n8813 ;
  assign n9455 = n9454 ^ n6907 ;
  assign n9456 = n9436 ^ n8820 ;
  assign n9457 = n9456 ^ n6913 ;
  assign n9458 = n9428 ^ n8826 ;
  assign n9459 = n9458 ^ n6981 ;
  assign n9485 = n9484 ^ n9483 ;
  assign n9487 = n9485 & ~n9486 ;
  assign n9488 = n9487 ^ n6967 ;
  assign n9460 = n9423 ^ n9421 ;
  assign n9461 = n9460 ^ n9418 ;
  assign n9489 = n9488 ^ n9461 ;
  assign n9490 = n9488 ^ n6854 ;
  assign n9491 = n9489 & n9490 ;
  assign n9492 = n9491 ^ n6854 ;
  assign n9493 = n9492 ^ n9458 ;
  assign n9494 = ~n9459 & ~n9493 ;
  assign n9495 = n9494 ^ n6981 ;
  assign n9496 = n9495 ^ n9456 ;
  assign n9497 = n9457 & ~n9496 ;
  assign n9498 = n9497 ^ n6913 ;
  assign n9499 = n9498 ^ n9454 ;
  assign n9500 = n9455 & ~n9499 ;
  assign n9501 = n9500 ^ n6907 ;
  assign n9502 = n9501 ^ n9452 ;
  assign n9503 = n9453 & n9502 ;
  assign n9504 = n9503 ^ n6905 ;
  assign n9450 = n9449 ^ n9448 ;
  assign n9530 = n9504 ^ n9450 ;
  assign n9531 = n9504 ^ n6900 ;
  assign n9532 = ~n9530 & n9531 ;
  assign n9533 = n9532 ^ n6900 ;
  assign n9774 = n9544 ^ n9533 ;
  assign n9775 = ~n9545 & n9774 ;
  assign n9776 = n9775 ^ n6898 ;
  assign n9777 = n9776 ^ n9772 ;
  assign n9778 = ~n9773 & n9777 ;
  assign n9779 = n9778 ^ n6890 ;
  assign n9771 = n9671 ^ n9659 ;
  assign n9780 = n9779 ^ n9771 ;
  assign n9781 = n9779 ^ n6887 ;
  assign n9782 = n9780 & n9781 ;
  assign n9783 = n9782 ^ n6887 ;
  assign n9784 = n9783 ^ n9769 ;
  assign n9785 = n9770 & n9784 ;
  assign n9786 = n9785 ^ n6879 ;
  assign n9768 = n9685 ^ n9677 ;
  assign n9787 = n9786 ^ n9768 ;
  assign n9788 = n9786 ^ n6873 ;
  assign n9789 = ~n9787 & ~n9788 ;
  assign n9790 = n9789 ^ n6873 ;
  assign n9791 = n9790 ^ n9766 ;
  assign n9792 = ~n9767 & n9791 ;
  assign n9793 = n9792 ^ n6868 ;
  assign n9795 = n9794 ^ n9793 ;
  assign n9796 = n9794 ^ n6861 ;
  assign n9797 = n9795 & ~n9796 ;
  assign n9798 = n9797 ^ n6861 ;
  assign n9799 = n9798 ^ n9763 ;
  assign n9800 = n9764 & ~n9799 ;
  assign n9801 = n9800 ^ n7121 ;
  assign n9802 = n9801 ^ n9761 ;
  assign n9803 = n9762 & n9802 ;
  assign n9804 = n9803 ^ n7182 ;
  assign n9760 = n9714 ^ n9634 ;
  assign n9805 = n9804 ^ n9760 ;
  assign n9806 = n9804 ^ n7306 ;
  assign n9807 = n9805 & n9806 ;
  assign n9808 = n9807 ^ n7306 ;
  assign n9810 = n9809 ^ n9808 ;
  assign n9811 = n9758 ^ n7336 ;
  assign n9812 = n9811 ^ n9758 ;
  assign n9813 = n9812 ^ n9808 ;
  assign n9814 = ~n9810 & ~n9813 ;
  assign n9815 = n9814 ^ n9811 ;
  assign n9816 = n9759 & ~n9815 ;
  assign n9817 = n9816 ^ n7421 ;
  assign n9819 = n9818 ^ n9817 ;
  assign n9820 = n9818 ^ n7453 ;
  assign n9821 = ~n9819 & n9820 ;
  assign n9822 = n9821 ^ n7453 ;
  assign n9823 = n9822 ^ n9756 ;
  assign n9824 = ~n9757 & n9823 ;
  assign n9825 = n9824 ^ n6715 ;
  assign n9826 = n9825 ^ n9754 ;
  assign n9827 = ~n9755 & n9826 ;
  assign n9828 = n9827 ^ n6714 ;
  assign n9829 = n9828 ^ n6729 ;
  assign n9830 = n9743 ^ n9609 ;
  assign n9831 = n9830 ^ n9828 ;
  assign n9832 = n9829 & ~n9831 ;
  assign n9833 = n9832 ^ n6729 ;
  assign n9753 = n9752 ^ n9750 ;
  assign n9834 = n9833 ^ n9753 ;
  assign n9835 = n9833 ^ n6711 ;
  assign n9836 = n9834 & n9835 ;
  assign n9837 = n9836 ^ n6711 ;
  assign n9838 = n9837 ^ n6705 ;
  assign n9848 = n9847 ^ n9841 ;
  assign n9980 = n9848 ^ n9837 ;
  assign n9981 = n9838 & ~n9980 ;
  assign n9982 = n9981 ^ n6705 ;
  assign n9983 = n9982 ^ n6744 ;
  assign n9995 = n9994 ^ n9983 ;
  assign n9849 = n9848 ^ n9838 ;
  assign n9850 = n9830 ^ n9829 ;
  assign n9851 = n9760 ^ n7306 ;
  assign n9852 = n9851 ^ n9804 ;
  assign n9853 = n9801 ^ n9762 ;
  assign n9854 = n9798 ^ n9764 ;
  assign n9855 = n9796 ^ n9793 ;
  assign n9856 = n9768 ^ n6873 ;
  assign n9857 = n9856 ^ n9786 ;
  assign n9858 = n9783 ^ n9770 ;
  assign n9859 = n9771 ^ n6887 ;
  assign n9860 = n9859 ^ n9779 ;
  assign n9451 = n9450 ^ n6900 ;
  assign n9505 = n9504 ^ n9451 ;
  assign n9506 = n9492 ^ n9459 ;
  assign n9507 = n9461 ^ n6854 ;
  assign n9508 = n9507 ^ n9488 ;
  assign n9519 = ~n9517 & ~n9518 ;
  assign n9520 = ~n9508 & n9519 ;
  assign n9521 = n9506 & ~n9520 ;
  assign n9522 = n9495 ^ n9457 ;
  assign n9523 = n9521 & n9522 ;
  assign n9524 = n9498 ^ n9455 ;
  assign n9525 = ~n9523 & ~n9524 ;
  assign n9526 = n9501 ^ n6905 ;
  assign n9527 = n9526 ^ n9452 ;
  assign n9528 = n9525 & ~n9527 ;
  assign n9529 = ~n9505 & ~n9528 ;
  assign n9546 = n9545 ^ n9533 ;
  assign n9861 = n9529 & n9546 ;
  assign n9862 = n9776 ^ n6890 ;
  assign n9863 = n9862 ^ n9772 ;
  assign n9864 = n9861 & n9863 ;
  assign n9865 = n9860 & n9864 ;
  assign n9866 = n9858 & ~n9865 ;
  assign n9867 = n9857 & n9866 ;
  assign n9868 = n9790 ^ n9767 ;
  assign n9869 = ~n9867 & n9868 ;
  assign n9870 = ~n9855 & ~n9869 ;
  assign n9871 = n9854 & n9870 ;
  assign n9872 = n9853 & n9871 ;
  assign n9873 = n9852 & n9872 ;
  assign n9874 = n9809 ^ n7336 ;
  assign n9875 = n9874 ^ n9808 ;
  assign n9876 = n9873 & n9875 ;
  assign n9877 = n9815 ^ n7421 ;
  assign n9878 = ~n9876 & ~n9877 ;
  assign n9879 = n9820 ^ n9817 ;
  assign n9880 = ~n9878 & n9879 ;
  assign n9881 = n9822 ^ n9757 ;
  assign n9882 = ~n9880 & n9881 ;
  assign n9883 = n9825 ^ n9755 ;
  assign n9884 = ~n9882 & ~n9883 ;
  assign n9885 = ~n9850 & ~n9884 ;
  assign n9886 = n9835 ^ n9753 ;
  assign n9887 = n9885 & n9886 ;
  assign n9979 = n9849 & ~n9887 ;
  assign n9996 = n9995 ^ n9979 ;
  assign n9891 = n9883 ^ n9882 ;
  assign n9892 = n9891 ^ x357 ;
  assign n9893 = n9881 ^ n9880 ;
  assign n9894 = n9893 ^ x358 ;
  assign n9895 = n9879 ^ n9878 ;
  assign n9896 = n9895 ^ x359 ;
  assign n9897 = n9877 ^ n9876 ;
  assign n9898 = n9897 ^ x360 ;
  assign n9899 = n9875 ^ n9873 ;
  assign n9900 = n9899 ^ x361 ;
  assign n9901 = n9871 ^ n9853 ;
  assign n9902 = n9901 ^ x363 ;
  assign n9903 = n9869 ^ n9855 ;
  assign n9904 = n9903 ^ x365 ;
  assign n9905 = n9868 ^ n9867 ;
  assign n9906 = n9905 ^ x366 ;
  assign n9907 = n9866 ^ n9857 ;
  assign n9908 = n9907 ^ x367 ;
  assign n9910 = n9864 ^ n9860 ;
  assign n9911 = n9910 ^ x369 ;
  assign n9912 = n9863 ^ n9861 ;
  assign n9913 = n9912 ^ x370 ;
  assign n9549 = n9528 ^ n9505 ;
  assign n9550 = n9549 ^ x372 ;
  assign n9597 = n9527 ^ n9525 ;
  assign n9551 = n9524 ^ n9523 ;
  assign n9552 = n9551 ^ x374 ;
  assign n9553 = n9522 ^ n9521 ;
  assign n9554 = n9553 ^ x375 ;
  assign n9555 = n9519 ^ n9508 ;
  assign n9556 = n9555 ^ x377 ;
  assign n9558 = n9557 ^ x378 ;
  assign n9580 = n9579 ^ n9557 ;
  assign n9581 = n9558 & ~n9580 ;
  assign n9582 = n9581 ^ x378 ;
  assign n9583 = n9582 ^ n9555 ;
  assign n9584 = ~n9556 & n9583 ;
  assign n9585 = n9584 ^ x377 ;
  assign n9586 = n9585 ^ x376 ;
  assign n9587 = n9520 ^ n9506 ;
  assign n9588 = n9587 ^ n9585 ;
  assign n9589 = n9586 & ~n9588 ;
  assign n9590 = n9589 ^ x376 ;
  assign n9591 = n9590 ^ n9553 ;
  assign n9592 = ~n9554 & n9591 ;
  assign n9593 = n9592 ^ x375 ;
  assign n9594 = n9593 ^ n9551 ;
  assign n9595 = n9552 & ~n9594 ;
  assign n9596 = n9595 ^ x374 ;
  assign n9598 = n9597 ^ n9596 ;
  assign n9599 = n9597 ^ x373 ;
  assign n9600 = n9598 & ~n9599 ;
  assign n9601 = n9600 ^ x373 ;
  assign n9602 = n9601 ^ n9549 ;
  assign n9603 = ~n9550 & n9602 ;
  assign n9604 = n9603 ^ x372 ;
  assign n9547 = n9546 ^ n9529 ;
  assign n9914 = n9604 ^ n9547 ;
  assign n9915 = n9604 ^ x371 ;
  assign n9916 = n9914 & n9915 ;
  assign n9917 = n9916 ^ x371 ;
  assign n9918 = n9917 ^ n9912 ;
  assign n9919 = ~n9913 & n9918 ;
  assign n9920 = n9919 ^ x370 ;
  assign n9921 = n9920 ^ n9910 ;
  assign n9922 = ~n9911 & n9921 ;
  assign n9923 = n9922 ^ x369 ;
  assign n9909 = n9865 ^ n9858 ;
  assign n9924 = n9923 ^ n9909 ;
  assign n9925 = n9907 ^ x368 ;
  assign n9926 = n9925 ^ n9907 ;
  assign n9927 = n9926 ^ n9909 ;
  assign n9928 = n9924 & ~n9927 ;
  assign n9929 = n9928 ^ n9925 ;
  assign n9930 = n9908 & ~n9929 ;
  assign n9931 = n9930 ^ x367 ;
  assign n9932 = n9931 ^ n9905 ;
  assign n9933 = n9906 & ~n9932 ;
  assign n9934 = n9933 ^ x366 ;
  assign n9935 = n9934 ^ n9903 ;
  assign n9936 = n9904 & ~n9935 ;
  assign n9937 = n9936 ^ x365 ;
  assign n9938 = n9937 ^ x364 ;
  assign n9939 = n9870 ^ n9854 ;
  assign n9940 = n9939 ^ n9937 ;
  assign n9941 = n9938 & ~n9940 ;
  assign n9942 = n9941 ^ x364 ;
  assign n9943 = n9942 ^ n9901 ;
  assign n9944 = n9902 & ~n9943 ;
  assign n9945 = n9944 ^ x363 ;
  assign n9946 = n9945 ^ x362 ;
  assign n9947 = n9872 ^ n9852 ;
  assign n9948 = n9947 ^ n9945 ;
  assign n9949 = n9946 & ~n9948 ;
  assign n9950 = n9949 ^ x362 ;
  assign n9951 = n9950 ^ n9899 ;
  assign n9952 = n9900 & ~n9951 ;
  assign n9953 = n9952 ^ x361 ;
  assign n9954 = n9953 ^ n9897 ;
  assign n9955 = ~n9898 & n9954 ;
  assign n9956 = n9955 ^ x360 ;
  assign n9957 = n9956 ^ n9895 ;
  assign n9958 = ~n9896 & n9957 ;
  assign n9959 = n9958 ^ x359 ;
  assign n9960 = n9959 ^ n9893 ;
  assign n9961 = n9894 & ~n9960 ;
  assign n9962 = n9961 ^ x358 ;
  assign n9963 = n9962 ^ n9891 ;
  assign n9964 = n9892 & ~n9963 ;
  assign n9965 = n9964 ^ x357 ;
  assign n9890 = n9884 ^ n9850 ;
  assign n9966 = n9965 ^ n9890 ;
  assign n9967 = n9965 ^ x356 ;
  assign n9968 = n9966 & n9967 ;
  assign n9969 = n9968 ^ x356 ;
  assign n9889 = n9886 ^ n9885 ;
  assign n9970 = n9969 ^ n9889 ;
  assign n9971 = n9969 ^ x355 ;
  assign n9972 = n9970 & n9971 ;
  assign n9973 = n9972 ^ x355 ;
  assign n9888 = n9887 ^ n9849 ;
  assign n9974 = n9973 ^ n9888 ;
  assign n9975 = n9973 ^ x354 ;
  assign n9976 = n9974 & n9975 ;
  assign n9977 = n9976 ^ x354 ;
  assign n9978 = n9977 ^ x353 ;
  assign n9997 = n9996 ^ n9978 ;
  assign n9998 = n9997 ^ n8185 ;
  assign n9999 = n9998 ^ n8829 ;
  assign n10000 = n9999 ^ n9997 ;
  assign n10001 = n8820 & ~n10000 ;
  assign n10002 = n10001 ^ n9998 ;
  assign n10009 = n8835 ^ n8156 ;
  assign n10010 = ~n8826 & ~n10009 ;
  assign n10011 = n10010 ^ n8156 ;
  assign n10008 = n9975 ^ n9888 ;
  assign n10012 = n10011 ^ n10008 ;
  assign n10018 = n9971 ^ n9889 ;
  assign n10026 = n10018 ^ n10011 ;
  assign n10013 = n9967 ^ n9890 ;
  assign n10014 = n8931 ^ n8095 ;
  assign n10015 = n8833 & n10014 ;
  assign n10016 = n10015 ^ n8095 ;
  assign n10017 = ~n10013 & n10016 ;
  assign n10019 = n10018 ^ n10017 ;
  assign n10020 = n10017 ^ n8104 ;
  assign n10021 = n10020 ^ n8926 ;
  assign n10022 = n10021 ^ n10017 ;
  assign n10023 = n9423 & ~n10022 ;
  assign n10024 = n10023 ^ n10020 ;
  assign n10025 = ~n10019 & ~n10024 ;
  assign n10027 = n10026 ^ n10025 ;
  assign n10028 = ~n10012 & ~n10027 ;
  assign n10029 = n10028 ^ n10011 ;
  assign n10003 = n8908 ^ n8308 ;
  assign n10004 = ~n8813 & ~n10003 ;
  assign n10005 = n10004 ^ n8308 ;
  assign n10006 = n10005 ^ n9997 ;
  assign n10007 = n10006 ^ n10005 ;
  assign n10030 = n10029 ^ n10007 ;
  assign n10031 = ~n10002 & ~n10030 ;
  assign n10032 = n10031 ^ n10006 ;
  assign n10033 = n8822 ^ n8306 ;
  assign n10034 = ~n8807 & ~n10033 ;
  assign n10035 = n10034 ^ n8306 ;
  assign n10059 = n10035 ^ n10005 ;
  assign n10051 = n7334 ^ n7325 ;
  assign n10052 = ~n8737 & ~n10051 ;
  assign n10046 = n9341 ^ n9338 ;
  assign n10047 = n10046 ^ n9371 ;
  assign n10048 = n10047 ^ n9993 ;
  assign n10049 = n10048 ^ n6744 ;
  assign n10045 = x353 ^ x352 ;
  assign n10050 = n10049 ^ n10045 ;
  assign n10053 = n10052 ^ n10050 ;
  assign n10043 = n9993 ^ n9985 ;
  assign n10044 = ~n9990 & n10043 ;
  assign n10054 = n10053 ^ n10044 ;
  assign n10042 = ~n9979 & ~n9995 ;
  assign n10055 = n10054 ^ n10042 ;
  assign n10039 = n9996 ^ n9977 ;
  assign n10040 = n9996 ^ x353 ;
  assign n10041 = n10039 & ~n10040 ;
  assign n10056 = n10055 ^ n10041 ;
  assign n10036 = n9994 ^ n9982 ;
  assign n10037 = n9994 ^ n6744 ;
  assign n10038 = n10036 & n10037 ;
  assign n10057 = n10056 ^ n10038 ;
  assign n10058 = n10057 ^ n10035 ;
  assign n10060 = n10059 ^ n10058 ;
  assign n10061 = ~n10032 & n10060 ;
  assign n10062 = n10061 ^ n10059 ;
  assign n10064 = n9565 ^ n9562 ;
  assign n10066 = n10064 ^ n10035 ;
  assign n10063 = n9510 ^ x383 ;
  assign n10065 = n10064 ^ n10063 ;
  assign n10067 = n10066 ^ n10065 ;
  assign n10068 = ~n10062 & n10067 ;
  assign n10069 = n10068 ^ n10066 ;
  assign n10118 = n8815 ^ n8332 ;
  assign n10119 = ~n9538 & ~n10118 ;
  assign n10120 = n10119 ^ n8332 ;
  assign n10122 = n10120 ^ n10064 ;
  assign n10070 = n8962 ^ n8323 ;
  assign n10071 = ~n9449 & ~n10070 ;
  assign n10072 = n10071 ^ n8323 ;
  assign n10121 = n10120 ^ n10072 ;
  assign n10123 = n10122 ^ n10121 ;
  assign n10124 = ~n10069 & ~n10123 ;
  assign n10125 = n10124 ^ n10122 ;
  assign n10126 = n9561 ^ x381 ;
  assign n10127 = n10126 ^ n9567 ;
  assign n10294 = n10127 ^ n10120 ;
  assign n10295 = ~n10125 & ~n10294 ;
  assign n10296 = n10295 ^ n10120 ;
  assign n10290 = n8893 ^ n8291 ;
  assign n10291 = ~n9654 & ~n10290 ;
  assign n10292 = n10291 ^ n8291 ;
  assign n10293 = n10292 ^ n10284 ;
  assign n10297 = n10296 ^ n10293 ;
  assign n10298 = n10297 ^ n10292 ;
  assign n10299 = ~n10289 & n10298 ;
  assign n10300 = n10299 ^ n10293 ;
  assign n10301 = n9577 ^ n9574 ;
  assign n10302 = n10301 ^ n10292 ;
  assign n10303 = n10300 & ~n10302 ;
  assign n10304 = n10303 ^ n10301 ;
  assign n10306 = n10305 ^ n10304 ;
  assign n10307 = n10306 ^ n10277 ;
  assign n10308 = ~n10282 & ~n10307 ;
  assign n10309 = n10308 ^ n10305 ;
  assign n10200 = n9582 ^ n9556 ;
  assign n10444 = n10309 ^ n10200 ;
  assign n10445 = n10444 ^ n7569 ;
  assign n10447 = n10296 ^ n10289 ;
  assign n10448 = n10447 ^ n7547 ;
  assign n10074 = n10063 ^ n10062 ;
  assign n10075 = n10074 ^ n6851 ;
  assign n10076 = n10029 ^ n10002 ;
  assign n10077 = n10076 ^ n7328 ;
  assign n10085 = n10027 ^ n10008 ;
  assign n10078 = n10016 ^ n10013 ;
  assign n10079 = n7386 & ~n10078 ;
  assign n10080 = n10079 ^ n7377 ;
  assign n10081 = n10024 ^ n10018 ;
  assign n10082 = n10081 ^ n10079 ;
  assign n10083 = n10080 & n10082 ;
  assign n10084 = n10083 ^ n7377 ;
  assign n10086 = n10085 ^ n10084 ;
  assign n10087 = n10085 ^ n7506 ;
  assign n10088 = ~n10086 & n10087 ;
  assign n10089 = n10088 ^ n7506 ;
  assign n10090 = n10089 ^ n10076 ;
  assign n10091 = n10077 & n10090 ;
  assign n10092 = n10091 ^ n7328 ;
  assign n10093 = n10092 ^ n6852 ;
  assign n10094 = n10057 ^ n10032 ;
  assign n10095 = n10094 ^ n10092 ;
  assign n10096 = ~n10093 & ~n10095 ;
  assign n10097 = n10096 ^ n6852 ;
  assign n10098 = n10097 ^ n10074 ;
  assign n10099 = ~n10075 & ~n10098 ;
  assign n10100 = n10099 ^ n6851 ;
  assign n10101 = n10100 ^ n7535 ;
  assign n10073 = n10072 ^ n10069 ;
  assign n10130 = n10100 ^ n10073 ;
  assign n10131 = n10101 & n10130 ;
  assign n10132 = n10131 ^ n7535 ;
  assign n10128 = n10127 ^ n10125 ;
  assign n10449 = n10132 ^ n10128 ;
  assign n10450 = n10132 ^ n7370 ;
  assign n10451 = ~n10449 & n10450 ;
  assign n10452 = n10451 ^ n7370 ;
  assign n10453 = n10452 ^ n10447 ;
  assign n10454 = ~n10448 & n10453 ;
  assign n10455 = n10454 ^ n7547 ;
  assign n10456 = n10455 ^ n7368 ;
  assign n10457 = n10301 ^ n10300 ;
  assign n10458 = n10457 ^ n10455 ;
  assign n10459 = n10456 & n10458 ;
  assign n10460 = n10459 ^ n7368 ;
  assign n10446 = n10304 ^ n10282 ;
  assign n10461 = n10460 ^ n10446 ;
  assign n10462 = n10460 ^ n7559 ;
  assign n10463 = n10461 & ~n10462 ;
  assign n10464 = n10463 ^ n7559 ;
  assign n10465 = n10464 ^ n10444 ;
  assign n10466 = ~n10445 & n10465 ;
  assign n10467 = n10466 ^ n7569 ;
  assign n10278 = n10277 ^ n10200 ;
  assign n10310 = ~n10278 & ~n10309 ;
  assign n10311 = n10310 ^ n10200 ;
  assign n10193 = n9587 ^ n9586 ;
  assign n10266 = n10193 ^ n8278 ;
  assign n10267 = n10266 ^ n8888 ;
  assign n10268 = n10267 ^ n10193 ;
  assign n10269 = ~n9692 & ~n10268 ;
  assign n10270 = n10269 ^ n10266 ;
  assign n10443 = n10311 ^ n10270 ;
  assign n10468 = n10467 ^ n10443 ;
  assign n10469 = n10467 ^ n7363 ;
  assign n10470 = n10468 & n10469 ;
  assign n10471 = n10470 ^ n7363 ;
  assign n10316 = n9590 ^ x375 ;
  assign n10317 = n10316 ^ n9553 ;
  assign n10271 = n8883 ^ n8273 ;
  assign n10272 = ~n9701 & n10271 ;
  assign n10273 = n10272 ^ n8273 ;
  assign n10274 = n10273 ^ n10193 ;
  assign n10312 = n10311 ^ n10274 ;
  assign n10313 = n10312 ^ n10273 ;
  assign n10314 = n10270 & ~n10313 ;
  assign n10315 = n10314 ^ n10274 ;
  assign n10441 = n10317 ^ n10315 ;
  assign n10442 = n10441 ^ n7351 ;
  assign n10556 = n10471 ^ n10442 ;
  assign n10543 = n10452 ^ n10448 ;
  assign n10102 = n10101 ^ n10073 ;
  assign n10103 = n10089 ^ n7328 ;
  assign n10104 = n10103 ^ n10076 ;
  assign n10105 = n10084 ^ n7506 ;
  assign n10106 = n10105 ^ n10085 ;
  assign n10107 = n10078 ^ n7386 ;
  assign n10108 = n10081 ^ n10080 ;
  assign n10109 = ~n10107 & ~n10108 ;
  assign n10110 = n10106 & n10109 ;
  assign n10111 = ~n10104 & ~n10110 ;
  assign n10112 = n10094 ^ n10093 ;
  assign n10113 = n10111 & ~n10112 ;
  assign n10114 = n10097 ^ n6851 ;
  assign n10115 = n10114 ^ n10074 ;
  assign n10116 = ~n10113 & ~n10115 ;
  assign n10117 = n10102 & n10116 ;
  assign n10129 = n10128 ^ n7370 ;
  assign n10133 = n10132 ^ n10129 ;
  assign n10544 = ~n10117 & n10133 ;
  assign n10545 = ~n10543 & n10544 ;
  assign n10546 = n10457 ^ n10456 ;
  assign n10547 = ~n10545 & n10546 ;
  assign n10548 = n10446 ^ n7559 ;
  assign n10549 = n10548 ^ n10460 ;
  assign n10550 = n10547 & ~n10549 ;
  assign n10551 = n10464 ^ n10445 ;
  assign n10552 = ~n10550 & n10551 ;
  assign n10553 = n10443 ^ n7363 ;
  assign n10554 = n10553 ^ n10467 ;
  assign n10555 = n10552 & n10554 ;
  assign n10615 = n10556 ^ n10555 ;
  assign n10616 = n10615 ^ x402 ;
  assign n10617 = n10554 ^ n10552 ;
  assign n10618 = n10617 ^ x403 ;
  assign n10619 = n10551 ^ n10550 ;
  assign n10620 = n10619 ^ x404 ;
  assign n10621 = n10549 ^ n10547 ;
  assign n10622 = n10621 ^ x405 ;
  assign n10623 = n10546 ^ n10545 ;
  assign n10624 = n10623 ^ x406 ;
  assign n10625 = n10544 ^ n10543 ;
  assign n10626 = n10625 ^ x407 ;
  assign n10135 = n10116 ^ n10102 ;
  assign n10136 = n10135 ^ x409 ;
  assign n10137 = n10112 ^ n10111 ;
  assign n10138 = n10137 ^ x411 ;
  assign n10146 = n10109 ^ n10106 ;
  assign n10140 = x415 & n10107 ;
  assign n10141 = n10140 ^ x414 ;
  assign n10142 = n10108 ^ n10107 ;
  assign n10143 = n10142 ^ n10140 ;
  assign n10144 = n10141 & ~n10143 ;
  assign n10145 = n10144 ^ x414 ;
  assign n10147 = n10146 ^ n10145 ;
  assign n10148 = n10146 ^ x413 ;
  assign n10149 = ~n10147 & n10148 ;
  assign n10150 = n10149 ^ x413 ;
  assign n10139 = n10110 ^ n10104 ;
  assign n10151 = n10150 ^ n10139 ;
  assign n10152 = n10150 ^ x412 ;
  assign n10153 = n10151 & n10152 ;
  assign n10154 = n10153 ^ x412 ;
  assign n10155 = n10154 ^ n10137 ;
  assign n10156 = n10138 & ~n10155 ;
  assign n10157 = n10156 ^ x411 ;
  assign n10158 = n10157 ^ x410 ;
  assign n10159 = n10115 ^ n10113 ;
  assign n10160 = n10159 ^ n10157 ;
  assign n10161 = n10158 & ~n10160 ;
  assign n10162 = n10161 ^ x410 ;
  assign n10163 = n10162 ^ n10135 ;
  assign n10164 = n10136 & ~n10163 ;
  assign n10165 = n10164 ^ x409 ;
  assign n10166 = n10165 ^ x408 ;
  assign n10134 = n10133 ^ n10117 ;
  assign n10627 = n10165 ^ n10134 ;
  assign n10628 = n10166 & ~n10627 ;
  assign n10629 = n10628 ^ x408 ;
  assign n10630 = n10629 ^ n10625 ;
  assign n10631 = n10626 & ~n10630 ;
  assign n10632 = n10631 ^ x407 ;
  assign n10633 = n10632 ^ n10623 ;
  assign n10634 = ~n10624 & n10633 ;
  assign n10635 = n10634 ^ x406 ;
  assign n10636 = n10635 ^ n10621 ;
  assign n10637 = ~n10622 & n10636 ;
  assign n10638 = n10637 ^ x405 ;
  assign n10639 = n10638 ^ n10619 ;
  assign n10640 = n10620 & ~n10639 ;
  assign n10641 = n10640 ^ x404 ;
  assign n10642 = n10641 ^ n10617 ;
  assign n10643 = ~n10618 & n10642 ;
  assign n10644 = n10643 ^ x403 ;
  assign n10645 = n10644 ^ n10615 ;
  assign n10646 = n10616 & ~n10645 ;
  assign n10647 = n10646 ^ x402 ;
  assign n10472 = n10471 ^ n10441 ;
  assign n10473 = n10442 & ~n10472 ;
  assign n10474 = n10473 ^ n7351 ;
  assign n10318 = n10317 ^ n10273 ;
  assign n10319 = n10315 & n10318 ;
  assign n10320 = n10319 ^ n10317 ;
  assign n10187 = n9593 ^ n9552 ;
  assign n10260 = n10187 ^ n8267 ;
  assign n10261 = n10260 ^ n8877 ;
  assign n10262 = n10261 ^ n10187 ;
  assign n10263 = ~n9638 & n10262 ;
  assign n10264 = n10263 ^ n10260 ;
  assign n10439 = n10320 ^ n10264 ;
  assign n10440 = n10439 ^ n7357 ;
  assign n10558 = n10474 ^ n10440 ;
  assign n10557 = n10555 & ~n10556 ;
  assign n10613 = n10558 ^ n10557 ;
  assign n10614 = n10613 ^ x401 ;
  assign n11019 = n10647 ^ n10614 ;
  assign n10223 = n9939 ^ n9938 ;
  assign n11016 = n9739 ^ n8840 ;
  assign n11017 = n10223 & ~n11016 ;
  assign n11018 = n11017 ^ n8840 ;
  assign n11020 = n11019 ^ n11018 ;
  assign n10227 = n9934 ^ n9904 ;
  assign n11023 = n9730 ^ n8854 ;
  assign n11024 = n10227 & n11023 ;
  assign n11025 = n11024 ^ n8854 ;
  assign n11021 = n10644 ^ x402 ;
  assign n11022 = n11021 ^ n10615 ;
  assign n11026 = n11025 ^ n11022 ;
  assign n11048 = n10641 ^ n10618 ;
  assign n10350 = n9929 ^ x367 ;
  assign n11029 = n9627 ^ n8866 ;
  assign n11030 = n10350 & n11029 ;
  assign n11031 = n11030 ^ n8866 ;
  assign n11027 = n10638 ^ x404 ;
  assign n11028 = n11027 ^ n10619 ;
  assign n11032 = n11031 ^ n11028 ;
  assign n10245 = n9920 ^ n9911 ;
  assign n10962 = n9635 ^ n8877 ;
  assign n10963 = ~n10245 & n10962 ;
  assign n10964 = n10963 ^ n8877 ;
  assign n10961 = n10632 ^ n10624 ;
  assign n10965 = n10964 ^ n10961 ;
  assign n9548 = n9547 ^ x371 ;
  assign n9605 = n9604 ^ n9548 ;
  assign n10167 = n10166 ^ n10134 ;
  assign n10168 = n10167 ^ n9638 ;
  assign n10169 = n10168 ^ n8888 ;
  assign n10170 = n10169 ^ n10167 ;
  assign n10171 = n9605 & n10170 ;
  assign n10172 = n10171 ^ n10168 ;
  assign n10178 = n10162 ^ x409 ;
  assign n10179 = n10178 ^ n10135 ;
  assign n10173 = n9601 ^ x372 ;
  assign n10174 = n10173 ^ n9549 ;
  assign n10175 = n9701 ^ n8990 ;
  assign n10176 = n10174 & ~n10175 ;
  assign n10177 = n10176 ^ n9701 ;
  assign n10180 = n10179 ^ n10177 ;
  assign n10182 = n9599 ^ n9596 ;
  assign n10183 = n9692 ^ n8980 ;
  assign n10184 = ~n10182 & n10183 ;
  assign n10185 = n10184 ^ n8980 ;
  assign n10181 = n10159 ^ n10158 ;
  assign n10186 = n10185 ^ n10181 ;
  assign n10191 = n10154 ^ n10138 ;
  assign n10188 = n9679 ^ n8893 ;
  assign n10189 = n10187 & ~n10188 ;
  assign n10190 = n10189 ^ n8893 ;
  assign n10192 = n10191 ^ n10190 ;
  assign n10772 = n10152 ^ n10139 ;
  assign n10194 = n10148 ^ n10145 ;
  assign n10195 = n10194 ^ n8815 ;
  assign n10196 = n10195 ^ n9654 ;
  assign n10197 = n10196 ^ n10194 ;
  assign n10198 = n10193 & ~n10197 ;
  assign n10199 = n10198 ^ n10195 ;
  assign n10204 = n10142 ^ n10141 ;
  assign n10201 = n9661 ^ n8962 ;
  assign n10202 = ~n10200 & n10201 ;
  assign n10203 = n10202 ^ n8962 ;
  assign n10205 = n10204 ^ n10203 ;
  assign n10211 = n10107 ^ x415 ;
  assign n10208 = n9538 ^ n8822 ;
  assign n10209 = n10207 & ~n10208 ;
  assign n10210 = n10209 ^ n8822 ;
  assign n10212 = n10211 ^ n10210 ;
  assign n10725 = n9449 ^ n8908 ;
  assign n10726 = ~n10301 & n10725 ;
  assign n10727 = n10726 ^ n8908 ;
  assign n10762 = n10727 ^ n10210 ;
  assign n10413 = n9959 ^ n9894 ;
  assign n10410 = n8770 ^ n7332 ;
  assign n10411 = ~n9384 & n10410 ;
  assign n10412 = n10411 ^ n7332 ;
  assign n10414 = n10413 ^ n10412 ;
  assign n10216 = n9956 ^ n9896 ;
  assign n10213 = n8737 ^ n8079 ;
  assign n10214 = ~n9386 & n10213 ;
  assign n10215 = n10214 ^ n8079 ;
  assign n10217 = n10216 ^ n10215 ;
  assign n10219 = n8684 ^ n8021 ;
  assign n10220 = ~n9393 & ~n10219 ;
  assign n10221 = n10220 ^ n8021 ;
  assign n10218 = n9950 ^ n9900 ;
  assign n10222 = n10221 ^ n10218 ;
  assign n10224 = n9045 ^ n8564 ;
  assign n10225 = n9752 & ~n10224 ;
  assign n10226 = n10225 ^ n8564 ;
  assign n10228 = n10227 ^ n10226 ;
  assign n10231 = n9035 ^ n8546 ;
  assign n10232 = n9609 & ~n10231 ;
  assign n10233 = n10232 ^ n8546 ;
  assign n10229 = n9931 ^ n9906 ;
  assign n10234 = n10233 ^ n10229 ;
  assign n10235 = n9923 ^ x368 ;
  assign n10236 = n10235 ^ n9909 ;
  assign n10351 = n10350 ^ n10236 ;
  assign n10237 = n10236 ^ n8481 ;
  assign n10238 = n10237 ^ n9024 ;
  assign n10239 = n10238 ^ n10236 ;
  assign n10240 = ~n9730 & ~n10239 ;
  assign n10241 = n10240 ^ n10237 ;
  assign n10242 = n8840 ^ n8467 ;
  assign n10243 = ~n9612 & ~n10242 ;
  assign n10244 = n10243 ^ n8467 ;
  assign n10246 = n10245 ^ n10244 ;
  assign n10247 = n8857 ^ n8245 ;
  assign n10248 = n9630 & n10247 ;
  assign n10249 = n10248 ^ n8857 ;
  assign n10250 = n10249 ^ n9605 ;
  assign n10251 = n10174 ^ n8256 ;
  assign n10252 = n10251 ^ n8866 ;
  assign n10253 = n10252 ^ n10174 ;
  assign n10254 = ~n9635 & n10253 ;
  assign n10255 = n10254 ^ n10251 ;
  assign n10327 = n10249 ^ n10174 ;
  assign n10256 = n8872 ^ n8262 ;
  assign n10257 = ~n9709 & ~n10256 ;
  assign n10258 = n10257 ^ n8262 ;
  assign n10259 = n10258 ^ n10182 ;
  assign n10321 = n10320 ^ n10258 ;
  assign n10265 = n10258 ^ n10187 ;
  assign n10322 = n10321 ^ n10265 ;
  assign n10323 = ~n10264 & ~n10322 ;
  assign n10324 = n10323 ^ n10265 ;
  assign n10325 = n10259 & ~n10324 ;
  assign n10326 = n10325 ^ n10258 ;
  assign n10328 = n10327 ^ n10326 ;
  assign n10329 = n10328 ^ n10249 ;
  assign n10330 = ~n10255 & n10329 ;
  assign n10331 = n10330 ^ n10327 ;
  assign n10332 = ~n10250 & n10331 ;
  assign n10333 = n10332 ^ n9605 ;
  assign n10334 = n10333 ^ n8377 ;
  assign n10335 = n10334 ^ n8854 ;
  assign n10336 = n10335 ^ n10333 ;
  assign n10337 = n9627 & ~n10336 ;
  assign n10338 = n10337 ^ n10334 ;
  assign n10340 = n9917 ^ x370 ;
  assign n10341 = n10340 ^ n9912 ;
  assign n10342 = n10341 ^ n10244 ;
  assign n10339 = n10333 ^ n10244 ;
  assign n10343 = n10342 ^ n10339 ;
  assign n10344 = n10338 & n10343 ;
  assign n10345 = n10344 ^ n10342 ;
  assign n10346 = n10246 & ~n10345 ;
  assign n10347 = n10346 ^ n10245 ;
  assign n10348 = n10347 ^ n10236 ;
  assign n10349 = n10241 & n10348 ;
  assign n10352 = n10351 ^ n10349 ;
  assign n10355 = n9034 ^ n8497 ;
  assign n10356 = ~n9739 & ~n10355 ;
  assign n10357 = n10356 ^ n8497 ;
  assign n10353 = n10350 ^ n10229 ;
  assign n10354 = n10353 ^ n10229 ;
  assign n10358 = n10357 ^ n10354 ;
  assign n10359 = ~n10352 & ~n10358 ;
  assign n10360 = n10359 ^ n10353 ;
  assign n10361 = ~n10234 & n10360 ;
  assign n10230 = n10229 ^ n10226 ;
  assign n10362 = n10361 ^ n10230 ;
  assign n10363 = n10228 & ~n10362 ;
  assign n10364 = n10363 ^ n10227 ;
  assign n10365 = n10364 ^ n10223 ;
  assign n10366 = n10223 ^ n8722 ;
  assign n10367 = n10366 ^ n9366 ;
  assign n10368 = n10367 ^ n10223 ;
  assign n10369 = ~n9842 & ~n10368 ;
  assign n10370 = n10369 ^ n10366 ;
  assign n10371 = n10365 & n10370 ;
  assign n10372 = n10371 ^ n10364 ;
  assign n10373 = n10372 ^ n7955 ;
  assign n10374 = n10373 ^ n8696 ;
  assign n10375 = n10374 ^ n10372 ;
  assign n10376 = ~n9985 & n10375 ;
  assign n10377 = n10376 ^ n10373 ;
  assign n10382 = n9942 ^ x363 ;
  assign n10383 = n10382 ^ n9901 ;
  assign n10378 = n8691 ^ n7992 ;
  assign n10379 = ~n10046 & ~n10378 ;
  assign n10380 = n10379 ^ n7992 ;
  assign n10384 = n10383 ^ n10380 ;
  assign n10381 = n10380 ^ n10372 ;
  assign n10385 = n10384 ^ n10381 ;
  assign n10386 = n10377 & n10385 ;
  assign n10387 = n10386 ^ n10384 ;
  assign n10390 = n10380 ^ n10221 ;
  assign n10388 = n9947 ^ n9946 ;
  assign n10389 = n10388 ^ n10221 ;
  assign n10391 = n10390 ^ n10389 ;
  assign n10392 = ~n10387 & n10391 ;
  assign n10393 = n10392 ^ n10389 ;
  assign n10394 = n10222 & n10393 ;
  assign n10395 = n10394 ^ n10221 ;
  assign n10396 = n10395 ^ n8055 ;
  assign n10397 = n10396 ^ n8683 ;
  assign n10398 = n10397 ^ n10395 ;
  assign n10399 = n9398 & ~n10398 ;
  assign n10400 = n10399 ^ n10396 ;
  assign n10404 = n10395 ^ n10216 ;
  assign n10401 = n9953 ^ x360 ;
  assign n10402 = n10401 ^ n9897 ;
  assign n10403 = n10402 ^ n10216 ;
  assign n10405 = n10404 ^ n10403 ;
  assign n10406 = ~n10400 & ~n10405 ;
  assign n10407 = n10406 ^ n10404 ;
  assign n10408 = n10217 & ~n10407 ;
  assign n10409 = n10408 ^ n10216 ;
  assign n10719 = n10412 ^ n10409 ;
  assign n10720 = n10414 & ~n10719 ;
  assign n10716 = n8936 ^ n7325 ;
  assign n10717 = n9379 & n10716 ;
  assign n10712 = n10412 ^ n10051 ;
  assign n10711 = n9962 ^ n9892 ;
  assign n10713 = n10712 ^ n10711 ;
  assign n10714 = n10713 ^ n7401 ;
  assign n10710 = x385 ^ x384 ;
  assign n10715 = n10714 ^ n10710 ;
  assign n10718 = n10717 ^ n10715 ;
  assign n10721 = n10720 ^ n10718 ;
  assign n10423 = n10370 ^ n10364 ;
  assign n10534 = n10423 ^ n8066 ;
  assign n10424 = n10362 ^ n10227 ;
  assign n10425 = n10424 ^ n8034 ;
  assign n10427 = n10357 ^ n10352 ;
  assign n10428 = n10427 ^ n7988 ;
  assign n10429 = n10347 ^ n10241 ;
  assign n10430 = n10429 ^ n7947 ;
  assign n10431 = n10345 ^ n10245 ;
  assign n10432 = n10431 ^ n7746 ;
  assign n10433 = n10341 ^ n10338 ;
  assign n10434 = n10433 ^ n7731 ;
  assign n10436 = n10326 ^ n10255 ;
  assign n10437 = n10436 ^ n7599 ;
  assign n10475 = n10474 ^ n10439 ;
  assign n10476 = n10440 & ~n10475 ;
  assign n10477 = n10476 ^ n7357 ;
  assign n10438 = n10324 ^ n10182 ;
  assign n10478 = n10477 ^ n10438 ;
  assign n10479 = n10477 ^ n7345 ;
  assign n10480 = ~n10478 & n10479 ;
  assign n10481 = n10480 ^ n7345 ;
  assign n10482 = n10481 ^ n10436 ;
  assign n10483 = ~n10437 & ~n10482 ;
  assign n10484 = n10483 ^ n7599 ;
  assign n10435 = n10331 ^ n9605 ;
  assign n10485 = n10484 ^ n10435 ;
  assign n10486 = n10484 ^ n7338 ;
  assign n10487 = n10485 & ~n10486 ;
  assign n10488 = n10487 ^ n7338 ;
  assign n10489 = n10488 ^ n10433 ;
  assign n10490 = n10434 & ~n10489 ;
  assign n10491 = n10490 ^ n7731 ;
  assign n10492 = n10491 ^ n10431 ;
  assign n10493 = ~n10432 & n10492 ;
  assign n10494 = n10493 ^ n7746 ;
  assign n10495 = n10494 ^ n10429 ;
  assign n10496 = n10430 & n10495 ;
  assign n10497 = n10496 ^ n7947 ;
  assign n10498 = n10497 ^ n10427 ;
  assign n10499 = n10428 & n10498 ;
  assign n10500 = n10499 ^ n7988 ;
  assign n10426 = n10360 ^ n10233 ;
  assign n10501 = n10500 ^ n10426 ;
  assign n10502 = n10500 ^ n8011 ;
  assign n10503 = n10501 & ~n10502 ;
  assign n10504 = n10503 ^ n8011 ;
  assign n10505 = n10504 ^ n10424 ;
  assign n10506 = ~n10425 & n10505 ;
  assign n10507 = n10506 ^ n8034 ;
  assign n10535 = n10534 ^ n10507 ;
  assign n10536 = n10504 ^ n8034 ;
  assign n10537 = n10536 ^ n10424 ;
  assign n10538 = n10426 ^ n8011 ;
  assign n10539 = n10538 ^ n10500 ;
  assign n10540 = n10435 ^ n7338 ;
  assign n10541 = n10540 ^ n10484 ;
  assign n10542 = n10481 ^ n10437 ;
  assign n10559 = n10557 & ~n10558 ;
  assign n10560 = n10438 ^ n7345 ;
  assign n10561 = n10560 ^ n10477 ;
  assign n10562 = ~n10559 & n10561 ;
  assign n10563 = ~n10542 & n10562 ;
  assign n10564 = n10541 & ~n10563 ;
  assign n10565 = n10488 ^ n10434 ;
  assign n10566 = ~n10564 & n10565 ;
  assign n10567 = n10491 ^ n7746 ;
  assign n10568 = n10567 ^ n10431 ;
  assign n10569 = n10566 & ~n10568 ;
  assign n10570 = n10494 ^ n10430 ;
  assign n10571 = n10569 & n10570 ;
  assign n10572 = n10497 ^ n10428 ;
  assign n10573 = n10571 & ~n10572 ;
  assign n10574 = n10539 & n10573 ;
  assign n10575 = ~n10537 & ~n10574 ;
  assign n10576 = ~n10535 & ~n10575 ;
  assign n10508 = n10507 ^ n10423 ;
  assign n10509 = n10507 ^ n8066 ;
  assign n10510 = ~n10508 & n10509 ;
  assign n10511 = n10510 ^ n8066 ;
  assign n10421 = n10383 ^ n10377 ;
  assign n10422 = n10421 ^ n7286 ;
  assign n10577 = n10511 ^ n10422 ;
  assign n10578 = ~n10576 & n10577 ;
  assign n10515 = n10388 ^ n10387 ;
  assign n10517 = n10515 ^ n7315 ;
  assign n10512 = n10511 ^ n10421 ;
  assign n10513 = n10422 & ~n10512 ;
  assign n10514 = n10513 ^ n7286 ;
  assign n10579 = n10517 ^ n10514 ;
  assign n10580 = ~n10578 & n10579 ;
  assign n10516 = n10515 ^ n10514 ;
  assign n10518 = n10516 & ~n10517 ;
  assign n10519 = n10518 ^ n7315 ;
  assign n10521 = n10519 ^ n7475 ;
  assign n10420 = n10393 ^ n10218 ;
  assign n10581 = n10521 ^ n10420 ;
  assign n10582 = ~n10580 & ~n10581 ;
  assign n10520 = n10519 ^ n10420 ;
  assign n10522 = n10520 & n10521 ;
  assign n10523 = n10522 ^ n7475 ;
  assign n10583 = n10523 ^ n7473 ;
  assign n10419 = n10402 ^ n10400 ;
  assign n10584 = n10583 ^ n10419 ;
  assign n10585 = n10582 & ~n10584 ;
  assign n10524 = n10523 ^ n10419 ;
  assign n10527 = n10419 ^ n7473 ;
  assign n10528 = n10524 & ~n10527 ;
  assign n10525 = n7473 ^ n7464 ;
  assign n10529 = n10528 ^ n10525 ;
  assign n10417 = n10407 ^ n10215 ;
  assign n10586 = n10529 ^ n10417 ;
  assign n10587 = ~n10585 & n10586 ;
  assign n10418 = n10417 ^ n7464 ;
  assign n10530 = ~n10418 & n10529 ;
  assign n10531 = n10530 ^ n7464 ;
  assign n10588 = n10531 ^ n7401 ;
  assign n10415 = n10414 ^ n10409 ;
  assign n10589 = n10588 ^ n10415 ;
  assign n10709 = ~n10587 & n10589 ;
  assign n10722 = n10721 ^ n10709 ;
  assign n10593 = n10579 ^ n10578 ;
  assign n10594 = n10593 ^ x389 ;
  assign n10595 = n10577 ^ n10576 ;
  assign n10596 = n10595 ^ x390 ;
  assign n10597 = n10575 ^ n10535 ;
  assign n10598 = n10597 ^ x391 ;
  assign n10600 = n10573 ^ n10539 ;
  assign n10601 = n10600 ^ x393 ;
  assign n10602 = n10572 ^ n10571 ;
  assign n10603 = n10602 ^ x394 ;
  assign n10604 = n10570 ^ n10569 ;
  assign n10605 = n10604 ^ x395 ;
  assign n10606 = n10568 ^ n10566 ;
  assign n10607 = n10606 ^ x396 ;
  assign n10608 = n10565 ^ n10564 ;
  assign n10609 = n10608 ^ x397 ;
  assign n10610 = n10562 ^ n10542 ;
  assign n10611 = n10610 ^ x399 ;
  assign n10648 = n10647 ^ n10613 ;
  assign n10649 = n10614 & ~n10648 ;
  assign n10650 = n10649 ^ x401 ;
  assign n10612 = n10561 ^ n10559 ;
  assign n10651 = n10650 ^ n10612 ;
  assign n10652 = n10610 ^ x400 ;
  assign n10653 = n10652 ^ n10612 ;
  assign n10654 = n10653 ^ n10610 ;
  assign n10655 = n10651 & ~n10654 ;
  assign n10656 = n10655 ^ n10652 ;
  assign n10657 = ~n10611 & n10656 ;
  assign n10658 = n10657 ^ x399 ;
  assign n10659 = n10658 ^ x398 ;
  assign n10660 = n10563 ^ n10541 ;
  assign n10661 = n10660 ^ n10658 ;
  assign n10662 = n10659 & ~n10661 ;
  assign n10663 = n10662 ^ x398 ;
  assign n10664 = n10663 ^ n10608 ;
  assign n10665 = ~n10609 & n10664 ;
  assign n10666 = n10665 ^ x397 ;
  assign n10667 = n10666 ^ n10606 ;
  assign n10668 = ~n10607 & n10667 ;
  assign n10669 = n10668 ^ x396 ;
  assign n10670 = n10669 ^ n10604 ;
  assign n10671 = n10605 & ~n10670 ;
  assign n10672 = n10671 ^ x395 ;
  assign n10673 = n10672 ^ n10602 ;
  assign n10674 = ~n10603 & n10673 ;
  assign n10675 = n10674 ^ x394 ;
  assign n10676 = n10675 ^ n10600 ;
  assign n10677 = n10601 & ~n10676 ;
  assign n10678 = n10677 ^ x393 ;
  assign n10599 = n10574 ^ n10537 ;
  assign n10679 = n10678 ^ n10599 ;
  assign n10680 = n10597 ^ x392 ;
  assign n10681 = n10680 ^ n10597 ;
  assign n10682 = n10681 ^ n10599 ;
  assign n10683 = n10679 & ~n10682 ;
  assign n10684 = n10683 ^ n10680 ;
  assign n10685 = n10598 & ~n10684 ;
  assign n10686 = n10685 ^ x391 ;
  assign n10687 = n10686 ^ n10595 ;
  assign n10688 = n10596 & ~n10687 ;
  assign n10689 = n10688 ^ x390 ;
  assign n10690 = n10689 ^ n10593 ;
  assign n10691 = ~n10594 & n10690 ;
  assign n10692 = n10691 ^ x389 ;
  assign n10693 = n10692 ^ x388 ;
  assign n10694 = n10581 ^ n10580 ;
  assign n10695 = n10694 ^ n10692 ;
  assign n10696 = n10693 & n10695 ;
  assign n10697 = n10696 ^ x388 ;
  assign n10592 = n10584 ^ n10582 ;
  assign n10698 = n10697 ^ n10592 ;
  assign n10699 = n10697 ^ x387 ;
  assign n10700 = ~n10698 & n10699 ;
  assign n10701 = n10700 ^ x387 ;
  assign n10591 = n10586 ^ n10585 ;
  assign n10702 = n10701 ^ n10591 ;
  assign n10703 = n10701 ^ x386 ;
  assign n10704 = n10702 & n10703 ;
  assign n10705 = n10704 ^ x386 ;
  assign n10590 = n10589 ^ n10587 ;
  assign n10706 = n10705 ^ n10590 ;
  assign n10707 = n10705 ^ x385 ;
  assign n10708 = ~n10706 & n10707 ;
  assign n10723 = n10722 ^ n10708 ;
  assign n10416 = n10415 ^ n7401 ;
  assign n10532 = n10531 ^ n10415 ;
  assign n10533 = n10416 & ~n10532 ;
  assign n10724 = n10723 ^ n10533 ;
  assign n10728 = n10727 ^ n10724 ;
  assign n10751 = n8829 ^ n8807 ;
  assign n10752 = ~n10284 & n10751 ;
  assign n10753 = n10752 ^ n8829 ;
  assign n10759 = n10753 ^ n10727 ;
  assign n10748 = n10703 ^ n10591 ;
  assign n10754 = n10753 ^ n10748 ;
  assign n10734 = n10699 ^ n10592 ;
  assign n10729 = n10694 ^ n10693 ;
  assign n10730 = n8931 ^ n8826 ;
  assign n10731 = ~n10063 & ~n10730 ;
  assign n10732 = n10731 ^ n8931 ;
  assign n10733 = ~n10729 & n10732 ;
  assign n10735 = n10734 ^ n10733 ;
  assign n10736 = n10733 ^ n8926 ;
  assign n10737 = n10736 ^ n8820 ;
  assign n10738 = n10737 ^ n10733 ;
  assign n10739 = n10064 & ~n10738 ;
  assign n10740 = n10739 ^ n10736 ;
  assign n10741 = n10735 & n10740 ;
  assign n10742 = n10741 ^ n10734 ;
  assign n10743 = n10742 ^ n8835 ;
  assign n10744 = n10743 ^ n8813 ;
  assign n10745 = n10744 ^ n10742 ;
  assign n10746 = n10127 & n10745 ;
  assign n10747 = n10746 ^ n10743 ;
  assign n10749 = n10748 ^ n10742 ;
  assign n10750 = n10747 & ~n10749 ;
  assign n10755 = n10754 ^ n10750 ;
  assign n10756 = n10707 ^ n10590 ;
  assign n10757 = n10756 ^ n10753 ;
  assign n10758 = n10755 & ~n10757 ;
  assign n10760 = n10759 ^ n10758 ;
  assign n10761 = n10728 & n10760 ;
  assign n10763 = n10762 ^ n10761 ;
  assign n10764 = n10212 & n10763 ;
  assign n10765 = n10764 ^ n10211 ;
  assign n10766 = n10765 ^ n10203 ;
  assign n10767 = n10205 & ~n10766 ;
  assign n10768 = n10767 ^ n10204 ;
  assign n10769 = n10768 ^ n10194 ;
  assign n10770 = n10199 & n10769 ;
  assign n10771 = n10770 ^ n10194 ;
  assign n10773 = n10772 ^ n10771 ;
  assign n10774 = n9649 ^ n8244 ;
  assign n10775 = n10317 & ~n10774 ;
  assign n10776 = n10775 ^ n9649 ;
  assign n10777 = n10776 ^ n10771 ;
  assign n10778 = ~n10773 & ~n10777 ;
  assign n10779 = n10778 ^ n10772 ;
  assign n10780 = n10779 ^ n10190 ;
  assign n10781 = ~n10192 & ~n10780 ;
  assign n10782 = n10781 ^ n10191 ;
  assign n10783 = n10782 ^ n10181 ;
  assign n10784 = ~n10186 & ~n10783 ;
  assign n10785 = n10784 ^ n10185 ;
  assign n10786 = n10785 ^ n10177 ;
  assign n10787 = ~n10180 & ~n10786 ;
  assign n10788 = n10787 ^ n10179 ;
  assign n10857 = n10788 ^ n10167 ;
  assign n10858 = ~n10172 & n10857 ;
  assign n10859 = n10858 ^ n10167 ;
  assign n10853 = n9709 ^ n8883 ;
  assign n10854 = ~n10341 & n10853 ;
  assign n10855 = n10854 ^ n8883 ;
  assign n10957 = n10859 ^ n10855 ;
  assign n10852 = n10629 ^ n10626 ;
  assign n10958 = n10859 ^ n10852 ;
  assign n10959 = ~n10957 & ~n10958 ;
  assign n10960 = n10959 ^ n10855 ;
  assign n11035 = n10961 ^ n10960 ;
  assign n11036 = n10965 & ~n11035 ;
  assign n11037 = n11036 ^ n10964 ;
  assign n11033 = n10635 ^ n10622 ;
  assign n11038 = n11037 ^ n11033 ;
  assign n11039 = n11033 ^ n8872 ;
  assign n11040 = n11039 ^ n9630 ;
  assign n11041 = n11040 ^ n11033 ;
  assign n11042 = ~n10236 & ~n11041 ;
  assign n11043 = n11042 ^ n11039 ;
  assign n11044 = n11038 & ~n11043 ;
  assign n11034 = n11033 ^ n11031 ;
  assign n11045 = n11044 ^ n11034 ;
  assign n11046 = n11032 & ~n11045 ;
  assign n11047 = n11046 ^ n11031 ;
  assign n11049 = n11048 ^ n11047 ;
  assign n11050 = n11048 ^ n8857 ;
  assign n11051 = n11050 ^ n9612 ;
  assign n11052 = n11051 ^ n11048 ;
  assign n11053 = n10229 & ~n11052 ;
  assign n11054 = n11053 ^ n11050 ;
  assign n11055 = ~n11049 & ~n11054 ;
  assign n11056 = n11055 ^ n11048 ;
  assign n11057 = n11056 ^ n11022 ;
  assign n11058 = ~n11026 & n11057 ;
  assign n11059 = n11058 ^ n11025 ;
  assign n11060 = n11059 ^ n11018 ;
  assign n11061 = n11020 & n11060 ;
  assign n11062 = n11061 ^ n11019 ;
  assign n11013 = n10650 ^ x400 ;
  assign n11014 = n11013 ^ n10612 ;
  assign n11010 = n9609 ^ n9024 ;
  assign n11011 = n10383 & n11010 ;
  assign n11012 = n11011 ^ n9024 ;
  assign n11015 = n11014 ^ n11012 ;
  assign n11132 = n11062 ^ n11015 ;
  assign n11134 = n11132 ^ n8481 ;
  assign n11127 = n11059 ^ n11020 ;
  assign n11118 = n11054 ^ n11047 ;
  assign n11105 = n11043 ^ n11037 ;
  assign n11106 = n11105 ^ n8262 ;
  assign n10856 = n10855 ^ n10852 ;
  assign n10860 = n10859 ^ n10856 ;
  assign n10861 = n10860 ^ n8273 ;
  assign n10789 = n10788 ^ n10172 ;
  assign n10790 = n10789 ^ n8278 ;
  assign n10791 = n10785 ^ n10180 ;
  assign n10792 = n10791 ^ n8355 ;
  assign n10794 = n10779 ^ n10192 ;
  assign n10795 = n10794 ^ n8291 ;
  assign n10796 = n10776 ^ n10772 ;
  assign n10797 = n10796 ^ n10771 ;
  assign n10798 = n10797 ^ n8294 ;
  assign n10831 = n10768 ^ n10199 ;
  assign n10799 = n10765 ^ n10205 ;
  assign n10800 = n10799 ^ n8323 ;
  assign n10801 = n10763 ^ n10211 ;
  assign n10802 = n10801 ^ n8306 ;
  assign n10803 = n10732 ^ n10729 ;
  assign n10804 = n8095 & ~n10803 ;
  assign n10805 = n10804 ^ n8104 ;
  assign n10806 = n10740 ^ n10734 ;
  assign n10807 = n10806 ^ n10804 ;
  assign n10808 = n10805 & n10807 ;
  assign n10809 = n10808 ^ n8104 ;
  assign n10810 = n10809 ^ n8156 ;
  assign n10811 = n10748 ^ n10747 ;
  assign n10812 = n10811 ^ n10809 ;
  assign n10813 = n10810 & ~n10812 ;
  assign n10814 = n10813 ^ n8156 ;
  assign n10815 = n10814 ^ n8185 ;
  assign n10816 = n10756 ^ n10755 ;
  assign n10817 = n10816 ^ n10814 ;
  assign n10818 = n10815 & ~n10817 ;
  assign n10819 = n10818 ^ n8185 ;
  assign n10820 = n10819 ^ n8308 ;
  assign n10821 = n10760 ^ n10724 ;
  assign n10822 = n10821 ^ n10819 ;
  assign n10823 = n10820 & n10822 ;
  assign n10824 = n10823 ^ n8308 ;
  assign n10825 = n10824 ^ n10801 ;
  assign n10826 = n10802 & n10825 ;
  assign n10827 = n10826 ^ n8306 ;
  assign n10828 = n10827 ^ n10799 ;
  assign n10829 = ~n10800 & n10828 ;
  assign n10830 = n10829 ^ n8323 ;
  assign n10832 = n10831 ^ n10830 ;
  assign n10833 = n10831 ^ n8332 ;
  assign n10834 = n10832 & ~n10833 ;
  assign n10835 = n10834 ^ n8332 ;
  assign n10836 = n10835 ^ n10797 ;
  assign n10837 = ~n10798 & ~n10836 ;
  assign n10838 = n10837 ^ n8294 ;
  assign n10839 = n10838 ^ n10794 ;
  assign n10840 = n10795 & ~n10839 ;
  assign n10841 = n10840 ^ n8291 ;
  assign n10793 = n10782 ^ n10186 ;
  assign n10842 = n10841 ^ n10793 ;
  assign n10843 = n10841 ^ n8286 ;
  assign n10844 = n10842 & ~n10843 ;
  assign n10845 = n10844 ^ n8286 ;
  assign n10846 = n10845 ^ n10791 ;
  assign n10847 = n10792 & n10846 ;
  assign n10848 = n10847 ^ n8355 ;
  assign n10849 = n10848 ^ n10789 ;
  assign n10850 = ~n10790 & n10849 ;
  assign n10851 = n10850 ^ n8278 ;
  assign n10968 = n10860 ^ n10851 ;
  assign n10969 = n10861 & n10968 ;
  assign n10970 = n10969 ^ n8273 ;
  assign n10966 = n10965 ^ n10960 ;
  assign n11107 = n10970 ^ n10966 ;
  assign n11108 = n10970 ^ n8267 ;
  assign n11109 = ~n11107 & n11108 ;
  assign n11110 = n11109 ^ n8267 ;
  assign n11111 = n11110 ^ n11105 ;
  assign n11112 = ~n11106 & n11111 ;
  assign n11113 = n11112 ^ n8262 ;
  assign n11104 = n11045 ^ n11028 ;
  assign n11114 = n11113 ^ n11104 ;
  assign n11115 = n11113 ^ n8256 ;
  assign n11116 = ~n11114 & ~n11115 ;
  assign n11117 = n11116 ^ n8256 ;
  assign n11119 = n11118 ^ n11117 ;
  assign n11120 = n11118 ^ n8245 ;
  assign n11121 = n11119 & ~n11120 ;
  assign n11122 = n11121 ^ n8245 ;
  assign n11103 = n11056 ^ n11026 ;
  assign n11123 = n11122 ^ n11103 ;
  assign n11124 = n11122 ^ n8377 ;
  assign n11125 = ~n11123 & n11124 ;
  assign n11126 = n11125 ^ n8377 ;
  assign n11128 = n11127 ^ n11126 ;
  assign n11129 = n11127 ^ n8467 ;
  assign n11130 = n11128 & n11129 ;
  assign n11131 = n11130 ^ n8467 ;
  assign n11206 = n11134 ^ n11131 ;
  assign n11192 = n11126 ^ n8467 ;
  assign n11193 = n11192 ^ n11127 ;
  assign n11194 = n11103 ^ n8377 ;
  assign n11195 = n11194 ^ n11122 ;
  assign n11196 = n11120 ^ n11117 ;
  assign n11197 = n11104 ^ n8256 ;
  assign n11198 = n11197 ^ n11113 ;
  assign n11199 = n11110 ^ n11106 ;
  assign n10862 = n10861 ^ n10851 ;
  assign n10863 = n10845 ^ n10792 ;
  assign n10864 = n10793 ^ n8286 ;
  assign n10865 = n10864 ^ n10841 ;
  assign n10866 = n10827 ^ n10800 ;
  assign n10867 = n10821 ^ n10820 ;
  assign n10868 = n10803 ^ n8095 ;
  assign n10869 = n10806 ^ n10805 ;
  assign n10870 = ~n10868 & ~n10869 ;
  assign n10871 = n10811 ^ n10810 ;
  assign n10872 = n10870 & n10871 ;
  assign n10873 = n10816 ^ n10815 ;
  assign n10874 = ~n10872 & ~n10873 ;
  assign n10875 = n10867 & n10874 ;
  assign n10876 = n10824 ^ n8306 ;
  assign n10877 = n10876 ^ n10801 ;
  assign n10878 = ~n10875 & n10877 ;
  assign n10879 = n10866 & n10878 ;
  assign n10880 = n10833 ^ n10830 ;
  assign n10881 = ~n10879 & ~n10880 ;
  assign n10882 = n10835 ^ n10798 ;
  assign n10883 = n10881 & ~n10882 ;
  assign n10884 = n10838 ^ n10795 ;
  assign n10885 = ~n10883 & n10884 ;
  assign n10886 = n10865 & n10885 ;
  assign n10887 = n10863 & ~n10886 ;
  assign n10888 = n10848 ^ n10790 ;
  assign n10889 = n10887 & n10888 ;
  assign n10956 = ~n10862 & n10889 ;
  assign n10967 = n10966 ^ n8267 ;
  assign n10971 = n10970 ^ n10967 ;
  assign n11200 = n10956 & n10971 ;
  assign n11201 = n11199 & ~n11200 ;
  assign n11202 = n11198 & n11201 ;
  assign n11203 = n11196 & ~n11202 ;
  assign n11204 = n11195 & ~n11203 ;
  assign n11205 = n11193 & n11204 ;
  assign n11268 = n11206 ^ n11205 ;
  assign n11269 = n11268 ^ x427 ;
  assign n11270 = n11203 ^ n11195 ;
  assign n11271 = n11270 ^ x429 ;
  assign n11272 = n11201 ^ n11198 ;
  assign n11273 = n11272 ^ x431 ;
  assign n10972 = n10971 ^ n10956 ;
  assign n10973 = n10972 ^ x433 ;
  assign n10890 = n10889 ^ n10862 ;
  assign n10891 = n10890 ^ x434 ;
  assign n10892 = n10888 ^ n10887 ;
  assign n10893 = n10892 ^ x435 ;
  assign n10894 = n10885 ^ n10865 ;
  assign n10895 = n10894 ^ x437 ;
  assign n10896 = n10884 ^ n10883 ;
  assign n10897 = n10896 ^ x438 ;
  assign n10898 = n10882 ^ n10881 ;
  assign n10899 = n10898 ^ x439 ;
  assign n10901 = n10878 ^ n10866 ;
  assign n10902 = n10901 ^ x441 ;
  assign n10903 = n10877 ^ n10875 ;
  assign n10904 = n10903 ^ x442 ;
  assign n10905 = n10874 ^ n10867 ;
  assign n10906 = n10905 ^ x443 ;
  assign n10907 = n10873 ^ n10872 ;
  assign n10908 = n10907 ^ x444 ;
  assign n10915 = n10871 ^ n10870 ;
  assign n10909 = x447 & n10868 ;
  assign n10910 = n10909 ^ x446 ;
  assign n10911 = n10869 ^ n10868 ;
  assign n10912 = n10911 ^ n10909 ;
  assign n10913 = n10910 & ~n10912 ;
  assign n10914 = n10913 ^ x446 ;
  assign n10916 = n10915 ^ n10914 ;
  assign n10917 = n10915 ^ x445 ;
  assign n10918 = ~n10916 & n10917 ;
  assign n10919 = n10918 ^ x445 ;
  assign n10920 = n10919 ^ n10907 ;
  assign n10921 = ~n10908 & n10920 ;
  assign n10922 = n10921 ^ x444 ;
  assign n10923 = n10922 ^ n10905 ;
  assign n10924 = ~n10906 & n10923 ;
  assign n10925 = n10924 ^ x443 ;
  assign n10926 = n10925 ^ n10903 ;
  assign n10927 = ~n10904 & n10926 ;
  assign n10928 = n10927 ^ x442 ;
  assign n10929 = n10928 ^ n10901 ;
  assign n10930 = n10902 & ~n10929 ;
  assign n10931 = n10930 ^ x441 ;
  assign n10900 = n10880 ^ n10879 ;
  assign n10932 = n10931 ^ n10900 ;
  assign n10933 = n10931 ^ x440 ;
  assign n10934 = n10932 & n10933 ;
  assign n10935 = n10934 ^ x440 ;
  assign n10936 = n10935 ^ n10898 ;
  assign n10937 = n10899 & ~n10936 ;
  assign n10938 = n10937 ^ x439 ;
  assign n10939 = n10938 ^ n10896 ;
  assign n10940 = ~n10897 & n10939 ;
  assign n10941 = n10940 ^ x438 ;
  assign n10942 = n10941 ^ n10894 ;
  assign n10943 = n10895 & ~n10942 ;
  assign n10944 = n10943 ^ x437 ;
  assign n10945 = n10944 ^ x436 ;
  assign n10946 = n10886 ^ n10863 ;
  assign n10947 = n10946 ^ n10944 ;
  assign n10948 = n10945 & ~n10947 ;
  assign n10949 = n10948 ^ x436 ;
  assign n10950 = n10949 ^ n10892 ;
  assign n10951 = ~n10893 & n10950 ;
  assign n10952 = n10951 ^ x435 ;
  assign n10953 = n10952 ^ n10890 ;
  assign n10954 = n10891 & ~n10953 ;
  assign n10955 = n10954 ^ x434 ;
  assign n11275 = n10972 ^ n10955 ;
  assign n11276 = ~n10973 & n11275 ;
  assign n11277 = n11276 ^ x433 ;
  assign n11274 = n11200 ^ n11199 ;
  assign n11278 = n11277 ^ n11274 ;
  assign n11279 = n11272 ^ x432 ;
  assign n11280 = n11279 ^ n11272 ;
  assign n11281 = n11280 ^ n11274 ;
  assign n11282 = n11278 & ~n11281 ;
  assign n11283 = n11282 ^ n11279 ;
  assign n11284 = n11273 & ~n11283 ;
  assign n11285 = n11284 ^ x431 ;
  assign n11286 = n11285 ^ x430 ;
  assign n11287 = n11202 ^ n11196 ;
  assign n11288 = n11287 ^ n11285 ;
  assign n11289 = n11286 & ~n11288 ;
  assign n11290 = n11289 ^ x430 ;
  assign n11291 = n11290 ^ n11270 ;
  assign n11292 = ~n11271 & n11291 ;
  assign n11293 = n11292 ^ x429 ;
  assign n11294 = n11293 ^ x428 ;
  assign n11295 = n11204 ^ n11193 ;
  assign n11296 = n11295 ^ n11293 ;
  assign n11297 = n11294 & ~n11296 ;
  assign n11298 = n11297 ^ x428 ;
  assign n11299 = n11298 ^ n11268 ;
  assign n11300 = ~n11269 & n11299 ;
  assign n11301 = n11300 ^ x427 ;
  assign n11712 = n11301 ^ x426 ;
  assign n11133 = n11132 ^ n11131 ;
  assign n11135 = ~n11133 & n11134 ;
  assign n11136 = n11135 ^ n8481 ;
  assign n11063 = n11062 ^ n11012 ;
  assign n11064 = ~n11015 & ~n11063 ;
  assign n11065 = n11064 ^ n11014 ;
  assign n10975 = n10656 ^ x399 ;
  assign n11002 = n10975 ^ n9034 ;
  assign n11003 = n11002 ^ n9752 ;
  assign n11004 = n11003 ^ n10975 ;
  assign n11005 = n10388 & n11004 ;
  assign n11006 = n11005 ^ n11002 ;
  assign n11101 = n11065 ^ n11006 ;
  assign n11102 = n11101 ^ n8497 ;
  assign n11208 = n11136 ^ n11102 ;
  assign n11207 = n11205 & ~n11206 ;
  assign n11266 = n11208 ^ n11207 ;
  assign n11713 = n11712 ^ n11266 ;
  assign n11226 = n10684 ^ x391 ;
  assign n11571 = n11295 ^ n11294 ;
  assign n11572 = n11571 ^ n10046 ;
  assign n11573 = n11572 ^ n10711 ;
  assign n11574 = n11573 ^ n11571 ;
  assign n11575 = n11226 & ~n11574 ;
  assign n11576 = n11575 ^ n11572 ;
  assign n11585 = n11290 ^ n11271 ;
  assign n11185 = n10678 ^ x392 ;
  assign n11186 = n11185 ^ n10599 ;
  assign n11582 = n10413 ^ n9985 ;
  assign n11583 = ~n11186 & ~n11582 ;
  assign n11584 = n11583 ^ n9985 ;
  assign n11586 = n11585 ^ n11584 ;
  assign n11593 = n11287 ^ n11286 ;
  assign n11693 = n11593 ^ n11584 ;
  assign n11095 = n10672 ^ x394 ;
  assign n11096 = n11095 ^ n10602 ;
  assign n11587 = n11283 ^ x431 ;
  assign n11588 = n11587 ^ n9752 ;
  assign n11589 = n11588 ^ n10402 ;
  assign n11590 = n11589 ^ n11587 ;
  assign n11591 = ~n11096 & ~n11590 ;
  assign n11592 = n11591 ^ n11588 ;
  assign n11684 = n11593 ^ n11587 ;
  assign n11597 = n11277 ^ x432 ;
  assign n11598 = n11597 ^ n11274 ;
  assign n10996 = n10669 ^ n10605 ;
  assign n11594 = n10218 ^ n9609 ;
  assign n11595 = n10996 & n11594 ;
  assign n11596 = n11595 ^ n9609 ;
  assign n11599 = n11598 ^ n11596 ;
  assign n11606 = n10952 ^ x434 ;
  assign n11607 = n11606 ^ n10890 ;
  assign n10997 = n10663 ^ n10609 ;
  assign n11603 = n10383 ^ n9730 ;
  assign n11604 = ~n10997 & ~n11603 ;
  assign n11605 = n11604 ^ n9730 ;
  assign n11608 = n11607 ^ n11605 ;
  assign n11612 = n10949 ^ n10893 ;
  assign n11007 = n10660 ^ n10659 ;
  assign n11609 = n10223 ^ n9612 ;
  assign n11610 = n11007 & ~n11609 ;
  assign n11611 = n11610 ^ n9612 ;
  assign n11613 = n11612 ^ n11611 ;
  assign n11614 = n10227 ^ n9627 ;
  assign n11615 = ~n10975 & n11614 ;
  assign n11616 = n11615 ^ n9627 ;
  assign n11533 = n10946 ^ n10945 ;
  assign n11617 = n11616 ^ n11533 ;
  assign n11651 = n10350 ^ n9635 ;
  assign n11652 = n11019 & ~n11651 ;
  assign n11653 = n11652 ^ n9635 ;
  assign n11618 = n10236 ^ n9709 ;
  assign n11619 = n11022 & n11618 ;
  assign n11620 = n11619 ^ n9709 ;
  assign n11546 = n10935 ^ n10899 ;
  assign n11621 = n11620 ^ n11546 ;
  assign n11622 = n10341 ^ n9701 ;
  assign n11623 = n11028 & n11622 ;
  assign n11624 = n11623 ^ n9701 ;
  assign n11557 = n10928 ^ n10902 ;
  assign n11625 = n11624 ^ n11557 ;
  assign n11521 = n10174 ^ n9679 ;
  assign n11522 = ~n10961 & ~n11521 ;
  assign n11523 = n11522 ^ n9679 ;
  assign n11520 = n10922 ^ n10906 ;
  assign n11524 = n11523 ^ n11520 ;
  assign n11452 = n10919 ^ x444 ;
  assign n11453 = n11452 ^ n10907 ;
  assign n11449 = n10182 ^ n9649 ;
  assign n11450 = n10852 & ~n11449 ;
  assign n11451 = n11450 ^ n9649 ;
  assign n11454 = n11453 ^ n11451 ;
  assign n11407 = n10917 ^ n10914 ;
  assign n11404 = n10187 ^ n9654 ;
  assign n11405 = n10167 & ~n11404 ;
  assign n11406 = n11405 ^ n9654 ;
  assign n11408 = n11407 ^ n11406 ;
  assign n10982 = n10911 ^ n10910 ;
  assign n10979 = n10317 ^ n9661 ;
  assign n10980 = n10179 & ~n10979 ;
  assign n10981 = n10980 ^ n9661 ;
  assign n10983 = n10982 ^ n10981 ;
  assign n10985 = n10193 ^ n9538 ;
  assign n10986 = n10181 & ~n10985 ;
  assign n10987 = n10986 ^ n9538 ;
  assign n10984 = n10868 ^ x447 ;
  assign n10988 = n10987 ^ n10984 ;
  assign n10989 = n10666 ^ x396 ;
  assign n10990 = n10989 ^ n10606 ;
  assign n10991 = n10990 ^ n9366 ;
  assign n10992 = n10991 ^ n10046 ;
  assign n10993 = n10992 ^ n10990 ;
  assign n10994 = ~n10216 & ~n10993 ;
  assign n10995 = n10994 ^ n10991 ;
  assign n11080 = n10996 ^ n10990 ;
  assign n10998 = n9985 ^ n9045 ;
  assign n10999 = ~n10402 & n10998 ;
  assign n11000 = n10999 ^ n9045 ;
  assign n11001 = n11000 ^ n10997 ;
  assign n11008 = n11007 ^ n10975 ;
  assign n11009 = n11008 ^ n11007 ;
  assign n11066 = n11065 ^ n11009 ;
  assign n11067 = ~n11006 & n11066 ;
  assign n11068 = n11067 ^ n11008 ;
  assign n11073 = n11007 ^ n11000 ;
  assign n11069 = n9842 ^ n9035 ;
  assign n11070 = n10218 & ~n11069 ;
  assign n11071 = n11070 ^ n9035 ;
  assign n11072 = n11071 ^ n11000 ;
  assign n11074 = n11073 ^ n11072 ;
  assign n11075 = ~n11068 & n11074 ;
  assign n11076 = n11075 ^ n11073 ;
  assign n11077 = n11001 & ~n11076 ;
  assign n11078 = n11077 ^ n11000 ;
  assign n11079 = n11078 ^ n10996 ;
  assign n11081 = n11080 ^ n11079 ;
  assign n11082 = n10995 & n11081 ;
  assign n11083 = n11082 ^ n11079 ;
  assign n11084 = n9398 ^ n8691 ;
  assign n11085 = n10711 & ~n11084 ;
  assign n11086 = n11085 ^ n8691 ;
  assign n11091 = n11086 ^ n10996 ;
  assign n11087 = n9393 ^ n8696 ;
  assign n11088 = n10413 & n11087 ;
  assign n11089 = n11088 ^ n8696 ;
  assign n11090 = n11089 ^ n11086 ;
  assign n11092 = n11091 ^ n11090 ;
  assign n11093 = ~n11083 & ~n11092 ;
  assign n11094 = n11093 ^ n11091 ;
  assign n11161 = n11096 ^ n11086 ;
  assign n11162 = ~n11094 & n11161 ;
  assign n11163 = n11162 ^ n11086 ;
  assign n11164 = n11163 ^ n8684 ;
  assign n11165 = n11164 ^ n9386 ;
  assign n11166 = n11165 ^ n11163 ;
  assign n11167 = ~n10013 & n11166 ;
  assign n11168 = n11167 ^ n11164 ;
  assign n11177 = n9384 ^ n8683 ;
  assign n11178 = ~n10018 & ~n11177 ;
  assign n11179 = n11178 ^ n8683 ;
  assign n11169 = n10675 ^ x393 ;
  assign n11170 = n11169 ^ n10600 ;
  assign n11181 = n11179 ^ n11170 ;
  assign n11180 = n11179 ^ n11163 ;
  assign n11182 = n11181 ^ n11180 ;
  assign n11183 = n11168 & ~n11182 ;
  assign n11184 = n11183 ^ n11180 ;
  assign n11228 = n11226 ^ n11186 ;
  assign n11227 = n11226 ^ n11179 ;
  assign n11229 = n11228 ^ n11227 ;
  assign n11230 = ~n11184 & ~n11229 ;
  assign n11231 = n11230 ^ n11227 ;
  assign n11240 = n10686 ^ x390 ;
  assign n11241 = n11240 ^ n10595 ;
  assign n11242 = n11241 ^ n11226 ;
  assign n11243 = n11242 ^ n11241 ;
  assign n11223 = n9379 ^ n8737 ;
  assign n11224 = n10008 & ~n11223 ;
  assign n11225 = n11224 ^ n9379 ;
  assign n11244 = n11243 ^ n11225 ;
  assign n11245 = n11231 & n11244 ;
  assign n11246 = n11245 ^ n11242 ;
  assign n11247 = n8833 ^ n8770 ;
  assign n11248 = ~n9997 & n11247 ;
  assign n11249 = n11248 ^ n8770 ;
  assign n11389 = n11249 ^ n11241 ;
  assign n11390 = ~n11246 & n11389 ;
  assign n11386 = n9423 ^ n8936 ;
  assign n11387 = n10057 & ~n11386 ;
  assign n11382 = n11249 ^ n10716 ;
  assign n11381 = n10689 ^ n10594 ;
  assign n11383 = n11382 ^ n11381 ;
  assign n11384 = n11383 ^ n7332 ;
  assign n11380 = x417 ^ x416 ;
  assign n11385 = n11384 ^ n11380 ;
  assign n11388 = n11387 ^ n11385 ;
  assign n11391 = n11390 ^ n11388 ;
  assign n11187 = n11186 ^ n11184 ;
  assign n11171 = n11170 ^ n11168 ;
  assign n11098 = n11089 ^ n11083 ;
  assign n11099 = n11098 ^ n7955 ;
  assign n11140 = n11071 ^ n11068 ;
  assign n11137 = n11136 ^ n11101 ;
  assign n11138 = ~n11102 & n11137 ;
  assign n11139 = n11138 ^ n8497 ;
  assign n11141 = n11140 ^ n11139 ;
  assign n11142 = n11140 ^ n8546 ;
  assign n11143 = ~n11141 & n11142 ;
  assign n11144 = n11143 ^ n8546 ;
  assign n11145 = n11144 ^ n8564 ;
  assign n11146 = n11076 ^ n10997 ;
  assign n11147 = n11146 ^ n11144 ;
  assign n11148 = ~n11145 & n11147 ;
  assign n11149 = n11148 ^ n8564 ;
  assign n11100 = n11078 ^ n10995 ;
  assign n11150 = n11149 ^ n11100 ;
  assign n11151 = n11149 ^ n8722 ;
  assign n11152 = ~n11150 & ~n11151 ;
  assign n11153 = n11152 ^ n8722 ;
  assign n11154 = n11153 ^ n11098 ;
  assign n11155 = ~n11099 & n11154 ;
  assign n11156 = n11155 ^ n7955 ;
  assign n11097 = n11096 ^ n11094 ;
  assign n11157 = n11156 ^ n11097 ;
  assign n11158 = n11156 ^ n7992 ;
  assign n11159 = n11157 & ~n11158 ;
  assign n11160 = n11159 ^ n7992 ;
  assign n11172 = n11171 ^ n11160 ;
  assign n11173 = n11171 ^ n8021 ;
  assign n11174 = ~n11172 & n11173 ;
  assign n11175 = n11174 ^ n8021 ;
  assign n11176 = n11175 ^ n8055 ;
  assign n11188 = n11187 ^ n11176 ;
  assign n11189 = n11160 ^ n8021 ;
  assign n11190 = n11189 ^ n11171 ;
  assign n11191 = n11146 ^ n11145 ;
  assign n11209 = n11207 & n11208 ;
  assign n11210 = n11142 ^ n11139 ;
  assign n11211 = n11209 & ~n11210 ;
  assign n11212 = n11191 & ~n11211 ;
  assign n11213 = n11100 ^ n8722 ;
  assign n11214 = n11213 ^ n11149 ;
  assign n11215 = ~n11212 & ~n11214 ;
  assign n11216 = n11153 ^ n11099 ;
  assign n11217 = ~n11215 & ~n11216 ;
  assign n11218 = n11097 ^ n7992 ;
  assign n11219 = n11218 ^ n11156 ;
  assign n11220 = ~n11217 & ~n11219 ;
  assign n11221 = ~n11190 & ~n11220 ;
  assign n11222 = n11188 & n11221 ;
  assign n11233 = n11187 ^ n11175 ;
  assign n11234 = n11187 ^ n8055 ;
  assign n11235 = ~n11233 & ~n11234 ;
  assign n11236 = n11235 ^ n8055 ;
  assign n11237 = n11236 ^ n8079 ;
  assign n11232 = n11231 ^ n11225 ;
  assign n11238 = n11237 ^ n11232 ;
  assign n11239 = ~n11222 & n11238 ;
  assign n11251 = n11236 ^ n11232 ;
  assign n11252 = n11232 ^ n8079 ;
  assign n11253 = n11251 & ~n11252 ;
  assign n11254 = n11253 ^ n8079 ;
  assign n11255 = n11254 ^ n7332 ;
  assign n11250 = n11249 ^ n11246 ;
  assign n11256 = n11255 ^ n11250 ;
  assign n11379 = ~n11239 & n11256 ;
  assign n11392 = n11391 ^ n11379 ;
  assign n11258 = n11219 ^ n11217 ;
  assign n11259 = n11258 ^ x421 ;
  assign n11260 = n11216 ^ n11215 ;
  assign n11261 = n11260 ^ x422 ;
  assign n11262 = n11214 ^ n11212 ;
  assign n11263 = n11262 ^ x423 ;
  assign n11264 = n11210 ^ n11209 ;
  assign n11265 = n11264 ^ x425 ;
  assign n11267 = n11266 ^ x426 ;
  assign n11302 = n11301 ^ n11266 ;
  assign n11303 = n11267 & ~n11302 ;
  assign n11304 = n11303 ^ x426 ;
  assign n11305 = n11304 ^ n11264 ;
  assign n11306 = ~n11265 & n11305 ;
  assign n11307 = n11306 ^ x425 ;
  assign n11308 = n11307 ^ x424 ;
  assign n11309 = n11211 ^ n11191 ;
  assign n11310 = n11309 ^ n11307 ;
  assign n11311 = n11308 & ~n11310 ;
  assign n11312 = n11311 ^ x424 ;
  assign n11313 = n11312 ^ n11262 ;
  assign n11314 = n11263 & ~n11313 ;
  assign n11315 = n11314 ^ x423 ;
  assign n11316 = n11315 ^ n11260 ;
  assign n11317 = ~n11261 & n11316 ;
  assign n11318 = n11317 ^ x422 ;
  assign n11319 = n11318 ^ n11258 ;
  assign n11320 = n11259 & ~n11319 ;
  assign n11321 = n11320 ^ x421 ;
  assign n11322 = n11321 ^ x420 ;
  assign n11323 = n11220 ^ n11190 ;
  assign n11324 = n11323 ^ n11321 ;
  assign n11325 = n11322 & n11324 ;
  assign n11326 = n11325 ^ x420 ;
  assign n11327 = n11326 ^ x419 ;
  assign n11328 = n11221 ^ n11188 ;
  assign n11329 = n11328 ^ n11326 ;
  assign n11330 = n11327 & n11329 ;
  assign n11331 = n11330 ^ x419 ;
  assign n11332 = n11331 ^ x418 ;
  assign n11333 = n11238 ^ n11222 ;
  assign n11334 = n11333 ^ n11331 ;
  assign n11335 = n11332 & n11334 ;
  assign n11336 = n11335 ^ x418 ;
  assign n11337 = n11336 ^ x417 ;
  assign n11257 = n11256 ^ n11239 ;
  assign n11377 = n11336 ^ n11257 ;
  assign n11378 = n11337 & ~n11377 ;
  assign n11393 = n11392 ^ n11378 ;
  assign n11375 = n11254 ^ n11250 ;
  assign n11376 = ~n11255 & n11375 ;
  assign n11394 = n11393 ^ n11376 ;
  assign n11397 = n11394 ^ n10987 ;
  assign n11340 = n11323 ^ n11322 ;
  assign n11341 = n10127 ^ n8826 ;
  assign n11342 = n10211 & ~n11341 ;
  assign n11343 = n11342 ^ n8826 ;
  assign n11344 = ~n11340 & ~n11343 ;
  assign n11339 = n11328 ^ n11327 ;
  assign n11345 = n11344 ^ n11339 ;
  assign n11346 = n11344 ^ n8820 ;
  assign n11347 = n11346 ^ n10284 ;
  assign n11348 = n11347 ^ n11344 ;
  assign n11349 = n10204 & ~n11348 ;
  assign n11350 = n11349 ^ n11346 ;
  assign n11351 = ~n11345 & n11350 ;
  assign n11352 = n11351 ^ n11344 ;
  assign n11353 = n11352 ^ n8813 ;
  assign n11354 = n11353 ^ n10301 ;
  assign n11355 = n11354 ^ n11352 ;
  assign n11356 = n10194 & n11355 ;
  assign n11357 = n11356 ^ n11353 ;
  assign n11358 = n11333 ^ n11332 ;
  assign n11359 = n11358 ^ n11352 ;
  assign n11360 = n11357 & ~n11359 ;
  assign n11361 = n11360 ^ n11358 ;
  assign n11338 = n11337 ^ n11257 ;
  assign n11362 = n11361 ^ n11338 ;
  assign n11363 = n11361 ^ n8807 ;
  assign n11364 = n11363 ^ n10207 ;
  assign n11365 = n11364 ^ n11361 ;
  assign n11366 = ~n10772 & ~n11365 ;
  assign n11367 = n11366 ^ n11363 ;
  assign n11368 = ~n11362 & n11367 ;
  assign n11369 = n11368 ^ n11361 ;
  assign n11370 = n11369 ^ n9449 ;
  assign n11371 = n11370 ^ n10200 ;
  assign n11372 = n11371 ^ n11369 ;
  assign n11373 = n10191 & n11372 ;
  assign n11374 = n11373 ^ n11370 ;
  assign n11395 = n11394 ^ n11369 ;
  assign n11396 = ~n11374 & ~n11395 ;
  assign n11398 = n11397 ^ n11396 ;
  assign n11399 = ~n10988 & ~n11398 ;
  assign n11400 = n11399 ^ n10987 ;
  assign n11401 = n11400 ^ n10981 ;
  assign n11402 = n10983 & n11401 ;
  assign n11403 = n11402 ^ n10982 ;
  assign n11446 = n11406 ^ n11403 ;
  assign n11447 = ~n11408 & n11446 ;
  assign n11448 = n11447 ^ n11407 ;
  assign n11517 = n11451 ^ n11448 ;
  assign n11518 = ~n11454 & ~n11517 ;
  assign n11519 = n11518 ^ n11453 ;
  assign n11626 = n11520 ^ n11519 ;
  assign n11627 = ~n11524 & ~n11626 ;
  assign n11628 = n11627 ^ n11523 ;
  assign n11564 = n10925 ^ x442 ;
  assign n11565 = n11564 ^ n10903 ;
  assign n11629 = n11628 ^ n11565 ;
  assign n11630 = n11565 ^ n9692 ;
  assign n11631 = n11630 ^ n9605 ;
  assign n11632 = n11631 ^ n11565 ;
  assign n11633 = ~n11033 & n11632 ;
  assign n11634 = n11633 ^ n11630 ;
  assign n11635 = ~n11629 & n11634 ;
  assign n11636 = n11635 ^ n11565 ;
  assign n11637 = n11636 ^ n11557 ;
  assign n11638 = ~n11625 & n11637 ;
  assign n11639 = n11638 ^ n11624 ;
  assign n11553 = n10933 ^ n10900 ;
  assign n11640 = n11639 ^ n11553 ;
  assign n11641 = n11553 ^ n9638 ;
  assign n11642 = n11641 ^ n10245 ;
  assign n11643 = n11642 ^ n11553 ;
  assign n11644 = ~n11048 & n11643 ;
  assign n11645 = n11644 ^ n11641 ;
  assign n11646 = n11640 & n11645 ;
  assign n11647 = n11646 ^ n11553 ;
  assign n11648 = n11647 ^ n11546 ;
  assign n11649 = ~n11621 & n11648 ;
  assign n11650 = n11649 ^ n11620 ;
  assign n11654 = n11653 ^ n11650 ;
  assign n11655 = n10938 ^ n10897 ;
  assign n11656 = n11655 ^ n11653 ;
  assign n11657 = ~n11654 & n11656 ;
  assign n11658 = n11657 ^ n11655 ;
  assign n11539 = n10941 ^ n10895 ;
  assign n11659 = n11658 ^ n11539 ;
  assign n11660 = n11539 ^ n9630 ;
  assign n11661 = n11660 ^ n10229 ;
  assign n11662 = n11661 ^ n11539 ;
  assign n11663 = ~n11014 & ~n11662 ;
  assign n11664 = n11663 ^ n11660 ;
  assign n11665 = ~n11659 & n11664 ;
  assign n11666 = n11665 ^ n11658 ;
  assign n11667 = n11666 ^ n11616 ;
  assign n11668 = n11617 & n11667 ;
  assign n11669 = n11668 ^ n11533 ;
  assign n11670 = n11669 ^ n11611 ;
  assign n11671 = n11613 & n11670 ;
  assign n11672 = n11671 ^ n11612 ;
  assign n11673 = n11672 ^ n11605 ;
  assign n11674 = ~n11608 & ~n11673 ;
  assign n11675 = n11674 ^ n11607 ;
  assign n11600 = n10388 ^ n9739 ;
  assign n11601 = n10990 & ~n11600 ;
  assign n11602 = n11601 ^ n10388 ;
  assign n11676 = n11675 ^ n11602 ;
  assign n10974 = n10973 ^ n10955 ;
  assign n11677 = n11675 ^ n10974 ;
  assign n11678 = ~n11676 & ~n11677 ;
  assign n11679 = n11678 ^ n10974 ;
  assign n11680 = n11679 ^ n11596 ;
  assign n11681 = ~n11599 & n11680 ;
  assign n11682 = n11681 ^ n11598 ;
  assign n11683 = n11682 ^ n11593 ;
  assign n11685 = n11684 ^ n11683 ;
  assign n11686 = n11592 & ~n11685 ;
  assign n11687 = n11686 ^ n11684 ;
  assign n11688 = n10216 ^ n9842 ;
  assign n11689 = n11170 & n11688 ;
  assign n11690 = n11689 ^ n9842 ;
  assign n11691 = n11690 ^ n11593 ;
  assign n11692 = n11687 & ~n11691 ;
  assign n11694 = n11693 ^ n11692 ;
  assign n11695 = n11586 & n11694 ;
  assign n11696 = n11695 ^ n11585 ;
  assign n11577 = n10013 ^ n9393 ;
  assign n11578 = n11241 & n11577 ;
  assign n11579 = n11578 ^ n9393 ;
  assign n11580 = n11579 ^ n11571 ;
  assign n11581 = n11580 ^ n11579 ;
  assign n11697 = n11696 ^ n11581 ;
  assign n11698 = ~n11576 & ~n11697 ;
  assign n11699 = n11698 ^ n11580 ;
  assign n11700 = n10018 ^ n9398 ;
  assign n11701 = ~n11381 & ~n11700 ;
  assign n11702 = n11701 ^ n9398 ;
  assign n11705 = n11702 ^ n11579 ;
  assign n11703 = n11298 ^ n11269 ;
  assign n11704 = n11703 ^ n11702 ;
  assign n11706 = n11705 ^ n11704 ;
  assign n11707 = n11699 & n11706 ;
  assign n11708 = n11707 ^ n11704 ;
  assign n11722 = n11713 ^ n11708 ;
  assign n11723 = n11722 ^ n8691 ;
  assign n11803 = n11703 ^ n11699 ;
  assign n11724 = n11696 ^ n11576 ;
  assign n11725 = n11724 ^ n9366 ;
  assign n11727 = n11690 ^ n11687 ;
  assign n11728 = n11727 ^ n9035 ;
  assign n11788 = n11682 ^ n11592 ;
  assign n11729 = n11679 ^ n11599 ;
  assign n11730 = n11729 ^ n9024 ;
  assign n11731 = n11602 ^ n10974 ;
  assign n11732 = n11731 ^ n11675 ;
  assign n11733 = n11732 ^ n8840 ;
  assign n11773 = n11669 ^ n11613 ;
  assign n11735 = n11666 ^ n11617 ;
  assign n11736 = n11735 ^ n8866 ;
  assign n11737 = n11664 ^ n11658 ;
  assign n11738 = n11737 ^ n8872 ;
  assign n11739 = n11656 ^ n11650 ;
  assign n11740 = n11739 ^ n8877 ;
  assign n11741 = n11647 ^ n11621 ;
  assign n11742 = n11741 ^ n8883 ;
  assign n11743 = n11645 ^ n11639 ;
  assign n11744 = n11743 ^ n8888 ;
  assign n11745 = n11636 ^ n11625 ;
  assign n11746 = n11745 ^ n8990 ;
  assign n11525 = n11524 ^ n11519 ;
  assign n11526 = n11525 ^ n8893 ;
  assign n11455 = n11454 ^ n11448 ;
  assign n11456 = n11455 ^ n8244 ;
  assign n11409 = n11408 ^ n11403 ;
  assign n11410 = n11409 ^ n8815 ;
  assign n11411 = n11400 ^ n10983 ;
  assign n11412 = n11411 ^ n8962 ;
  assign n11435 = n11398 ^ n10984 ;
  assign n11413 = n11394 ^ n11374 ;
  assign n11414 = n11413 ^ n8908 ;
  assign n11427 = n11367 ^ n11338 ;
  assign n11415 = n11343 ^ n11340 ;
  assign n11416 = n8931 & n11415 ;
  assign n11417 = n11416 ^ n8926 ;
  assign n11418 = n11350 ^ n11339 ;
  assign n11419 = n11418 ^ n11416 ;
  assign n11420 = ~n11417 & n11419 ;
  assign n11421 = n11420 ^ n8926 ;
  assign n11422 = n11421 ^ n8835 ;
  assign n11423 = n11358 ^ n11357 ;
  assign n11424 = n11423 ^ n11421 ;
  assign n11425 = n11422 & n11424 ;
  assign n11426 = n11425 ^ n8835 ;
  assign n11428 = n11427 ^ n11426 ;
  assign n11429 = n11427 ^ n8829 ;
  assign n11430 = n11428 & ~n11429 ;
  assign n11431 = n11430 ^ n8829 ;
  assign n11432 = n11431 ^ n11413 ;
  assign n11433 = ~n11414 & n11432 ;
  assign n11434 = n11433 ^ n8908 ;
  assign n11436 = n11435 ^ n11434 ;
  assign n11437 = n11435 ^ n8822 ;
  assign n11438 = ~n11436 & ~n11437 ;
  assign n11439 = n11438 ^ n8822 ;
  assign n11440 = n11439 ^ n11411 ;
  assign n11441 = ~n11412 & n11440 ;
  assign n11442 = n11441 ^ n8962 ;
  assign n11443 = n11442 ^ n11409 ;
  assign n11444 = ~n11410 & n11443 ;
  assign n11445 = n11444 ^ n8815 ;
  assign n11514 = n11455 ^ n11445 ;
  assign n11515 = n11456 & n11514 ;
  assign n11516 = n11515 ^ n8244 ;
  assign n11748 = n11525 ^ n11516 ;
  assign n11749 = ~n11526 & n11748 ;
  assign n11750 = n11749 ^ n8893 ;
  assign n11747 = n11634 ^ n11628 ;
  assign n11751 = n11750 ^ n11747 ;
  assign n11752 = n11750 ^ n8980 ;
  assign n11753 = n11751 & n11752 ;
  assign n11754 = n11753 ^ n8980 ;
  assign n11755 = n11754 ^ n11745 ;
  assign n11756 = n11746 & n11755 ;
  assign n11757 = n11756 ^ n8990 ;
  assign n11758 = n11757 ^ n11743 ;
  assign n11759 = n11744 & n11758 ;
  assign n11760 = n11759 ^ n8888 ;
  assign n11761 = n11760 ^ n11741 ;
  assign n11762 = ~n11742 & n11761 ;
  assign n11763 = n11762 ^ n8883 ;
  assign n11764 = n11763 ^ n11739 ;
  assign n11765 = n11740 & ~n11764 ;
  assign n11766 = n11765 ^ n8877 ;
  assign n11767 = n11766 ^ n11737 ;
  assign n11768 = n11738 & n11767 ;
  assign n11769 = n11768 ^ n8872 ;
  assign n11770 = n11769 ^ n11735 ;
  assign n11771 = ~n11736 & n11770 ;
  assign n11772 = n11771 ^ n8866 ;
  assign n11774 = n11773 ^ n11772 ;
  assign n11775 = n11773 ^ n8857 ;
  assign n11776 = ~n11774 & n11775 ;
  assign n11777 = n11776 ^ n8857 ;
  assign n11734 = n11672 ^ n11608 ;
  assign n11778 = n11777 ^ n11734 ;
  assign n11779 = n11777 ^ n8854 ;
  assign n11780 = ~n11778 & ~n11779 ;
  assign n11781 = n11780 ^ n8854 ;
  assign n11782 = n11781 ^ n11732 ;
  assign n11783 = ~n11733 & ~n11782 ;
  assign n11784 = n11783 ^ n8840 ;
  assign n11785 = n11784 ^ n11729 ;
  assign n11786 = n11730 & ~n11785 ;
  assign n11787 = n11786 ^ n9024 ;
  assign n11789 = n11788 ^ n11787 ;
  assign n11790 = n11788 ^ n9034 ;
  assign n11791 = n11789 & ~n11790 ;
  assign n11792 = n11791 ^ n9034 ;
  assign n11793 = n11792 ^ n11727 ;
  assign n11794 = ~n11728 & n11793 ;
  assign n11795 = n11794 ^ n9035 ;
  assign n11726 = n11694 ^ n11585 ;
  assign n11796 = n11795 ^ n11726 ;
  assign n11797 = n11795 ^ n9045 ;
  assign n11798 = ~n11796 & ~n11797 ;
  assign n11799 = n11798 ^ n9045 ;
  assign n11800 = n11799 ^ n11724 ;
  assign n11801 = n11725 & n11800 ;
  assign n11802 = n11801 ^ n9366 ;
  assign n11804 = n11803 ^ n11802 ;
  assign n11805 = n11803 ^ n8696 ;
  assign n11806 = ~n11804 & ~n11805 ;
  assign n11807 = n11806 ^ n8696 ;
  assign n11808 = n11807 ^ n11722 ;
  assign n11809 = n11723 & ~n11808 ;
  assign n11810 = n11809 ^ n8691 ;
  assign n11719 = n11304 ^ n11265 ;
  assign n11709 = n10008 ^ n9386 ;
  assign n11710 = ~n10729 & n11709 ;
  assign n11711 = n11710 ^ n9386 ;
  assign n11715 = n11711 ^ n11702 ;
  assign n11714 = n11713 ^ n11711 ;
  assign n11716 = n11715 ^ n11714 ;
  assign n11717 = n11708 & n11716 ;
  assign n11718 = n11717 ^ n11714 ;
  assign n11720 = n11719 ^ n11718 ;
  assign n11721 = n11720 ^ n8684 ;
  assign n11981 = n11810 ^ n11721 ;
  assign n11855 = n11807 ^ n11723 ;
  assign n11856 = n11781 ^ n11733 ;
  assign n11857 = n11734 ^ n8854 ;
  assign n11858 = n11857 ^ n11777 ;
  assign n11859 = n11775 ^ n11772 ;
  assign n11860 = n11757 ^ n11744 ;
  assign n11861 = n11747 ^ n8980 ;
  assign n11862 = n11861 ^ n11750 ;
  assign n11527 = n11526 ^ n11516 ;
  assign n11457 = n11456 ^ n11445 ;
  assign n11458 = n11415 ^ n8931 ;
  assign n11459 = n11418 ^ n11417 ;
  assign n11460 = n11458 & n11459 ;
  assign n11461 = n11423 ^ n11422 ;
  assign n11462 = n11460 & n11461 ;
  assign n11463 = n11429 ^ n11426 ;
  assign n11464 = ~n11462 & ~n11463 ;
  assign n11465 = n11431 ^ n11414 ;
  assign n11466 = n11464 & ~n11465 ;
  assign n11467 = n11437 ^ n11434 ;
  assign n11468 = ~n11466 & n11467 ;
  assign n11469 = n11439 ^ n11412 ;
  assign n11470 = n11468 & ~n11469 ;
  assign n11471 = n11442 ^ n11410 ;
  assign n11472 = ~n11470 & n11471 ;
  assign n11528 = ~n11457 & n11472 ;
  assign n11863 = n11527 & ~n11528 ;
  assign n11864 = n11862 & n11863 ;
  assign n11865 = n11754 ^ n11746 ;
  assign n11866 = ~n11864 & n11865 ;
  assign n11867 = ~n11860 & n11866 ;
  assign n11868 = n11760 ^ n11742 ;
  assign n11869 = n11867 & ~n11868 ;
  assign n11870 = n11763 ^ n11740 ;
  assign n11871 = n11869 & n11870 ;
  assign n11872 = n11766 ^ n11738 ;
  assign n11873 = ~n11871 & ~n11872 ;
  assign n11874 = n11769 ^ n11736 ;
  assign n11875 = n11873 & ~n11874 ;
  assign n11876 = ~n11859 & ~n11875 ;
  assign n11877 = ~n11858 & ~n11876 ;
  assign n11878 = n11856 & n11877 ;
  assign n11879 = n11784 ^ n11730 ;
  assign n11880 = n11878 & n11879 ;
  assign n11881 = n11790 ^ n11787 ;
  assign n11882 = n11880 & ~n11881 ;
  assign n11883 = n11792 ^ n11728 ;
  assign n11884 = n11882 & ~n11883 ;
  assign n11885 = n11797 ^ n11726 ;
  assign n11886 = ~n11884 & n11885 ;
  assign n11887 = n11799 ^ n11725 ;
  assign n11888 = ~n11886 & ~n11887 ;
  assign n11889 = n11805 ^ n11802 ;
  assign n11890 = ~n11888 & n11889 ;
  assign n11982 = ~n11855 & ~n11890 ;
  assign n11989 = ~n11981 & ~n11982 ;
  assign n11822 = n11309 ^ n11308 ;
  assign n11814 = n11719 ^ n11711 ;
  assign n11815 = n11718 & n11814 ;
  assign n11816 = n11815 ^ n11719 ;
  assign n11817 = n11816 ^ n9384 ;
  assign n11818 = n11817 ^ n9997 ;
  assign n11819 = n11818 ^ n11816 ;
  assign n11820 = n10734 & n11819 ;
  assign n11821 = n11820 ^ n11817 ;
  assign n11823 = n11822 ^ n11821 ;
  assign n11825 = n11823 ^ n8683 ;
  assign n11811 = n11810 ^ n11720 ;
  assign n11812 = ~n11721 & n11811 ;
  assign n11813 = n11812 ^ n8684 ;
  assign n11988 = n11825 ^ n11813 ;
  assign n11990 = n11989 ^ n11988 ;
  assign n11891 = n11890 ^ n11855 ;
  assign n11892 = n11891 ^ x453 ;
  assign n11893 = n11889 ^ n11888 ;
  assign n11894 = n11893 ^ x454 ;
  assign n11895 = n11887 ^ n11886 ;
  assign n11896 = n11895 ^ x455 ;
  assign n11897 = n11885 ^ n11884 ;
  assign n11898 = n11897 ^ x456 ;
  assign n11963 = n11883 ^ n11882 ;
  assign n11899 = n11881 ^ n11880 ;
  assign n11900 = n11899 ^ x458 ;
  assign n11901 = n11879 ^ n11878 ;
  assign n11902 = n11901 ^ x459 ;
  assign n11903 = n11876 ^ n11858 ;
  assign n11904 = n11903 ^ x461 ;
  assign n11905 = n11875 ^ n11859 ;
  assign n11906 = n11905 ^ x462 ;
  assign n11907 = n11874 ^ n11873 ;
  assign n11908 = n11907 ^ x463 ;
  assign n11910 = n11870 ^ n11869 ;
  assign n11911 = n11910 ^ x465 ;
  assign n11912 = n11868 ^ n11867 ;
  assign n11913 = n11912 ^ x466 ;
  assign n11927 = n11866 ^ n11860 ;
  assign n11914 = n11863 ^ n11862 ;
  assign n11915 = n11914 ^ x469 ;
  assign n11529 = n11528 ^ n11527 ;
  assign n11530 = n11529 ^ x470 ;
  assign n11473 = n11472 ^ n11457 ;
  assign n11474 = n11473 ^ x471 ;
  assign n11475 = n11471 ^ n11470 ;
  assign n11476 = n11475 ^ x472 ;
  assign n11477 = n11469 ^ n11468 ;
  assign n11478 = n11477 ^ x473 ;
  assign n11479 = n11467 ^ n11466 ;
  assign n11480 = n11479 ^ x474 ;
  assign n11497 = n11465 ^ n11464 ;
  assign n11481 = n11463 ^ n11462 ;
  assign n11482 = n11481 ^ x476 ;
  assign n11489 = n11461 ^ n11460 ;
  assign n11483 = x479 & ~n11458 ;
  assign n11484 = n11483 ^ x478 ;
  assign n11485 = n11459 ^ n11458 ;
  assign n11486 = n11485 ^ n11483 ;
  assign n11487 = n11484 & ~n11486 ;
  assign n11488 = n11487 ^ x478 ;
  assign n11490 = n11489 ^ n11488 ;
  assign n11491 = n11489 ^ x477 ;
  assign n11492 = ~n11490 & n11491 ;
  assign n11493 = n11492 ^ x477 ;
  assign n11494 = n11493 ^ n11481 ;
  assign n11495 = ~n11482 & n11494 ;
  assign n11496 = n11495 ^ x476 ;
  assign n11498 = n11497 ^ n11496 ;
  assign n11499 = n11497 ^ x475 ;
  assign n11500 = ~n11498 & n11499 ;
  assign n11501 = n11500 ^ x475 ;
  assign n11502 = n11501 ^ n11479 ;
  assign n11503 = ~n11480 & n11502 ;
  assign n11504 = n11503 ^ x474 ;
  assign n11505 = n11504 ^ n11477 ;
  assign n11506 = ~n11478 & n11505 ;
  assign n11507 = n11506 ^ x473 ;
  assign n11508 = n11507 ^ n11475 ;
  assign n11509 = n11476 & ~n11508 ;
  assign n11510 = n11509 ^ x472 ;
  assign n11511 = n11510 ^ n11473 ;
  assign n11512 = n11474 & ~n11511 ;
  assign n11513 = n11512 ^ x471 ;
  assign n11916 = n11529 ^ n11513 ;
  assign n11917 = ~n11530 & n11916 ;
  assign n11918 = n11917 ^ x470 ;
  assign n11919 = n11918 ^ n11914 ;
  assign n11920 = n11915 & ~n11919 ;
  assign n11921 = n11920 ^ x469 ;
  assign n11922 = n11921 ^ x468 ;
  assign n11923 = n11865 ^ n11864 ;
  assign n11924 = n11923 ^ n11921 ;
  assign n11925 = n11922 & ~n11924 ;
  assign n11926 = n11925 ^ x468 ;
  assign n11928 = n11927 ^ n11926 ;
  assign n11929 = n11927 ^ x467 ;
  assign n11930 = ~n11928 & n11929 ;
  assign n11931 = n11930 ^ x467 ;
  assign n11932 = n11931 ^ n11912 ;
  assign n11933 = n11913 & ~n11932 ;
  assign n11934 = n11933 ^ x466 ;
  assign n11935 = n11934 ^ n11910 ;
  assign n11936 = ~n11911 & n11935 ;
  assign n11937 = n11936 ^ x465 ;
  assign n11909 = n11872 ^ n11871 ;
  assign n11938 = n11937 ^ n11909 ;
  assign n11939 = n11907 ^ x464 ;
  assign n11940 = n11939 ^ n11907 ;
  assign n11941 = n11940 ^ n11909 ;
  assign n11942 = ~n11938 & n11941 ;
  assign n11943 = n11942 ^ n11939 ;
  assign n11944 = ~n11908 & n11943 ;
  assign n11945 = n11944 ^ x463 ;
  assign n11946 = n11945 ^ n11905 ;
  assign n11947 = ~n11906 & n11946 ;
  assign n11948 = n11947 ^ x462 ;
  assign n11949 = n11948 ^ n11903 ;
  assign n11950 = n11904 & ~n11949 ;
  assign n11951 = n11950 ^ x461 ;
  assign n11952 = n11951 ^ x460 ;
  assign n11953 = n11877 ^ n11856 ;
  assign n11954 = n11953 ^ n11951 ;
  assign n11955 = n11952 & ~n11954 ;
  assign n11956 = n11955 ^ x460 ;
  assign n11957 = n11956 ^ n11901 ;
  assign n11958 = n11902 & ~n11957 ;
  assign n11959 = n11958 ^ x459 ;
  assign n11960 = n11959 ^ n11899 ;
  assign n11961 = ~n11900 & n11960 ;
  assign n11962 = n11961 ^ x458 ;
  assign n11964 = n11963 ^ n11962 ;
  assign n11965 = n11963 ^ x457 ;
  assign n11966 = n11964 & ~n11965 ;
  assign n11967 = n11966 ^ x457 ;
  assign n11968 = n11967 ^ n11897 ;
  assign n11969 = n11898 & ~n11968 ;
  assign n11970 = n11969 ^ x456 ;
  assign n11971 = n11970 ^ n11895 ;
  assign n11972 = n11896 & ~n11971 ;
  assign n11973 = n11972 ^ x455 ;
  assign n11974 = n11973 ^ n11893 ;
  assign n11975 = n11894 & ~n11974 ;
  assign n11976 = n11975 ^ x454 ;
  assign n11977 = n11976 ^ n11891 ;
  assign n11978 = n11892 & ~n11977 ;
  assign n11979 = n11978 ^ x453 ;
  assign n11980 = n11979 ^ x452 ;
  assign n11983 = n11982 ^ n11981 ;
  assign n11984 = n11983 ^ n11979 ;
  assign n11985 = n11980 & n11984 ;
  assign n11986 = n11985 ^ x452 ;
  assign n11987 = n11986 ^ x451 ;
  assign n12050 = n11990 ^ n11987 ;
  assign n12040 = n11983 ^ n11980 ;
  assign n12041 = n10194 ^ n10127 ;
  assign n12042 = n10984 & n12041 ;
  assign n12043 = n12042 ^ n10127 ;
  assign n12044 = ~n12040 & n12043 ;
  assign n12045 = n12044 ^ n10284 ;
  assign n12046 = n12045 ^ n10772 ;
  assign n12047 = n12046 ^ n12044 ;
  assign n12048 = n10982 & n12047 ;
  assign n12049 = n12048 ^ n12045 ;
  assign n12142 = n12050 ^ n12049 ;
  assign n12140 = n12043 ^ n12040 ;
  assign n12141 = ~n8826 & ~n12140 ;
  assign n12143 = n12142 ^ n12141 ;
  assign n12144 = n12142 ^ n8820 ;
  assign n12145 = ~n12143 & n12144 ;
  assign n12146 = n12145 ^ n8820 ;
  assign n12034 = n10301 ^ n10191 ;
  assign n12035 = n11407 & ~n12034 ;
  assign n12036 = n12035 ^ n10301 ;
  assign n12052 = n12044 ^ n12036 ;
  assign n12051 = n12050 ^ n12036 ;
  assign n12053 = n12052 ^ n12051 ;
  assign n12054 = ~n12049 & ~n12053 ;
  assign n12055 = n12054 ^ n12052 ;
  assign n11997 = n11988 & n11989 ;
  assign n11833 = n10057 ^ n9379 ;
  assign n11834 = ~n10748 & n11833 ;
  assign n11835 = n11834 ^ n9379 ;
  assign n11830 = n11312 ^ n11263 ;
  assign n11831 = n11830 ^ n11822 ;
  assign n11828 = n11822 ^ n11816 ;
  assign n11829 = ~n11821 & ~n11828 ;
  assign n11832 = n11831 ^ n11829 ;
  assign n11836 = n11835 ^ n11832 ;
  assign n11995 = n11836 ^ n8737 ;
  assign n11824 = n11823 ^ n11813 ;
  assign n11826 = n11824 & n11825 ;
  assign n11827 = n11826 ^ n8683 ;
  assign n11996 = n11995 ^ n11827 ;
  assign n11998 = n11997 ^ n11996 ;
  assign n11991 = n11990 ^ n11986 ;
  assign n11992 = n11987 & n11991 ;
  assign n11993 = n11992 ^ x451 ;
  assign n11994 = n11993 ^ x450 ;
  assign n12038 = n11998 ^ n11994 ;
  assign n12138 = n12055 ^ n12038 ;
  assign n12139 = n12138 ^ n8813 ;
  assign n12215 = n12146 ^ n12139 ;
  assign n12216 = n12140 ^ n8826 ;
  assign n12217 = n12141 ^ n8820 ;
  assign n12218 = n12217 ^ n12142 ;
  assign n12219 = n12216 & n12218 ;
  assign n12220 = n12215 & n12219 ;
  assign n12039 = n12038 ^ n12036 ;
  assign n12056 = ~n12039 & ~n12055 ;
  assign n12030 = n10207 ^ n10181 ;
  assign n12031 = ~n11453 & n12030 ;
  assign n12032 = n12031 ^ n10207 ;
  assign n12037 = n12036 ^ n12032 ;
  assign n12057 = n12056 ^ n12037 ;
  assign n12005 = ~n11996 & ~n11997 ;
  assign n11837 = n11836 ^ n11827 ;
  assign n11838 = n11827 ^ n8737 ;
  assign n11839 = n11837 & n11838 ;
  assign n11840 = n11839 ^ n11836 ;
  assign n12003 = n11840 ^ n8770 ;
  assign n11848 = n10063 ^ n8833 ;
  assign n11849 = n10756 & ~n11848 ;
  assign n11850 = n11849 ^ n8833 ;
  assign n11841 = n11315 ^ x422 ;
  assign n11842 = n11841 ^ n11260 ;
  assign n11844 = n11842 ^ n11830 ;
  assign n11843 = n11842 ^ n11835 ;
  assign n11845 = n11844 ^ n11843 ;
  assign n11846 = n11832 & n11845 ;
  assign n11847 = n11846 ^ n11844 ;
  assign n11851 = n11850 ^ n11847 ;
  assign n12004 = n12003 ^ n11851 ;
  assign n12006 = n12005 ^ n12004 ;
  assign n11999 = n11998 ^ n11993 ;
  assign n12000 = n11994 & ~n11999 ;
  assign n12001 = n12000 ^ x450 ;
  assign n12002 = n12001 ^ x449 ;
  assign n12029 = n12006 ^ n12002 ;
  assign n12137 = n12057 ^ n12029 ;
  assign n12213 = n12137 ^ n8807 ;
  assign n12147 = n12146 ^ n12138 ;
  assign n12148 = n12139 & n12147 ;
  assign n12149 = n12148 ^ n8813 ;
  assign n12214 = n12213 ^ n12149 ;
  assign n12276 = n12220 ^ n12214 ;
  assign n12264 = x511 & ~n12216 ;
  assign n12265 = n12264 ^ x510 ;
  assign n12266 = n12218 ^ n12216 ;
  assign n12267 = n12266 ^ n12264 ;
  assign n12268 = n12265 & ~n12267 ;
  assign n12269 = n12268 ^ x510 ;
  assign n12270 = n12269 ^ x509 ;
  assign n12271 = n12219 ^ n12215 ;
  assign n12272 = n12271 ^ n12269 ;
  assign n12273 = n12270 & ~n12272 ;
  assign n12274 = n12273 ^ x509 ;
  assign n12275 = n12274 ^ x508 ;
  assign n12356 = n12276 ^ n12275 ;
  assign n12337 = n11929 ^ n11926 ;
  assign n12197 = n11923 ^ n11922 ;
  assign n12198 = n12197 ^ n10227 ;
  assign n12199 = n12198 ^ n10997 ;
  assign n12200 = n12199 ^ n12197 ;
  assign n12201 = n11587 & ~n12200 ;
  assign n12202 = n12201 ^ n12198 ;
  assign n12329 = n10990 ^ n10223 ;
  assign n12330 = n11593 & ~n12329 ;
  assign n12331 = n12330 ^ n10223 ;
  assign n12333 = n12331 ^ n12197 ;
  assign n12118 = n11918 ^ n11915 ;
  assign n12115 = n11007 ^ n10229 ;
  assign n12116 = n11598 & n12115 ;
  assign n12117 = n12116 ^ n11007 ;
  assign n12119 = n12118 ^ n12117 ;
  assign n11531 = n11530 ^ n11513 ;
  assign n10976 = n10975 ^ n10350 ;
  assign n10977 = n10974 & ~n10976 ;
  assign n10978 = n10977 ^ n10975 ;
  assign n11532 = n11531 ^ n10978 ;
  assign n12102 = n11510 ^ x471 ;
  assign n12103 = n12102 ^ n11473 ;
  assign n12092 = n11507 ^ x472 ;
  assign n12093 = n12092 ^ n11475 ;
  assign n11537 = n11504 ^ n11478 ;
  assign n11534 = n11022 ^ n10341 ;
  assign n11535 = ~n11533 & ~n11534 ;
  assign n11536 = n11535 ^ n11022 ;
  assign n11538 = n11537 ^ n11536 ;
  assign n11543 = n11501 ^ x474 ;
  assign n11544 = n11543 ^ n11479 ;
  assign n11540 = n11048 ^ n9605 ;
  assign n11541 = n11539 & n11540 ;
  assign n11542 = n11541 ^ n9605 ;
  assign n11545 = n11544 ^ n11542 ;
  assign n12077 = n11499 ^ n11496 ;
  assign n11550 = n11493 ^ x476 ;
  assign n11551 = n11550 ^ n11481 ;
  assign n11547 = n11033 ^ n10182 ;
  assign n11548 = n11546 & n11547 ;
  assign n11549 = n11548 ^ n10182 ;
  assign n11552 = n11551 ^ n11549 ;
  assign n11558 = n11485 ^ n11484 ;
  assign n11559 = n11558 ^ n10317 ;
  assign n11560 = n11559 ^ n10852 ;
  assign n11561 = n11560 ^ n11558 ;
  assign n11562 = n11557 & ~n11561 ;
  assign n11563 = n11562 ^ n11559 ;
  assign n11569 = n11458 ^ x479 ;
  assign n11566 = n10193 ^ n10167 ;
  assign n11567 = ~n11565 & n11566 ;
  assign n11568 = n11567 ^ n10193 ;
  assign n11570 = n11569 ^ n11568 ;
  assign n12025 = n10200 ^ n10179 ;
  assign n12026 = ~n11520 & ~n12025 ;
  assign n12027 = n12026 ^ n10200 ;
  assign n12019 = n11850 ^ n11842 ;
  assign n12020 = n11847 & ~n12019 ;
  assign n12016 = n10064 ^ n9423 ;
  assign n12017 = ~n10724 & n12016 ;
  assign n12012 = n11850 ^ n11386 ;
  assign n12011 = n11318 ^ n11259 ;
  assign n12013 = n12012 ^ n12011 ;
  assign n12014 = n12013 ^ n8770 ;
  assign n12010 = x449 ^ x448 ;
  assign n12015 = n12014 ^ n12010 ;
  assign n12018 = n12017 ^ n12015 ;
  assign n12021 = n12020 ^ n12018 ;
  assign n12009 = n12004 & ~n12005 ;
  assign n12022 = n12021 ^ n12009 ;
  assign n12007 = n12006 ^ n12001 ;
  assign n12008 = n12002 & ~n12007 ;
  assign n12023 = n12022 ^ n12008 ;
  assign n11852 = n11851 ^ n11840 ;
  assign n11853 = n11851 ^ n8770 ;
  assign n11854 = n11852 & ~n11853 ;
  assign n12024 = n12023 ^ n11854 ;
  assign n12028 = n12027 ^ n12024 ;
  assign n12033 = n12032 ^ n12029 ;
  assign n12058 = n12033 & ~n12057 ;
  assign n12059 = n12058 ^ n12032 ;
  assign n12060 = n12059 ^ n12024 ;
  assign n12061 = ~n12028 & ~n12060 ;
  assign n12062 = n12061 ^ n12027 ;
  assign n12063 = n12062 ^ n11568 ;
  assign n12064 = ~n11570 & n12063 ;
  assign n12065 = n12064 ^ n11569 ;
  assign n12066 = n12065 ^ n11558 ;
  assign n12067 = ~n11563 & ~n12066 ;
  assign n12068 = n12067 ^ n11558 ;
  assign n11554 = n10961 ^ n10187 ;
  assign n11555 = ~n11553 & ~n11554 ;
  assign n11556 = n11555 ^ n10187 ;
  assign n12069 = n12068 ^ n11556 ;
  assign n12070 = n11491 ^ n11488 ;
  assign n12071 = n12070 ^ n11556 ;
  assign n12072 = n12069 & ~n12071 ;
  assign n12073 = n12072 ^ n12068 ;
  assign n12074 = n12073 ^ n11549 ;
  assign n12075 = n11552 & n12074 ;
  assign n12076 = n12075 ^ n11551 ;
  assign n12078 = n12077 ^ n12076 ;
  assign n12079 = n12077 ^ n10174 ;
  assign n12080 = n12079 ^ n11028 ;
  assign n12081 = n12080 ^ n12077 ;
  assign n12082 = ~n11655 & ~n12081 ;
  assign n12083 = n12082 ^ n12079 ;
  assign n12084 = ~n12078 & ~n12083 ;
  assign n12085 = n12084 ^ n12077 ;
  assign n12086 = n12085 ^ n11542 ;
  assign n12087 = n11545 & n12086 ;
  assign n12088 = n12087 ^ n11544 ;
  assign n12089 = n12088 ^ n11536 ;
  assign n12090 = ~n11538 & n12089 ;
  assign n12091 = n12090 ^ n11537 ;
  assign n12094 = n12093 ^ n12091 ;
  assign n12095 = n12093 ^ n10245 ;
  assign n12096 = n12095 ^ n11019 ;
  assign n12097 = n12096 ^ n12093 ;
  assign n12098 = ~n11612 & ~n12097 ;
  assign n12099 = n12098 ^ n12095 ;
  assign n12100 = ~n12094 & ~n12099 ;
  assign n12101 = n12100 ^ n12093 ;
  assign n12104 = n12103 ^ n12101 ;
  assign n12105 = n12103 ^ n11014 ;
  assign n12106 = n12105 ^ n10236 ;
  assign n12107 = n12106 ^ n12103 ;
  assign n12108 = ~n11607 & n12107 ;
  assign n12109 = n12108 ^ n12105 ;
  assign n12110 = n12104 & ~n12109 ;
  assign n12111 = n12110 ^ n12103 ;
  assign n12112 = n12111 ^ n10978 ;
  assign n12113 = n11532 & n12112 ;
  assign n12114 = n12113 ^ n11531 ;
  assign n12203 = n12117 ^ n12114 ;
  assign n12204 = n12119 & n12203 ;
  assign n12205 = n12204 ^ n12118 ;
  assign n12332 = n12331 ^ n12205 ;
  assign n12334 = n12333 ^ n12332 ;
  assign n12335 = n12202 & n12334 ;
  assign n12336 = n12335 ^ n12333 ;
  assign n12338 = n12337 ^ n12336 ;
  assign n12339 = n12338 ^ n9612 ;
  assign n12206 = n12205 ^ n12202 ;
  assign n12207 = n12206 ^ n9627 ;
  assign n12120 = n12119 ^ n12114 ;
  assign n12121 = n12120 ^ n9630 ;
  assign n12189 = n12111 ^ n11532 ;
  assign n12122 = n12109 ^ n12101 ;
  assign n12123 = n12122 ^ n9709 ;
  assign n12181 = n12099 ^ n12091 ;
  assign n12124 = n12088 ^ n11538 ;
  assign n12125 = n12124 ^ n9701 ;
  assign n12126 = n12085 ^ n11545 ;
  assign n12127 = n12126 ^ n9692 ;
  assign n12170 = n12083 ^ n12076 ;
  assign n12128 = n12073 ^ n11552 ;
  assign n12129 = n12128 ^ n9649 ;
  assign n12130 = n12071 ^ n12068 ;
  assign n12131 = n12130 ^ n9654 ;
  assign n12133 = n12062 ^ n11570 ;
  assign n12134 = n12133 ^ n9538 ;
  assign n12135 = n12059 ^ n12028 ;
  assign n12136 = n12135 ^ n9449 ;
  assign n12150 = n12149 ^ n12137 ;
  assign n12151 = n12149 ^ n8807 ;
  assign n12152 = ~n12150 & n12151 ;
  assign n12153 = n12152 ^ n8807 ;
  assign n12154 = n12153 ^ n12135 ;
  assign n12155 = n12136 & ~n12154 ;
  assign n12156 = n12155 ^ n9449 ;
  assign n12157 = n12156 ^ n12133 ;
  assign n12158 = ~n12134 & n12157 ;
  assign n12159 = n12158 ^ n9538 ;
  assign n12132 = n12065 ^ n11563 ;
  assign n12160 = n12159 ^ n12132 ;
  assign n12161 = n12159 ^ n9661 ;
  assign n12162 = n12160 & ~n12161 ;
  assign n12163 = n12162 ^ n9661 ;
  assign n12164 = n12163 ^ n12130 ;
  assign n12165 = ~n12131 & ~n12164 ;
  assign n12166 = n12165 ^ n9654 ;
  assign n12167 = n12166 ^ n12128 ;
  assign n12168 = n12129 & n12167 ;
  assign n12169 = n12168 ^ n9649 ;
  assign n12171 = n12170 ^ n12169 ;
  assign n12172 = n12170 ^ n9679 ;
  assign n12173 = ~n12171 & n12172 ;
  assign n12174 = n12173 ^ n9679 ;
  assign n12175 = n12174 ^ n12126 ;
  assign n12176 = ~n12127 & ~n12175 ;
  assign n12177 = n12176 ^ n9692 ;
  assign n12178 = n12177 ^ n12124 ;
  assign n12179 = ~n12125 & n12178 ;
  assign n12180 = n12179 ^ n9701 ;
  assign n12182 = n12181 ^ n12180 ;
  assign n12183 = n12181 ^ n9638 ;
  assign n12184 = n12182 & ~n12183 ;
  assign n12185 = n12184 ^ n9638 ;
  assign n12186 = n12185 ^ n12122 ;
  assign n12187 = n12123 & ~n12186 ;
  assign n12188 = n12187 ^ n9709 ;
  assign n12190 = n12189 ^ n12188 ;
  assign n12191 = n12189 ^ n9635 ;
  assign n12192 = n12190 & ~n12191 ;
  assign n12193 = n12192 ^ n9635 ;
  assign n12194 = n12193 ^ n12120 ;
  assign n12195 = n12121 & ~n12194 ;
  assign n12196 = n12195 ^ n9630 ;
  assign n12326 = n12206 ^ n12196 ;
  assign n12327 = n12207 & n12326 ;
  assign n12328 = n12327 ^ n9627 ;
  assign n12494 = n12338 ^ n12328 ;
  assign n12495 = ~n12339 & ~n12494 ;
  assign n12496 = n12495 ^ n9612 ;
  assign n12432 = n11931 ^ x466 ;
  assign n12433 = n12432 ^ n11912 ;
  assign n12424 = n10996 ^ n10383 ;
  assign n12425 = ~n11585 & n12424 ;
  assign n12426 = n12425 ^ n10383 ;
  assign n12428 = n12426 ^ n12331 ;
  assign n12427 = n12426 ^ n12337 ;
  assign n12429 = n12428 ^ n12427 ;
  assign n12430 = n12336 & n12429 ;
  assign n12431 = n12430 ^ n12428 ;
  assign n12493 = n12433 ^ n12431 ;
  assign n12497 = n12496 ^ n12493 ;
  assign n12498 = n12496 ^ n9730 ;
  assign n12499 = n12497 & n12498 ;
  assign n12500 = n12499 ^ n9730 ;
  assign n12418 = n11096 ^ n10388 ;
  assign n12419 = n11571 & ~n12418 ;
  assign n12420 = n12419 ^ n10388 ;
  assign n12435 = n12426 ^ n12420 ;
  assign n12434 = n12433 ^ n12420 ;
  assign n12436 = n12435 ^ n12434 ;
  assign n12437 = n12431 & n12436 ;
  assign n12438 = n12437 ^ n12435 ;
  assign n12422 = n11934 ^ n11911 ;
  assign n12491 = n12438 ^ n12422 ;
  assign n12492 = n12491 ^ n9739 ;
  assign n12540 = n12500 ^ n12492 ;
  assign n12541 = n12493 ^ n9730 ;
  assign n12542 = n12541 ^ n12496 ;
  assign n12340 = n12339 ^ n12328 ;
  assign n12208 = n12207 ^ n12196 ;
  assign n12209 = n12174 ^ n12127 ;
  assign n12210 = n12172 ^ n12169 ;
  assign n12211 = n12132 ^ n9661 ;
  assign n12212 = n12211 ^ n12159 ;
  assign n12221 = n12214 & ~n12220 ;
  assign n12222 = n12153 ^ n12136 ;
  assign n12223 = n12221 & n12222 ;
  assign n12224 = n12156 ^ n12134 ;
  assign n12225 = ~n12223 & n12224 ;
  assign n12226 = ~n12212 & n12225 ;
  assign n12227 = n12163 ^ n12131 ;
  assign n12228 = ~n12226 & n12227 ;
  assign n12229 = n12166 ^ n12129 ;
  assign n12230 = n12228 & n12229 ;
  assign n12231 = n12210 & ~n12230 ;
  assign n12232 = ~n12209 & n12231 ;
  assign n12233 = n12177 ^ n12125 ;
  assign n12234 = ~n12232 & ~n12233 ;
  assign n12235 = n12183 ^ n12180 ;
  assign n12236 = n12234 & ~n12235 ;
  assign n12237 = n12185 ^ n12123 ;
  assign n12238 = n12236 & n12237 ;
  assign n12239 = n12191 ^ n12188 ;
  assign n12240 = n12238 & ~n12239 ;
  assign n12241 = n12193 ^ n12121 ;
  assign n12242 = ~n12240 & ~n12241 ;
  assign n12341 = ~n12208 & n12242 ;
  assign n12543 = n12340 & ~n12341 ;
  assign n12544 = n12542 & ~n12543 ;
  assign n12545 = ~n12540 & n12544 ;
  assign n12501 = n12500 ^ n12491 ;
  assign n12502 = n12492 & ~n12501 ;
  assign n12503 = n12502 ^ n9739 ;
  assign n12423 = n12422 ^ n12420 ;
  assign n12439 = ~n12423 & n12438 ;
  assign n12414 = n11170 ^ n10218 ;
  assign n12415 = ~n11703 & n12414 ;
  assign n12416 = n12415 ^ n10218 ;
  assign n12421 = n12420 ^ n12416 ;
  assign n12440 = n12439 ^ n12421 ;
  assign n12412 = n11937 ^ x464 ;
  assign n12413 = n12412 ^ n11909 ;
  assign n12489 = n12440 ^ n12413 ;
  assign n12490 = n12489 ^ n9609 ;
  assign n12546 = n12503 ^ n12490 ;
  assign n12547 = n12545 & ~n12546 ;
  assign n12417 = n12416 ^ n12413 ;
  assign n12441 = n12417 & n12440 ;
  assign n12442 = n12441 ^ n12416 ;
  assign n12408 = n11186 ^ n10402 ;
  assign n12409 = n11713 & n12408 ;
  assign n12410 = n12409 ^ n10402 ;
  assign n12407 = n11943 ^ x463 ;
  assign n12411 = n12410 ^ n12407 ;
  assign n12488 = n12442 ^ n12411 ;
  assign n12538 = n12488 ^ n9752 ;
  assign n12504 = n12503 ^ n12489 ;
  assign n12505 = n12490 & n12504 ;
  assign n12506 = n12505 ^ n9609 ;
  assign n12539 = n12538 ^ n12506 ;
  assign n12569 = n12547 ^ n12539 ;
  assign n12570 = n12569 ^ x490 ;
  assign n12571 = n12546 ^ n12545 ;
  assign n12572 = n12571 ^ x491 ;
  assign n12573 = n12543 ^ n12542 ;
  assign n12574 = n12573 ^ x493 ;
  assign n12342 = n12341 ^ n12340 ;
  assign n12575 = n12342 ^ x494 ;
  assign n12243 = n12242 ^ n12208 ;
  assign n12244 = n12243 ^ x495 ;
  assign n12246 = n12239 ^ n12238 ;
  assign n12247 = n12246 ^ x497 ;
  assign n12248 = n12235 ^ n12234 ;
  assign n12249 = n12248 ^ x499 ;
  assign n12250 = n12233 ^ n12232 ;
  assign n12251 = n12250 ^ x500 ;
  assign n12298 = n12231 ^ n12209 ;
  assign n12252 = n12230 ^ n12210 ;
  assign n12253 = n12252 ^ x502 ;
  assign n12254 = n12229 ^ n12228 ;
  assign n12255 = n12254 ^ x503 ;
  assign n12256 = n12227 ^ n12226 ;
  assign n12257 = n12256 ^ x504 ;
  assign n12258 = n12225 ^ n12212 ;
  assign n12259 = n12258 ^ x505 ;
  assign n12260 = n12224 ^ n12223 ;
  assign n12261 = n12260 ^ x506 ;
  assign n12262 = n12222 ^ n12221 ;
  assign n12263 = n12262 ^ x507 ;
  assign n12277 = n12276 ^ n12274 ;
  assign n12278 = n12275 & ~n12277 ;
  assign n12279 = n12278 ^ x508 ;
  assign n12280 = n12279 ^ n12262 ;
  assign n12281 = ~n12263 & n12280 ;
  assign n12282 = n12281 ^ x507 ;
  assign n12283 = n12282 ^ n12260 ;
  assign n12284 = ~n12261 & n12283 ;
  assign n12285 = n12284 ^ x506 ;
  assign n12286 = n12285 ^ n12258 ;
  assign n12287 = ~n12259 & n12286 ;
  assign n12288 = n12287 ^ x505 ;
  assign n12289 = n12288 ^ n12256 ;
  assign n12290 = n12257 & ~n12289 ;
  assign n12291 = n12290 ^ x504 ;
  assign n12292 = n12291 ^ n12254 ;
  assign n12293 = ~n12255 & n12292 ;
  assign n12294 = n12293 ^ x503 ;
  assign n12295 = n12294 ^ n12252 ;
  assign n12296 = ~n12253 & n12295 ;
  assign n12297 = n12296 ^ x502 ;
  assign n12299 = n12298 ^ n12297 ;
  assign n12300 = n12298 ^ x501 ;
  assign n12301 = n12299 & ~n12300 ;
  assign n12302 = n12301 ^ x501 ;
  assign n12303 = n12302 ^ n12250 ;
  assign n12304 = ~n12251 & n12303 ;
  assign n12305 = n12304 ^ x500 ;
  assign n12306 = n12305 ^ n12248 ;
  assign n12307 = n12249 & ~n12306 ;
  assign n12308 = n12307 ^ x499 ;
  assign n12309 = n12308 ^ x498 ;
  assign n12310 = n12237 ^ n12236 ;
  assign n12311 = n12310 ^ n12308 ;
  assign n12312 = n12309 & n12311 ;
  assign n12313 = n12312 ^ x498 ;
  assign n12314 = n12313 ^ n12246 ;
  assign n12315 = n12247 & ~n12314 ;
  assign n12316 = n12315 ^ x497 ;
  assign n12245 = n12241 ^ n12240 ;
  assign n12317 = n12316 ^ n12245 ;
  assign n12318 = n12243 ^ x496 ;
  assign n12319 = n12318 ^ n12243 ;
  assign n12320 = n12319 ^ n12245 ;
  assign n12321 = ~n12317 & n12320 ;
  assign n12322 = n12321 ^ n12318 ;
  assign n12323 = ~n12244 & n12322 ;
  assign n12324 = n12323 ^ x495 ;
  assign n12576 = n12342 ^ n12324 ;
  assign n12577 = n12575 & ~n12576 ;
  assign n12578 = n12577 ^ x494 ;
  assign n12579 = n12578 ^ n12573 ;
  assign n12580 = ~n12574 & n12579 ;
  assign n12581 = n12580 ^ x493 ;
  assign n12582 = n12581 ^ x492 ;
  assign n12583 = n12544 ^ n12540 ;
  assign n12584 = n12583 ^ n12581 ;
  assign n12585 = n12582 & n12584 ;
  assign n12586 = n12585 ^ x492 ;
  assign n12587 = n12586 ^ n12571 ;
  assign n12588 = ~n12572 & n12587 ;
  assign n12589 = n12588 ^ x491 ;
  assign n12590 = n12589 ^ n12569 ;
  assign n12591 = n12570 & ~n12590 ;
  assign n12592 = n12591 ^ x490 ;
  assign n12548 = n12539 & n12547 ;
  assign n12507 = n12506 ^ n12488 ;
  assign n12508 = n12506 ^ n9752 ;
  assign n12509 = ~n12507 & n12508 ;
  assign n12510 = n12509 ^ n9752 ;
  assign n12443 = n12442 ^ n12407 ;
  assign n12444 = n12411 & n12443 ;
  assign n12445 = n12444 ^ n12410 ;
  assign n12403 = n11226 ^ n10216 ;
  assign n12404 = ~n11719 & ~n12403 ;
  assign n12405 = n12404 ^ n10216 ;
  assign n12401 = n11945 ^ x462 ;
  assign n12402 = n12401 ^ n11905 ;
  assign n12406 = n12405 ^ n12402 ;
  assign n12486 = n12445 ^ n12406 ;
  assign n12487 = n12486 ^ n9842 ;
  assign n12537 = n12510 ^ n12487 ;
  assign n12568 = n12548 ^ n12537 ;
  assign n12593 = n12592 ^ n12568 ;
  assign n12594 = n12592 ^ x489 ;
  assign n12595 = ~n12593 & n12594 ;
  assign n12596 = n12595 ^ x489 ;
  assign n13170 = n12596 ^ x488 ;
  assign n12511 = n12510 ^ n12486 ;
  assign n12512 = n12487 & n12511 ;
  assign n12513 = n12512 ^ n9842 ;
  assign n12446 = n12445 ^ n12402 ;
  assign n12447 = n12406 & ~n12446 ;
  assign n12448 = n12447 ^ n12405 ;
  assign n12399 = n11948 ^ n11904 ;
  assign n12396 = n11241 ^ n10413 ;
  assign n12397 = n11822 & n12396 ;
  assign n12398 = n12397 ^ n10413 ;
  assign n12400 = n12399 ^ n12398 ;
  assign n12484 = n12448 ^ n12400 ;
  assign n12485 = n12484 ^ n9985 ;
  assign n12550 = n12513 ^ n12485 ;
  assign n12549 = n12537 & n12548 ;
  assign n12566 = n12550 ^ n12549 ;
  assign n13171 = n13170 ^ n12566 ;
  assign n12645 = n11973 ^ x454 ;
  assign n12646 = n12645 ^ n11893 ;
  assign n12959 = n12586 ^ x491 ;
  assign n12960 = n12959 ^ n12571 ;
  assign n12961 = n12960 ^ n10729 ;
  assign n12962 = n12961 ^ n11340 ;
  assign n12963 = n12962 ^ n12960 ;
  assign n12964 = n12646 & n12963 ;
  assign n12965 = n12964 ^ n12961 ;
  assign n12464 = n11970 ^ n11896 ;
  assign n12972 = n12011 ^ n11381 ;
  assign n12973 = n12464 & ~n12972 ;
  assign n12974 = n12973 ^ n11381 ;
  assign n12971 = n12583 ^ n12582 ;
  assign n12975 = n12974 ^ n12971 ;
  assign n12369 = n11967 ^ x456 ;
  assign n12370 = n12369 ^ n11897 ;
  assign n12977 = n11842 ^ n11241 ;
  assign n12978 = n12370 & ~n12977 ;
  assign n12979 = n12978 ^ n11241 ;
  assign n12976 = n12578 ^ n12574 ;
  assign n12980 = n12979 ^ n12976 ;
  assign n13046 = n12322 ^ x495 ;
  assign n12390 = n11956 ^ n11902 ;
  assign n12983 = n11719 ^ n11170 ;
  assign n12984 = n12390 & ~n12983 ;
  assign n12985 = n12984 ^ n11170 ;
  assign n12981 = n12316 ^ x496 ;
  assign n12982 = n12981 ^ n12245 ;
  assign n12986 = n12985 ^ n12982 ;
  assign n12344 = n11953 ^ n11952 ;
  assign n12987 = n11713 ^ n11096 ;
  assign n12988 = n12344 & ~n12987 ;
  assign n12989 = n12988 ^ n11096 ;
  assign n12899 = n12313 ^ n12247 ;
  assign n12990 = n12989 ^ n12899 ;
  assign n12991 = n11571 ^ n10990 ;
  assign n12992 = ~n12402 & ~n12991 ;
  assign n12993 = n12992 ^ n10990 ;
  assign n12913 = n12305 ^ n12249 ;
  assign n12994 = n12993 ^ n12913 ;
  assign n13018 = n11585 ^ n10997 ;
  assign n13019 = ~n12407 & n13018 ;
  assign n13020 = n13019 ^ n10997 ;
  assign n13028 = n13020 ^ n12993 ;
  assign n12940 = n12294 ^ n12253 ;
  assign n12995 = n12940 ^ n10975 ;
  assign n12996 = n12995 ^ n11587 ;
  assign n12997 = n12996 ^ n12940 ;
  assign n12998 = ~n12422 & ~n12997 ;
  assign n12999 = n12998 ^ n12995 ;
  assign n13010 = n11593 ^ n11007 ;
  assign n13011 = n12413 & n13010 ;
  assign n13012 = n13011 ^ n11007 ;
  assign n13014 = n13012 ^ n12940 ;
  assign n13003 = n11598 ^ n11014 ;
  assign n13004 = n12433 & n13003 ;
  assign n13005 = n13004 ^ n11014 ;
  assign n12887 = n11019 ^ n10974 ;
  assign n12888 = n12337 & ~n12887 ;
  assign n12889 = n12888 ^ n11019 ;
  assign n12885 = n12288 ^ x504 ;
  assign n12886 = n12885 ^ n12256 ;
  assign n12890 = n12889 ^ n12886 ;
  assign n12789 = n11607 ^ n11022 ;
  assign n12790 = n12197 & n12789 ;
  assign n12791 = n12790 ^ n11022 ;
  assign n12788 = n12285 ^ n12259 ;
  assign n12792 = n12791 ^ n12788 ;
  assign n12726 = n11612 ^ n11048 ;
  assign n12727 = n12118 & n12726 ;
  assign n12728 = n12727 ^ n11048 ;
  assign n12724 = n12282 ^ x506 ;
  assign n12725 = n12724 ^ n12260 ;
  assign n12729 = n12728 ^ n12725 ;
  assign n12349 = n11533 ^ n11028 ;
  assign n12350 = ~n11531 & n12349 ;
  assign n12351 = n12350 ^ n11028 ;
  assign n12348 = n12279 ^ n12263 ;
  assign n12352 = n12351 ^ n12348 ;
  assign n12353 = n11539 ^ n11033 ;
  assign n12354 = n12103 & ~n12353 ;
  assign n12355 = n12354 ^ n11033 ;
  assign n12357 = n12356 ^ n12355 ;
  assign n12709 = n12271 ^ n12270 ;
  assign n12359 = n11546 ^ n10852 ;
  assign n12360 = ~n11537 & n12359 ;
  assign n12361 = n12360 ^ n10852 ;
  assign n12358 = n12266 ^ n12265 ;
  assign n12362 = n12361 ^ n12358 ;
  assign n12673 = n11557 ^ n10179 ;
  assign n12674 = n12077 & n12673 ;
  assign n12675 = n12674 ^ n10179 ;
  assign n12622 = n11520 ^ n10191 ;
  assign n12623 = n12070 & ~n12622 ;
  assign n12624 = n12623 ^ n10191 ;
  assign n12387 = n10729 ^ n10013 ;
  assign n12388 = ~n11842 & n12387 ;
  assign n12389 = n12388 ^ n10013 ;
  assign n12391 = n12390 ^ n12389 ;
  assign n12392 = n11381 ^ n10711 ;
  assign n12393 = n11830 & ~n12392 ;
  assign n12394 = n12393 ^ n10711 ;
  assign n12395 = n12394 ^ n12344 ;
  assign n12449 = n12448 ^ n12398 ;
  assign n12450 = n12400 & n12449 ;
  assign n12451 = n12450 ^ n12399 ;
  assign n12452 = n12451 ^ n12394 ;
  assign n12453 = n12395 & ~n12452 ;
  assign n12454 = n12453 ^ n12344 ;
  assign n12455 = n12454 ^ n12389 ;
  assign n12456 = ~n12391 & n12455 ;
  assign n12457 = n12456 ^ n12390 ;
  assign n12384 = n11959 ^ x458 ;
  assign n12385 = n12384 ^ n11899 ;
  assign n12381 = n10734 ^ n10018 ;
  assign n12382 = n12011 & ~n12381 ;
  assign n12383 = n12382 ^ n10018 ;
  assign n12386 = n12385 ^ n12383 ;
  assign n12479 = n12457 ^ n12386 ;
  assign n12555 = n12479 ^ n9398 ;
  assign n12480 = n12454 ^ n12391 ;
  assign n12481 = n12480 ^ n9393 ;
  assign n12482 = n12451 ^ n12395 ;
  assign n12483 = n12482 ^ n10046 ;
  assign n12514 = n12513 ^ n12484 ;
  assign n12515 = n12485 & ~n12514 ;
  assign n12516 = n12515 ^ n9985 ;
  assign n12517 = n12516 ^ n12482 ;
  assign n12518 = ~n12483 & n12517 ;
  assign n12519 = n12518 ^ n10046 ;
  assign n12520 = n12519 ^ n12480 ;
  assign n12521 = n12481 & ~n12520 ;
  assign n12522 = n12521 ^ n9393 ;
  assign n12556 = n12555 ^ n12522 ;
  assign n12536 = n12519 ^ n12481 ;
  assign n12551 = ~n12549 & n12550 ;
  assign n12552 = n12516 ^ n12483 ;
  assign n12553 = ~n12551 & n12552 ;
  assign n12554 = n12536 & ~n12553 ;
  assign n12606 = n12556 ^ n12554 ;
  assign n12562 = n12553 ^ n12536 ;
  assign n12563 = n12562 ^ x486 ;
  assign n12564 = n12552 ^ n12551 ;
  assign n12565 = n12564 ^ x487 ;
  assign n12567 = n12566 ^ x488 ;
  assign n12597 = n12596 ^ n12566 ;
  assign n12598 = n12567 & ~n12597 ;
  assign n12599 = n12598 ^ x488 ;
  assign n12600 = n12599 ^ n12564 ;
  assign n12601 = ~n12565 & n12600 ;
  assign n12602 = n12601 ^ x487 ;
  assign n12603 = n12602 ^ n12562 ;
  assign n12604 = n12563 & ~n12603 ;
  assign n12605 = n12604 ^ x486 ;
  assign n12607 = n12606 ^ n12605 ;
  assign n12608 = n12606 ^ x485 ;
  assign n12609 = ~n12607 & n12608 ;
  assign n12610 = n12609 ^ x485 ;
  assign n12611 = n12610 ^ x484 ;
  assign n12557 = ~n12554 & ~n12556 ;
  assign n12523 = n12522 ^ n12479 ;
  assign n12524 = n12522 ^ n9398 ;
  assign n12525 = n12523 & ~n12524 ;
  assign n12526 = n12525 ^ n9398 ;
  assign n12458 = n12457 ^ n12383 ;
  assign n12459 = n12386 & n12458 ;
  assign n12460 = n12459 ^ n12385 ;
  assign n12379 = n11965 ^ n11962 ;
  assign n12376 = n10748 ^ n10008 ;
  assign n12377 = ~n11340 & n12376 ;
  assign n12378 = n12377 ^ n10008 ;
  assign n12380 = n12379 ^ n12378 ;
  assign n12477 = n12460 ^ n12380 ;
  assign n12478 = n12477 ^ n9386 ;
  assign n12535 = n12526 ^ n12478 ;
  assign n12612 = n12557 ^ n12535 ;
  assign n12613 = n12612 ^ n12610 ;
  assign n12614 = n12611 & n12613 ;
  assign n12615 = n12614 ^ x484 ;
  assign n12558 = ~n12535 & ~n12557 ;
  assign n12527 = n12526 ^ n12477 ;
  assign n12528 = n12478 & n12527 ;
  assign n12529 = n12528 ^ n9386 ;
  assign n12461 = n12460 ^ n12378 ;
  assign n12462 = n12380 & ~n12461 ;
  assign n12463 = n12462 ^ n12379 ;
  assign n12371 = n12370 ^ n9997 ;
  assign n12372 = n12371 ^ n10756 ;
  assign n12373 = n12372 ^ n12370 ;
  assign n12374 = ~n11339 & ~n12373 ;
  assign n12375 = n12374 ^ n12371 ;
  assign n12475 = n12463 ^ n12375 ;
  assign n12476 = n12475 ^ n9384 ;
  assign n12534 = n12529 ^ n12476 ;
  assign n12561 = n12558 ^ n12534 ;
  assign n12616 = n12615 ^ n12561 ;
  assign n12617 = n12615 ^ x483 ;
  assign n12618 = ~n12616 & n12617 ;
  assign n12619 = n12618 ^ x483 ;
  assign n12620 = n12619 ^ x482 ;
  assign n12559 = ~n12534 & n12558 ;
  assign n12530 = n12529 ^ n12475 ;
  assign n12531 = ~n12476 & n12530 ;
  assign n12532 = n12531 ^ n9384 ;
  assign n12470 = n10724 ^ n10057 ;
  assign n12471 = ~n11358 & ~n12470 ;
  assign n12472 = n12471 ^ n10057 ;
  assign n12466 = n12464 ^ n12370 ;
  assign n12465 = n12464 ^ n12463 ;
  assign n12467 = n12466 ^ n12465 ;
  assign n12468 = ~n12375 & ~n12467 ;
  assign n12469 = n12468 ^ n12466 ;
  assign n12473 = n12472 ^ n12469 ;
  assign n12474 = n12473 ^ n9379 ;
  assign n12533 = n12532 ^ n12474 ;
  assign n12560 = n12559 ^ n12533 ;
  assign n12621 = n12620 ^ n12560 ;
  assign n12625 = n12624 ^ n12621 ;
  assign n12628 = n11407 ^ n10194 ;
  assign n12629 = ~n11569 & n12628 ;
  assign n12630 = n12629 ^ n10194 ;
  assign n12631 = n12612 ^ n12611 ;
  assign n12632 = n12630 & ~n12631 ;
  assign n12626 = n12561 ^ x483 ;
  assign n12627 = n12626 ^ n12615 ;
  assign n12633 = n12632 ^ n12627 ;
  assign n12634 = n12632 ^ n10772 ;
  assign n12635 = n12634 ^ n11453 ;
  assign n12636 = n12635 ^ n12632 ;
  assign n12637 = n11558 & n12636 ;
  assign n12638 = n12637 ^ n12634 ;
  assign n12639 = n12633 & ~n12638 ;
  assign n12640 = n12639 ^ n12632 ;
  assign n12641 = n12640 ^ n12621 ;
  assign n12642 = n12625 & ~n12641 ;
  assign n12643 = n12642 ^ n12624 ;
  assign n12366 = n11565 ^ n10181 ;
  assign n12367 = ~n11551 & ~n12366 ;
  assign n12368 = n12367 ^ n10181 ;
  assign n12644 = n12643 ^ n12368 ;
  assign n12664 = n12560 ^ x482 ;
  assign n12665 = n12619 ^ n12560 ;
  assign n12666 = n12664 & ~n12665 ;
  assign n12667 = n12666 ^ x482 ;
  assign n12668 = n12667 ^ x481 ;
  assign n12662 = ~n12533 & ~n12559 ;
  assign n12656 = n12532 ^ n12473 ;
  assign n12657 = n12532 ^ n9379 ;
  assign n12658 = n12656 & ~n12657 ;
  assign n12659 = n12658 ^ n9379 ;
  assign n12660 = n12659 ^ n8833 ;
  assign n12652 = n10211 ^ n10063 ;
  assign n12653 = n11338 & ~n12652 ;
  assign n12654 = n12653 ^ n10063 ;
  assign n12648 = n12646 ^ n12464 ;
  assign n12647 = n12646 ^ n12472 ;
  assign n12649 = n12648 ^ n12647 ;
  assign n12650 = n12469 & n12649 ;
  assign n12651 = n12650 ^ n12648 ;
  assign n12655 = n12654 ^ n12651 ;
  assign n12661 = n12660 ^ n12655 ;
  assign n12663 = n12662 ^ n12661 ;
  assign n12669 = n12668 ^ n12663 ;
  assign n12670 = n12669 ^ n12643 ;
  assign n12671 = ~n12644 & n12670 ;
  assign n12672 = n12671 ^ n12669 ;
  assign n12676 = n12675 ^ n12672 ;
  assign n12691 = n10204 ^ n10064 ;
  assign n12692 = n11394 & n12691 ;
  assign n12687 = n12654 ^ n12016 ;
  assign n12686 = n11976 ^ n11892 ;
  assign n12688 = n12687 ^ n12686 ;
  assign n12689 = n12688 ^ n8833 ;
  assign n12685 = x481 ^ x480 ;
  assign n12690 = n12689 ^ n12685 ;
  assign n12693 = n12692 ^ n12690 ;
  assign n12683 = n12654 ^ n12646 ;
  assign n12684 = ~n12651 & ~n12683 ;
  assign n12694 = n12693 ^ n12684 ;
  assign n12682 = n12661 & ~n12662 ;
  assign n12695 = n12694 ^ n12682 ;
  assign n12680 = n12667 ^ n12663 ;
  assign n12681 = n12668 & ~n12680 ;
  assign n12696 = n12695 ^ n12681 ;
  assign n12677 = n12659 ^ n12655 ;
  assign n12678 = n12655 ^ n8833 ;
  assign n12679 = n12677 & ~n12678 ;
  assign n12697 = n12696 ^ n12679 ;
  assign n12698 = n12697 ^ n12672 ;
  assign n12699 = n12676 & ~n12698 ;
  assign n12700 = n12699 ^ n12675 ;
  assign n12363 = n11553 ^ n10167 ;
  assign n12364 = ~n11544 & ~n12363 ;
  assign n12365 = n12364 ^ n10167 ;
  assign n12701 = n12700 ^ n12365 ;
  assign n12702 = n12216 ^ x511 ;
  assign n12703 = n12702 ^ n12700 ;
  assign n12704 = ~n12701 & ~n12703 ;
  assign n12705 = n12704 ^ n12702 ;
  assign n12706 = n12705 ^ n12358 ;
  assign n12707 = n12362 & n12706 ;
  assign n12708 = n12707 ^ n12361 ;
  assign n12710 = n12709 ^ n12708 ;
  assign n12711 = n12709 ^ n10961 ;
  assign n12712 = n12711 ^ n11655 ;
  assign n12713 = n12712 ^ n12709 ;
  assign n12714 = n12093 & n12713 ;
  assign n12715 = n12714 ^ n12711 ;
  assign n12716 = n12710 & ~n12715 ;
  assign n12717 = n12716 ^ n12709 ;
  assign n12718 = n12717 ^ n12355 ;
  assign n12719 = ~n12357 & n12718 ;
  assign n12720 = n12719 ^ n12356 ;
  assign n12721 = n12720 ^ n12348 ;
  assign n12722 = ~n12352 & n12721 ;
  assign n12723 = n12722 ^ n12351 ;
  assign n12785 = n12725 ^ n12723 ;
  assign n12786 = n12729 & n12785 ;
  assign n12787 = n12786 ^ n12728 ;
  assign n12882 = n12788 ^ n12787 ;
  assign n12883 = ~n12792 & ~n12882 ;
  assign n12884 = n12883 ^ n12791 ;
  assign n13000 = n12886 ^ n12884 ;
  assign n13001 = n12890 & ~n13000 ;
  assign n13002 = n13001 ^ n12889 ;
  assign n13006 = n13005 ^ n13002 ;
  assign n12935 = n12291 ^ x503 ;
  assign n12936 = n12935 ^ n12254 ;
  assign n13007 = n13005 ^ n12936 ;
  assign n13008 = n13006 & n13007 ;
  assign n13009 = n13008 ^ n12936 ;
  assign n13013 = n13012 ^ n13009 ;
  assign n13015 = n13014 ^ n13013 ;
  assign n13016 = n12999 & n13015 ;
  assign n13017 = n13016 ^ n13014 ;
  assign n12928 = n12300 ^ n12297 ;
  assign n13022 = n13020 ^ n12928 ;
  assign n13021 = n13020 ^ n13012 ;
  assign n13023 = n13022 ^ n13021 ;
  assign n13024 = ~n13017 & ~n13023 ;
  assign n13025 = n13024 ^ n13021 ;
  assign n12919 = n12302 ^ x500 ;
  assign n12920 = n12919 ^ n12250 ;
  assign n13026 = n13020 ^ n12920 ;
  assign n13027 = ~n13025 & n13026 ;
  assign n13029 = n13028 ^ n13027 ;
  assign n13030 = ~n12994 & n13029 ;
  assign n13031 = n13030 ^ n12993 ;
  assign n12906 = n12310 ^ n12309 ;
  assign n13032 = n13031 ^ n12906 ;
  assign n13033 = n12906 ^ n10996 ;
  assign n13034 = n13033 ^ n11703 ;
  assign n13035 = n13034 ^ n12906 ;
  assign n13036 = n12399 & ~n13035 ;
  assign n13037 = n13036 ^ n13033 ;
  assign n13038 = n13032 & ~n13037 ;
  assign n13039 = n13038 ^ n12906 ;
  assign n13040 = n13039 ^ n12899 ;
  assign n13041 = ~n12990 & n13040 ;
  assign n13042 = n13041 ^ n12989 ;
  assign n13043 = n13042 ^ n12982 ;
  assign n13044 = n12986 & n13043 ;
  assign n13045 = n13044 ^ n12985 ;
  assign n13047 = n13046 ^ n13045 ;
  assign n13048 = n13046 ^ n11186 ;
  assign n13049 = n13048 ^ n11822 ;
  assign n13050 = n13049 ^ n13046 ;
  assign n13051 = ~n12385 & ~n13050 ;
  assign n13052 = n13051 ^ n13048 ;
  assign n13053 = ~n13047 & n13052 ;
  assign n13054 = n13053 ^ n13046 ;
  assign n12325 = n12324 ^ x494 ;
  assign n12343 = n12342 ^ n12325 ;
  assign n13055 = n13054 ^ n12343 ;
  assign n13056 = n12343 ^ n11226 ;
  assign n13057 = n13056 ^ n11830 ;
  assign n13058 = n13057 ^ n12343 ;
  assign n13059 = ~n12379 & n13058 ;
  assign n13060 = n13059 ^ n13056 ;
  assign n13061 = ~n13055 & n13060 ;
  assign n13062 = n13061 ^ n12343 ;
  assign n13063 = n13062 ^ n12976 ;
  assign n13064 = ~n12980 & n13063 ;
  assign n13065 = n13064 ^ n12979 ;
  assign n13066 = n13065 ^ n12971 ;
  assign n13067 = n12975 & n13066 ;
  assign n13068 = n13067 ^ n12974 ;
  assign n12966 = n11339 ^ n10734 ;
  assign n12967 = n12686 & ~n12966 ;
  assign n12968 = n12967 ^ n10734 ;
  assign n12969 = n12968 ^ n12960 ;
  assign n12970 = n12969 ^ n12968 ;
  assign n13069 = n13068 ^ n12970 ;
  assign n13070 = n12965 & n13069 ;
  assign n13071 = n13070 ^ n12969 ;
  assign n13072 = n11358 ^ n10748 ;
  assign n13073 = ~n12040 & n13072 ;
  assign n13074 = n13073 ^ n10748 ;
  assign n13078 = n13074 ^ n12968 ;
  assign n13075 = n12589 ^ x490 ;
  assign n13076 = n13075 ^ n12569 ;
  assign n13077 = n13076 ^ n13074 ;
  assign n13079 = n13078 ^ n13077 ;
  assign n13080 = ~n13071 & n13079 ;
  assign n13081 = n13080 ^ n13078 ;
  assign n13082 = n12568 ^ x489 ;
  assign n13083 = n13082 ^ n12592 ;
  assign n13162 = n13083 ^ n13074 ;
  assign n13163 = ~n13081 & ~n13162 ;
  assign n13164 = n13163 ^ n13074 ;
  assign n13165 = n13164 ^ n10756 ;
  assign n13166 = n13165 ^ n11338 ;
  assign n13167 = n13166 ^ n13164 ;
  assign n13168 = ~n12050 & n13167 ;
  assign n13169 = n13168 ^ n13165 ;
  assign n13172 = n13171 ^ n13169 ;
  assign n13173 = n13172 ^ n9997 ;
  assign n13084 = n13083 ^ n13081 ;
  assign n13085 = n13084 ^ n10008 ;
  assign n13086 = n13076 ^ n13071 ;
  assign n13087 = n13086 ^ n10018 ;
  assign n13088 = n13068 ^ n12965 ;
  assign n13089 = n13088 ^ n10013 ;
  assign n13091 = n13062 ^ n12980 ;
  assign n13092 = n13091 ^ n10413 ;
  assign n13093 = n13060 ^ n13054 ;
  assign n13094 = n13093 ^ n10216 ;
  assign n13138 = n13052 ^ n13045 ;
  assign n13129 = n13039 ^ n12990 ;
  assign n13096 = n13037 ^ n13031 ;
  assign n13097 = n13096 ^ n10383 ;
  assign n13098 = n13029 ^ n12913 ;
  assign n13099 = n13098 ^ n10223 ;
  assign n13100 = n13025 ^ n12920 ;
  assign n13101 = n13100 ^ n10227 ;
  assign n13115 = n13017 ^ n12928 ;
  assign n13102 = n13009 ^ n12999 ;
  assign n13103 = n13102 ^ n10350 ;
  assign n13104 = n13007 ^ n13002 ;
  assign n13105 = n13104 ^ n10236 ;
  assign n12891 = n12890 ^ n12884 ;
  assign n12892 = n12891 ^ n10245 ;
  assign n12793 = n12792 ^ n12787 ;
  assign n12794 = n12793 ^ n10341 ;
  assign n12730 = n12729 ^ n12723 ;
  assign n12731 = n12730 ^ n9605 ;
  assign n12732 = n12720 ^ n12352 ;
  assign n12733 = n12732 ^ n10174 ;
  assign n12774 = n12717 ^ n12357 ;
  assign n12734 = n12715 ^ n12708 ;
  assign n12735 = n12734 ^ n10187 ;
  assign n12737 = n12702 ^ n12365 ;
  assign n12738 = n12737 ^ n12700 ;
  assign n12739 = n12738 ^ n10193 ;
  assign n12740 = n12697 ^ n12675 ;
  assign n12741 = n12740 ^ n12672 ;
  assign n12742 = n12741 ^ n10200 ;
  assign n12745 = n12640 ^ n12625 ;
  assign n12746 = n12745 ^ n10301 ;
  assign n12749 = n12638 ^ n12627 ;
  assign n12747 = n12631 ^ n12630 ;
  assign n12748 = n10127 & ~n12747 ;
  assign n12750 = n12749 ^ n12748 ;
  assign n12751 = n12749 ^ n10284 ;
  assign n12752 = n12750 & n12751 ;
  assign n12753 = n12752 ^ n10284 ;
  assign n12754 = n12753 ^ n12745 ;
  assign n12755 = ~n12746 & n12754 ;
  assign n12756 = n12755 ^ n10301 ;
  assign n12743 = n12669 ^ n12368 ;
  assign n12744 = n12743 ^ n12643 ;
  assign n12757 = n12756 ^ n12744 ;
  assign n12758 = n12756 ^ n10207 ;
  assign n12759 = n12757 & ~n12758 ;
  assign n12760 = n12759 ^ n10207 ;
  assign n12761 = n12760 ^ n12741 ;
  assign n12762 = ~n12742 & ~n12761 ;
  assign n12763 = n12762 ^ n10200 ;
  assign n12764 = n12763 ^ n12738 ;
  assign n12765 = ~n12739 & ~n12764 ;
  assign n12766 = n12765 ^ n10193 ;
  assign n12736 = n12705 ^ n12362 ;
  assign n12767 = n12766 ^ n12736 ;
  assign n12768 = n12766 ^ n10317 ;
  assign n12769 = n12767 & ~n12768 ;
  assign n12770 = n12769 ^ n10317 ;
  assign n12771 = n12770 ^ n12734 ;
  assign n12772 = ~n12735 & ~n12771 ;
  assign n12773 = n12772 ^ n10187 ;
  assign n12775 = n12774 ^ n12773 ;
  assign n12776 = n12774 ^ n10182 ;
  assign n12777 = n12775 & n12776 ;
  assign n12778 = n12777 ^ n10182 ;
  assign n12779 = n12778 ^ n12732 ;
  assign n12780 = n12733 & ~n12779 ;
  assign n12781 = n12780 ^ n10174 ;
  assign n12782 = n12781 ^ n12730 ;
  assign n12783 = ~n12731 & n12782 ;
  assign n12784 = n12783 ^ n9605 ;
  assign n12879 = n12793 ^ n12784 ;
  assign n12880 = ~n12794 & n12879 ;
  assign n12881 = n12880 ^ n10341 ;
  assign n13106 = n12891 ^ n12881 ;
  assign n13107 = ~n12892 & n13106 ;
  assign n13108 = n13107 ^ n10245 ;
  assign n13109 = n13108 ^ n13104 ;
  assign n13110 = ~n13105 & n13109 ;
  assign n13111 = n13110 ^ n10236 ;
  assign n13112 = n13111 ^ n13102 ;
  assign n13113 = ~n13103 & ~n13112 ;
  assign n13114 = n13113 ^ n10350 ;
  assign n13116 = n13115 ^ n13114 ;
  assign n13117 = n13115 ^ n10229 ;
  assign n13118 = ~n13116 & n13117 ;
  assign n13119 = n13118 ^ n10229 ;
  assign n13120 = n13119 ^ n13100 ;
  assign n13121 = n13101 & ~n13120 ;
  assign n13122 = n13121 ^ n10227 ;
  assign n13123 = n13122 ^ n13098 ;
  assign n13124 = n13099 & ~n13123 ;
  assign n13125 = n13124 ^ n10223 ;
  assign n13126 = n13125 ^ n13096 ;
  assign n13127 = n13097 & ~n13126 ;
  assign n13128 = n13127 ^ n10383 ;
  assign n13130 = n13129 ^ n13128 ;
  assign n13131 = n13129 ^ n10388 ;
  assign n13132 = ~n13130 & n13131 ;
  assign n13133 = n13132 ^ n10388 ;
  assign n13095 = n13042 ^ n12986 ;
  assign n13134 = n13133 ^ n13095 ;
  assign n13135 = n13133 ^ n10218 ;
  assign n13136 = n13134 & n13135 ;
  assign n13137 = n13136 ^ n10218 ;
  assign n13139 = n13138 ^ n13137 ;
  assign n13140 = n13138 ^ n10402 ;
  assign n13141 = ~n13139 & ~n13140 ;
  assign n13142 = n13141 ^ n10402 ;
  assign n13143 = n13142 ^ n13093 ;
  assign n13144 = n13094 & ~n13143 ;
  assign n13145 = n13144 ^ n10216 ;
  assign n13146 = n13145 ^ n13091 ;
  assign n13147 = ~n13092 & ~n13146 ;
  assign n13148 = n13147 ^ n10413 ;
  assign n13090 = n13065 ^ n12975 ;
  assign n13149 = n13148 ^ n13090 ;
  assign n13150 = n13148 ^ n10711 ;
  assign n13151 = ~n13149 & n13150 ;
  assign n13152 = n13151 ^ n10711 ;
  assign n13153 = n13152 ^ n13088 ;
  assign n13154 = n13089 & n13153 ;
  assign n13155 = n13154 ^ n10013 ;
  assign n13156 = n13155 ^ n13086 ;
  assign n13157 = n13087 & ~n13156 ;
  assign n13158 = n13157 ^ n10018 ;
  assign n13159 = n13158 ^ n13084 ;
  assign n13160 = n13085 & ~n13159 ;
  assign n13161 = n13160 ^ n10008 ;
  assign n13306 = n13172 ^ n13161 ;
  assign n13307 = n13173 & ~n13306 ;
  assign n13308 = n13307 ^ n9997 ;
  assign n13301 = n11394 ^ n10724 ;
  assign n13302 = n12038 & ~n13301 ;
  assign n13303 = n13302 ^ n10724 ;
  assign n13295 = n12599 ^ n12565 ;
  assign n13297 = n13295 ^ n13164 ;
  assign n13296 = n13295 ^ n13171 ;
  assign n13298 = n13297 ^ n13296 ;
  assign n13299 = ~n13169 & ~n13298 ;
  assign n13300 = n13299 ^ n13297 ;
  assign n13304 = n13303 ^ n13300 ;
  assign n13305 = n13304 ^ n10057 ;
  assign n13309 = n13308 ^ n13305 ;
  assign n13174 = n13173 ^ n13161 ;
  assign n13175 = n13158 ^ n13085 ;
  assign n13176 = n13142 ^ n13094 ;
  assign n13177 = n13140 ^ n13137 ;
  assign n13178 = n13095 ^ n10218 ;
  assign n13179 = n13178 ^ n13133 ;
  assign n13180 = n13131 ^ n13128 ;
  assign n13181 = n13111 ^ n13103 ;
  assign n13182 = n13108 ^ n13105 ;
  assign n12795 = n12794 ^ n12784 ;
  assign n12796 = n12778 ^ n12733 ;
  assign n12797 = n12776 ^ n12773 ;
  assign n12798 = n12736 ^ n10317 ;
  assign n12799 = n12798 ^ n12766 ;
  assign n12800 = n12747 ^ n10127 ;
  assign n12801 = n12748 ^ n10284 ;
  assign n12802 = n12801 ^ n12749 ;
  assign n12803 = ~n12800 & n12802 ;
  assign n12804 = n12753 ^ n12746 ;
  assign n12805 = n12803 & n12804 ;
  assign n12806 = n12744 ^ n10207 ;
  assign n12807 = n12806 ^ n12756 ;
  assign n12808 = ~n12805 & n12807 ;
  assign n12809 = n12760 ^ n12742 ;
  assign n12810 = n12808 & n12809 ;
  assign n12811 = n12763 ^ n12739 ;
  assign n12812 = ~n12810 & n12811 ;
  assign n12813 = n12799 & n12812 ;
  assign n12814 = n12770 ^ n12735 ;
  assign n12815 = ~n12813 & ~n12814 ;
  assign n12816 = ~n12797 & n12815 ;
  assign n12817 = ~n12796 & ~n12816 ;
  assign n12818 = n12781 ^ n12731 ;
  assign n12819 = n12817 & n12818 ;
  assign n12878 = ~n12795 & ~n12819 ;
  assign n12893 = n12892 ^ n12881 ;
  assign n13183 = n12878 & ~n12893 ;
  assign n13184 = ~n13182 & n13183 ;
  assign n13185 = ~n13181 & n13184 ;
  assign n13186 = n13117 ^ n13114 ;
  assign n13187 = ~n13185 & n13186 ;
  assign n13188 = n13119 ^ n13101 ;
  assign n13189 = n13187 & n13188 ;
  assign n13190 = n13122 ^ n13099 ;
  assign n13191 = ~n13189 & ~n13190 ;
  assign n13192 = n13125 ^ n13097 ;
  assign n13193 = ~n13191 & n13192 ;
  assign n13194 = n13180 & n13193 ;
  assign n13195 = ~n13179 & n13194 ;
  assign n13196 = ~n13177 & n13195 ;
  assign n13197 = ~n13176 & n13196 ;
  assign n13198 = n13145 ^ n13092 ;
  assign n13199 = ~n13197 & ~n13198 ;
  assign n13200 = n13090 ^ n10711 ;
  assign n13201 = n13200 ^ n13148 ;
  assign n13202 = ~n13199 & n13201 ;
  assign n13203 = n13152 ^ n13089 ;
  assign n13204 = ~n13202 & ~n13203 ;
  assign n13205 = n13155 ^ n13087 ;
  assign n13206 = ~n13204 & ~n13205 ;
  assign n13207 = n13175 & ~n13206 ;
  assign n13294 = n13174 & n13207 ;
  assign n13310 = n13309 ^ n13294 ;
  assign n13311 = n13310 ^ n1796 ;
  assign n13348 = ~n13294 & n13309 ;
  assign n13342 = n12602 ^ x486 ;
  assign n13343 = n13342 ^ n12562 ;
  assign n13344 = n13343 ^ n13295 ;
  assign n13340 = n13303 ^ n13295 ;
  assign n13341 = n13300 & n13340 ;
  assign n13345 = n13344 ^ n13341 ;
  assign n13337 = n10984 ^ n10211 ;
  assign n13338 = n12029 & n13337 ;
  assign n13339 = n13338 ^ n10211 ;
  assign n13346 = n13345 ^ n13339 ;
  assign n13332 = n13308 ^ n13304 ;
  assign n13333 = n13308 ^ n10057 ;
  assign n13334 = ~n13332 & ~n13333 ;
  assign n13335 = n13334 ^ n10057 ;
  assign n13336 = n13335 ^ n10063 ;
  assign n13347 = n13346 ^ n13336 ;
  assign n13349 = n13348 ^ n13347 ;
  assign n13350 = n13349 ^ n1796 ;
  assign n13351 = n13350 ^ n13349 ;
  assign n13209 = n13206 ^ n13175 ;
  assign n13210 = n13209 ^ n2459 ;
  assign n13211 = n13205 ^ n13204 ;
  assign n13212 = n13211 ^ n2444 ;
  assign n13214 = n13201 ^ n13199 ;
  assign n13215 = n13214 ^ n2557 ;
  assign n13216 = n13198 ^ n13197 ;
  assign n13217 = n13216 ^ n2551 ;
  assign n13218 = n13196 ^ n13176 ;
  assign n13219 = n13218 ^ n1395 ;
  assign n13221 = n13194 ^ n13179 ;
  assign n13222 = n13221 ^ n1154 ;
  assign n13224 = n13192 ^ n13191 ;
  assign n13225 = n13224 ^ n974 ;
  assign n13226 = n13190 ^ n13189 ;
  assign n828 = x431 ^ x79 ;
  assign n829 = n828 ^ x271 ;
  assign n830 = n829 ^ x15 ;
  assign n13227 = n13226 ^ n830 ;
  assign n13228 = n13188 ^ n13187 ;
  assign n13229 = n13228 ^ n833 ;
  assign n13247 = n13228 ^ n737 ;
  assign n13230 = n13186 ^ n13185 ;
  assign n13231 = n13230 ^ n737 ;
  assign n13232 = n13184 ^ n13181 ;
  assign n13233 = n13232 ^ n678 ;
  assign n13241 = n13232 ^ n666 ;
  assign n13234 = n13183 ^ n13182 ;
  assign n13235 = n13234 ^ n666 ;
  assign n12894 = n12893 ^ n12878 ;
  assign n12895 = n12894 ^ n1511 ;
  assign n12820 = n12819 ^ n12795 ;
  assign n12821 = n12820 ^ n1511 ;
  assign n12822 = n12818 ^ n12817 ;
  assign n12823 = n12822 ^ n1505 ;
  assign n12824 = n12816 ^ n12796 ;
  assign n12825 = n12824 ^ n515 ;
  assign n12828 = n12815 ^ n12797 ;
  assign n12829 = n12828 ^ n2914 ;
  assign n12830 = n12814 ^ n12813 ;
  assign n12831 = n12830 ^ n566 ;
  assign n12835 = n12809 ^ n12808 ;
  assign n12836 = n12835 ^ n2154 ;
  assign n12837 = n12807 ^ n12805 ;
  assign n12838 = n12837 ^ n2062 ;
  assign n12839 = n12804 ^ n12803 ;
  assign n12840 = n12839 ^ n2042 ;
  assign n1869 = x416 ^ x64 ;
  assign n1870 = n1869 ^ x256 ;
  assign n1871 = n1870 ^ x0 ;
  assign n12843 = n1871 & n12800 ;
  assign n12844 = n12843 ^ n2046 ;
  assign n12845 = n12802 ^ n12800 ;
  assign n12846 = n12845 ^ n12843 ;
  assign n12847 = n12844 & n12846 ;
  assign n12848 = n12847 ^ n2046 ;
  assign n12841 = n12837 ^ n2042 ;
  assign n12842 = n12841 ^ n12837 ;
  assign n12849 = n12848 ^ n12842 ;
  assign n12850 = n12840 & n12849 ;
  assign n12851 = n12850 ^ n12841 ;
  assign n12852 = n12838 & ~n12851 ;
  assign n12853 = n12852 ^ n2062 ;
  assign n12854 = n12853 ^ n2154 ;
  assign n12855 = ~n12836 & n12854 ;
  assign n12856 = n12855 ^ n2154 ;
  assign n12857 = n12856 ^ n1457 ;
  assign n12858 = n12811 ^ n12810 ;
  assign n12859 = n12858 ^ n12856 ;
  assign n12860 = n12857 & n12859 ;
  assign n12861 = n12860 ^ n1457 ;
  assign n12834 = n12812 ^ n12799 ;
  assign n12862 = n12861 ^ n12834 ;
  assign n12863 = n12861 ^ n2291 ;
  assign n12864 = ~n12862 & n12863 ;
  assign n12865 = n12864 ^ n2291 ;
  assign n12832 = n12828 ^ n566 ;
  assign n12833 = n12832 ^ n12828 ;
  assign n12866 = n12865 ^ n12833 ;
  assign n12867 = ~n12831 & n12866 ;
  assign n12868 = n12867 ^ n12832 ;
  assign n12869 = n12829 & ~n12868 ;
  assign n12870 = n12869 ^ n2914 ;
  assign n12826 = n12822 ^ n515 ;
  assign n12827 = n12826 ^ n12822 ;
  assign n12871 = n12870 ^ n12827 ;
  assign n12872 = n12825 & n12871 ;
  assign n12873 = n12872 ^ n12826 ;
  assign n12874 = n12823 & ~n12873 ;
  assign n12875 = n12874 ^ n1505 ;
  assign n12876 = n12875 ^ n1511 ;
  assign n12877 = ~n12821 & n12876 ;
  assign n12896 = n12895 ^ n12877 ;
  assign n13236 = n12894 ^ n660 ;
  assign n13237 = ~n12896 & n13236 ;
  assign n13238 = n13237 ^ n660 ;
  assign n13239 = n13238 ^ n666 ;
  assign n13240 = n13235 & n13239 ;
  assign n13242 = n13241 ^ n13240 ;
  assign n13243 = n13233 & n13242 ;
  assign n13244 = n13243 ^ n13232 ;
  assign n13245 = n13244 ^ n737 ;
  assign n13246 = ~n13231 & n13245 ;
  assign n13248 = n13247 ^ n13246 ;
  assign n13249 = n13229 & ~n13248 ;
  assign n13250 = n13249 ^ n833 ;
  assign n13251 = n13250 ^ n13226 ;
  assign n13252 = ~n13227 & n13251 ;
  assign n13253 = n13252 ^ n830 ;
  assign n13254 = n13253 ^ n13224 ;
  assign n13255 = ~n13225 & n13254 ;
  assign n13256 = n13255 ^ n974 ;
  assign n13223 = n13193 ^ n13180 ;
  assign n13257 = n13256 ^ n13223 ;
  assign n13258 = n13221 ^ n1203 ;
  assign n13259 = n13258 ^ n13221 ;
  assign n13260 = n13259 ^ n13223 ;
  assign n13261 = ~n13257 & n13260 ;
  assign n13262 = n13261 ^ n13258 ;
  assign n13263 = ~n13222 & n13262 ;
  assign n13264 = n13263 ^ n1154 ;
  assign n13220 = n13195 ^ n13177 ;
  assign n13265 = n13264 ^ n13220 ;
  assign n13266 = n13218 ^ n1359 ;
  assign n13267 = n13266 ^ n13218 ;
  assign n13268 = n13267 ^ n13220 ;
  assign n13269 = n13265 & ~n13268 ;
  assign n13270 = n13269 ^ n13266 ;
  assign n13271 = ~n13219 & n13270 ;
  assign n13272 = n13271 ^ n1395 ;
  assign n13273 = n13272 ^ n13216 ;
  assign n13274 = ~n13217 & n13273 ;
  assign n13275 = n13274 ^ n2551 ;
  assign n13276 = n13275 ^ n13214 ;
  assign n13277 = ~n13215 & n13276 ;
  assign n13278 = n13277 ^ n2557 ;
  assign n13213 = n13203 ^ n13202 ;
  assign n13279 = n13278 ^ n13213 ;
  assign n13280 = n13211 ^ n2484 ;
  assign n13281 = n13280 ^ n13211 ;
  assign n13282 = n13281 ^ n13213 ;
  assign n13283 = n13279 & ~n13282 ;
  assign n13284 = n13283 ^ n13280 ;
  assign n13285 = n13212 & ~n13284 ;
  assign n13286 = n13285 ^ n2444 ;
  assign n13287 = n13286 ^ n13209 ;
  assign n13288 = n13210 & ~n13287 ;
  assign n13289 = n13288 ^ n2459 ;
  assign n13208 = n13207 ^ n13174 ;
  assign n13290 = n13289 ^ n13208 ;
  assign n13291 = n13289 ^ n1805 ;
  assign n13292 = n13290 & n13291 ;
  assign n13293 = n13292 ^ n1805 ;
  assign n13352 = n13351 ^ n13293 ;
  assign n13353 = ~n13311 & n13352 ;
  assign n13354 = n13353 ^ n13350 ;
  assign n13355 = n13354 ^ n1785 ;
  assign n13357 = n13355 ^ n11565 ;
  assign n13358 = n13357 ^ n11544 ;
  assign n13359 = n13358 ^ n13355 ;
  assign n13360 = n12356 & n13359 ;
  assign n13361 = n13360 ^ n13357 ;
  assign n13312 = n13311 ^ n13293 ;
  assign n12956 = n12077 ^ n11520 ;
  assign n12957 = n12709 & ~n12956 ;
  assign n12958 = n12957 ^ n11520 ;
  assign n13313 = n13312 ^ n12958 ;
  assign n13316 = n13286 ^ n13210 ;
  assign n13317 = n12070 ^ n11407 ;
  assign n13318 = ~n12702 & n13317 ;
  assign n13319 = n13318 ^ n11407 ;
  assign n13320 = n13316 & n13319 ;
  assign n13314 = n13208 ^ n1805 ;
  assign n13315 = n13314 ^ n13289 ;
  assign n13321 = n13320 ^ n13315 ;
  assign n13322 = n13320 ^ n11453 ;
  assign n13323 = n13322 ^ n11551 ;
  assign n13324 = n13323 ^ n13320 ;
  assign n13325 = n12358 & n13324 ;
  assign n13326 = n13325 ^ n13322 ;
  assign n13327 = ~n13321 & ~n13326 ;
  assign n13328 = n13327 ^ n13320 ;
  assign n13329 = n13328 ^ n12958 ;
  assign n13330 = n13313 & n13329 ;
  assign n13331 = n13330 ^ n13312 ;
  assign n13482 = n13361 ^ n13331 ;
  assign n13483 = n13482 ^ n10181 ;
  assign n13491 = n13328 ^ n13313 ;
  assign n13486 = n13326 ^ n13315 ;
  assign n13484 = n13319 ^ n13316 ;
  assign n13485 = n10194 & n13484 ;
  assign n13487 = n13486 ^ n13485 ;
  assign n13488 = n13486 ^ n10772 ;
  assign n13489 = ~n13487 & ~n13488 ;
  assign n13490 = n13489 ^ n10772 ;
  assign n13492 = n13491 ^ n13490 ;
  assign n13493 = n13491 ^ n10191 ;
  assign n13494 = n13492 & n13493 ;
  assign n13495 = n13494 ^ n10191 ;
  assign n13496 = n13495 ^ n13482 ;
  assign n13497 = ~n13483 & n13496 ;
  assign n13498 = n13497 ^ n10181 ;
  assign n13381 = n13347 & n13348 ;
  assign n13374 = n12608 ^ n12605 ;
  assign n13375 = n13374 ^ n12691 ;
  assign n13376 = n13375 ^ n13339 ;
  assign n13377 = n13376 ^ n10063 ;
  assign n3066 = x417 ^ x65 ;
  assign n3067 = n3066 ^ x257 ;
  assign n3068 = n3067 ^ x1 ;
  assign n13378 = n13377 ^ n3068 ;
  assign n13372 = n10982 ^ n10204 ;
  assign n13373 = n12024 & n13372 ;
  assign n13379 = n13378 ^ n13373 ;
  assign n13370 = n13343 ^ n13339 ;
  assign n13371 = n13345 & n13370 ;
  assign n13380 = n13379 ^ n13371 ;
  assign n13382 = n13381 ^ n13380 ;
  assign n13368 = n13349 ^ n1785 ;
  assign n13369 = ~n13354 & ~n13368 ;
  assign n13383 = n13382 ^ n13369 ;
  assign n13365 = n13346 ^ n10063 ;
  assign n13366 = n13346 ^ n13335 ;
  assign n13367 = n13365 & n13366 ;
  assign n13384 = n13383 ^ n13367 ;
  assign n12952 = n11557 ^ n11537 ;
  assign n12953 = ~n12348 & ~n12952 ;
  assign n12954 = n12953 ^ n11557 ;
  assign n13363 = n13355 ^ n12954 ;
  assign n13356 = n13355 ^ n13331 ;
  assign n13362 = n13356 & n13361 ;
  assign n13364 = n13363 ^ n13362 ;
  assign n13480 = n13384 ^ n13364 ;
  assign n13481 = n13480 ^ n10179 ;
  assign n13556 = n13498 ^ n13481 ;
  assign n13557 = n13485 ^ n10772 ;
  assign n13558 = n13557 ^ n13486 ;
  assign n13559 = n13484 ^ n10194 ;
  assign n13560 = ~n13558 & n13559 ;
  assign n13561 = n13493 ^ n13490 ;
  assign n13562 = n13560 & ~n13561 ;
  assign n13563 = n13495 ^ n13483 ;
  assign n13564 = ~n13562 & n13563 ;
  assign n13565 = n13556 & n13564 ;
  assign n13385 = n13384 ^ n12954 ;
  assign n13386 = ~n13364 & n13385 ;
  assign n12947 = n12093 ^ n11553 ;
  assign n12948 = ~n12725 & ~n12947 ;
  assign n12949 = n12948 ^ n11553 ;
  assign n12955 = n12954 ^ n12949 ;
  assign n13387 = n13386 ^ n12955 ;
  assign n12950 = n12800 ^ n1871 ;
  assign n13479 = n13387 ^ n12950 ;
  assign n13554 = n13479 ^ n10167 ;
  assign n13499 = n13498 ^ n13480 ;
  assign n13500 = ~n13481 & n13499 ;
  assign n13501 = n13500 ^ n10179 ;
  assign n13555 = n13554 ^ n13501 ;
  assign n13657 = n13565 ^ n13555 ;
  assign n13743 = n13657 ^ n2258 ;
  assign n13658 = n13564 ^ n13556 ;
  assign n13659 = n13658 ^ n2075 ;
  assign n13660 = n13563 ^ n13562 ;
  assign n13661 = n13660 ^ n2244 ;
  assign n1972 = x478 ^ x126 ;
  assign n1973 = n1972 ^ x318 ;
  assign n1974 = n1973 ^ x62 ;
  assign n13672 = n13660 ^ n1974 ;
  assign n13662 = n13561 ^ n13560 ;
  assign n13663 = n13662 ^ n1974 ;
  assign n1901 = x448 ^ x96 ;
  assign n1902 = n1901 ^ x288 ;
  assign n1903 = n1902 ^ x32 ;
  assign n13664 = n1903 & ~n13559 ;
  assign n1907 = x479 ^ x127 ;
  assign n1908 = n1907 ^ x319 ;
  assign n1909 = n1908 ^ x63 ;
  assign n13665 = n13664 ^ n1909 ;
  assign n13666 = n13559 ^ n13558 ;
  assign n13667 = n13666 ^ n13664 ;
  assign n13668 = ~n13665 & ~n13667 ;
  assign n13669 = n13668 ^ n13666 ;
  assign n13670 = n13669 ^ n1974 ;
  assign n13671 = ~n13663 & ~n13670 ;
  assign n13673 = n13672 ^ n13671 ;
  assign n13674 = n13661 & ~n13673 ;
  assign n13675 = n13674 ^ n2244 ;
  assign n13676 = n13675 ^ n2075 ;
  assign n13677 = ~n13659 & n13676 ;
  assign n13678 = n13677 ^ n2075 ;
  assign n13744 = n13743 ^ n13678 ;
  assign n13769 = n13223 ^ n1203 ;
  assign n13770 = n13769 ^ n13256 ;
  assign n13765 = n12040 ^ n11340 ;
  assign n13766 = n13343 & n13765 ;
  assign n13767 = n13766 ^ n11340 ;
  assign n13808 = n13770 ^ n13767 ;
  assign n13771 = n13770 ^ n12011 ;
  assign n13772 = n13771 ^ n12686 ;
  assign n13773 = n13772 ^ n13770 ;
  assign n13774 = ~n13295 & n13773 ;
  assign n13775 = n13774 ^ n13771 ;
  assign n13776 = n13253 ^ n13225 ;
  assign n13777 = n13776 ^ n11842 ;
  assign n13778 = n13777 ^ n12646 ;
  assign n13779 = n13778 ^ n13776 ;
  assign n13780 = n13171 & ~n13779 ;
  assign n13781 = n13780 ^ n13777 ;
  assign n13794 = n13250 ^ n13227 ;
  assign n13785 = n13248 ^ n833 ;
  assign n13594 = n13242 ^ n678 ;
  assign n13595 = n13594 ^ n11713 ;
  assign n13596 = n13595 ^ n12385 ;
  assign n13597 = n13596 ^ n13594 ;
  assign n13598 = ~n12971 & ~n13597 ;
  assign n13599 = n13598 ^ n13595 ;
  assign n13455 = n12390 ^ n11703 ;
  assign n13456 = ~n12976 & ~n13455 ;
  assign n13457 = n13456 ^ n11703 ;
  assign n13454 = n13238 ^ n13235 ;
  assign n13458 = n13457 ^ n13454 ;
  assign n12897 = n12896 ^ n660 ;
  assign n12345 = n12344 ^ n11571 ;
  assign n12346 = ~n12343 & n12345 ;
  assign n12347 = n12346 ^ n12344 ;
  assign n12898 = n12897 ^ n12347 ;
  assign n12900 = n12870 ^ n12825 ;
  assign n12901 = n12900 ^ n12407 ;
  assign n12902 = n12901 ^ n11587 ;
  assign n12903 = n12902 ^ n12900 ;
  assign n12904 = ~n12899 & ~n12903 ;
  assign n12905 = n12904 ^ n12901 ;
  assign n13429 = n12402 ^ n11593 ;
  assign n13430 = ~n12982 & ~n13429 ;
  assign n13431 = n13430 ^ n12402 ;
  assign n13432 = n13431 ^ n12900 ;
  assign n12907 = n12868 ^ n2914 ;
  assign n12908 = n12907 ^ n12413 ;
  assign n12909 = n12908 ^ n11598 ;
  assign n12910 = n12909 ^ n12907 ;
  assign n12911 = n12906 & ~n12910 ;
  assign n12912 = n12911 ^ n12908 ;
  assign n12917 = n12865 ^ n12831 ;
  assign n12914 = n12422 ^ n10974 ;
  assign n12915 = n12913 & n12914 ;
  assign n12916 = n12915 ^ n10974 ;
  assign n12918 = n12917 ^ n12916 ;
  assign n12921 = n12834 ^ n2291 ;
  assign n12922 = n12921 ^ n12861 ;
  assign n12924 = n12922 ^ n11607 ;
  assign n12923 = n12922 ^ n12433 ;
  assign n12925 = n12924 ^ n12923 ;
  assign n12926 = ~n12920 & n12925 ;
  assign n12927 = n12926 ^ n12924 ;
  assign n13420 = n12922 ^ n12916 ;
  assign n12932 = n12858 ^ n1457 ;
  assign n12933 = n12932 ^ n12856 ;
  assign n12929 = n12337 ^ n11612 ;
  assign n12930 = ~n12928 & ~n12929 ;
  assign n12931 = n12930 ^ n11612 ;
  assign n12934 = n12933 ^ n12931 ;
  assign n12945 = n12851 ^ n2062 ;
  assign n12937 = n12118 ^ n11539 ;
  assign n12938 = ~n12936 & n12937 ;
  assign n12939 = n12938 ^ n11539 ;
  assign n12946 = n12945 ^ n12939 ;
  assign n13389 = n12845 ^ n12844 ;
  assign n13390 = n13389 ^ n12950 ;
  assign n12951 = n12950 ^ n12949 ;
  assign n13388 = ~n12951 & n13387 ;
  assign n13391 = n13390 ^ n13388 ;
  assign n13397 = n12103 ^ n11546 ;
  assign n13398 = ~n12788 & n13397 ;
  assign n13399 = n13398 ^ n11546 ;
  assign n13392 = n11655 ^ n11531 ;
  assign n13393 = n12886 & n13392 ;
  assign n13394 = n13393 ^ n11655 ;
  assign n13395 = n13394 ^ n13389 ;
  assign n13396 = n13395 ^ n13394 ;
  assign n13400 = n13399 ^ n13396 ;
  assign n13401 = ~n13391 & ~n13400 ;
  assign n13402 = n13401 ^ n13395 ;
  assign n13405 = n13394 ^ n12939 ;
  assign n13403 = n12848 ^ n12840 ;
  assign n13404 = n13403 ^ n12939 ;
  assign n13406 = n13405 ^ n13404 ;
  assign n13407 = n13402 & ~n13406 ;
  assign n13408 = n13407 ^ n13405 ;
  assign n13409 = n12946 & ~n13408 ;
  assign n12941 = n12197 ^ n11533 ;
  assign n12942 = ~n12940 & n12941 ;
  assign n12943 = n12942 ^ n11533 ;
  assign n12944 = n12943 ^ n12939 ;
  assign n13410 = n13409 ^ n12944 ;
  assign n13413 = n12943 ^ n12931 ;
  assign n13411 = n12853 ^ n12836 ;
  assign n13412 = n13411 ^ n12931 ;
  assign n13414 = n13413 ^ n13412 ;
  assign n13415 = ~n13410 & ~n13414 ;
  assign n13416 = n13415 ^ n13412 ;
  assign n13417 = n12934 & ~n13416 ;
  assign n13418 = n13417 ^ n12933 ;
  assign n13419 = n13418 ^ n12916 ;
  assign n13421 = n13420 ^ n13419 ;
  assign n13422 = n12927 & ~n13421 ;
  assign n13423 = n13422 ^ n13420 ;
  assign n13424 = n12918 & n13423 ;
  assign n13425 = n13424 ^ n12917 ;
  assign n13426 = n13425 ^ n12907 ;
  assign n13427 = n12912 & ~n13426 ;
  assign n13428 = n13427 ^ n12907 ;
  assign n13433 = n13432 ^ n13428 ;
  assign n13434 = n13433 ^ n13431 ;
  assign n13435 = ~n12905 & n13434 ;
  assign n13436 = n13435 ^ n13432 ;
  assign n13440 = n12873 ^ n1505 ;
  assign n13437 = n12399 ^ n11585 ;
  assign n13438 = n13046 & ~n13437 ;
  assign n13439 = n13438 ^ n12399 ;
  assign n13441 = n13440 ^ n13439 ;
  assign n13442 = n13441 ^ n13431 ;
  assign n13443 = n13442 ^ n13439 ;
  assign n13444 = n13436 & ~n13443 ;
  assign n13445 = n13444 ^ n13441 ;
  assign n13447 = n12875 ^ n12821 ;
  assign n13448 = n13447 ^ n12347 ;
  assign n13446 = n13439 ^ n12347 ;
  assign n13449 = n13448 ^ n13446 ;
  assign n13450 = ~n13445 & ~n13449 ;
  assign n13451 = n13450 ^ n13448 ;
  assign n13452 = n12898 & n13451 ;
  assign n13453 = n13452 ^ n12897 ;
  assign n13591 = n13454 ^ n13453 ;
  assign n13592 = ~n13458 & ~n13591 ;
  assign n13593 = n13592 ^ n13457 ;
  assign n13613 = n13594 ^ n13593 ;
  assign n13614 = n13599 & ~n13613 ;
  assign n13609 = n12379 ^ n11719 ;
  assign n13610 = ~n12960 & n13609 ;
  assign n13611 = n13610 ^ n11719 ;
  assign n13612 = n13611 ^ n13594 ;
  assign n13615 = n13614 ^ n13612 ;
  assign n13616 = n13244 ^ n13231 ;
  assign n13782 = n13616 ^ n13611 ;
  assign n13783 = n13615 & n13782 ;
  assign n13784 = n13783 ^ n13616 ;
  assign n13786 = n13785 ^ n13784 ;
  assign n13787 = n13785 ^ n11822 ;
  assign n13788 = n13787 ^ n12370 ;
  assign n13789 = n13788 ^ n13785 ;
  assign n13790 = n13076 & n13789 ;
  assign n13791 = n13790 ^ n13787 ;
  assign n13792 = ~n13786 & n13791 ;
  assign n13793 = n13792 ^ n13785 ;
  assign n13795 = n13794 ^ n13793 ;
  assign n13796 = n13794 ^ n11830 ;
  assign n13797 = n13796 ^ n12464 ;
  assign n13798 = n13797 ^ n13794 ;
  assign n13799 = n13083 & n13798 ;
  assign n13800 = n13799 ^ n13796 ;
  assign n13801 = ~n13795 & ~n13800 ;
  assign n13802 = n13801 ^ n13794 ;
  assign n13803 = n13802 ^ n13776 ;
  assign n13804 = n13781 & n13803 ;
  assign n13805 = n13804 ^ n13776 ;
  assign n13806 = n13805 ^ n13770 ;
  assign n13807 = n13775 & ~n13806 ;
  assign n13809 = n13808 ^ n13807 ;
  assign n13726 = n13262 ^ n1154 ;
  assign n13864 = n13809 ^ n13726 ;
  assign n13865 = n13864 ^ n10729 ;
  assign n13867 = n13802 ^ n13781 ;
  assign n13868 = n13867 ^ n11241 ;
  assign n13873 = n13791 ^ n13784 ;
  assign n13617 = n13616 ^ n13615 ;
  assign n13618 = n13617 ^ n11170 ;
  assign n13600 = n13599 ^ n13593 ;
  assign n13601 = n13600 ^ n11096 ;
  assign n13543 = n13451 ^ n12897 ;
  assign n13461 = n13447 ^ n13445 ;
  assign n13462 = n13461 ^ n10997 ;
  assign n13535 = n13440 ^ n13436 ;
  assign n13463 = n13428 ^ n12905 ;
  assign n13464 = n13463 ^ n10975 ;
  assign n13465 = n13425 ^ n12912 ;
  assign n13466 = n13465 ^ n11014 ;
  assign n13524 = n13423 ^ n12917 ;
  assign n13467 = n13418 ^ n12927 ;
  assign n13468 = n13467 ^ n11022 ;
  assign n13469 = n13416 ^ n12933 ;
  assign n13470 = n13469 ^ n11048 ;
  assign n13471 = n13411 ^ n13410 ;
  assign n13472 = n13471 ^ n11028 ;
  assign n13473 = n13408 ^ n12945 ;
  assign n13474 = n13473 ^ n11033 ;
  assign n13475 = n13403 ^ n13402 ;
  assign n13476 = n13475 ^ n10961 ;
  assign n13477 = n13399 ^ n13391 ;
  assign n13478 = n13477 ^ n10852 ;
  assign n13502 = n13501 ^ n13479 ;
  assign n13503 = n13501 ^ n10167 ;
  assign n13504 = n13502 & n13503 ;
  assign n13505 = n13504 ^ n10167 ;
  assign n13506 = n13505 ^ n13477 ;
  assign n13507 = ~n13478 & n13506 ;
  assign n13508 = n13507 ^ n10852 ;
  assign n13509 = n13508 ^ n13475 ;
  assign n13510 = ~n13476 & ~n13509 ;
  assign n13511 = n13510 ^ n10961 ;
  assign n13512 = n13511 ^ n13473 ;
  assign n13513 = n13474 & ~n13512 ;
  assign n13514 = n13513 ^ n11033 ;
  assign n13515 = n13514 ^ n13471 ;
  assign n13516 = ~n13472 & ~n13515 ;
  assign n13517 = n13516 ^ n11028 ;
  assign n13518 = n13517 ^ n13469 ;
  assign n13519 = n13470 & n13518 ;
  assign n13520 = n13519 ^ n11048 ;
  assign n13521 = n13520 ^ n13467 ;
  assign n13522 = ~n13468 & ~n13521 ;
  assign n13523 = n13522 ^ n11022 ;
  assign n13525 = n13524 ^ n13523 ;
  assign n13526 = n13524 ^ n11019 ;
  assign n13527 = ~n13525 & n13526 ;
  assign n13528 = n13527 ^ n11019 ;
  assign n13529 = n13528 ^ n13465 ;
  assign n13530 = n13466 & n13529 ;
  assign n13531 = n13530 ^ n11014 ;
  assign n13532 = n13531 ^ n13463 ;
  assign n13533 = n13464 & ~n13532 ;
  assign n13534 = n13533 ^ n10975 ;
  assign n13536 = n13535 ^ n13534 ;
  assign n13537 = n13535 ^ n11007 ;
  assign n13538 = ~n13536 & ~n13537 ;
  assign n13539 = n13538 ^ n11007 ;
  assign n13540 = n13539 ^ n13461 ;
  assign n13541 = n13462 & n13540 ;
  assign n13542 = n13541 ^ n10997 ;
  assign n13544 = n13543 ^ n13542 ;
  assign n13545 = n13543 ^ n10990 ;
  assign n13546 = ~n13544 & n13545 ;
  assign n13547 = n13546 ^ n10990 ;
  assign n13459 = n13458 ^ n13453 ;
  assign n13587 = n13547 ^ n13459 ;
  assign n13588 = n13547 ^ n10996 ;
  assign n13589 = ~n13587 & ~n13588 ;
  assign n13590 = n13589 ^ n10996 ;
  assign n13606 = n13600 ^ n13590 ;
  assign n13607 = n13601 & n13606 ;
  assign n13608 = n13607 ^ n11096 ;
  assign n13870 = n13617 ^ n13608 ;
  assign n13871 = n13618 & n13870 ;
  assign n13872 = n13871 ^ n11170 ;
  assign n13874 = n13873 ^ n13872 ;
  assign n13875 = n13873 ^ n11186 ;
  assign n13876 = n13874 & n13875 ;
  assign n13877 = n13876 ^ n11186 ;
  assign n13869 = n13800 ^ n13793 ;
  assign n13878 = n13877 ^ n13869 ;
  assign n13879 = n13877 ^ n11226 ;
  assign n13880 = ~n13878 & ~n13879 ;
  assign n13881 = n13880 ^ n11226 ;
  assign n13882 = n13881 ^ n13867 ;
  assign n13883 = ~n13868 & n13882 ;
  assign n13884 = n13883 ^ n11241 ;
  assign n13866 = n13805 ^ n13775 ;
  assign n13885 = n13884 ^ n13866 ;
  assign n13886 = n13884 ^ n11381 ;
  assign n13887 = n13885 & ~n13886 ;
  assign n13888 = n13887 ^ n11381 ;
  assign n13889 = n13888 ^ n13864 ;
  assign n13890 = ~n13865 & n13889 ;
  assign n13891 = n13890 ^ n10729 ;
  assign n13821 = n13220 ^ n1359 ;
  assign n13822 = n13821 ^ n13264 ;
  assign n13768 = n13767 ^ n13726 ;
  assign n13810 = n13768 & ~n13809 ;
  assign n13811 = n13810 ^ n13767 ;
  assign n13812 = n13811 ^ n11339 ;
  assign n13813 = n13812 ^ n12050 ;
  assign n13814 = n13813 ^ n13811 ;
  assign n13815 = n13374 & n13814 ;
  assign n13816 = n13815 ^ n13812 ;
  assign n13863 = n13822 ^ n13816 ;
  assign n13892 = n13891 ^ n13863 ;
  assign n13893 = n13891 ^ n10734 ;
  assign n13894 = ~n13892 & ~n13893 ;
  assign n13895 = n13894 ^ n10734 ;
  assign n13830 = n13270 ^ n1395 ;
  assign n13817 = n12038 ^ n11358 ;
  assign n13818 = ~n12631 & ~n13817 ;
  assign n13819 = n13818 ^ n11358 ;
  assign n13823 = n13822 ^ n13819 ;
  assign n13820 = n13819 ^ n13811 ;
  assign n13824 = n13823 ^ n13820 ;
  assign n13825 = ~n13816 & n13824 ;
  assign n13826 = n13825 ^ n13823 ;
  assign n13861 = n13830 ^ n13826 ;
  assign n13862 = n13861 ^ n10748 ;
  assign n13927 = n13895 ^ n13862 ;
  assign n13910 = n13869 ^ n11226 ;
  assign n13911 = n13910 ^ n13877 ;
  assign n13912 = n13875 ^ n13872 ;
  assign n13460 = n13459 ^ n10996 ;
  assign n13548 = n13547 ^ n13460 ;
  assign n13549 = n13545 ^ n13542 ;
  assign n13550 = n13539 ^ n13462 ;
  assign n13551 = n13537 ^ n13534 ;
  assign n13552 = n13528 ^ n13466 ;
  assign n13553 = n13526 ^ n13523 ;
  assign n13566 = ~n13555 & ~n13565 ;
  assign n13567 = n13505 ^ n13478 ;
  assign n13568 = n13566 & ~n13567 ;
  assign n13569 = n13508 ^ n13476 ;
  assign n13570 = ~n13568 & n13569 ;
  assign n13571 = n13511 ^ n13474 ;
  assign n13572 = n13570 & n13571 ;
  assign n13573 = n13514 ^ n13472 ;
  assign n13574 = ~n13572 & n13573 ;
  assign n13575 = n13517 ^ n13470 ;
  assign n13576 = n13574 & n13575 ;
  assign n13577 = n13520 ^ n13468 ;
  assign n13578 = ~n13576 & ~n13577 ;
  assign n13579 = ~n13553 & n13578 ;
  assign n13580 = ~n13552 & n13579 ;
  assign n13581 = n13531 ^ n13464 ;
  assign n13582 = n13580 & n13581 ;
  assign n13583 = n13551 & ~n13582 ;
  assign n13584 = n13550 & n13583 ;
  assign n13585 = n13549 & ~n13584 ;
  assign n13586 = n13548 & ~n13585 ;
  assign n13602 = n13601 ^ n13590 ;
  assign n13605 = n13586 & n13602 ;
  assign n13619 = n13618 ^ n13608 ;
  assign n13913 = n13605 & ~n13619 ;
  assign n13914 = n13912 & n13913 ;
  assign n13915 = n13911 & n13914 ;
  assign n13916 = n13881 ^ n11241 ;
  assign n13917 = n13916 ^ n13867 ;
  assign n13918 = ~n13915 & n13917 ;
  assign n13919 = n13866 ^ n11381 ;
  assign n13920 = n13919 ^ n13884 ;
  assign n13921 = ~n13918 & n13920 ;
  assign n13922 = n13888 ^ n13865 ;
  assign n13923 = ~n13921 & ~n13922 ;
  assign n13924 = n13863 ^ n10734 ;
  assign n13925 = n13924 ^ n13891 ;
  assign n13926 = ~n13923 & n13925 ;
  assign n13974 = n13927 ^ n13926 ;
  assign n14024 = n13974 ^ n2528 ;
  assign n13939 = n13925 ^ n13923 ;
  assign n13940 = n13939 ^ n2586 ;
  assign n13942 = n13920 ^ n13918 ;
  assign n13943 = n13942 ^ n3109 ;
  assign n13958 = n13917 ^ n13915 ;
  assign n13944 = n13914 ^ n13911 ;
  assign n13945 = n13944 ^ n2501 ;
  assign n13603 = n13602 ^ n13586 ;
  assign n13604 = n13603 ^ n1053 ;
  assign n13623 = n13585 ^ n13548 ;
  assign n13624 = n13623 ^ n907 ;
  assign n13625 = n13584 ^ n13549 ;
  assign n13626 = n13625 ^ n901 ;
  assign n13629 = n13583 ^ n13550 ;
  assign n13715 = n13629 ^ n13625 ;
  assign n13627 = n13582 ^ n13551 ;
  assign n13628 = n13627 ^ n805 ;
  assign n13632 = n13581 ^ n13580 ;
  assign n13633 = n13632 ^ n799 ;
  assign n13701 = n13579 ^ n13552 ;
  assign n13634 = n13578 ^ n13553 ;
  assign n13635 = n13634 ^ n1565 ;
  assign n13636 = n13577 ^ n13576 ;
  assign n13637 = n13636 ^ n525 ;
  assign n13640 = n13575 ^ n13574 ;
  assign n13641 = n13640 ^ n545 ;
  assign n13642 = n13573 ^ n13572 ;
  assign n13643 = n13642 ^ n560 ;
  assign n13646 = n13571 ^ n13570 ;
  assign n13650 = n13649 ^ n13646 ;
  assign n13651 = n13569 ^ n13568 ;
  assign n13652 = n13651 ^ n1451 ;
  assign n13655 = n13567 ^ n13566 ;
  assign n13656 = n13655 ^ n2274 ;
  assign n13679 = n13678 ^ n13657 ;
  assign n13680 = n13678 ^ n2258 ;
  assign n13681 = ~n13679 & n13680 ;
  assign n13682 = n13681 ^ n2258 ;
  assign n13683 = n13682 ^ n13655 ;
  assign n13684 = ~n13656 & n13683 ;
  assign n13685 = n13684 ^ n2274 ;
  assign n13653 = n13646 ^ n1451 ;
  assign n13654 = n13653 ^ n13646 ;
  assign n13686 = n13685 ^ n13654 ;
  assign n13687 = n13652 & n13686 ;
  assign n13688 = n13687 ^ n13653 ;
  assign n13689 = ~n13650 & n13688 ;
  assign n13690 = n13689 ^ n13649 ;
  assign n13644 = n13640 ^ n560 ;
  assign n13645 = n13644 ^ n13640 ;
  assign n13691 = n13690 ^ n13645 ;
  assign n13692 = ~n13643 & n13691 ;
  assign n13693 = n13692 ^ n13644 ;
  assign n13694 = n13641 & ~n13693 ;
  assign n13695 = n13694 ^ n545 ;
  assign n13638 = n13634 ^ n525 ;
  assign n13639 = n13638 ^ n13634 ;
  assign n13696 = n13695 ^ n13639 ;
  assign n13697 = ~n13637 & n13696 ;
  assign n13698 = n13697 ^ n13638 ;
  assign n13699 = n13635 & n13698 ;
  assign n13700 = n13699 ^ n13634 ;
  assign n13702 = n13701 ^ n13700 ;
  assign n13703 = n13632 ^ n536 ;
  assign n13704 = n13703 ^ n13632 ;
  assign n13705 = n13704 ^ n13700 ;
  assign n13706 = ~n13702 & n13705 ;
  assign n13707 = n13706 ^ n13703 ;
  assign n13708 = ~n13633 & ~n13707 ;
  assign n13709 = n13708 ^ n13632 ;
  assign n13630 = n13629 ^ n805 ;
  assign n13631 = n13630 ^ n13629 ;
  assign n13710 = n13709 ^ n13631 ;
  assign n13711 = ~n13628 & ~n13710 ;
  assign n13712 = n13711 ^ n13630 ;
  assign n13713 = n13629 ^ n817 ;
  assign n13714 = n13712 & n13713 ;
  assign n13716 = n13715 ^ n13714 ;
  assign n13717 = n13626 & n13716 ;
  assign n13718 = n13717 ^ n13625 ;
  assign n13719 = n13718 ^ n13623 ;
  assign n13720 = ~n13624 & n13719 ;
  assign n13721 = n13720 ^ n907 ;
  assign n13620 = n13619 ^ n13605 ;
  assign n13621 = n13620 ^ n1053 ;
  assign n13622 = n13621 ^ n13620 ;
  assign n13722 = n13721 ^ n13622 ;
  assign n13723 = n13604 & n13722 ;
  assign n13724 = n13723 ^ n13621 ;
  assign n13947 = n13620 ^ n1244 ;
  assign n13948 = n13724 & ~n13947 ;
  assign n13949 = n13948 ^ n1244 ;
  assign n13946 = n13913 ^ n13912 ;
  assign n13950 = n13949 ^ n13946 ;
  assign n13951 = n13944 ^ n1238 ;
  assign n13952 = n13951 ^ n13944 ;
  assign n13953 = n13952 ^ n13946 ;
  assign n13954 = ~n13950 & n13953 ;
  assign n13955 = n13954 ^ n13951 ;
  assign n13956 = n13945 & ~n13955 ;
  assign n13957 = n13956 ^ n2501 ;
  assign n13959 = n13958 ^ n13957 ;
  assign n13960 = n13958 ^ n2848 ;
  assign n13961 = ~n13959 & n13960 ;
  assign n13962 = n13961 ^ n2848 ;
  assign n13963 = n13962 ^ n13942 ;
  assign n13964 = ~n13943 & n13963 ;
  assign n13965 = n13964 ^ n3109 ;
  assign n13941 = n13922 ^ n13921 ;
  assign n13966 = n13965 ^ n13941 ;
  assign n13967 = n13939 ^ n1829 ;
  assign n13968 = n13967 ^ n13939 ;
  assign n13969 = n13968 ^ n13941 ;
  assign n13970 = n13966 & ~n13969 ;
  assign n13971 = n13970 ^ n13967 ;
  assign n13972 = ~n13940 & n13971 ;
  assign n13973 = n13972 ^ n2586 ;
  assign n14025 = n14024 ^ n13973 ;
  assign n14021 = n12709 ^ n12070 ;
  assign n14022 = n12950 & n14021 ;
  assign n14023 = n14022 ^ n12070 ;
  assign n14116 = n14025 ^ n14023 ;
  assign n14207 = n14116 ^ n11407 ;
  assign n1947 = x480 ^ x128 ;
  assign n1948 = n1947 ^ x64 ;
  assign n1949 = n1948 ^ x320 ;
  assign n14377 = n14207 ^ n1949 ;
  assign n14378 = n14377 ^ n12886 ;
  assign n14379 = n14378 ^ n12917 ;
  assign n14380 = n14379 ^ n14377 ;
  assign n14381 = n13744 & ~n14380 ;
  assign n14382 = n14381 ^ n14378 ;
  assign n14067 = n13675 ^ n13659 ;
  assign n14652 = n12922 ^ n12788 ;
  assign n14653 = n14067 & ~n14652 ;
  assign n14654 = n14653 ^ n12922 ;
  assign n14475 = n12697 ^ n12024 ;
  assign n14476 = ~n13312 & n14475 ;
  assign n14477 = n14476 ^ n12024 ;
  assign n14468 = n13962 ^ n13943 ;
  assign n14465 = n13960 ^ n13957 ;
  assign n14469 = n14468 ^ n14465 ;
  assign n14384 = n12621 ^ n12038 ;
  assign n14385 = n13316 & n14384 ;
  assign n14386 = n14385 ^ n12038 ;
  assign n14383 = n13955 ^ n2501 ;
  assign n14387 = n14386 ^ n14383 ;
  assign n14388 = n13946 ^ n1238 ;
  assign n14389 = n14388 ^ n13949 ;
  assign n14456 = n14389 ^ n14386 ;
  assign n13988 = n13284 ^ n2444 ;
  assign n14390 = n14389 ^ n12050 ;
  assign n14391 = n14390 ^ n12627 ;
  assign n14392 = n14391 ^ n14389 ;
  assign n14393 = n13988 & ~n14392 ;
  assign n14394 = n14393 ^ n14390 ;
  assign n13846 = n13213 ^ n2484 ;
  assign n13847 = n13846 ^ n13278 ;
  assign n14395 = n12631 ^ n12040 ;
  assign n14396 = ~n13847 & n14395 ;
  assign n14397 = n14396 ^ n12040 ;
  assign n13725 = n13724 ^ n1244 ;
  assign n14398 = n14397 ^ n13725 ;
  assign n13837 = n13272 ^ n13217 ;
  assign n14402 = n13718 ^ n13624 ;
  assign n14403 = n14402 ^ n12646 ;
  assign n14404 = n14403 ^ n13343 ;
  assign n14405 = n14404 ^ n14402 ;
  assign n14406 = ~n13837 & n14405 ;
  assign n14407 = n14406 ^ n14403 ;
  assign n14409 = n13295 ^ n12464 ;
  assign n14410 = ~n13830 & ~n14409 ;
  assign n14411 = n14410 ^ n12464 ;
  assign n14408 = n13716 ^ n901 ;
  assign n14412 = n14411 ^ n14408 ;
  assign n14416 = n13712 ^ n817 ;
  assign n14413 = n13171 ^ n12370 ;
  assign n14414 = ~n13822 & n14413 ;
  assign n14415 = n14414 ^ n12370 ;
  assign n14417 = n14416 ^ n14415 ;
  assign n14419 = n13083 ^ n12379 ;
  assign n14420 = ~n13726 & ~n14419 ;
  assign n14421 = n14420 ^ n12379 ;
  assign n14418 = n13709 ^ n13628 ;
  assign n14422 = n14421 ^ n14418 ;
  assign n14426 = n13707 ^ n799 ;
  assign n14423 = n13076 ^ n12385 ;
  assign n14424 = n13770 & ~n14423 ;
  assign n14425 = n14424 ^ n12385 ;
  assign n14427 = n14426 ^ n14425 ;
  assign n14332 = n13701 ^ n536 ;
  assign n14333 = n14332 ^ n13700 ;
  assign n14334 = n14333 ^ n12390 ;
  assign n14335 = n14334 ^ n12960 ;
  assign n14336 = n14335 ^ n14333 ;
  assign n14337 = ~n13776 & ~n14336 ;
  assign n14338 = n14337 ^ n14334 ;
  assign n14190 = n13698 ^ n1565 ;
  assign n14191 = n14190 ^ n12344 ;
  assign n14192 = n14191 ^ n12971 ;
  assign n14193 = n14192 ^ n14190 ;
  assign n14194 = ~n13794 & ~n14193 ;
  assign n14195 = n14194 ^ n14191 ;
  assign n14176 = n13695 ^ n13637 ;
  assign n14177 = n14176 ^ n12399 ;
  assign n14178 = n14177 ^ n12976 ;
  assign n14179 = n14178 ^ n14176 ;
  assign n14180 = n13785 & ~n14179 ;
  assign n14181 = n14180 ^ n14177 ;
  assign n14092 = n12402 ^ n12343 ;
  assign n14093 = ~n13616 & ~n14092 ;
  assign n14094 = n14093 ^ n12402 ;
  assign n14084 = n13690 ^ n13643 ;
  assign n14095 = n14094 ^ n14084 ;
  assign n13729 = n12982 ^ n12413 ;
  assign n13730 = n13454 & n13729 ;
  assign n13731 = n13730 ^ n12413 ;
  assign n13728 = n13688 ^ n13649 ;
  assign n13732 = n13731 ^ n13728 ;
  assign n13736 = n13685 ^ n13652 ;
  assign n13733 = n12899 ^ n12422 ;
  assign n13734 = n12897 & ~n13733 ;
  assign n13735 = n13734 ^ n12422 ;
  assign n13737 = n13736 ^ n13735 ;
  assign n13739 = n12906 ^ n12433 ;
  assign n13740 = ~n13447 & ~n13739 ;
  assign n13741 = n13740 ^ n12433 ;
  assign n13738 = n13682 ^ n13656 ;
  assign n13742 = n13741 ^ n13738 ;
  assign n13745 = n12913 ^ n12337 ;
  assign n13746 = n13440 & n13745 ;
  assign n13747 = n13746 ^ n12337 ;
  assign n13748 = n13747 ^ n13744 ;
  assign n13749 = n13669 ^ n13663 ;
  assign n13750 = n13749 ^ n11531 ;
  assign n13751 = n13750 ^ n12940 ;
  assign n13752 = n13751 ^ n13749 ;
  assign n13753 = ~n12917 & n13752 ;
  assign n13754 = n13753 ^ n13750 ;
  assign n14050 = n12928 ^ n12118 ;
  assign n14051 = n12907 & ~n14050 ;
  assign n14052 = n14051 ^ n12118 ;
  assign n14054 = n14052 ^ n13749 ;
  assign n13756 = n12936 ^ n12103 ;
  assign n13757 = n12922 & ~n13756 ;
  assign n13758 = n13757 ^ n12103 ;
  assign n13755 = n13666 ^ n13665 ;
  assign n13759 = n13758 ^ n13755 ;
  assign n13761 = n12886 ^ n12093 ;
  assign n13762 = ~n12933 & n13761 ;
  assign n13763 = n13762 ^ n12093 ;
  assign n14046 = n13763 ^ n13755 ;
  assign n13760 = n13559 ^ n1903 ;
  assign n13764 = n13763 ^ n13760 ;
  assign n14005 = n12788 ^ n11537 ;
  assign n14006 = ~n13411 & n14005 ;
  assign n14007 = n14006 ^ n11537 ;
  assign n14043 = n14007 ^ n13763 ;
  assign n13843 = n12024 ^ n11394 ;
  assign n13844 = n12621 & n13843 ;
  assign n13845 = n13844 ^ n11394 ;
  assign n13827 = n12029 ^ n11338 ;
  assign n13828 = n12627 & n13827 ;
  assign n13829 = n13828 ^ n11338 ;
  assign n13832 = n13829 ^ n13819 ;
  assign n13831 = n13830 ^ n13829 ;
  assign n13833 = n13832 ^ n13831 ;
  assign n13834 = n13826 & n13833 ;
  assign n13835 = n13834 ^ n13832 ;
  assign n13836 = n13275 ^ n13215 ;
  assign n13839 = n13836 ^ n13829 ;
  assign n13838 = n13837 ^ n13836 ;
  assign n13840 = n13839 ^ n13838 ;
  assign n13841 = ~n13835 & ~n13840 ;
  assign n13842 = n13841 ^ n13839 ;
  assign n13858 = n13845 ^ n13842 ;
  assign n13859 = n13858 ^ n10724 ;
  assign n13896 = n13895 ^ n13861 ;
  assign n13897 = n13862 & n13896 ;
  assign n13898 = n13897 ^ n10748 ;
  assign n13860 = n13837 ^ n13835 ;
  assign n13899 = n13898 ^ n13860 ;
  assign n13900 = n13898 ^ n10756 ;
  assign n13901 = n13899 & ~n13900 ;
  assign n13902 = n13901 ^ n10756 ;
  assign n13903 = n13902 ^ n13858 ;
  assign n13904 = n13859 & n13903 ;
  assign n13905 = n13904 ^ n10724 ;
  assign n13932 = n13905 ^ n10211 ;
  assign n13853 = n11569 ^ n10984 ;
  assign n13854 = ~n12669 & ~n13853 ;
  assign n13855 = n13854 ^ n11569 ;
  assign n13849 = n13847 ^ n13836 ;
  assign n13848 = n13847 ^ n13845 ;
  assign n13850 = n13849 ^ n13848 ;
  assign n13851 = ~n13842 & ~n13850 ;
  assign n13852 = n13851 ^ n13849 ;
  assign n13856 = n13855 ^ n13852 ;
  assign n13933 = n13932 ^ n13856 ;
  assign n13908 = n13860 ^ n10756 ;
  assign n13909 = n13908 ^ n13898 ;
  assign n13928 = ~n13926 & ~n13927 ;
  assign n13929 = n13909 & n13928 ;
  assign n13930 = n13902 ^ n13859 ;
  assign n13931 = ~n13929 & n13930 ;
  assign n13999 = n13933 ^ n13931 ;
  assign n14000 = n13999 ^ n1856 ;
  assign n13935 = n13930 ^ n13929 ;
  assign n13936 = n13935 ^ n2742 ;
  assign n13937 = n13928 ^ n13909 ;
  assign n13938 = n13937 ^ n2454 ;
  assign n13975 = n13974 ^ n13973 ;
  assign n13976 = n13937 ^ n2528 ;
  assign n13977 = n13976 ^ n13937 ;
  assign n13978 = n13977 ^ n13973 ;
  assign n13979 = n13975 & n13978 ;
  assign n13980 = n13979 ^ n13976 ;
  assign n13981 = ~n13938 & n13980 ;
  assign n13982 = n13981 ^ n2454 ;
  assign n13983 = n13982 ^ n13935 ;
  assign n13984 = ~n13936 & n13983 ;
  assign n13985 = n13984 ^ n2742 ;
  assign n14001 = n13985 ^ n1856 ;
  assign n14002 = n14000 & n14001 ;
  assign n13995 = n13855 ^ n13847 ;
  assign n13996 = ~n13852 & n13995 ;
  assign n13992 = n11558 ^ n10982 ;
  assign n13993 = n12697 & n13992 ;
  assign n13987 = n13855 ^ n13372 ;
  assign n13989 = n13988 ^ n13987 ;
  assign n13990 = n13989 ^ n10211 ;
  assign n13986 = n13985 ^ n1862 ;
  assign n13991 = n13990 ^ n13986 ;
  assign n13994 = n13993 ^ n13991 ;
  assign n13997 = n13996 ^ n13994 ;
  assign n13934 = ~n13931 & ~n13933 ;
  assign n13998 = n13997 ^ n13934 ;
  assign n14003 = n14002 ^ n13998 ;
  assign n13857 = n13856 ^ n10211 ;
  assign n13906 = n13905 ^ n13856 ;
  assign n13907 = ~n13857 & ~n13906 ;
  assign n14004 = n14003 ^ n13907 ;
  assign n14008 = n14007 ^ n14004 ;
  assign n14009 = n14000 ^ n13985 ;
  assign n14040 = n14009 ^ n14007 ;
  assign n14010 = n14009 ^ n11544 ;
  assign n14011 = n14010 ^ n12725 ;
  assign n14012 = n14011 ^ n14009 ;
  assign n14013 = n12945 & n14012 ;
  assign n14014 = n14013 ^ n14010 ;
  assign n14018 = n13982 ^ n13936 ;
  assign n14015 = n12348 ^ n12077 ;
  assign n14016 = n13403 & ~n14015 ;
  assign n14017 = n14016 ^ n12077 ;
  assign n14019 = n14018 ^ n14017 ;
  assign n14026 = n14023 & ~n14025 ;
  assign n14020 = n13980 ^ n2454 ;
  assign n14027 = n14026 ^ n14020 ;
  assign n14028 = n14026 ^ n11551 ;
  assign n14029 = n14028 ^ n12356 ;
  assign n14030 = n14029 ^ n14026 ;
  assign n14031 = ~n13389 & ~n14030 ;
  assign n14032 = n14031 ^ n14028 ;
  assign n14033 = ~n14027 & ~n14032 ;
  assign n14034 = n14033 ^ n14026 ;
  assign n14035 = n14034 ^ n14017 ;
  assign n14036 = ~n14019 & ~n14035 ;
  assign n14037 = n14036 ^ n14018 ;
  assign n14038 = n14037 ^ n14009 ;
  assign n14039 = n14014 & n14038 ;
  assign n14041 = n14040 ^ n14039 ;
  assign n14042 = ~n14008 & n14041 ;
  assign n14044 = n14043 ^ n14042 ;
  assign n14045 = ~n13764 & ~n14044 ;
  assign n14047 = n14046 ^ n14045 ;
  assign n14048 = ~n13759 & n14047 ;
  assign n14049 = n14048 ^ n13758 ;
  assign n14053 = n14052 ^ n14049 ;
  assign n14055 = n14054 ^ n14053 ;
  assign n14056 = ~n13754 & n14055 ;
  assign n14057 = n14056 ^ n14054 ;
  assign n14058 = n12920 ^ n12197 ;
  assign n14059 = n12900 & ~n14058 ;
  assign n14060 = n14059 ^ n12197 ;
  assign n14063 = n14060 ^ n14052 ;
  assign n14061 = n13673 ^ n2244 ;
  assign n14062 = n14061 ^ n14060 ;
  assign n14064 = n14063 ^ n14062 ;
  assign n14065 = n14057 & n14064 ;
  assign n14066 = n14065 ^ n14063 ;
  assign n14069 = n14060 ^ n13747 ;
  assign n14068 = n14067 ^ n13747 ;
  assign n14070 = n14069 ^ n14068 ;
  assign n14071 = n14066 & ~n14070 ;
  assign n14072 = n14071 ^ n14069 ;
  assign n14073 = n13748 & n14072 ;
  assign n14074 = n14073 ^ n13747 ;
  assign n14075 = n14074 ^ n13741 ;
  assign n14076 = n13742 & n14075 ;
  assign n14077 = n14076 ^ n14074 ;
  assign n14078 = n14077 ^ n13735 ;
  assign n14079 = ~n13737 & n14078 ;
  assign n14080 = n14079 ^ n13736 ;
  assign n14081 = n14080 ^ n13728 ;
  assign n14082 = ~n13732 & n14081 ;
  assign n14083 = n14082 ^ n13731 ;
  assign n14085 = n14084 ^ n14083 ;
  assign n14086 = n14084 ^ n12407 ;
  assign n14087 = n14086 ^ n13046 ;
  assign n14088 = n14087 ^ n14084 ;
  assign n14089 = n13594 & n14088 ;
  assign n14090 = n14089 ^ n14086 ;
  assign n14091 = ~n14085 & n14090 ;
  assign n14096 = n14095 ^ n14091 ;
  assign n14097 = n13693 ^ n545 ;
  assign n14182 = n14097 ^ n14094 ;
  assign n14183 = n14096 & ~n14182 ;
  assign n14184 = n14183 ^ n14094 ;
  assign n14196 = n14184 ^ n14176 ;
  assign n14197 = ~n14181 & n14196 ;
  assign n14198 = n14197 ^ n14176 ;
  assign n14339 = n14198 ^ n14190 ;
  assign n14340 = ~n14195 & ~n14339 ;
  assign n14341 = n14340 ^ n14198 ;
  assign n14428 = n14341 ^ n14333 ;
  assign n14429 = n14338 & ~n14428 ;
  assign n14430 = n14429 ^ n14333 ;
  assign n14431 = n14430 ^ n14425 ;
  assign n14432 = n14427 & n14431 ;
  assign n14433 = n14432 ^ n14426 ;
  assign n14434 = n14433 ^ n14418 ;
  assign n14435 = ~n14422 & n14434 ;
  assign n14436 = n14435 ^ n14421 ;
  assign n14437 = n14436 ^ n14415 ;
  assign n14438 = n14417 & n14437 ;
  assign n14439 = n14438 ^ n14416 ;
  assign n14440 = n14439 ^ n14408 ;
  assign n14441 = n14412 & ~n14440 ;
  assign n14442 = n14441 ^ n14411 ;
  assign n14443 = n14442 ^ n14402 ;
  assign n14444 = ~n14407 & ~n14443 ;
  assign n14445 = n14444 ^ n14402 ;
  assign n14399 = n13374 ^ n12686 ;
  assign n14400 = ~n13836 & n14399 ;
  assign n14401 = n14400 ^ n12686 ;
  assign n14446 = n14445 ^ n14401 ;
  assign n14447 = n13721 ^ n13604 ;
  assign n14448 = n14447 ^ n14401 ;
  assign n14449 = ~n14446 & ~n14448 ;
  assign n14450 = n14449 ^ n14445 ;
  assign n14451 = n14450 ^ n14397 ;
  assign n14452 = n14398 & ~n14451 ;
  assign n14453 = n14452 ^ n13725 ;
  assign n14454 = n14453 ^ n14389 ;
  assign n14455 = ~n14394 & ~n14454 ;
  assign n14457 = n14456 ^ n14455 ;
  assign n14458 = n14387 & n14457 ;
  assign n14459 = n14458 ^ n14386 ;
  assign n14460 = n14459 ^ n12029 ;
  assign n14461 = n14460 ^ n12669 ;
  assign n14462 = n14461 ^ n14459 ;
  assign n14463 = ~n13315 & n14462 ;
  assign n14464 = n14463 ^ n14460 ;
  assign n14466 = n14465 ^ n14459 ;
  assign n14467 = ~n14464 & n14466 ;
  assign n14470 = n14469 ^ n14467 ;
  assign n14486 = n14477 ^ n14470 ;
  assign n14487 = n14486 ^ n11394 ;
  assign n14488 = n14465 ^ n14464 ;
  assign n14489 = n14488 ^ n11338 ;
  assign n14490 = n14457 ^ n14383 ;
  assign n14491 = n14490 ^ n11358 ;
  assign n14530 = n14453 ^ n14394 ;
  assign n14492 = n14450 ^ n14398 ;
  assign n14493 = n14492 ^ n11340 ;
  assign n14522 = n14448 ^ n14445 ;
  assign n14494 = n14442 ^ n14407 ;
  assign n14495 = n14494 ^ n11842 ;
  assign n14514 = n14439 ^ n14412 ;
  assign n14496 = n14436 ^ n14417 ;
  assign n14497 = n14496 ^ n11822 ;
  assign n14498 = n14433 ^ n14422 ;
  assign n14499 = n14498 ^ n11719 ;
  assign n14500 = n14430 ^ n14427 ;
  assign n14501 = n14500 ^ n11713 ;
  assign n14342 = n14341 ^ n14338 ;
  assign n14343 = n14342 ^ n11703 ;
  assign n14199 = n14198 ^ n14195 ;
  assign n14200 = n14199 ^ n11571 ;
  assign n14185 = n14184 ^ n14181 ;
  assign n14098 = n14097 ^ n14096 ;
  assign n14099 = n14098 ^ n11593 ;
  assign n14168 = n14090 ^ n14083 ;
  assign n14100 = n14080 ^ n13732 ;
  assign n14101 = n14100 ^ n11598 ;
  assign n14102 = n14077 ^ n13737 ;
  assign n14103 = n14102 ^ n10974 ;
  assign n14104 = n14074 ^ n13742 ;
  assign n14105 = n14104 ^ n11607 ;
  assign n14107 = n14067 ^ n14066 ;
  assign n14108 = n14107 ^ n11533 ;
  assign n14143 = n14049 ^ n13754 ;
  assign n14110 = n14047 ^ n13758 ;
  assign n14111 = n14110 ^ n11546 ;
  assign n14112 = n14044 ^ n13760 ;
  assign n14113 = n14112 ^ n11553 ;
  assign n14131 = n14041 ^ n14004 ;
  assign n14114 = n14037 ^ n14014 ;
  assign n14115 = n14114 ^ n11565 ;
  assign n14123 = n14034 ^ n14019 ;
  assign n14117 = n11407 & ~n14116 ;
  assign n14118 = n14117 ^ n11453 ;
  assign n14119 = n14032 ^ n14020 ;
  assign n14120 = n14119 ^ n14117 ;
  assign n14121 = ~n14118 & ~n14120 ;
  assign n14122 = n14121 ^ n11453 ;
  assign n14124 = n14123 ^ n14122 ;
  assign n14125 = n14123 ^ n11520 ;
  assign n14126 = ~n14124 & n14125 ;
  assign n14127 = n14126 ^ n11520 ;
  assign n14128 = n14127 ^ n14114 ;
  assign n14129 = n14115 & ~n14128 ;
  assign n14130 = n14129 ^ n11565 ;
  assign n14132 = n14131 ^ n14130 ;
  assign n14133 = n14112 ^ n11557 ;
  assign n14134 = n14133 ^ n14112 ;
  assign n14135 = n14134 ^ n14130 ;
  assign n14136 = n14132 & ~n14135 ;
  assign n14137 = n14136 ^ n14133 ;
  assign n14138 = ~n14113 & ~n14137 ;
  assign n14139 = n14138 ^ n11553 ;
  assign n14140 = n14139 ^ n14110 ;
  assign n14141 = ~n14111 & ~n14140 ;
  assign n14142 = n14141 ^ n11546 ;
  assign n14144 = n14143 ^ n14142 ;
  assign n14145 = n14143 ^ n11655 ;
  assign n14146 = n14144 & n14145 ;
  assign n14147 = n14146 ^ n11655 ;
  assign n14109 = n14061 ^ n14057 ;
  assign n14148 = n14147 ^ n14109 ;
  assign n14149 = n14147 ^ n11539 ;
  assign n14150 = n14148 & ~n14149 ;
  assign n14151 = n14150 ^ n11539 ;
  assign n14152 = n14151 ^ n14107 ;
  assign n14153 = ~n14108 & n14152 ;
  assign n14154 = n14153 ^ n11533 ;
  assign n14106 = n14072 ^ n13744 ;
  assign n14155 = n14154 ^ n14106 ;
  assign n14156 = n14154 ^ n11612 ;
  assign n14157 = ~n14155 & ~n14156 ;
  assign n14158 = n14157 ^ n11612 ;
  assign n14159 = n14158 ^ n14104 ;
  assign n14160 = ~n14105 & ~n14159 ;
  assign n14161 = n14160 ^ n11607 ;
  assign n14162 = n14161 ^ n14102 ;
  assign n14163 = n14103 & n14162 ;
  assign n14164 = n14163 ^ n10974 ;
  assign n14165 = n14164 ^ n14100 ;
  assign n14166 = n14101 & ~n14165 ;
  assign n14167 = n14166 ^ n11598 ;
  assign n14169 = n14168 ^ n14167 ;
  assign n14170 = n14168 ^ n11587 ;
  assign n14171 = n14169 & n14170 ;
  assign n14172 = n14171 ^ n11587 ;
  assign n14173 = n14172 ^ n14098 ;
  assign n14174 = n14099 & ~n14173 ;
  assign n14175 = n14174 ^ n11593 ;
  assign n14186 = n14185 ^ n14175 ;
  assign n14187 = n14185 ^ n11585 ;
  assign n14188 = ~n14186 & ~n14187 ;
  assign n14189 = n14188 ^ n11585 ;
  assign n14344 = n14199 ^ n14189 ;
  assign n14345 = ~n14200 & ~n14344 ;
  assign n14346 = n14345 ^ n11571 ;
  assign n14502 = n14346 ^ n14342 ;
  assign n14503 = n14343 & n14502 ;
  assign n14504 = n14503 ^ n11703 ;
  assign n14505 = n14504 ^ n14500 ;
  assign n14506 = n14501 & n14505 ;
  assign n14507 = n14506 ^ n11713 ;
  assign n14508 = n14507 ^ n14498 ;
  assign n14509 = ~n14499 & ~n14508 ;
  assign n14510 = n14509 ^ n11719 ;
  assign n14511 = n14510 ^ n14496 ;
  assign n14512 = ~n14497 & ~n14511 ;
  assign n14513 = n14512 ^ n11822 ;
  assign n14515 = n14514 ^ n14513 ;
  assign n14516 = n14514 ^ n11830 ;
  assign n14517 = ~n14515 & n14516 ;
  assign n14518 = n14517 ^ n11830 ;
  assign n14519 = n14518 ^ n14494 ;
  assign n14520 = n14495 & n14519 ;
  assign n14521 = n14520 ^ n11842 ;
  assign n14523 = n14522 ^ n14521 ;
  assign n14524 = n14522 ^ n12011 ;
  assign n14525 = ~n14523 & ~n14524 ;
  assign n14526 = n14525 ^ n12011 ;
  assign n14527 = n14526 ^ n14492 ;
  assign n14528 = n14493 & n14527 ;
  assign n14529 = n14528 ^ n11340 ;
  assign n14531 = n14530 ^ n14529 ;
  assign n14532 = n14530 ^ n11339 ;
  assign n14533 = n14531 & ~n14532 ;
  assign n14534 = n14533 ^ n11339 ;
  assign n14535 = n14534 ^ n14490 ;
  assign n14536 = ~n14491 & n14535 ;
  assign n14537 = n14536 ^ n11358 ;
  assign n14538 = n14537 ^ n14488 ;
  assign n14539 = n14489 & n14538 ;
  assign n14540 = n14539 ^ n11338 ;
  assign n14541 = n14540 ^ n11394 ;
  assign n14542 = ~n14487 & n14541 ;
  assign n14543 = n14542 ^ n11394 ;
  assign n14569 = n14543 ^ n10984 ;
  assign n14481 = n12702 ^ n11569 ;
  assign n14482 = ~n13355 & n14481 ;
  assign n14483 = n14482 ^ n11569 ;
  assign n14471 = n13941 ^ n1829 ;
  assign n14472 = n14471 ^ n13965 ;
  assign n14473 = n14472 ^ n14468 ;
  assign n14474 = n14473 ^ n14472 ;
  assign n14478 = n14477 ^ n14474 ;
  assign n14479 = ~n14470 & ~n14478 ;
  assign n14480 = n14479 ^ n14473 ;
  assign n14484 = n14483 ^ n14480 ;
  assign n14570 = n14569 ^ n14484 ;
  assign n14546 = n14540 ^ n14487 ;
  assign n14547 = n14537 ^ n14489 ;
  assign n14548 = n14532 ^ n14529 ;
  assign n14549 = n14507 ^ n14499 ;
  assign n14550 = n14504 ^ n14501 ;
  assign n14347 = n14346 ^ n14343 ;
  assign n14201 = n14200 ^ n14189 ;
  assign n14202 = n14161 ^ n14103 ;
  assign n14203 = n14158 ^ n14105 ;
  assign n14204 = n14109 ^ n11539 ;
  assign n14205 = n14204 ^ n14147 ;
  assign n14206 = n14145 ^ n14142 ;
  assign n14208 = n14119 ^ n14118 ;
  assign n14209 = ~n14207 & ~n14208 ;
  assign n14210 = n14125 ^ n14122 ;
  assign n14211 = n14209 & ~n14210 ;
  assign n14212 = n14127 ^ n14115 ;
  assign n14213 = ~n14211 & n14212 ;
  assign n14214 = n14131 ^ n11557 ;
  assign n14215 = n14214 ^ n14130 ;
  assign n14216 = n14213 & n14215 ;
  assign n14217 = n14137 ^ n11553 ;
  assign n14218 = ~n14216 & ~n14217 ;
  assign n14219 = n14139 ^ n14111 ;
  assign n14220 = n14218 & n14219 ;
  assign n14221 = ~n14206 & ~n14220 ;
  assign n14222 = n14205 & n14221 ;
  assign n14223 = n14151 ^ n14108 ;
  assign n14224 = ~n14222 & ~n14223 ;
  assign n14225 = n14106 ^ n11612 ;
  assign n14226 = n14225 ^ n14154 ;
  assign n14227 = n14224 & ~n14226 ;
  assign n14228 = ~n14203 & ~n14227 ;
  assign n14229 = ~n14202 & n14228 ;
  assign n14230 = n14164 ^ n14101 ;
  assign n14231 = n14229 & n14230 ;
  assign n14232 = n14170 ^ n14167 ;
  assign n14233 = n14231 & n14232 ;
  assign n14234 = n14172 ^ n14099 ;
  assign n14235 = ~n14233 & n14234 ;
  assign n14236 = n14187 ^ n14175 ;
  assign n14237 = n14235 & ~n14236 ;
  assign n14348 = ~n14201 & ~n14237 ;
  assign n14551 = n14347 & ~n14348 ;
  assign n14552 = ~n14550 & n14551 ;
  assign n14553 = ~n14549 & n14552 ;
  assign n14554 = n14510 ^ n14497 ;
  assign n14555 = n14553 & n14554 ;
  assign n14556 = n14516 ^ n14513 ;
  assign n14557 = n14555 & n14556 ;
  assign n14558 = n14518 ^ n14495 ;
  assign n14559 = ~n14557 & ~n14558 ;
  assign n14560 = n14524 ^ n14521 ;
  assign n14561 = ~n14559 & n14560 ;
  assign n14562 = n14526 ^ n14493 ;
  assign n14563 = ~n14561 & ~n14562 ;
  assign n14564 = n14548 & ~n14563 ;
  assign n14565 = n14534 ^ n14491 ;
  assign n14566 = ~n14564 & ~n14565 ;
  assign n14567 = n14547 & n14566 ;
  assign n14568 = ~n14546 & ~n14567 ;
  assign n14584 = n14570 ^ n14568 ;
  assign n14585 = n14584 ^ n3009 ;
  assign n14586 = n14567 ^ n14546 ;
  assign n14587 = n14586 ^ n1778 ;
  assign n14590 = n14566 ^ n14547 ;
  assign n14591 = n14590 ^ n2711 ;
  assign n14592 = n14565 ^ n14564 ;
  assign n14593 = n14592 ^ n1814 ;
  assign n14596 = n14563 ^ n14548 ;
  assign n14597 = n14596 ^ n2462 ;
  assign n14599 = n14560 ^ n14559 ;
  assign n14600 = n14599 ^ n2478 ;
  assign n14601 = n14558 ^ n14557 ;
  assign n14602 = n14601 ^ n2618 ;
  assign n14603 = n14556 ^ n14555 ;
  assign n14604 = n14603 ^ n1373 ;
  assign n14606 = n14552 ^ n14549 ;
  assign n14607 = n14606 ^ n1174 ;
  assign n14349 = n14348 ^ n14347 ;
  assign n14350 = n14349 ^ n1028 ;
  assign n14238 = n14237 ^ n14201 ;
  assign n14239 = n14238 ^ n839 ;
  assign n14320 = n14236 ^ n14235 ;
  assign n14328 = n14320 ^ n14238 ;
  assign n14318 = n14234 ^ n14233 ;
  assign n14240 = n14232 ^ n14231 ;
  assign n14241 = n14240 ^ n652 ;
  assign n14314 = n14240 ^ n646 ;
  assign n14242 = n14230 ^ n14229 ;
  assign n14243 = n14242 ^ n646 ;
  assign n14244 = n14228 ^ n14202 ;
  assign n14245 = n14244 ^ n555 ;
  assign n14246 = n14227 ^ n14203 ;
  assign n14247 = n14246 ^ n613 ;
  assign n14249 = n14226 ^ n14224 ;
  assign n14250 = n14249 ^ n1486 ;
  assign n14251 = n14223 ^ n14222 ;
  assign n14252 = n14251 ^ n1480 ;
  assign n14255 = n14221 ^ n14205 ;
  assign n14256 = n14255 ^ n2906 ;
  assign n14257 = n14220 ^ n14206 ;
  assign n14261 = n14260 ^ n14257 ;
  assign n14264 = n14219 ^ n14218 ;
  assign n14265 = n14264 ^ n581 ;
  assign n14266 = n14217 ^ n14216 ;
  assign n14267 = n14266 ^ n2146 ;
  assign n14268 = n14215 ^ n14213 ;
  assign n14269 = n14268 ^ n2140 ;
  assign n14270 = n14212 ^ n14211 ;
  assign n14271 = n14270 ^ n2030 ;
  assign n14272 = n14210 ^ n14209 ;
  assign n14273 = n14272 ^ n1968 ;
  assign n14276 = n1949 & n14207 ;
  assign n14277 = n14276 ^ n1956 ;
  assign n14278 = n14208 ^ n14207 ;
  assign n14279 = n14278 ^ n1956 ;
  assign n14280 = n14277 & ~n14279 ;
  assign n14281 = n14280 ^ n14276 ;
  assign n14274 = n14270 ^ n1968 ;
  assign n14275 = n14274 ^ n14270 ;
  assign n14282 = n14281 ^ n14275 ;
  assign n14283 = ~n14273 & n14282 ;
  assign n14284 = n14283 ^ n14274 ;
  assign n14285 = n14271 & n14284 ;
  assign n14286 = n14285 ^ n14270 ;
  assign n14287 = n14286 ^ n2140 ;
  assign n14288 = ~n14269 & n14287 ;
  assign n14289 = n14288 ^ n2140 ;
  assign n14290 = n14289 ^ n14266 ;
  assign n14291 = n14267 & ~n14290 ;
  assign n14292 = n14291 ^ n2146 ;
  assign n14293 = n14292 ^ n14264 ;
  assign n14294 = n14265 & ~n14293 ;
  assign n14295 = n14294 ^ n581 ;
  assign n14262 = n14260 ^ n14255 ;
  assign n14263 = n14262 ^ n14255 ;
  assign n14296 = n14295 ^ n14263 ;
  assign n14297 = ~n14261 & n14296 ;
  assign n14298 = n14297 ^ n14262 ;
  assign n14299 = ~n14256 & n14298 ;
  assign n14300 = n14299 ^ n2906 ;
  assign n14253 = n14249 ^ n1480 ;
  assign n14254 = n14253 ^ n14249 ;
  assign n14301 = n14300 ^ n14254 ;
  assign n14302 = n14252 & n14301 ;
  assign n14303 = n14302 ^ n14253 ;
  assign n14304 = ~n14250 & n14303 ;
  assign n14305 = n14304 ^ n1486 ;
  assign n14248 = n14244 ^ n613 ;
  assign n14306 = n14305 ^ n14248 ;
  assign n14307 = n14306 ^ n14244 ;
  assign n14308 = ~n14247 & n14307 ;
  assign n14309 = n14308 ^ n14248 ;
  assign n14310 = n14245 & ~n14309 ;
  assign n14311 = n14310 ^ n555 ;
  assign n14312 = n14311 ^ n646 ;
  assign n14313 = ~n14243 & n14312 ;
  assign n14315 = n14314 ^ n14313 ;
  assign n14316 = ~n14241 & ~n14315 ;
  assign n14317 = n14316 ^ n14240 ;
  assign n14319 = n14318 ^ n14317 ;
  assign n14321 = n14320 ^ n725 ;
  assign n14322 = n14321 ^ n14320 ;
  assign n14323 = n14322 ^ n14317 ;
  assign n14324 = ~n14319 & ~n14323 ;
  assign n14325 = n14324 ^ n14321 ;
  assign n14326 = n14320 ^ n1013 ;
  assign n14327 = ~n14325 & ~n14326 ;
  assign n14329 = n14328 ^ n14327 ;
  assign n14330 = ~n14239 & ~n14329 ;
  assign n14331 = n14330 ^ n839 ;
  assign n14609 = n14349 ^ n14331 ;
  assign n14610 = ~n14350 & n14609 ;
  assign n14611 = n14610 ^ n1028 ;
  assign n14615 = n14611 ^ n14606 ;
  assign n14608 = n14551 ^ n14550 ;
  assign n14612 = n14611 ^ n14608 ;
  assign n14613 = n14608 ^ n1046 ;
  assign n14614 = ~n14612 & n14613 ;
  assign n14616 = n14615 ^ n14614 ;
  assign n14617 = ~n14607 & n14616 ;
  assign n14618 = n14617 ^ n1174 ;
  assign n14605 = n14554 ^ n14553 ;
  assign n14619 = n14618 ^ n14605 ;
  assign n14620 = n14603 ^ n1338 ;
  assign n14621 = n14620 ^ n14603 ;
  assign n14622 = n14621 ^ n14605 ;
  assign n14623 = ~n14619 & n14622 ;
  assign n14624 = n14623 ^ n14620 ;
  assign n14625 = n14604 & ~n14624 ;
  assign n14626 = n14625 ^ n1373 ;
  assign n14627 = n14626 ^ n14601 ;
  assign n14628 = ~n14602 & n14627 ;
  assign n14629 = n14628 ^ n2618 ;
  assign n14630 = n14629 ^ n14599 ;
  assign n14631 = ~n14600 & n14630 ;
  assign n14632 = n14631 ^ n2478 ;
  assign n14598 = n14562 ^ n14561 ;
  assign n14633 = n14632 ^ n14598 ;
  assign n14634 = n14596 ^ n3096 ;
  assign n14635 = n14634 ^ n14596 ;
  assign n14636 = n14635 ^ n14598 ;
  assign n14637 = n14633 & ~n14636 ;
  assign n14638 = n14637 ^ n14634 ;
  assign n14639 = ~n14597 & n14638 ;
  assign n14640 = n14639 ^ n2462 ;
  assign n14594 = n14590 ^ n1814 ;
  assign n14595 = n14594 ^ n14590 ;
  assign n14641 = n14640 ^ n14595 ;
  assign n14642 = ~n14593 & n14641 ;
  assign n14643 = n14642 ^ n14594 ;
  assign n14644 = ~n14591 & n14643 ;
  assign n14645 = n14644 ^ n2711 ;
  assign n14588 = n14584 ^ n1778 ;
  assign n14589 = n14588 ^ n14584 ;
  assign n14646 = n14645 ^ n14589 ;
  assign n14647 = n14587 & n14646 ;
  assign n14648 = n14647 ^ n14588 ;
  assign n14649 = n14585 & n14648 ;
  assign n14580 = n14483 ^ n14472 ;
  assign n14581 = ~n14480 & n14580 ;
  assign n14577 = n12358 ^ n11558 ;
  assign n14578 = n13384 & n14577 ;
  assign n14572 = n13971 ^ n2586 ;
  assign n14573 = n14572 ^ n13992 ;
  assign n14574 = n14573 ^ n14483 ;
  assign n14575 = n14574 ^ n10984 ;
  assign n14576 = n14575 ^ n3021 ;
  assign n14579 = n14578 ^ n14576 ;
  assign n14582 = n14581 ^ n14579 ;
  assign n14571 = n14568 & ~n14570 ;
  assign n14583 = n14582 ^ n14571 ;
  assign n14650 = n14649 ^ n14583 ;
  assign n14485 = n14484 ^ n10984 ;
  assign n14544 = n14543 ^ n14484 ;
  assign n14545 = ~n14485 & n14544 ;
  assign n14651 = n14650 ^ n14545 ;
  assign n14655 = n14654 ^ n14651 ;
  assign n14662 = n14645 ^ n14587 ;
  assign n14659 = n13411 ^ n12348 ;
  assign n14660 = n13749 & n14659 ;
  assign n14661 = n14660 ^ n12348 ;
  assign n14663 = n14662 ^ n14661 ;
  assign n14669 = n14643 ^ n2711 ;
  assign n14664 = n13403 ^ n12709 ;
  assign n14665 = ~n13760 & n14664 ;
  assign n14666 = n14665 ^ n12709 ;
  assign n14667 = n14640 ^ n14593 ;
  assign n14668 = n14666 & ~n14667 ;
  assign n14670 = n14669 ^ n14668 ;
  assign n14671 = n14668 ^ n12356 ;
  assign n14672 = n14671 ^ n12945 ;
  assign n14673 = n14672 ^ n14668 ;
  assign n14674 = ~n13755 & n14673 ;
  assign n14675 = n14674 ^ n14671 ;
  assign n14676 = ~n14670 & ~n14675 ;
  assign n14677 = n14676 ^ n14669 ;
  assign n14678 = n14677 ^ n14661 ;
  assign n14679 = ~n14663 & ~n14678 ;
  assign n14680 = n14679 ^ n14662 ;
  assign n14656 = n12933 ^ n12725 ;
  assign n14657 = n14061 & n14656 ;
  assign n14658 = n14657 ^ n12725 ;
  assign n14681 = n14680 ^ n14658 ;
  assign n14682 = n14648 ^ n3009 ;
  assign n14683 = n14682 ^ n14680 ;
  assign n14684 = n14681 & n14683 ;
  assign n14685 = n14684 ^ n14682 ;
  assign n14686 = n14685 ^ n14651 ;
  assign n14687 = ~n14655 & n14686 ;
  assign n14688 = n14687 ^ n14654 ;
  assign n14689 = n14688 ^ n14377 ;
  assign n14690 = n14382 & n14689 ;
  assign n14691 = n14690 ^ n14377 ;
  assign n14375 = n14278 ^ n14277 ;
  assign n14372 = n12936 ^ n12907 ;
  assign n14373 = ~n13738 & ~n14372 ;
  assign n14374 = n14373 ^ n12936 ;
  assign n14376 = n14375 ^ n14374 ;
  assign n14734 = n14691 ^ n14376 ;
  assign n14802 = n14734 ^ n12103 ;
  assign n14735 = n14688 ^ n14382 ;
  assign n14736 = n14735 ^ n12093 ;
  assign n14738 = n14682 ^ n14658 ;
  assign n14739 = n14738 ^ n14680 ;
  assign n14740 = n14739 ^ n11544 ;
  assign n14748 = n14677 ^ n14663 ;
  assign n14743 = n14675 ^ n14669 ;
  assign n14741 = n14667 ^ n14666 ;
  assign n14742 = n12070 & ~n14741 ;
  assign n14744 = n14743 ^ n14742 ;
  assign n14745 = n14743 ^ n11551 ;
  assign n14746 = n14744 & n14745 ;
  assign n14747 = n14746 ^ n11551 ;
  assign n14749 = n14748 ^ n14747 ;
  assign n14750 = n14748 ^ n12077 ;
  assign n14751 = n14749 & n14750 ;
  assign n14752 = n14751 ^ n12077 ;
  assign n14753 = n14752 ^ n14739 ;
  assign n14754 = n14740 & n14753 ;
  assign n14755 = n14754 ^ n11544 ;
  assign n14737 = n14685 ^ n14655 ;
  assign n14756 = n14755 ^ n14737 ;
  assign n14757 = n14755 ^ n11537 ;
  assign n14758 = ~n14756 & n14757 ;
  assign n14759 = n14758 ^ n11537 ;
  assign n14760 = n14759 ^ n14735 ;
  assign n14761 = n14736 & n14760 ;
  assign n14762 = n14761 ^ n12093 ;
  assign n14803 = n14802 ^ n14762 ;
  assign n14789 = n14759 ^ n14736 ;
  assign n14790 = n14737 ^ n11537 ;
  assign n14791 = n14790 ^ n14755 ;
  assign n14792 = n14750 ^ n14747 ;
  assign n14793 = n14741 ^ n12070 ;
  assign n14794 = n14742 ^ n11551 ;
  assign n14795 = n14794 ^ n14743 ;
  assign n14796 = ~n14793 & n14795 ;
  assign n14797 = ~n14792 & n14796 ;
  assign n14798 = n14752 ^ n14740 ;
  assign n14799 = ~n14797 & ~n14798 ;
  assign n14800 = n14791 & n14799 ;
  assign n14801 = ~n14789 & ~n14800 ;
  assign n14830 = n14803 ^ n14801 ;
  assign n14831 = n14830 ^ n1460 ;
  assign n14832 = n14800 ^ n14789 ;
  assign n14833 = n14832 ^ n2223 ;
  assign n14834 = n14799 ^ n14791 ;
  assign n14835 = n14834 ^ n2122 ;
  assign n14836 = n14798 ^ n14797 ;
  assign n14837 = n14836 ^ n2102 ;
  assign n14838 = n14796 ^ n14792 ;
  assign n14839 = n14838 ^ n2106 ;
  assign n14842 = n3068 ^ x160 ;
  assign n14843 = n14842 ^ x352 ;
  assign n14844 = n14843 ^ x96 ;
  assign n14845 = n14793 & n14844 ;
  assign n1896 = n1871 ^ x191 ;
  assign n1897 = n1896 ^ x383 ;
  assign n1898 = n1897 ^ x127 ;
  assign n14846 = n14845 ^ n1898 ;
  assign n14847 = n14795 ^ n14793 ;
  assign n14848 = n14847 ^ n1898 ;
  assign n14849 = n14846 & n14848 ;
  assign n14850 = n14849 ^ n14845 ;
  assign n14840 = n14836 ^ n2106 ;
  assign n14841 = n14840 ^ n14836 ;
  assign n14851 = n14850 ^ n14841 ;
  assign n14852 = ~n14839 & n14851 ;
  assign n14853 = n14852 ^ n14840 ;
  assign n14854 = ~n14837 & n14853 ;
  assign n14855 = n14854 ^ n2102 ;
  assign n14856 = n14855 ^ n2122 ;
  assign n14857 = ~n14835 & n14856 ;
  assign n14858 = n14857 ^ n2122 ;
  assign n14859 = n14858 ^ n2223 ;
  assign n14860 = n14833 & ~n14859 ;
  assign n14861 = n14860 ^ n14832 ;
  assign n14862 = n14861 ^ n1460 ;
  assign n14863 = ~n14831 & n14862 ;
  assign n14864 = n14863 ^ n1460 ;
  assign n14804 = n14801 & ~n14803 ;
  assign n14763 = n14762 ^ n14734 ;
  assign n14764 = n14762 ^ n12103 ;
  assign n14765 = n14763 & n14764 ;
  assign n14766 = n14765 ^ n12103 ;
  assign n14696 = n14281 ^ n14273 ;
  assign n14369 = n12940 ^ n12900 ;
  assign n14370 = n13736 & ~n14369 ;
  assign n14371 = n14370 ^ n12940 ;
  assign n14731 = n14696 ^ n14371 ;
  assign n14692 = n14691 ^ n14374 ;
  assign n14693 = ~n14376 & n14692 ;
  assign n14694 = n14693 ^ n14375 ;
  assign n14732 = n14731 ^ n14694 ;
  assign n14733 = n14732 ^ n11531 ;
  assign n14788 = n14766 ^ n14733 ;
  assign n14826 = n14804 ^ n14788 ;
  assign n14827 = n14826 ^ n2372 ;
  assign n14932 = n14864 ^ n14827 ;
  assign n14718 = n14295 ^ n14261 ;
  assign n16276 = n14932 ^ n14718 ;
  assign n15340 = n14067 ^ n13411 ;
  assign n15341 = n15340 ^ n14696 ;
  assign n14983 = n13726 ^ n12960 ;
  assign n14984 = ~n14402 & n14983 ;
  assign n14985 = n14984 ^ n12960 ;
  assign n14930 = n14309 ^ n555 ;
  assign n15020 = n14985 ^ n14930 ;
  assign n14987 = n14930 ^ n12971 ;
  assign n14988 = n14987 ^ n13770 ;
  assign n14989 = n14988 ^ n14930 ;
  assign n14990 = n14408 & ~n14989 ;
  assign n14991 = n14990 ^ n14987 ;
  assign n14992 = n13794 ^ n12343 ;
  assign n14993 = n14418 & ~n14992 ;
  assign n14994 = n14993 ^ n12343 ;
  assign n14942 = n14303 ^ n1486 ;
  assign n14995 = n14994 ^ n14942 ;
  assign n14947 = n14300 ^ n14252 ;
  assign n14996 = n14947 ^ n13046 ;
  assign n14997 = n14996 ^ n13785 ;
  assign n14998 = n14997 ^ n14947 ;
  assign n14999 = ~n14426 & ~n14998 ;
  assign n15000 = n14999 ^ n14996 ;
  assign n14719 = n14718 ^ n12899 ;
  assign n14720 = n14719 ^ n13594 ;
  assign n14721 = n14720 ^ n14718 ;
  assign n14722 = n14190 & n14721 ;
  assign n14723 = n14722 ^ n14719 ;
  assign n14356 = n14292 ^ n14265 ;
  assign n14353 = n13454 ^ n12906 ;
  assign n14354 = ~n14176 & ~n14353 ;
  assign n14355 = n14354 ^ n12906 ;
  assign n14357 = n14356 ^ n14355 ;
  assign n14358 = n14289 ^ n14267 ;
  assign n14714 = n14358 ^ n14355 ;
  assign n14359 = n14358 ^ n12913 ;
  assign n14360 = n14359 ^ n12897 ;
  assign n14361 = n14360 ^ n14358 ;
  assign n14362 = n14097 & n14361 ;
  assign n14363 = n14362 ^ n14359 ;
  assign n14365 = n13447 ^ n12920 ;
  assign n14366 = ~n14084 & n14365 ;
  assign n14367 = n14366 ^ n12920 ;
  assign n14364 = n14286 ^ n14269 ;
  assign n14368 = n14367 ^ n14364 ;
  assign n14700 = n14284 ^ n2030 ;
  assign n14695 = n14694 ^ n14371 ;
  assign n14697 = n14696 ^ n14694 ;
  assign n14698 = n14695 & ~n14697 ;
  assign n14699 = n14698 ^ n14696 ;
  assign n14701 = n14700 ^ n14699 ;
  assign n14702 = n14700 ^ n12928 ;
  assign n14703 = n14702 ^ n13440 ;
  assign n14704 = n14703 ^ n14700 ;
  assign n14705 = ~n13728 & ~n14704 ;
  assign n14706 = n14705 ^ n14702 ;
  assign n14707 = ~n14701 & ~n14706 ;
  assign n14708 = n14707 ^ n14700 ;
  assign n14709 = n14708 ^ n14367 ;
  assign n14710 = ~n14368 & ~n14709 ;
  assign n14711 = n14710 ^ n14708 ;
  assign n14712 = n14711 ^ n14358 ;
  assign n14713 = n14363 & n14712 ;
  assign n14715 = n14714 ^ n14713 ;
  assign n14716 = ~n14357 & n14715 ;
  assign n14717 = n14716 ^ n14356 ;
  assign n14888 = n14718 ^ n14717 ;
  assign n14889 = ~n14723 & ~n14888 ;
  assign n14884 = n13616 ^ n12982 ;
  assign n14885 = n14333 & ~n14884 ;
  assign n14886 = n14885 ^ n12982 ;
  assign n14887 = n14886 ^ n14718 ;
  assign n14890 = n14889 ^ n14887 ;
  assign n14891 = n14298 ^ n2906 ;
  assign n15001 = n14891 ^ n14886 ;
  assign n15002 = n14890 & ~n15001 ;
  assign n15003 = n15002 ^ n14891 ;
  assign n15004 = n15003 ^ n14947 ;
  assign n15005 = ~n15000 & ~n15004 ;
  assign n15006 = n15005 ^ n14947 ;
  assign n15007 = n15006 ^ n14994 ;
  assign n15008 = ~n14995 & ~n15007 ;
  assign n15009 = n15008 ^ n14942 ;
  assign n14935 = n14305 ^ n14247 ;
  assign n15010 = n15009 ^ n14935 ;
  assign n15012 = n14935 ^ n12976 ;
  assign n15011 = n14935 ^ n13776 ;
  assign n15013 = n15012 ^ n15011 ;
  assign n15014 = n14416 & n15013 ;
  assign n15015 = n15014 ^ n15012 ;
  assign n15016 = n15010 & n15015 ;
  assign n15017 = n15016 ^ n14935 ;
  assign n15018 = n15017 ^ n14930 ;
  assign n15019 = ~n14991 & ~n15018 ;
  assign n15021 = n15020 ^ n15019 ;
  assign n14925 = n14311 ^ n14243 ;
  assign n15077 = n15021 ^ n14925 ;
  assign n15079 = n15077 ^ n12390 ;
  assign n15054 = n15017 ^ n14991 ;
  assign n15055 = n15054 ^ n12344 ;
  assign n15056 = n15015 ^ n15009 ;
  assign n15057 = n15056 ^ n12399 ;
  assign n15062 = n15003 ^ n15000 ;
  assign n14892 = n14891 ^ n14890 ;
  assign n14893 = n14892 ^ n12413 ;
  assign n14724 = n14723 ^ n14717 ;
  assign n14725 = n14724 ^ n12422 ;
  assign n14726 = n14715 ^ n14356 ;
  assign n14727 = n14726 ^ n12433 ;
  assign n14777 = n14711 ^ n14363 ;
  assign n14728 = n14708 ^ n14368 ;
  assign n14729 = n14728 ^ n12197 ;
  assign n14767 = n14766 ^ n14732 ;
  assign n14768 = ~n14733 & ~n14767 ;
  assign n14769 = n14768 ^ n11531 ;
  assign n14730 = n14706 ^ n14699 ;
  assign n14770 = n14769 ^ n14730 ;
  assign n14771 = n14769 ^ n12118 ;
  assign n14772 = n14770 & ~n14771 ;
  assign n14773 = n14772 ^ n12118 ;
  assign n14774 = n14773 ^ n14728 ;
  assign n14775 = n14729 & ~n14774 ;
  assign n14776 = n14775 ^ n12197 ;
  assign n14778 = n14777 ^ n14776 ;
  assign n14779 = n14777 ^ n12337 ;
  assign n14780 = ~n14778 & n14779 ;
  assign n14781 = n14780 ^ n12337 ;
  assign n14782 = n14781 ^ n14726 ;
  assign n14783 = ~n14727 & n14782 ;
  assign n14784 = n14783 ^ n12433 ;
  assign n14881 = n14784 ^ n14724 ;
  assign n14882 = n14725 & n14881 ;
  assign n14883 = n14882 ^ n12422 ;
  assign n15059 = n14892 ^ n14883 ;
  assign n15060 = n14893 & n15059 ;
  assign n15061 = n15060 ^ n12413 ;
  assign n15063 = n15062 ^ n15061 ;
  assign n15064 = n15062 ^ n12407 ;
  assign n15065 = ~n15063 & ~n15064 ;
  assign n15066 = n15065 ^ n12407 ;
  assign n15058 = n15006 ^ n14995 ;
  assign n15067 = n15066 ^ n15058 ;
  assign n15068 = n15066 ^ n12402 ;
  assign n15069 = ~n15067 & n15068 ;
  assign n15070 = n15069 ^ n12402 ;
  assign n15071 = n15070 ^ n15056 ;
  assign n15072 = ~n15057 & ~n15071 ;
  assign n15073 = n15072 ^ n12399 ;
  assign n15074 = n15073 ^ n15054 ;
  assign n15075 = n15055 & ~n15074 ;
  assign n15076 = n15075 ^ n12344 ;
  assign n15111 = n15079 ^ n15076 ;
  assign n15112 = n15073 ^ n15055 ;
  assign n15113 = n15058 ^ n12402 ;
  assign n15114 = n15113 ^ n15066 ;
  assign n14894 = n14893 ^ n14883 ;
  assign n14785 = n14784 ^ n14725 ;
  assign n14786 = n14730 ^ n12118 ;
  assign n14787 = n14786 ^ n14769 ;
  assign n14805 = n14788 & ~n14804 ;
  assign n14806 = n14787 & n14805 ;
  assign n14807 = n14773 ^ n14729 ;
  assign n14808 = ~n14806 & n14807 ;
  assign n14809 = n14779 ^ n14776 ;
  assign n14810 = n14808 & n14809 ;
  assign n14811 = n14781 ^ n14727 ;
  assign n14812 = ~n14810 & n14811 ;
  assign n14895 = ~n14785 & n14812 ;
  assign n15115 = n14894 & n14895 ;
  assign n15116 = n15064 ^ n15061 ;
  assign n15117 = n15115 & n15116 ;
  assign n15118 = ~n15114 & ~n15117 ;
  assign n15119 = n15070 ^ n15057 ;
  assign n15120 = n15118 & n15119 ;
  assign n15121 = ~n15112 & ~n15120 ;
  assign n15122 = n15111 & ~n15121 ;
  assign n15078 = n15077 ^ n15076 ;
  assign n15080 = ~n15078 & n15079 ;
  assign n15081 = n15080 ^ n12390 ;
  assign n14917 = n14315 ^ n652 ;
  assign n15025 = n14917 ^ n13076 ;
  assign n15026 = n15025 ^ n13822 ;
  assign n15027 = n15026 ^ n14917 ;
  assign n15028 = n14447 & ~n15027 ;
  assign n15029 = n15028 ^ n15025 ;
  assign n14986 = n14985 ^ n14925 ;
  assign n15022 = n14986 & n15021 ;
  assign n15023 = n15022 ^ n14925 ;
  assign n15052 = n15029 ^ n15023 ;
  assign n15053 = n15052 ^ n12385 ;
  assign n15123 = n15081 ^ n15053 ;
  assign n15124 = n15122 & ~n15123 ;
  assign n14913 = n14318 ^ n725 ;
  assign n14914 = n14913 ^ n14317 ;
  assign n15033 = n14914 ^ n13083 ;
  assign n15034 = n15033 ^ n13830 ;
  assign n15035 = n15034 ^ n14914 ;
  assign n15036 = ~n13725 & ~n15035 ;
  assign n15037 = n15036 ^ n15033 ;
  assign n15024 = n15023 ^ n14917 ;
  assign n15030 = n15024 & ~n15029 ;
  assign n15031 = n15030 ^ n14917 ;
  assign n15085 = n15037 ^ n15031 ;
  assign n15087 = n15085 ^ n12379 ;
  assign n15082 = n15081 ^ n15052 ;
  assign n15083 = ~n15053 & ~n15082 ;
  assign n15084 = n15083 ^ n12385 ;
  assign n15125 = n15087 ^ n15084 ;
  assign n15126 = n15124 & ~n15125 ;
  assign n15086 = n15085 ^ n15084 ;
  assign n15088 = ~n15086 & n15087 ;
  assign n15089 = n15088 ^ n12379 ;
  assign n15032 = n15031 ^ n14914 ;
  assign n15038 = ~n15032 & ~n15037 ;
  assign n15039 = n15038 ^ n15031 ;
  assign n14907 = n14325 ^ n1013 ;
  assign n14978 = n14907 ^ n13171 ;
  assign n14979 = n14978 ^ n13837 ;
  assign n14980 = n14979 ^ n14907 ;
  assign n14981 = n14389 & ~n14980 ;
  assign n14982 = n14981 ^ n14978 ;
  assign n15050 = n15039 ^ n14982 ;
  assign n15051 = n15050 ^ n12370 ;
  assign n15127 = n15089 ^ n15051 ;
  assign n15128 = n15126 & ~n15127 ;
  assign n15090 = n15089 ^ n15050 ;
  assign n15091 = n15051 & n15090 ;
  assign n15092 = n15091 ^ n12370 ;
  assign n15129 = n15092 ^ n12464 ;
  assign n14903 = n14329 ^ n839 ;
  assign n15042 = n14907 ^ n14903 ;
  assign n15040 = n15039 ^ n14907 ;
  assign n15041 = ~n14982 & n15040 ;
  assign n15043 = n15042 ^ n15041 ;
  assign n14974 = n13836 ^ n13295 ;
  assign n14975 = n14383 & n14974 ;
  assign n14976 = n14975 ^ n13295 ;
  assign n15048 = n15043 ^ n14976 ;
  assign n15130 = n15129 ^ n15048 ;
  assign n15131 = n15128 & n15130 ;
  assign n15049 = n15048 ^ n12464 ;
  assign n15093 = n15092 ^ n15048 ;
  assign n15094 = n15049 & ~n15093 ;
  assign n15095 = n15094 ^ n12464 ;
  assign n14977 = n14976 ^ n14903 ;
  assign n15044 = ~n14977 & n15043 ;
  assign n15045 = n15044 ^ n14976 ;
  assign n14351 = n14350 ^ n14331 ;
  assign n14969 = n14351 ^ n13343 ;
  assign n14970 = n14969 ^ n13847 ;
  assign n14971 = n14970 ^ n14351 ;
  assign n14972 = n14465 & ~n14971 ;
  assign n14973 = n14972 ^ n14969 ;
  assign n15046 = n15045 ^ n14973 ;
  assign n15047 = n15046 ^ n12646 ;
  assign n15132 = n15095 ^ n15047 ;
  assign n15133 = ~n15131 & ~n15132 ;
  assign n15105 = n15045 ^ n14351 ;
  assign n15106 = ~n14973 & n15105 ;
  assign n15107 = n15106 ^ n14351 ;
  assign n15099 = n14613 ^ n14611 ;
  assign n15100 = n15099 ^ n13374 ;
  assign n15101 = n15100 ^ n13988 ;
  assign n15102 = n15101 ^ n15099 ;
  assign n15103 = ~n14468 & n15102 ;
  assign n15104 = n15103 ^ n15100 ;
  assign n15108 = n15107 ^ n15104 ;
  assign n15109 = n15108 ^ n12686 ;
  assign n15096 = n15095 ^ n15046 ;
  assign n15097 = n15047 & ~n15096 ;
  assign n15098 = n15097 ^ n12646 ;
  assign n15110 = n15109 ^ n15098 ;
  assign n15153 = n15133 ^ n15110 ;
  assign n15154 = n15153 ^ n2563 ;
  assign n15155 = n15132 ^ n15131 ;
  assign n15156 = n15155 ^ n2821 ;
  assign n15157 = n15130 ^ n15128 ;
  assign n15158 = n15157 ^ n2796 ;
  assign n15160 = n15125 ^ n15124 ;
  assign n15161 = n15160 ^ n1305 ;
  assign n15187 = n15121 ^ n15111 ;
  assign n15163 = n15120 ^ n15112 ;
  assign n15164 = n15163 ^ n912 ;
  assign n15167 = n15119 ^ n15118 ;
  assign n15183 = n15167 ^ n15163 ;
  assign n15165 = n15117 ^ n15114 ;
  assign n15166 = n15165 ^ n720 ;
  assign n15170 = n15116 ^ n15115 ;
  assign n15171 = n15170 ^ n708 ;
  assign n15174 = n15170 ^ n702 ;
  assign n14896 = n14895 ^ n14894 ;
  assign n14897 = n14896 ^ n702 ;
  assign n14813 = n14812 ^ n14785 ;
  assign n14814 = n14813 ^ n1529 ;
  assign n14815 = n14811 ^ n14810 ;
  assign n14816 = n14815 ^ n1523 ;
  assign n14819 = n14809 ^ n14808 ;
  assign n14820 = n14819 ^ n518 ;
  assign n14821 = n14807 ^ n14806 ;
  assign n14822 = n14821 ^ n2920 ;
  assign n14824 = n14805 ^ n14787 ;
  assign n14825 = n14824 ^ n569 ;
  assign n14828 = n14824 ^ n2372 ;
  assign n14829 = n14828 ^ n14824 ;
  assign n14865 = n14864 ^ n14829 ;
  assign n14866 = n14827 & n14865 ;
  assign n14867 = n14866 ^ n14828 ;
  assign n14868 = ~n14825 & n14867 ;
  assign n14869 = n14868 ^ n569 ;
  assign n14823 = n14819 ^ n2920 ;
  assign n14870 = n14869 ^ n14823 ;
  assign n14871 = n14870 ^ n14819 ;
  assign n14872 = ~n14822 & n14871 ;
  assign n14873 = n14872 ^ n14823 ;
  assign n14874 = n14820 & ~n14873 ;
  assign n14875 = n14874 ^ n518 ;
  assign n14817 = n14813 ^ n1523 ;
  assign n14818 = n14817 ^ n14813 ;
  assign n14876 = n14875 ^ n14818 ;
  assign n14877 = n14816 & n14876 ;
  assign n14878 = n14877 ^ n14817 ;
  assign n14879 = n14814 & n14878 ;
  assign n14880 = n14879 ^ n14813 ;
  assign n15172 = n14880 ^ n702 ;
  assign n15173 = ~n14897 & n15172 ;
  assign n15175 = n15174 ^ n15173 ;
  assign n15176 = ~n15171 & ~n15175 ;
  assign n15177 = n15176 ^ n15170 ;
  assign n15168 = n15167 ^ n720 ;
  assign n15169 = n15168 ^ n15167 ;
  assign n15178 = n15177 ^ n15169 ;
  assign n15179 = n15166 & ~n15178 ;
  assign n15180 = n15179 ^ n15168 ;
  assign n15181 = n15167 ^ n785 ;
  assign n15182 = n15180 & n15181 ;
  assign n15184 = n15183 ^ n15182 ;
  assign n15185 = ~n15164 & n15184 ;
  assign n15186 = n15185 ^ n912 ;
  assign n15188 = n15187 ^ n15186 ;
  assign n894 = n830 ^ x174 ;
  assign n895 = n894 ^ x366 ;
  assign n896 = n895 ^ x110 ;
  assign n15189 = n15187 ^ n896 ;
  assign n15190 = n15188 & ~n15189 ;
  assign n15191 = n15190 ^ n896 ;
  assign n15162 = n15123 ^ n15122 ;
  assign n15192 = n15191 ^ n15162 ;
  assign n15193 = n15160 ^ n1061 ;
  assign n15194 = n15193 ^ n15160 ;
  assign n15195 = n15194 ^ n15162 ;
  assign n15196 = n15192 & ~n15195 ;
  assign n15197 = n15196 ^ n15193 ;
  assign n15198 = ~n15161 & n15197 ;
  assign n15199 = n15198 ^ n1305 ;
  assign n15159 = n15127 ^ n15126 ;
  assign n15200 = n15199 ^ n15159 ;
  assign n15201 = n15157 ^ n1256 ;
  assign n15202 = n15201 ^ n15157 ;
  assign n15203 = n15202 ^ n15159 ;
  assign n15204 = n15200 & ~n15203 ;
  assign n15205 = n15204 ^ n15201 ;
  assign n15206 = n15158 & ~n15205 ;
  assign n15207 = n15206 ^ n2796 ;
  assign n15208 = n15207 ^ n15155 ;
  assign n15209 = ~n15156 & n15208 ;
  assign n15210 = n15209 ^ n2821 ;
  assign n15211 = n15210 ^ n15153 ;
  assign n15212 = ~n15154 & n15211 ;
  assign n15213 = n15212 ^ n2563 ;
  assign n15135 = n15108 ^ n15098 ;
  assign n15144 = n14616 ^ n1174 ;
  assign n15136 = n15107 ^ n15099 ;
  assign n15137 = ~n15104 & n15136 ;
  assign n15138 = n15137 ^ n15099 ;
  assign n15139 = n15138 ^ n12631 ;
  assign n15140 = n15139 ^ n13316 ;
  assign n15141 = n15140 ^ n15138 ;
  assign n15142 = ~n14472 & ~n15141 ;
  assign n15143 = n15142 ^ n15139 ;
  assign n15145 = n15144 ^ n15143 ;
  assign n15146 = n15145 ^ n12686 ;
  assign n15147 = n15146 ^ n15098 ;
  assign n15148 = n15147 ^ n15145 ;
  assign n15149 = ~n15135 & n15148 ;
  assign n15150 = n15149 ^ n15146 ;
  assign n15151 = n15150 ^ n12040 ;
  assign n15134 = n15110 & ~n15133 ;
  assign n15152 = n15151 ^ n15134 ;
  assign n15214 = n15213 ^ n15152 ;
  assign n15227 = n14605 ^ n1338 ;
  assign n15228 = n15227 ^ n14618 ;
  assign n15219 = n13315 ^ n12627 ;
  assign n15220 = ~n14572 & ~n15219 ;
  assign n15221 = n15220 ^ n12627 ;
  assign n15223 = n15221 ^ n15138 ;
  assign n15222 = n15221 ^ n15144 ;
  assign n15224 = n15223 ^ n15222 ;
  assign n15225 = n15143 & n15224 ;
  assign n15226 = n15225 ^ n15223 ;
  assign n15229 = n15228 ^ n15226 ;
  assign n15230 = n15229 ^ n12050 ;
  assign n15216 = n15145 ^ n12040 ;
  assign n15217 = n15150 & n15216 ;
  assign n15218 = n15217 ^ n12040 ;
  assign n15231 = n15230 ^ n15218 ;
  assign n15215 = ~n15134 & ~n15151 ;
  assign n15232 = n15231 ^ n15215 ;
  assign n15233 = n15232 ^ n2569 ;
  assign n15234 = n15233 ^ n15152 ;
  assign n15235 = n15234 ^ n15232 ;
  assign n15236 = n15214 & ~n15235 ;
  assign n15237 = n15236 ^ n15233 ;
  assign n15250 = n15229 ^ n15218 ;
  assign n15251 = n15230 & ~n15250 ;
  assign n15252 = n15251 ^ n12050 ;
  assign n15247 = n14624 ^ n1373 ;
  assign n15239 = n13312 ^ n12621 ;
  assign n15240 = ~n14025 & ~n15239 ;
  assign n15241 = n15240 ^ n12621 ;
  assign n15243 = n15241 ^ n15221 ;
  assign n15242 = n15241 ^ n15228 ;
  assign n15244 = n15243 ^ n15242 ;
  assign n15245 = ~n15226 & n15244 ;
  assign n15246 = n15245 ^ n15243 ;
  assign n15248 = n15247 ^ n15246 ;
  assign n15249 = n15248 ^ n12038 ;
  assign n15253 = n15252 ^ n15249 ;
  assign n15238 = ~n15215 & ~n15231 ;
  assign n15254 = n15253 ^ n15238 ;
  assign n15256 = n15254 ^ n2490 ;
  assign n15255 = n15254 ^ n15232 ;
  assign n15257 = n15256 ^ n15255 ;
  assign n15258 = ~n15237 & n15257 ;
  assign n15259 = n15258 ^ n15256 ;
  assign n15260 = n15259 ^ n2447 ;
  assign n15261 = n14377 ^ n13403 ;
  assign n15262 = n15261 ^ n13749 ;
  assign n15263 = n15260 & n15262 ;
  assign n14967 = n14061 ^ n12945 ;
  assign n14968 = n14967 ^ n14375 ;
  assign n15264 = n15263 ^ n14968 ;
  assign n15278 = n14626 ^ n14602 ;
  assign n15270 = n13355 ^ n12669 ;
  assign n15271 = ~n14020 & ~n15270 ;
  assign n15272 = n15271 ^ n12669 ;
  assign n15274 = n15272 ^ n15241 ;
  assign n15273 = n15272 ^ n15247 ;
  assign n15275 = n15274 ^ n15273 ;
  assign n15276 = n15246 & n15275 ;
  assign n15277 = n15276 ^ n15274 ;
  assign n15279 = n15278 ^ n15277 ;
  assign n15280 = n15279 ^ n12029 ;
  assign n15266 = n15252 ^ n15248 ;
  assign n15267 = n15252 ^ n12038 ;
  assign n15268 = n15266 & ~n15267 ;
  assign n15269 = n15268 ^ n12038 ;
  assign n15281 = n15280 ^ n15269 ;
  assign n15265 = ~n15238 & n15253 ;
  assign n15282 = n15281 ^ n15265 ;
  assign n15285 = n15282 ^ n2447 ;
  assign n15284 = n15282 ^ n15254 ;
  assign n15286 = n15285 ^ n15284 ;
  assign n15287 = ~n15259 & n15286 ;
  assign n15288 = n15287 ^ n15285 ;
  assign n15312 = n15288 ^ n2472 ;
  assign n15303 = n15279 ^ n15269 ;
  assign n15304 = ~n15280 & n15303 ;
  assign n15305 = n15304 ^ n12029 ;
  assign n15295 = n14629 ^ n14600 ;
  assign n15297 = n15295 ^ n15272 ;
  assign n15296 = n15295 ^ n15278 ;
  assign n15298 = n15297 ^ n15296 ;
  assign n15299 = n15277 & ~n15298 ;
  assign n15300 = n15299 ^ n15297 ;
  assign n15292 = n13384 ^ n12697 ;
  assign n15293 = n14018 & n15292 ;
  assign n15294 = n15293 ^ n13384 ;
  assign n15301 = n15300 ^ n15294 ;
  assign n15302 = n15301 ^ n12024 ;
  assign n15306 = n15305 ^ n15302 ;
  assign n15291 = n15265 & n15281 ;
  assign n15307 = n15306 ^ n15291 ;
  assign n15308 = n15307 ^ n1808 ;
  assign n15283 = n15282 ^ n2472 ;
  assign n15289 = ~n15283 & n15288 ;
  assign n15290 = n15289 ^ n2472 ;
  assign n15309 = n15308 ^ n15290 ;
  assign n15310 = n15309 ^ n14968 ;
  assign n15311 = n15310 ^ n15309 ;
  assign n15313 = n15312 ^ n15311 ;
  assign n15314 = n15264 & ~n15313 ;
  assign n15315 = n15314 ^ n15310 ;
  assign n15452 = n15341 ^ n15315 ;
  assign n15538 = n15452 ^ n12348 ;
  assign n15454 = n15262 ^ n15260 ;
  assign n15455 = n12709 & n15454 ;
  assign n15453 = n15312 ^ n15264 ;
  assign n15456 = n15455 ^ n15453 ;
  assign n15457 = n15455 ^ n12356 ;
  assign n15458 = n15456 & n15457 ;
  assign n15459 = n15458 ^ n12356 ;
  assign n15539 = n15538 ^ n15459 ;
  assign n15535 = n15457 ^ n15453 ;
  assign n15536 = n15454 ^ n12709 ;
  assign n15537 = ~n15535 & n15536 ;
  assign n15608 = n15539 ^ n15537 ;
  assign n1940 = n1909 ^ x222 ;
  assign n1941 = n1940 ^ x414 ;
  assign n1942 = n1941 ^ x158 ;
  assign n15609 = n15608 ^ n1942 ;
  assign n15610 = n15536 ^ n15535 ;
  assign n1934 = n1903 ^ x223 ;
  assign n1935 = n1934 ^ x415 ;
  assign n1936 = n1935 ^ x159 ;
  assign n15611 = n15610 ^ n1936 ;
  assign n1887 = n1862 ^ x192 ;
  assign n1888 = n1887 ^ x384 ;
  assign n1889 = n1888 ^ x128 ;
  assign n15612 = n1889 & ~n15536 ;
  assign n15613 = n15612 ^ n1936 ;
  assign n15614 = ~n15611 & ~n15613 ;
  assign n15615 = n15614 ^ n15610 ;
  assign n15616 = n15615 ^ n1942 ;
  assign n15617 = n15609 & ~n15616 ;
  assign n15618 = n15617 ^ n1942 ;
  assign n15622 = n15618 ^ n2325 ;
  assign n15460 = n15459 ^ n15452 ;
  assign n15461 = n15459 ^ n12348 ;
  assign n15462 = n15460 & ~n15461 ;
  assign n15463 = n15462 ^ n12348 ;
  assign n15368 = n13744 ^ n12933 ;
  assign n15369 = n15368 ^ n14700 ;
  assign n15328 = n15305 ^ n12024 ;
  assign n15329 = n15302 & n15328 ;
  assign n15330 = n15329 ^ n15305 ;
  assign n15331 = n15330 ^ n11569 ;
  assign n15324 = n12950 ^ n12702 ;
  assign n15325 = ~n14009 & ~n15324 ;
  assign n15326 = n15325 ^ n12702 ;
  assign n15317 = n14598 ^ n3096 ;
  assign n15318 = n15317 ^ n14632 ;
  assign n15319 = n15318 ^ n15295 ;
  assign n15320 = n15319 ^ n15318 ;
  assign n15321 = n15320 ^ n15294 ;
  assign n15322 = ~n15300 & ~n15321 ;
  assign n15323 = n15322 ^ n15319 ;
  assign n15327 = n15326 ^ n15323 ;
  assign n15332 = n15331 ^ n15327 ;
  assign n15316 = ~n15291 & ~n15306 ;
  assign n15333 = n15332 ^ n15316 ;
  assign n15334 = n15333 ^ n1808 ;
  assign n15335 = n15334 ^ n15290 ;
  assign n15336 = n15335 ^ n15333 ;
  assign n15337 = n15308 & n15336 ;
  assign n15338 = n15337 ^ n15334 ;
  assign n15339 = n15338 ^ n1799 ;
  assign n15343 = n15339 ^ n15309 ;
  assign n15342 = n15341 ^ n15339 ;
  assign n15344 = n15343 ^ n15342 ;
  assign n15345 = n15315 & ~n15344 ;
  assign n15346 = n15345 ^ n15343 ;
  assign n15450 = n15369 ^ n15346 ;
  assign n15451 = n15450 ^ n12725 ;
  assign n15541 = n15463 ^ n15451 ;
  assign n15540 = n15537 & n15539 ;
  assign n15607 = n15541 ^ n15540 ;
  assign n15619 = n15618 ^ n15607 ;
  assign n2017 = n1974 ^ x221 ;
  assign n2018 = n2017 ^ x413 ;
  assign n2019 = n2018 ^ x157 ;
  assign n15620 = n15607 ^ n2019 ;
  assign n15621 = n15619 & ~n15620 ;
  assign n15623 = n15622 ^ n15621 ;
  assign n15464 = n15463 ^ n15450 ;
  assign n15465 = ~n15451 & n15464 ;
  assign n15466 = n15465 ^ n12725 ;
  assign n15376 = n13738 ^ n12922 ;
  assign n15377 = n15376 ^ n14364 ;
  assign n15364 = n15316 & n15332 ;
  assign n15357 = n14638 ^ n2462 ;
  assign n15358 = n15357 ^ n12358 ;
  assign n15356 = n15318 ^ n11558 ;
  assign n15359 = n15358 ^ n15356 ;
  assign n15360 = n15359 ^ n11569 ;
  assign n15361 = n15360 ^ n1791 ;
  assign n15354 = n15326 ^ n15318 ;
  assign n15355 = n15323 & n15354 ;
  assign n15362 = n15361 ^ n15355 ;
  assign n15352 = n13389 ^ n12358 ;
  assign n15353 = n14004 & ~n15352 ;
  assign n15363 = n15362 ^ n15353 ;
  assign n15365 = n15364 ^ n15363 ;
  assign n15350 = n15333 ^ n1799 ;
  assign n15351 = ~n15338 & ~n15350 ;
  assign n15366 = n15365 ^ n15351 ;
  assign n15347 = n15327 ^ n11569 ;
  assign n15348 = n15330 ^ n15327 ;
  assign n15349 = n15347 & n15348 ;
  assign n15367 = n15366 ^ n15349 ;
  assign n15371 = n15367 ^ n15339 ;
  assign n15370 = n15369 ^ n15367 ;
  assign n15372 = n15371 ^ n15370 ;
  assign n15373 = ~n15346 & n15372 ;
  assign n15374 = n15373 ^ n15371 ;
  assign n15449 = n15377 ^ n15374 ;
  assign n15467 = n15466 ^ n15449 ;
  assign n15468 = n15466 ^ n12788 ;
  assign n15469 = ~n15467 & n15468 ;
  assign n15470 = n15469 ^ n12788 ;
  assign n14962 = n14844 ^ n14793 ;
  assign n15378 = n15377 ^ n14962 ;
  assign n15375 = n15367 ^ n14962 ;
  assign n15379 = n15378 ^ n15375 ;
  assign n15380 = ~n15374 & n15379 ;
  assign n15381 = n15380 ^ n15375 ;
  assign n14964 = n13736 ^ n12917 ;
  assign n14965 = n14964 ^ n14358 ;
  assign n15447 = n15381 ^ n14965 ;
  assign n15448 = n15447 ^ n12886 ;
  assign n15544 = n15470 ^ n15448 ;
  assign n15533 = n15449 ^ n12788 ;
  assign n15534 = n15533 ^ n15466 ;
  assign n15542 = n15540 & n15541 ;
  assign n15543 = ~n15534 & n15542 ;
  assign n15605 = n15544 ^ n15543 ;
  assign n15626 = n15605 ^ n2325 ;
  assign n15624 = n15542 ^ n15534 ;
  assign n15625 = n15624 ^ n15605 ;
  assign n15627 = n15626 ^ n15625 ;
  assign n15628 = n15623 & ~n15627 ;
  assign n15629 = n15628 ^ n15626 ;
  assign n15689 = n15629 ^ n2135 ;
  assign n16277 = n16276 ^ n15689 ;
  assign n15744 = n14572 ^ n13988 ;
  assign n15745 = n15744 ^ n15295 ;
  assign n15717 = n15184 ^ n912 ;
  assign n15715 = n14468 ^ n13836 ;
  assign n15716 = n15715 ^ n15247 ;
  assign n15718 = n15717 ^ n15716 ;
  assign n15724 = n15180 ^ n785 ;
  assign n15722 = n14465 ^ n13837 ;
  assign n15723 = n15722 ^ n15228 ;
  assign n15725 = n15724 ^ n15723 ;
  assign n15420 = n14389 ^ n13822 ;
  assign n15421 = n15420 ^ n15099 ;
  assign n15419 = n15175 ^ n708 ;
  assign n15422 = n15421 ^ n15419 ;
  assign n14898 = n14897 ^ n14880 ;
  assign n13727 = n13726 ^ n13725 ;
  assign n14352 = n14351 ^ n13727 ;
  assign n14899 = n14898 ^ n14352 ;
  assign n14902 = n14447 ^ n13770 ;
  assign n14904 = n14903 ^ n14902 ;
  assign n14900 = n14878 ^ n1529 ;
  assign n14905 = n14904 ^ n14900 ;
  assign n14909 = n14875 ^ n14816 ;
  assign n14906 = n14402 ^ n13776 ;
  assign n14908 = n14907 ^ n14906 ;
  assign n14910 = n14909 ^ n14908 ;
  assign n14912 = n14408 ^ n13794 ;
  assign n14915 = n14914 ^ n14912 ;
  assign n14911 = n14873 ^ n518 ;
  assign n14916 = n14915 ^ n14911 ;
  assign n14920 = n14869 ^ n14822 ;
  assign n14918 = n14917 ^ n13785 ;
  assign n14919 = n14918 ^ n14416 ;
  assign n14921 = n14920 ^ n14919 ;
  assign n14927 = n14867 ^ n569 ;
  assign n14924 = n14418 ^ n13616 ;
  assign n14926 = n14925 ^ n14924 ;
  assign n14928 = n14927 ^ n14926 ;
  assign n15402 = n14932 ^ n14927 ;
  assign n14929 = n14426 ^ n13594 ;
  assign n14931 = n14930 ^ n14929 ;
  assign n14933 = n14932 ^ n14931 ;
  assign n14937 = n14861 ^ n14831 ;
  assign n14934 = n14333 ^ n13454 ;
  assign n14936 = n14935 ^ n14934 ;
  assign n14938 = n14937 ^ n14936 ;
  assign n14941 = n14190 ^ n12897 ;
  assign n14943 = n14942 ^ n14941 ;
  assign n14939 = n14858 ^ n14833 ;
  assign n14944 = n14943 ^ n14939 ;
  assign n14946 = n14176 ^ n13447 ;
  assign n14948 = n14947 ^ n14946 ;
  assign n14945 = n14855 ^ n14835 ;
  assign n14949 = n14948 ^ n14945 ;
  assign n14952 = n14853 ^ n2102 ;
  assign n15391 = n14952 ^ n14945 ;
  assign n14950 = n14097 ^ n13440 ;
  assign n14951 = n14950 ^ n14891 ;
  assign n14953 = n14952 ^ n14951 ;
  assign n14955 = n14084 ^ n12900 ;
  assign n14956 = n14955 ^ n14718 ;
  assign n15388 = n14956 ^ n14952 ;
  assign n14954 = n14850 ^ n14839 ;
  assign n14957 = n14956 ^ n14954 ;
  assign n14959 = n13728 ^ n12907 ;
  assign n14960 = n14959 ^ n14356 ;
  assign n15385 = n14960 ^ n14954 ;
  assign n14958 = n14847 ^ n14846 ;
  assign n14961 = n14960 ^ n14958 ;
  assign n14966 = n14965 ^ n14962 ;
  assign n15382 = ~n14966 & n15381 ;
  assign n14963 = n14962 ^ n14958 ;
  assign n15383 = n15382 ^ n14963 ;
  assign n15384 = n14961 & n15383 ;
  assign n15386 = n15385 ^ n15384 ;
  assign n15387 = ~n14957 & ~n15386 ;
  assign n15389 = n15388 ^ n15387 ;
  assign n15390 = n14953 & ~n15389 ;
  assign n15392 = n15391 ^ n15390 ;
  assign n15393 = ~n14949 & ~n15392 ;
  assign n15394 = n15393 ^ n14948 ;
  assign n15395 = n15394 ^ n14939 ;
  assign n15396 = ~n14944 & n15395 ;
  assign n14940 = n14939 ^ n14937 ;
  assign n15397 = n15396 ^ n14940 ;
  assign n15398 = n14938 & ~n15397 ;
  assign n15399 = n15398 ^ n14937 ;
  assign n15400 = n15399 ^ n14931 ;
  assign n15401 = ~n14933 & ~n15400 ;
  assign n15403 = n15402 ^ n15401 ;
  assign n15404 = ~n14928 & ~n15403 ;
  assign n15405 = n15404 ^ n14927 ;
  assign n14922 = n14920 ^ n14911 ;
  assign n14923 = n14922 ^ n14911 ;
  assign n15406 = n15405 ^ n14923 ;
  assign n15407 = n14921 & n15406 ;
  assign n15408 = n15407 ^ n14922 ;
  assign n15409 = ~n14916 & n15408 ;
  assign n15410 = n15409 ^ n14915 ;
  assign n15411 = n15410 ^ n14908 ;
  assign n15412 = ~n14910 & ~n15411 ;
  assign n15413 = n15412 ^ n14909 ;
  assign n15414 = n15413 ^ n14900 ;
  assign n15415 = n14905 & n15414 ;
  assign n14901 = n14900 ^ n14898 ;
  assign n15416 = n15415 ^ n14901 ;
  assign n15417 = n14899 & ~n15416 ;
  assign n15418 = n15417 ^ n14898 ;
  assign n15523 = n15419 ^ n15418 ;
  assign n15524 = ~n15422 & n15523 ;
  assign n15520 = n14383 ^ n13830 ;
  assign n15521 = n15520 ^ n15144 ;
  assign n15522 = n15521 ^ n15419 ;
  assign n15525 = n15524 ^ n15522 ;
  assign n15526 = n15177 ^ n15166 ;
  assign n15726 = n15526 ^ n15521 ;
  assign n15727 = n15525 & ~n15726 ;
  assign n15728 = n15727 ^ n15526 ;
  assign n15729 = n15728 ^ n15723 ;
  assign n15730 = ~n15725 & ~n15729 ;
  assign n15731 = n15730 ^ n15724 ;
  assign n15719 = n15189 ^ n15186 ;
  assign n15720 = n15719 ^ n15717 ;
  assign n15721 = n15720 ^ n15719 ;
  assign n15732 = n15731 ^ n15721 ;
  assign n15733 = ~n15718 & ~n15732 ;
  assign n15734 = n15733 ^ n15720 ;
  assign n15737 = n15162 ^ n1061 ;
  assign n15738 = n15737 ^ n15191 ;
  assign n15740 = n15738 ^ n15719 ;
  assign n15735 = n14472 ^ n13847 ;
  assign n15736 = n15735 ^ n15278 ;
  assign n15739 = n15738 ^ n15736 ;
  assign n15741 = n15740 ^ n15739 ;
  assign n15742 = n15734 & n15741 ;
  assign n15743 = n15742 ^ n15740 ;
  assign n15786 = n15745 ^ n15743 ;
  assign n15787 = n15786 ^ n13374 ;
  assign n15788 = n15736 ^ n15734 ;
  assign n15789 = n15788 ^ n13343 ;
  assign n15798 = n15731 ^ n15718 ;
  assign n15790 = n15728 ^ n15725 ;
  assign n15791 = n15790 ^ n13171 ;
  assign n15527 = n15526 ^ n15525 ;
  assign n15528 = n15527 ^ n13083 ;
  assign n15423 = n15422 ^ n15418 ;
  assign n15424 = n15423 ^ n13076 ;
  assign n15425 = n15416 ^ n14352 ;
  assign n15426 = n15425 ^ n12960 ;
  assign n15427 = n15413 ^ n14905 ;
  assign n15428 = n15427 ^ n12971 ;
  assign n15429 = n15410 ^ n14910 ;
  assign n15430 = n15429 ^ n12976 ;
  assign n15503 = n15408 ^ n14915 ;
  assign n15431 = n15405 ^ n14921 ;
  assign n15432 = n15431 ^ n13046 ;
  assign n15495 = n15403 ^ n14926 ;
  assign n15433 = n15399 ^ n14933 ;
  assign n15434 = n15433 ^ n12899 ;
  assign n15435 = n15397 ^ n14936 ;
  assign n15436 = n15435 ^ n12906 ;
  assign n15437 = n15394 ^ n14944 ;
  assign n15438 = n15437 ^ n12913 ;
  assign n15439 = n15392 ^ n14948 ;
  assign n15440 = n15439 ^ n12920 ;
  assign n15441 = n15389 ^ n14951 ;
  assign n15442 = n15441 ^ n12928 ;
  assign n15443 = n15386 ^ n14956 ;
  assign n15444 = n15443 ^ n12940 ;
  assign n15445 = n15383 ^ n14960 ;
  assign n15446 = n15445 ^ n12936 ;
  assign n15471 = n15470 ^ n15447 ;
  assign n15472 = ~n15448 & ~n15471 ;
  assign n15473 = n15472 ^ n12886 ;
  assign n15474 = n15473 ^ n15445 ;
  assign n15475 = ~n15446 & ~n15474 ;
  assign n15476 = n15475 ^ n12936 ;
  assign n15477 = n15476 ^ n15443 ;
  assign n15478 = ~n15444 & n15477 ;
  assign n15479 = n15478 ^ n12940 ;
  assign n15480 = n15479 ^ n15441 ;
  assign n15481 = ~n15442 & n15480 ;
  assign n15482 = n15481 ^ n12928 ;
  assign n15483 = n15482 ^ n15439 ;
  assign n15484 = ~n15440 & n15483 ;
  assign n15485 = n15484 ^ n12920 ;
  assign n15486 = n15485 ^ n15437 ;
  assign n15487 = ~n15438 & ~n15486 ;
  assign n15488 = n15487 ^ n12913 ;
  assign n15489 = n15488 ^ n15435 ;
  assign n15490 = ~n15436 & ~n15489 ;
  assign n15491 = n15490 ^ n12906 ;
  assign n15492 = n15491 ^ n15433 ;
  assign n15493 = n15434 & n15492 ;
  assign n15494 = n15493 ^ n12899 ;
  assign n15496 = n15495 ^ n15494 ;
  assign n15497 = n15495 ^ n12982 ;
  assign n15498 = n15496 & ~n15497 ;
  assign n15499 = n15498 ^ n12982 ;
  assign n15500 = n15499 ^ n15431 ;
  assign n15501 = n15432 & n15500 ;
  assign n15502 = n15501 ^ n13046 ;
  assign n15504 = n15503 ^ n15502 ;
  assign n15505 = n15503 ^ n12343 ;
  assign n15506 = n15504 & n15505 ;
  assign n15507 = n15506 ^ n12343 ;
  assign n15508 = n15507 ^ n15429 ;
  assign n15509 = ~n15430 & ~n15508 ;
  assign n15510 = n15509 ^ n12976 ;
  assign n15511 = n15510 ^ n15427 ;
  assign n15512 = ~n15428 & n15511 ;
  assign n15513 = n15512 ^ n12971 ;
  assign n15514 = n15513 ^ n15425 ;
  assign n15515 = ~n15426 & n15514 ;
  assign n15516 = n15515 ^ n12960 ;
  assign n15517 = n15516 ^ n15423 ;
  assign n15518 = n15424 & n15517 ;
  assign n15519 = n15518 ^ n13076 ;
  assign n15792 = n15527 ^ n15519 ;
  assign n15793 = n15528 & ~n15792 ;
  assign n15794 = n15793 ^ n13083 ;
  assign n15795 = n15794 ^ n15790 ;
  assign n15796 = n15791 & ~n15795 ;
  assign n15797 = n15796 ^ n13171 ;
  assign n15799 = n15798 ^ n15797 ;
  assign n15800 = n15798 ^ n13295 ;
  assign n15801 = n15799 & n15800 ;
  assign n15802 = n15801 ^ n13295 ;
  assign n15803 = n15802 ^ n15788 ;
  assign n15804 = ~n15789 & ~n15803 ;
  assign n15805 = n15804 ^ n13343 ;
  assign n15806 = n15805 ^ n15786 ;
  assign n15807 = n15787 & ~n15806 ;
  assign n15808 = n15807 ^ n13374 ;
  assign n15753 = n14025 ^ n13316 ;
  assign n15754 = n15753 ^ n15318 ;
  assign n15676 = n15197 ^ n1305 ;
  assign n15747 = n15738 ^ n15676 ;
  assign n15746 = n15745 ^ n15676 ;
  assign n15748 = n15747 ^ n15746 ;
  assign n15749 = n15743 & ~n15748 ;
  assign n15750 = n15749 ^ n15747 ;
  assign n15784 = n15754 ^ n15750 ;
  assign n15785 = n15784 ^ n12631 ;
  assign n15857 = n15808 ^ n15785 ;
  assign n15848 = n15800 ^ n15797 ;
  assign n15529 = n15528 ^ n15519 ;
  assign n15530 = n15516 ^ n15424 ;
  assign n15531 = n15510 ^ n15428 ;
  assign n15532 = n15491 ^ n15434 ;
  assign n15545 = ~n15543 & ~n15544 ;
  assign n15546 = n15473 ^ n15446 ;
  assign n15547 = ~n15545 & ~n15546 ;
  assign n15548 = n15476 ^ n15444 ;
  assign n15549 = ~n15547 & ~n15548 ;
  assign n15550 = n15479 ^ n15442 ;
  assign n15551 = n15549 & ~n15550 ;
  assign n15552 = n15482 ^ n15440 ;
  assign n15553 = n15551 & ~n15552 ;
  assign n15554 = n15485 ^ n15438 ;
  assign n15555 = ~n15553 & n15554 ;
  assign n15556 = n15488 ^ n15436 ;
  assign n15557 = ~n15555 & n15556 ;
  assign n15558 = ~n15532 & ~n15557 ;
  assign n15559 = n15497 ^ n15494 ;
  assign n15560 = ~n15558 & n15559 ;
  assign n15561 = n15499 ^ n15432 ;
  assign n15562 = n15560 & ~n15561 ;
  assign n15563 = n15505 ^ n15502 ;
  assign n15564 = n15562 & n15563 ;
  assign n15565 = n15507 ^ n15430 ;
  assign n15566 = n15564 & n15565 ;
  assign n15567 = n15531 & ~n15566 ;
  assign n15568 = n15513 ^ n15426 ;
  assign n15569 = n15567 & n15568 ;
  assign n15570 = n15530 & ~n15569 ;
  assign n15849 = ~n15529 & n15570 ;
  assign n15850 = n15794 ^ n15791 ;
  assign n15851 = ~n15849 & n15850 ;
  assign n15852 = ~n15848 & ~n15851 ;
  assign n15853 = n15802 ^ n15789 ;
  assign n15854 = n15852 & ~n15853 ;
  assign n15855 = n15805 ^ n15787 ;
  assign n15856 = ~n15854 & n15855 ;
  assign n15886 = n15857 ^ n15856 ;
  assign n3113 = n3109 ^ x199 ;
  assign n3114 = n3113 ^ x391 ;
  assign n3115 = n3114 ^ x135 ;
  assign n15887 = n15886 ^ n3115 ;
  assign n15891 = n15855 ^ n15854 ;
  assign n15892 = n15891 ^ n2893 ;
  assign n15893 = n15853 ^ n15852 ;
  assign n15894 = n15893 ^ n2504 ;
  assign n15896 = n15850 ^ n15849 ;
  assign n15897 = n15896 ^ n1343 ;
  assign n15573 = n15569 ^ n15530 ;
  assign n15574 = n15573 ^ n1002 ;
  assign n15671 = n15573 ^ n990 ;
  assign n15575 = n15568 ^ n15567 ;
  assign n15576 = n15575 ^ n990 ;
  assign n15577 = n15566 ^ n15531 ;
  assign n15578 = n15577 ^ n883 ;
  assign n15579 = n15563 ^ n15562 ;
  assign n15580 = n15579 ^ n865 ;
  assign n15581 = n15561 ^ n15560 ;
  assign n15582 = n15581 ^ n641 ;
  assign n15584 = n15557 ^ n15532 ;
  assign n15585 = n15584 ^ n531 ;
  assign n15586 = n15556 ^ n15555 ;
  assign n15587 = n15586 ^ n548 ;
  assign n15588 = n15554 ^ n15553 ;
  assign n15589 = n15588 ^ n563 ;
  assign n15590 = n15552 ^ n15551 ;
  assign n15594 = n15593 ^ n15590 ;
  assign n15597 = n15550 ^ n15549 ;
  assign n15598 = n15597 ^ n1454 ;
  assign n15599 = n15548 ^ n15547 ;
  assign n15600 = n15599 ^ n2353 ;
  assign n15603 = n15546 ^ n15545 ;
  assign n15604 = n15603 ^ n2339 ;
  assign n15606 = n15605 ^ n2135 ;
  assign n15630 = ~n15606 & n15629 ;
  assign n15631 = n15630 ^ n2135 ;
  assign n15632 = n15631 ^ n15603 ;
  assign n15633 = n15604 & ~n15632 ;
  assign n15634 = n15633 ^ n2339 ;
  assign n15601 = n15597 ^ n2353 ;
  assign n15602 = n15601 ^ n15597 ;
  assign n15635 = n15634 ^ n15602 ;
  assign n15636 = ~n15600 & n15635 ;
  assign n15637 = n15636 ^ n15601 ;
  assign n15638 = n15598 & ~n15637 ;
  assign n15639 = n15638 ^ n1454 ;
  assign n15640 = n15639 ^ n15593 ;
  assign n15641 = n15594 & n15640 ;
  assign n15595 = n15593 ^ n15588 ;
  assign n15642 = n15641 ^ n15595 ;
  assign n15643 = ~n15589 & n15642 ;
  assign n15644 = n15643 ^ n563 ;
  assign n15645 = n15644 ^ n15586 ;
  assign n15646 = n15587 & ~n15645 ;
  assign n15647 = n15646 ^ n548 ;
  assign n15648 = n15647 ^ n15584 ;
  assign n15649 = n15585 & ~n15648 ;
  assign n15650 = n15649 ^ n531 ;
  assign n15654 = n15650 ^ n15581 ;
  assign n15583 = n15559 ^ n15558 ;
  assign n15651 = n15650 ^ n15583 ;
  assign n15652 = n15583 ^ n1581 ;
  assign n15653 = n15651 & ~n15652 ;
  assign n15655 = n15654 ^ n15653 ;
  assign n15656 = n15582 & ~n15655 ;
  assign n15657 = n15656 ^ n641 ;
  assign n15658 = n15657 ^ n865 ;
  assign n15659 = ~n15580 & ~n15658 ;
  assign n15660 = n15659 ^ n15579 ;
  assign n15661 = n15660 ^ n871 ;
  assign n15662 = n15565 ^ n15564 ;
  assign n15663 = n15662 ^ n871 ;
  assign n15664 = ~n15661 & ~n15663 ;
  assign n15665 = n15664 ^ n871 ;
  assign n15666 = n15665 ^ n883 ;
  assign n15667 = ~n15578 & ~n15666 ;
  assign n15668 = n15667 ^ n15577 ;
  assign n15669 = n15668 ^ n990 ;
  assign n15670 = n15576 & ~n15669 ;
  assign n15672 = n15671 ^ n15670 ;
  assign n15673 = n15574 & ~n15672 ;
  assign n15674 = n15673 ^ n1002 ;
  assign n15571 = n15570 ^ n15529 ;
  assign n15898 = n15674 ^ n15571 ;
  assign n15899 = n15896 ^ n1140 ;
  assign n15900 = n15899 ^ n15896 ;
  assign n15901 = n15900 ^ n15571 ;
  assign n15902 = ~n15898 & n15901 ;
  assign n15903 = n15902 ^ n15899 ;
  assign n15904 = ~n15897 & n15903 ;
  assign n15905 = n15904 ^ n1343 ;
  assign n15895 = n15851 ^ n15848 ;
  assign n15906 = n15905 ^ n15895 ;
  assign n15907 = n15893 ^ n1376 ;
  assign n15908 = n15907 ^ n15893 ;
  assign n15909 = n15908 ^ n15895 ;
  assign n15910 = n15906 & ~n15909 ;
  assign n15911 = n15910 ^ n15907 ;
  assign n15912 = n15894 & ~n15911 ;
  assign n15913 = n15912 ^ n2504 ;
  assign n15914 = n15913 ^ n15891 ;
  assign n15915 = ~n15892 & n15914 ;
  assign n15916 = n15915 ^ n2893 ;
  assign n15809 = n15808 ^ n15784 ;
  assign n15810 = ~n15785 & ~n15809 ;
  assign n15811 = n15810 ^ n12631 ;
  assign n15760 = n14020 ^ n13315 ;
  assign n15761 = n15760 ^ n15357 ;
  assign n15751 = n15159 ^ n1256 ;
  assign n15752 = n15751 ^ n15199 ;
  assign n15756 = n15752 ^ n15676 ;
  assign n15755 = n15754 ^ n15752 ;
  assign n15757 = n15756 ^ n15755 ;
  assign n15758 = n15750 & ~n15757 ;
  assign n15759 = n15758 ^ n15756 ;
  assign n15782 = n15761 ^ n15759 ;
  assign n15783 = n15782 ^ n12627 ;
  assign n15859 = n15811 ^ n15783 ;
  assign n15858 = ~n15856 & n15857 ;
  assign n15888 = n15859 ^ n15858 ;
  assign n15889 = n15888 ^ n3115 ;
  assign n15890 = n15889 ^ n15888 ;
  assign n15917 = n15916 ^ n15890 ;
  assign n15918 = n15887 & n15917 ;
  assign n15919 = n15918 ^ n15889 ;
  assign n15812 = n15811 ^ n15782 ;
  assign n15813 = ~n15783 & ~n15812 ;
  assign n15814 = n15813 ^ n12627 ;
  assign n15768 = n14018 ^ n13312 ;
  assign n15769 = n15768 ^ n14667 ;
  assign n15762 = n15205 ^ n2796 ;
  assign n15764 = n15762 ^ n15752 ;
  assign n15763 = n15762 ^ n15761 ;
  assign n15765 = n15764 ^ n15763 ;
  assign n15766 = n15759 & n15765 ;
  assign n15767 = n15766 ^ n15764 ;
  assign n15780 = n15769 ^ n15767 ;
  assign n15781 = n15780 ^ n12621 ;
  assign n15861 = n15814 ^ n15781 ;
  assign n15860 = n15858 & ~n15859 ;
  assign n15920 = n15861 ^ n15860 ;
  assign n15922 = n15920 ^ n1832 ;
  assign n15921 = n15920 ^ n15888 ;
  assign n15923 = n15922 ^ n15921 ;
  assign n15924 = ~n15919 & n15923 ;
  assign n15925 = n15924 ^ n15922 ;
  assign n15956 = n15925 ^ n2601 ;
  assign n15954 = n14696 ^ n13749 ;
  assign n15955 = n15954 ^ n14962 ;
  assign n16017 = n15956 ^ n15955 ;
  assign n16081 = n16017 ^ n13403 ;
  assign n3049 = n3021 ^ x224 ;
  assign n3050 = n3049 ^ x416 ;
  assign n3051 = n3050 ^ x160 ;
  assign n16275 = n16081 ^ n3051 ;
  assign n16278 = n16277 ^ n16275 ;
  assign n3035 = x417 ^ x225 ;
  assign n3036 = n3035 ^ n3009 ;
  assign n3037 = n3036 ^ x161 ;
  assign n16541 = n3037 ^ n1781 ;
  assign n16428 = n14377 ^ n13760 ;
  assign n16429 = n16428 ^ n15339 ;
  assign n16281 = n14667 ^ n14025 ;
  assign n15835 = n15152 ^ n2569 ;
  assign n15836 = n15835 ^ n15213 ;
  assign n16282 = n16281 ^ n15836 ;
  assign n15572 = n15571 ^ n1140 ;
  assign n15675 = n15674 ^ n15572 ;
  assign n16283 = n16282 ^ n15675 ;
  assign n16288 = n15357 ^ n14572 ;
  assign n15821 = n15210 ^ n15154 ;
  assign n16289 = n16288 ^ n15821 ;
  assign n16287 = n15672 ^ n1002 ;
  assign n16290 = n16289 ^ n16287 ;
  assign n16293 = n15668 ^ n15576 ;
  assign n15770 = n15207 ^ n15156 ;
  assign n16291 = n15770 ^ n14472 ;
  assign n16292 = n16291 ^ n15318 ;
  assign n16294 = n16293 ^ n16292 ;
  assign n16297 = n15295 ^ n14468 ;
  assign n16298 = n16297 ^ n15762 ;
  assign n16295 = n15665 ^ n15578 ;
  assign n16299 = n16298 ^ n16295 ;
  assign n16301 = n15278 ^ n14465 ;
  assign n16302 = n16301 ^ n15752 ;
  assign n16300 = n15663 ^ n15660 ;
  assign n16303 = n16302 ^ n16300 ;
  assign n16305 = n15247 ^ n14383 ;
  assign n16306 = n16305 ^ n15676 ;
  assign n16304 = n15657 ^ n15580 ;
  assign n16307 = n16306 ^ n16304 ;
  assign n16310 = n15655 ^ n641 ;
  assign n16308 = n15228 ^ n14389 ;
  assign n16309 = n16308 ^ n15738 ;
  assign n16311 = n16310 ^ n16309 ;
  assign n16246 = n15652 ^ n15650 ;
  assign n16231 = n15647 ^ n15585 ;
  assign n16247 = n16246 ^ n16231 ;
  assign n16229 = n15099 ^ n14447 ;
  assign n16230 = n16229 ^ n15717 ;
  assign n16232 = n16231 ^ n16230 ;
  assign n16127 = n14402 ^ n14351 ;
  assign n16128 = n16127 ^ n15724 ;
  assign n16126 = n15644 ^ n15587 ;
  assign n16129 = n16128 ^ n16126 ;
  assign n16070 = n15639 ^ n15594 ;
  assign n16068 = n14907 ^ n14416 ;
  assign n16069 = n16068 ^ n15419 ;
  assign n16071 = n16070 ^ n16069 ;
  assign n16111 = n15642 ^ n563 ;
  assign n15679 = n14917 ^ n14426 ;
  assign n15680 = n15679 ^ n14900 ;
  assign n15678 = n15634 ^ n15600 ;
  assign n15681 = n15680 ^ n15678 ;
  assign n15685 = n15631 ^ n15604 ;
  assign n15683 = n14925 ^ n14333 ;
  assign n15684 = n15683 ^ n14909 ;
  assign n15686 = n15685 ^ n15684 ;
  assign n15687 = n14930 ^ n14190 ;
  assign n15688 = n15687 ^ n14911 ;
  assign n15690 = n15689 ^ n15688 ;
  assign n15694 = n14935 ^ n14176 ;
  assign n15695 = n15694 ^ n14920 ;
  assign n15693 = n15624 ^ n15623 ;
  assign n15696 = n15695 ^ n15693 ;
  assign n15699 = n15620 ^ n15618 ;
  assign n15985 = n15699 ^ n15693 ;
  assign n15697 = n14942 ^ n14097 ;
  assign n15698 = n15697 ^ n14927 ;
  assign n15700 = n15699 ^ n15698 ;
  assign n15702 = n14947 ^ n14084 ;
  assign n15703 = n15702 ^ n14932 ;
  assign n15701 = n15615 ^ n15609 ;
  assign n15704 = n15703 ^ n15701 ;
  assign n15707 = n15613 ^ n15610 ;
  assign n15979 = n15707 ^ n15701 ;
  assign n15705 = n14891 ^ n13728 ;
  assign n15706 = n15705 ^ n14937 ;
  assign n15708 = n15707 ^ n15706 ;
  assign n15711 = n15536 ^ n1889 ;
  assign n15709 = n14718 ^ n13736 ;
  assign n15710 = n15709 ^ n14939 ;
  assign n15712 = n15711 ^ n15710 ;
  assign n15827 = n14004 ^ n13384 ;
  assign n15828 = n15827 ^ n14662 ;
  assign n15772 = n15770 ^ n15762 ;
  assign n15771 = n15770 ^ n15769 ;
  assign n15773 = n15772 ^ n15771 ;
  assign n15774 = ~n15767 & ~n15773 ;
  assign n15775 = n15774 ^ n15772 ;
  assign n15823 = n15821 ^ n15770 ;
  assign n15776 = n14009 ^ n13355 ;
  assign n15777 = n15776 ^ n14669 ;
  assign n15822 = n15821 ^ n15777 ;
  assign n15824 = n15823 ^ n15822 ;
  assign n15825 = ~n15775 & n15824 ;
  assign n15826 = n15825 ^ n15823 ;
  assign n15829 = n15828 ^ n15826 ;
  assign n15846 = n15829 ^ n12697 ;
  assign n15778 = n15777 ^ n15775 ;
  assign n15779 = n15778 ^ n12669 ;
  assign n15815 = n15814 ^ n15780 ;
  assign n15816 = n15781 & ~n15815 ;
  assign n15817 = n15816 ^ n12621 ;
  assign n15818 = n15817 ^ n15778 ;
  assign n15819 = n15779 & ~n15818 ;
  assign n15820 = n15819 ^ n12669 ;
  assign n15847 = n15846 ^ n15820 ;
  assign n15862 = n15860 & ~n15861 ;
  assign n15863 = n15817 ^ n15779 ;
  assign n15864 = ~n15862 & n15863 ;
  assign n15865 = ~n15847 & ~n15864 ;
  assign n15842 = n13760 ^ n12950 ;
  assign n15843 = n15842 ^ n14682 ;
  assign n15838 = n15836 ^ n15821 ;
  assign n15837 = n15836 ^ n15828 ;
  assign n15839 = n15838 ^ n15837 ;
  assign n15840 = n15826 & ~n15839 ;
  assign n15841 = n15840 ^ n15838 ;
  assign n15844 = n15843 ^ n15841 ;
  assign n15830 = n15829 ^ n15820 ;
  assign n15831 = n15820 ^ n12697 ;
  assign n15832 = n15830 & ~n15831 ;
  assign n15833 = n15832 ^ n15829 ;
  assign n15834 = n15833 ^ n12702 ;
  assign n15845 = n15844 ^ n15834 ;
  assign n15884 = n15865 ^ n15845 ;
  assign n15885 = n15884 ^ n2998 ;
  assign n15926 = n15863 ^ n15862 ;
  assign n15928 = n15926 ^ n2601 ;
  assign n15927 = n15926 ^ n15920 ;
  assign n15929 = n15928 ^ n15927 ;
  assign n15930 = ~n15925 & n15929 ;
  assign n15931 = n15930 ^ n15928 ;
  assign n15932 = n15864 ^ n15847 ;
  assign n15934 = n15932 ^ n15926 ;
  assign n15933 = n15932 ^ n2615 ;
  assign n15935 = n15934 ^ n15933 ;
  assign n15936 = n15931 & ~n15935 ;
  assign n15937 = n15936 ^ n15933 ;
  assign n15939 = n2998 ^ n2688 ;
  assign n15938 = n15932 ^ n2998 ;
  assign n15940 = n15939 ^ n15938 ;
  assign n15941 = n15937 & ~n15940 ;
  assign n15942 = n15941 ^ n15939 ;
  assign n15943 = n15885 & n15942 ;
  assign n15880 = n15843 ^ n15836 ;
  assign n15881 = ~n15841 & n15880 ;
  assign n15877 = n2998 ^ n1883 ;
  assign n15875 = n12702 ^ n12358 ;
  assign n15871 = n13755 ^ n13389 ;
  assign n15872 = n15871 ^ n14651 ;
  assign n15873 = n15872 ^ n15843 ;
  assign n15870 = n15237 ^ n2490 ;
  assign n15874 = n15873 ^ n15870 ;
  assign n15876 = n15875 ^ n15874 ;
  assign n15878 = n15877 ^ n15876 ;
  assign n15867 = n15844 ^ n12702 ;
  assign n15868 = n15844 ^ n15833 ;
  assign n15869 = n15867 & n15868 ;
  assign n15879 = n15878 ^ n15869 ;
  assign n15882 = n15881 ^ n15879 ;
  assign n15866 = ~n15845 & n15865 ;
  assign n15883 = n15882 ^ n15866 ;
  assign n15944 = n15943 ^ n15883 ;
  assign n15973 = n15944 ^ n15711 ;
  assign n15713 = n14356 ^ n13738 ;
  assign n15714 = n15713 ^ n14945 ;
  assign n15945 = n15944 ^ n15714 ;
  assign n15948 = n15942 ^ n15884 ;
  assign n15946 = n14358 ^ n13744 ;
  assign n15947 = n15946 ^ n14952 ;
  assign n15949 = n15948 ^ n15947 ;
  assign n15952 = n15937 ^ n2688 ;
  assign n15967 = n15952 ^ n15948 ;
  assign n15950 = n14954 ^ n14067 ;
  assign n15951 = n15950 ^ n14364 ;
  assign n15953 = n15952 ^ n15951 ;
  assign n15958 = n14700 ^ n14061 ;
  assign n15959 = n15958 ^ n14958 ;
  assign n15964 = n15959 ^ n15952 ;
  assign n15957 = ~n15955 & n15956 ;
  assign n15960 = n15959 ^ n15957 ;
  assign n15961 = n15931 ^ n2615 ;
  assign n15962 = n15961 ^ n15959 ;
  assign n15963 = ~n15960 & n15962 ;
  assign n15965 = n15964 ^ n15963 ;
  assign n15966 = n15953 & n15965 ;
  assign n15968 = n15967 ^ n15966 ;
  assign n15969 = ~n15949 & ~n15968 ;
  assign n15970 = n15969 ^ n15948 ;
  assign n15971 = n15970 ^ n15714 ;
  assign n15972 = n15945 & ~n15971 ;
  assign n15974 = n15973 ^ n15972 ;
  assign n15975 = n15712 & ~n15974 ;
  assign n15976 = n15975 ^ n15711 ;
  assign n15977 = n15976 ^ n15706 ;
  assign n15978 = n15708 & ~n15977 ;
  assign n15980 = n15979 ^ n15978 ;
  assign n15981 = n15704 & ~n15980 ;
  assign n15982 = n15981 ^ n15703 ;
  assign n15983 = n15982 ^ n15699 ;
  assign n15984 = n15700 & ~n15983 ;
  assign n15986 = n15985 ^ n15984 ;
  assign n15987 = n15696 & n15986 ;
  assign n15988 = n15987 ^ n15695 ;
  assign n15989 = n15988 ^ n15689 ;
  assign n15990 = ~n15690 & n15989 ;
  assign n15691 = n15689 ^ n15685 ;
  assign n15991 = n15990 ^ n15691 ;
  assign n15992 = ~n15686 & ~n15991 ;
  assign n15993 = n15992 ^ n15685 ;
  assign n15682 = n15637 ^ n1454 ;
  assign n15994 = n15993 ^ n15682 ;
  assign n15995 = n15994 ^ n15678 ;
  assign n15996 = n15995 ^ n15682 ;
  assign n15997 = n15681 & ~n15996 ;
  assign n15998 = n15997 ^ n15994 ;
  assign n15999 = n14914 ^ n14418 ;
  assign n16000 = n15999 ^ n14898 ;
  assign n16072 = n16000 ^ n15682 ;
  assign n16073 = n15998 & ~n16072 ;
  assign n16074 = n16073 ^ n15682 ;
  assign n16112 = n16111 ^ n16074 ;
  assign n16113 = n16112 ^ n16069 ;
  assign n16114 = n16113 ^ n16111 ;
  assign n16115 = ~n16071 & n16114 ;
  assign n16116 = n16115 ^ n16112 ;
  assign n16117 = n14903 ^ n14408 ;
  assign n16118 = n16117 ^ n15526 ;
  assign n16123 = n16118 ^ n16111 ;
  assign n16124 = n16116 & n16123 ;
  assign n16125 = n16124 ^ n16118 ;
  assign n16226 = n16126 ^ n16125 ;
  assign n16227 = n16129 & ~n16226 ;
  assign n16228 = n16227 ^ n16126 ;
  assign n16244 = n16230 ^ n16228 ;
  assign n16245 = n16232 & ~n16244 ;
  assign n16248 = n16247 ^ n16245 ;
  assign n16249 = n15144 ^ n13725 ;
  assign n16250 = n16249 ^ n15719 ;
  assign n16314 = n16250 ^ n16246 ;
  assign n16315 = n16248 & ~n16314 ;
  assign n16316 = n16315 ^ n16246 ;
  assign n16317 = n16316 ^ n16310 ;
  assign n16318 = ~n16311 & n16317 ;
  assign n16312 = n16310 ^ n16304 ;
  assign n16319 = n16318 ^ n16312 ;
  assign n16320 = n16307 & n16319 ;
  assign n16321 = n16320 ^ n16306 ;
  assign n16322 = n16321 ^ n16300 ;
  assign n16323 = n16303 & n16322 ;
  assign n16324 = n16323 ^ n16302 ;
  assign n16325 = n16324 ^ n16295 ;
  assign n16326 = ~n16299 & ~n16325 ;
  assign n16296 = n16295 ^ n16293 ;
  assign n16327 = n16326 ^ n16296 ;
  assign n16328 = n16294 & n16327 ;
  assign n16329 = n16328 ^ n16293 ;
  assign n16330 = n16329 ^ n16287 ;
  assign n16331 = ~n16290 & n16330 ;
  assign n16332 = n16331 ^ n16289 ;
  assign n16284 = n15903 ^ n1343 ;
  assign n16285 = n16284 ^ n15675 ;
  assign n16286 = n16285 ^ n16284 ;
  assign n16333 = n16332 ^ n16286 ;
  assign n16334 = ~n16283 & ~n16333 ;
  assign n16335 = n16334 ^ n16285 ;
  assign n16338 = n15895 ^ n1376 ;
  assign n16339 = n16338 ^ n15905 ;
  assign n16341 = n16339 ^ n16284 ;
  assign n16336 = n14669 ^ n14020 ;
  assign n16337 = n16336 ^ n15870 ;
  assign n16340 = n16339 ^ n16337 ;
  assign n16342 = n16341 ^ n16340 ;
  assign n16343 = ~n16335 & ~n16342 ;
  assign n16344 = n16343 ^ n16341 ;
  assign n16347 = n15911 ^ n2504 ;
  assign n16349 = n16347 ^ n16339 ;
  assign n16345 = n14662 ^ n14018 ;
  assign n16346 = n16345 ^ n15260 ;
  assign n16348 = n16347 ^ n16346 ;
  assign n16350 = n16349 ^ n16348 ;
  assign n16351 = n16344 & n16350 ;
  assign n16352 = n16351 ^ n16349 ;
  assign n16353 = n15913 ^ n15892 ;
  assign n16357 = n16353 ^ n16347 ;
  assign n16354 = n14682 ^ n14009 ;
  assign n16355 = n16354 ^ n15312 ;
  assign n16356 = n16355 ^ n16353 ;
  assign n16358 = n16357 ^ n16356 ;
  assign n16359 = ~n16352 & n16358 ;
  assign n16360 = n16359 ^ n16357 ;
  assign n16422 = n15916 ^ n15887 ;
  assign n16424 = n16422 ^ n16353 ;
  assign n16361 = n14651 ^ n14004 ;
  assign n16362 = n16361 ^ n15309 ;
  assign n16423 = n16422 ^ n16362 ;
  assign n16425 = n16424 ^ n16423 ;
  assign n16426 = ~n16360 & n16425 ;
  assign n16427 = n16426 ^ n16424 ;
  assign n16430 = n16429 ^ n16427 ;
  assign n16363 = n16362 ^ n16360 ;
  assign n16364 = n16363 ^ n13384 ;
  assign n16366 = n16337 ^ n16335 ;
  assign n16367 = n16366 ^ n13315 ;
  assign n16368 = n16332 ^ n16283 ;
  assign n16369 = n16368 ^ n13316 ;
  assign n16398 = n16329 ^ n16290 ;
  assign n16371 = n16324 ^ n16299 ;
  assign n16372 = n16371 ^ n13836 ;
  assign n16374 = n16319 ^ n16306 ;
  assign n16375 = n16374 ^ n13830 ;
  assign n16376 = n16316 ^ n16311 ;
  assign n16377 = n16376 ^ n13822 ;
  assign n16251 = n16250 ^ n16248 ;
  assign n16252 = n16251 ^ n13726 ;
  assign n16233 = n16232 ^ n16228 ;
  assign n16234 = n16233 ^ n13770 ;
  assign n16130 = n16129 ^ n16125 ;
  assign n16131 = n16130 ^ n13776 ;
  assign n16119 = n16118 ^ n16116 ;
  assign n16120 = n16119 ^ n13794 ;
  assign n16075 = n16074 ^ n16071 ;
  assign n16076 = n16075 ^ n13785 ;
  assign n16002 = n15993 ^ n15681 ;
  assign n16003 = n16002 ^ n13594 ;
  assign n16005 = n15988 ^ n15690 ;
  assign n16006 = n16005 ^ n12897 ;
  assign n16007 = n15986 ^ n15695 ;
  assign n16008 = n16007 ^ n13447 ;
  assign n16046 = n15982 ^ n15700 ;
  assign n16009 = n15980 ^ n15703 ;
  assign n16010 = n16009 ^ n12900 ;
  assign n16011 = n15976 ^ n15708 ;
  assign n16012 = n16011 ^ n12907 ;
  assign n16013 = n15974 ^ n15710 ;
  assign n16014 = n16013 ^ n12917 ;
  assign n16032 = n15970 ^ n15945 ;
  assign n16015 = n15968 ^ n15947 ;
  assign n16016 = n16015 ^ n12933 ;
  assign n16024 = n15965 ^ n15951 ;
  assign n16018 = n13403 & ~n16017 ;
  assign n16019 = n16018 ^ n12945 ;
  assign n16020 = n15961 ^ n15960 ;
  assign n16021 = n16020 ^ n16018 ;
  assign n16022 = n16019 & ~n16021 ;
  assign n16023 = n16022 ^ n12945 ;
  assign n16025 = n16024 ^ n16023 ;
  assign n16026 = n16024 ^ n13411 ;
  assign n16027 = n16025 & n16026 ;
  assign n16028 = n16027 ^ n13411 ;
  assign n16029 = n16028 ^ n16015 ;
  assign n16030 = ~n16016 & n16029 ;
  assign n16031 = n16030 ^ n12933 ;
  assign n16033 = n16032 ^ n16031 ;
  assign n16034 = n16032 ^ n12922 ;
  assign n16035 = n16033 & n16034 ;
  assign n16036 = n16035 ^ n12922 ;
  assign n16037 = n16036 ^ n16013 ;
  assign n16038 = ~n16014 & ~n16037 ;
  assign n16039 = n16038 ^ n12917 ;
  assign n16040 = n16039 ^ n16011 ;
  assign n16041 = ~n16012 & ~n16040 ;
  assign n16042 = n16041 ^ n12907 ;
  assign n16043 = n16042 ^ n16009 ;
  assign n16044 = ~n16010 & n16043 ;
  assign n16045 = n16044 ^ n12900 ;
  assign n16047 = n16046 ^ n16045 ;
  assign n16048 = n16046 ^ n13440 ;
  assign n16049 = n16047 & ~n16048 ;
  assign n16050 = n16049 ^ n13440 ;
  assign n16051 = n16050 ^ n16007 ;
  assign n16052 = ~n16008 & ~n16051 ;
  assign n16053 = n16052 ^ n13447 ;
  assign n16054 = n16053 ^ n16005 ;
  assign n16055 = n16006 & n16054 ;
  assign n16056 = n16055 ^ n12897 ;
  assign n16004 = n15991 ^ n15684 ;
  assign n16057 = n16056 ^ n16004 ;
  assign n16058 = n16056 ^ n13454 ;
  assign n16059 = ~n16057 & n16058 ;
  assign n16060 = n16059 ^ n13454 ;
  assign n16061 = n16060 ^ n16002 ;
  assign n16062 = ~n16003 & n16061 ;
  assign n16063 = n16062 ^ n13594 ;
  assign n16001 = n16000 ^ n15998 ;
  assign n16064 = n16063 ^ n16001 ;
  assign n16065 = n16063 ^ n13616 ;
  assign n16066 = n16064 & ~n16065 ;
  assign n16067 = n16066 ^ n13616 ;
  assign n16108 = n16075 ^ n16067 ;
  assign n16109 = n16076 & n16108 ;
  assign n16110 = n16109 ^ n13785 ;
  assign n16132 = n16119 ^ n16110 ;
  assign n16133 = ~n16120 & ~n16132 ;
  assign n16134 = n16133 ^ n13794 ;
  assign n16223 = n16134 ^ n16130 ;
  assign n16224 = n16131 & ~n16223 ;
  assign n16225 = n16224 ^ n13776 ;
  assign n16241 = n16233 ^ n16225 ;
  assign n16242 = n16234 & n16241 ;
  assign n16243 = n16242 ^ n13770 ;
  assign n16378 = n16251 ^ n16243 ;
  assign n16379 = n16252 & n16378 ;
  assign n16380 = n16379 ^ n13726 ;
  assign n16381 = n16380 ^ n16376 ;
  assign n16382 = n16377 & ~n16381 ;
  assign n16383 = n16382 ^ n13822 ;
  assign n16384 = n16383 ^ n16374 ;
  assign n16385 = ~n16375 & n16384 ;
  assign n16386 = n16385 ^ n13830 ;
  assign n16373 = n16321 ^ n16303 ;
  assign n16387 = n16386 ^ n16373 ;
  assign n16388 = n16386 ^ n13837 ;
  assign n16389 = ~n16387 & n16388 ;
  assign n16390 = n16389 ^ n13837 ;
  assign n16391 = n16390 ^ n16371 ;
  assign n16392 = n16372 & ~n16391 ;
  assign n16393 = n16392 ^ n13836 ;
  assign n16370 = n16327 ^ n16292 ;
  assign n16394 = n16393 ^ n16370 ;
  assign n16395 = n16393 ^ n13847 ;
  assign n16396 = ~n16394 & n16395 ;
  assign n16397 = n16396 ^ n13847 ;
  assign n16399 = n16398 ^ n16397 ;
  assign n16400 = n16398 ^ n13988 ;
  assign n16401 = n16399 & n16400 ;
  assign n16402 = n16401 ^ n13988 ;
  assign n16403 = n16402 ^ n16368 ;
  assign n16404 = n16369 & ~n16403 ;
  assign n16405 = n16404 ^ n13316 ;
  assign n16406 = n16405 ^ n16366 ;
  assign n16407 = n16367 & n16406 ;
  assign n16408 = n16407 ^ n13315 ;
  assign n16409 = n16408 ^ n13312 ;
  assign n16410 = n16346 ^ n16344 ;
  assign n16411 = n16410 ^ n16408 ;
  assign n16412 = n16409 & ~n16411 ;
  assign n16413 = n16412 ^ n13312 ;
  assign n16365 = n16355 ^ n16352 ;
  assign n16414 = n16413 ^ n16365 ;
  assign n16415 = n16413 ^ n13355 ;
  assign n16416 = ~n16414 & n16415 ;
  assign n16417 = n16416 ^ n13355 ;
  assign n16418 = n16417 ^ n16363 ;
  assign n16419 = n16364 & n16418 ;
  assign n16420 = n16419 ^ n13384 ;
  assign n16534 = n16430 ^ n16420 ;
  assign n16432 = n16405 ^ n16367 ;
  assign n16433 = n16400 ^ n16397 ;
  assign n16434 = n16370 ^ n13847 ;
  assign n16435 = n16434 ^ n16393 ;
  assign n16436 = n16390 ^ n16372 ;
  assign n16437 = n16373 ^ n13837 ;
  assign n16438 = n16437 ^ n16386 ;
  assign n16253 = n16252 ^ n16243 ;
  assign n16077 = n16076 ^ n16067 ;
  assign n16078 = n16053 ^ n16006 ;
  assign n16079 = n16050 ^ n16008 ;
  assign n16080 = n16048 ^ n16045 ;
  assign n16082 = n16020 ^ n16019 ;
  assign n16083 = ~n16081 & n16082 ;
  assign n16084 = n16026 ^ n16023 ;
  assign n16085 = n16083 & n16084 ;
  assign n16086 = n16028 ^ n16016 ;
  assign n16087 = n16085 & n16086 ;
  assign n16088 = n16034 ^ n16031 ;
  assign n16089 = n16087 & ~n16088 ;
  assign n16090 = n16036 ^ n16014 ;
  assign n16091 = ~n16089 & n16090 ;
  assign n16092 = n16039 ^ n16012 ;
  assign n16093 = ~n16091 & n16092 ;
  assign n16094 = n16042 ^ n16010 ;
  assign n16095 = ~n16093 & n16094 ;
  assign n16096 = n16080 & n16095 ;
  assign n16097 = n16079 & n16096 ;
  assign n16098 = ~n16078 & ~n16097 ;
  assign n16099 = n16004 ^ n13454 ;
  assign n16100 = n16099 ^ n16056 ;
  assign n16101 = ~n16098 & ~n16100 ;
  assign n16102 = n16060 ^ n16003 ;
  assign n16103 = ~n16101 & ~n16102 ;
  assign n16104 = n16001 ^ n13616 ;
  assign n16105 = n16104 ^ n16063 ;
  assign n16106 = ~n16103 & ~n16105 ;
  assign n16107 = n16077 & n16106 ;
  assign n16121 = n16120 ^ n16110 ;
  assign n16122 = n16107 & n16121 ;
  assign n16135 = n16134 ^ n16131 ;
  assign n16222 = n16122 & n16135 ;
  assign n16235 = n16234 ^ n16225 ;
  assign n16254 = ~n16222 & ~n16235 ;
  assign n16439 = n16253 & n16254 ;
  assign n16440 = n16380 ^ n16377 ;
  assign n16441 = ~n16439 & n16440 ;
  assign n16442 = n16383 ^ n16375 ;
  assign n16443 = n16441 & ~n16442 ;
  assign n16444 = ~n16438 & ~n16443 ;
  assign n16445 = n16436 & ~n16444 ;
  assign n16446 = n16435 & n16445 ;
  assign n16447 = ~n16433 & ~n16446 ;
  assign n16448 = n16402 ^ n16369 ;
  assign n16449 = ~n16447 & ~n16448 ;
  assign n16450 = ~n16432 & n16449 ;
  assign n16451 = n16410 ^ n16409 ;
  assign n16452 = n16450 & n16451 ;
  assign n16453 = n16365 ^ n13355 ;
  assign n16454 = n16453 ^ n16413 ;
  assign n16455 = ~n16452 & ~n16454 ;
  assign n16456 = n16417 ^ n16364 ;
  assign n16457 = ~n16455 & n16456 ;
  assign n16537 = n16534 ^ n16457 ;
  assign n16538 = n12950 & n16537 ;
  assign n16535 = n16457 ^ n16420 ;
  assign n16536 = n16534 & n16535 ;
  assign n16539 = n16538 ^ n16536 ;
  assign n16531 = n16429 ^ n16422 ;
  assign n16532 = n16427 & n16531 ;
  assign n16528 = n15919 ^ n1832 ;
  assign n16525 = n14375 ^ n13755 ;
  assign n16526 = n16525 ^ n16429 ;
  assign n16527 = n16526 ^ n15367 ;
  assign n16529 = n16528 ^ n16527 ;
  assign n16530 = n16529 ^ n13390 ;
  assign n16533 = n16532 ^ n16530 ;
  assign n16540 = n16539 ^ n16533 ;
  assign n16542 = n16541 ^ n16540 ;
  assign n16421 = n16420 ^ n12950 ;
  assign n16431 = n16430 ^ n16421 ;
  assign n16458 = n16457 ^ n16431 ;
  assign n16459 = n16458 ^ n1781 ;
  assign n16517 = n16456 ^ n16455 ;
  assign n16460 = n16454 ^ n16452 ;
  assign n16461 = n16460 ^ n1817 ;
  assign n16463 = n16449 ^ n16432 ;
  assign n16464 = n16463 ^ n3133 ;
  assign n16466 = n16446 ^ n16433 ;
  assign n16467 = n16466 ^ n2621 ;
  assign n16468 = n16445 ^ n16435 ;
  assign n16469 = n16468 ^ n2544 ;
  assign n16471 = n16443 ^ n16438 ;
  assign n16472 = n16471 ^ n1276 ;
  assign n16474 = n16440 ^ n16439 ;
  assign n16475 = n16474 ^ n1102 ;
  assign n16255 = n16254 ^ n16253 ;
  assign n16256 = n16255 ^ n925 ;
  assign n16476 = n16474 ^ n925 ;
  assign n16477 = n16476 ^ n16474 ;
  assign n16236 = n16235 ^ n16222 ;
  assign n16136 = n16135 ^ n16122 ;
  assign n16137 = n16136 ^ n773 ;
  assign n16138 = n16121 ^ n16107 ;
  assign n16139 = n16138 ^ n694 ;
  assign n16140 = n16106 ^ n16077 ;
  assign n16141 = n16140 ^ n688 ;
  assign n16142 = n16105 ^ n16103 ;
  assign n16143 = n16142 ^ n632 ;
  assign n16146 = n16102 ^ n16101 ;
  assign n16147 = n16146 ^ n626 ;
  assign n16203 = n16100 ^ n16098 ;
  assign n16148 = n16097 ^ n16078 ;
  assign n16149 = n16148 ^ n1492 ;
  assign n16199 = n16148 ^ n2909 ;
  assign n16150 = n16096 ^ n16079 ;
  assign n16151 = n16150 ^ n2909 ;
  assign n16152 = n16095 ^ n16080 ;
  assign n16156 = n16155 ^ n16152 ;
  assign n16157 = n16094 ^ n16093 ;
  assign n16158 = n16157 ^ n584 ;
  assign n16161 = n16092 ^ n16091 ;
  assign n16162 = n16161 ^ n2215 ;
  assign n16163 = n16090 ^ n16089 ;
  assign n16164 = n16163 ^ n2209 ;
  assign n16185 = n16163 ^ n2090 ;
  assign n16165 = n16088 ^ n16087 ;
  assign n16166 = n16165 ^ n2090 ;
  assign n16167 = n16086 ^ n16085 ;
  assign n16168 = n16167 ^ n2013 ;
  assign n16169 = n3051 & n16081 ;
  assign n1992 = n1949 ^ x255 ;
  assign n1993 = n1992 ^ x447 ;
  assign n1994 = n1993 ^ x191 ;
  assign n16170 = n16169 ^ n1994 ;
  assign n16171 = n16082 ^ n16081 ;
  assign n16172 = n16171 ^ n16169 ;
  assign n16173 = n16170 & n16172 ;
  assign n16174 = n16173 ^ n1994 ;
  assign n16175 = n16174 ^ n2001 ;
  assign n16176 = n16084 ^ n16083 ;
  assign n16177 = n16176 ^ n2001 ;
  assign n16178 = n16175 & n16177 ;
  assign n16179 = n16178 ^ n2001 ;
  assign n16180 = n16179 ^ n16167 ;
  assign n16181 = n16168 & ~n16180 ;
  assign n16182 = n16181 ^ n2013 ;
  assign n16183 = n16182 ^ n2090 ;
  assign n16184 = ~n16166 & n16183 ;
  assign n16186 = n16185 ^ n16184 ;
  assign n16187 = n16164 & n16186 ;
  assign n16188 = n16187 ^ n16163 ;
  assign n16189 = n16188 ^ n16161 ;
  assign n16190 = ~n16162 & n16189 ;
  assign n16191 = n16190 ^ n2215 ;
  assign n16159 = n16152 ^ n584 ;
  assign n16160 = n16159 ^ n16152 ;
  assign n16192 = n16191 ^ n16160 ;
  assign n16193 = n16158 & n16192 ;
  assign n16194 = n16193 ^ n16159 ;
  assign n16195 = ~n16156 & n16194 ;
  assign n16196 = n16195 ^ n16155 ;
  assign n16197 = n16196 ^ n2909 ;
  assign n16198 = ~n16151 & n16197 ;
  assign n16200 = n16199 ^ n16198 ;
  assign n16201 = n16149 & ~n16200 ;
  assign n16202 = n16201 ^ n1492 ;
  assign n16204 = n16203 ^ n16202 ;
  assign n16205 = n16202 ^ n1498 ;
  assign n16206 = ~n16204 & ~n16205 ;
  assign n16207 = n16206 ^ n16203 ;
  assign n16208 = n16207 ^ n626 ;
  assign n16209 = n16147 & n16208 ;
  assign n16210 = n16209 ^ n16146 ;
  assign n16144 = n16140 ^ n632 ;
  assign n16145 = n16144 ^ n16140 ;
  assign n16211 = n16210 ^ n16145 ;
  assign n16212 = ~n16143 & n16211 ;
  assign n16213 = n16212 ^ n16144 ;
  assign n16214 = ~n16141 & ~n16213 ;
  assign n16215 = n16214 ^ n16140 ;
  assign n16216 = n16215 ^ n694 ;
  assign n16217 = ~n16139 & n16216 ;
  assign n16218 = n16217 ^ n16138 ;
  assign n16219 = n16218 ^ n16136 ;
  assign n16220 = ~n16137 & ~n16219 ;
  assign n16221 = n16220 ^ n773 ;
  assign n16237 = n16236 ^ n16221 ;
  assign n16238 = n16221 ^ n1110 ;
  assign n16239 = n16237 & ~n16238 ;
  assign n16240 = n16239 ^ n16236 ;
  assign n16478 = n16477 ^ n16240 ;
  assign n16479 = n16256 & n16478 ;
  assign n16480 = n16479 ^ n16476 ;
  assign n16481 = n16475 & ~n16480 ;
  assign n16482 = n16481 ^ n1102 ;
  assign n16486 = n16482 ^ n16471 ;
  assign n16473 = n16442 ^ n16441 ;
  assign n16483 = n16482 ^ n16473 ;
  assign n16484 = n16473 ^ n1133 ;
  assign n16485 = n16483 & ~n16484 ;
  assign n16487 = n16486 ^ n16485 ;
  assign n16488 = n16472 & ~n16487 ;
  assign n16489 = n16488 ^ n1276 ;
  assign n16470 = n16444 ^ n16436 ;
  assign n16490 = n16489 ^ n16470 ;
  assign n16491 = n16468 ^ n2788 ;
  assign n16492 = n16491 ^ n16468 ;
  assign n16493 = n16492 ^ n16470 ;
  assign n16494 = ~n16490 & n16493 ;
  assign n16495 = n16494 ^ n16491 ;
  assign n16496 = ~n16469 & n16495 ;
  assign n16497 = n16496 ^ n2544 ;
  assign n16498 = n16497 ^ n16466 ;
  assign n16499 = n16467 & ~n16498 ;
  assign n16500 = n16499 ^ n2621 ;
  assign n16465 = n16448 ^ n16447 ;
  assign n16501 = n16500 ^ n16465 ;
  assign n16502 = n16463 ^ n2480 ;
  assign n16503 = n16502 ^ n16463 ;
  assign n16504 = n16503 ^ n16465 ;
  assign n16505 = n16501 & ~n16504 ;
  assign n16506 = n16505 ^ n16502 ;
  assign n16507 = n16464 & ~n16506 ;
  assign n16508 = n16507 ^ n3133 ;
  assign n16462 = n16451 ^ n16450 ;
  assign n16509 = n16508 ^ n16462 ;
  assign n16510 = n16460 ^ n2465 ;
  assign n16511 = n16510 ^ n16460 ;
  assign n16512 = n16511 ^ n16462 ;
  assign n16513 = n16509 & ~n16512 ;
  assign n16514 = n16513 ^ n16510 ;
  assign n16515 = n16461 & ~n16514 ;
  assign n16516 = n16515 ^ n1817 ;
  assign n16518 = n16517 ^ n16516 ;
  assign n16519 = n16458 ^ n2763 ;
  assign n16520 = n16519 ^ n16458 ;
  assign n16521 = n16520 ^ n16516 ;
  assign n16522 = ~n16518 & n16521 ;
  assign n16523 = n16522 ^ n16519 ;
  assign n16524 = ~n16459 & n16523 ;
  assign n16543 = n16542 ^ n16524 ;
  assign n16574 = n16543 ^ n16275 ;
  assign n16279 = n14937 ^ n14356 ;
  assign n16280 = n16279 ^ n15693 ;
  assign n16544 = n16543 ^ n16280 ;
  assign n16547 = n16523 ^ n1781 ;
  assign n16545 = n15699 ^ n14939 ;
  assign n16546 = n16545 ^ n14358 ;
  assign n16548 = n16547 ^ n16546 ;
  assign n16552 = n14945 ^ n14364 ;
  assign n16553 = n16552 ^ n15701 ;
  assign n16549 = n16517 ^ n2763 ;
  assign n16550 = n16549 ^ n16516 ;
  assign n16554 = n16553 ^ n16550 ;
  assign n16557 = n14954 ^ n14696 ;
  assign n16558 = n16557 ^ n15711 ;
  assign n16559 = n16462 ^ n2465 ;
  assign n16560 = n16559 ^ n16508 ;
  assign n16561 = ~n16558 & ~n16560 ;
  assign n16555 = n14952 ^ n14700 ;
  assign n16556 = n16555 ^ n15707 ;
  assign n16562 = n16561 ^ n16556 ;
  assign n16563 = n16514 ^ n1817 ;
  assign n16564 = n16563 ^ n16556 ;
  assign n16565 = n16562 & ~n16564 ;
  assign n16566 = n16565 ^ n16561 ;
  assign n16567 = n16566 ^ n16550 ;
  assign n16568 = ~n16554 & n16567 ;
  assign n16551 = n16550 ^ n16547 ;
  assign n16569 = n16568 ^ n16551 ;
  assign n16570 = ~n16548 & ~n16569 ;
  assign n16571 = n16570 ^ n16547 ;
  assign n16572 = n16571 ^ n16543 ;
  assign n16573 = ~n16544 & n16572 ;
  assign n16575 = n16574 ^ n16573 ;
  assign n16576 = n16278 & n16575 ;
  assign n16577 = n16576 ^ n16277 ;
  assign n16272 = n14927 ^ n14891 ;
  assign n16273 = n16272 ^ n15685 ;
  assign n16270 = n16171 ^ n16170 ;
  assign n16274 = n16273 ^ n16270 ;
  assign n16641 = n16577 ^ n16274 ;
  assign n16643 = n16641 ^ n13728 ;
  assign n16614 = n16575 ^ n16277 ;
  assign n16615 = n16614 ^ n13736 ;
  assign n16633 = n16571 ^ n16544 ;
  assign n16616 = n16569 ^ n16546 ;
  assign n16617 = n16616 ^ n13744 ;
  assign n16625 = n16566 ^ n16554 ;
  assign n16618 = n16560 ^ n16558 ;
  assign n16619 = n13749 & n16618 ;
  assign n16620 = n16619 ^ n14061 ;
  assign n16621 = n16563 ^ n16562 ;
  assign n16622 = n16621 ^ n16619 ;
  assign n16623 = n16620 & ~n16622 ;
  assign n16624 = n16623 ^ n14061 ;
  assign n16626 = n16625 ^ n16624 ;
  assign n16627 = n16625 ^ n14067 ;
  assign n16628 = n16626 & n16627 ;
  assign n16629 = n16628 ^ n14067 ;
  assign n16630 = n16629 ^ n16616 ;
  assign n16631 = ~n16617 & ~n16630 ;
  assign n16632 = n16631 ^ n13744 ;
  assign n16634 = n16633 ^ n16632 ;
  assign n16635 = n16633 ^ n13738 ;
  assign n16636 = ~n16634 & ~n16635 ;
  assign n16637 = n16636 ^ n13738 ;
  assign n16638 = n16637 ^ n16614 ;
  assign n16639 = ~n16615 & ~n16638 ;
  assign n16640 = n16639 ^ n13736 ;
  assign n16660 = n16643 ^ n16640 ;
  assign n16661 = n16629 ^ n16617 ;
  assign n16662 = n16618 ^ n13749 ;
  assign n16663 = n16621 ^ n16620 ;
  assign n16664 = n16662 & n16663 ;
  assign n16665 = n16627 ^ n16624 ;
  assign n16666 = n16664 & n16665 ;
  assign n16667 = n16661 & n16666 ;
  assign n16668 = n16635 ^ n16632 ;
  assign n16669 = n16667 & ~n16668 ;
  assign n16670 = n16637 ^ n16615 ;
  assign n16671 = ~n16669 & ~n16670 ;
  assign n16672 = n16660 & ~n16671 ;
  assign n16642 = n16641 ^ n16640 ;
  assign n16644 = n16642 & n16643 ;
  assign n16645 = n16644 ^ n13728 ;
  assign n16578 = n16577 ^ n16270 ;
  assign n16579 = ~n16274 & ~n16578 ;
  assign n16266 = n16177 ^ n16174 ;
  assign n16271 = n16270 ^ n16266 ;
  assign n16580 = n16579 ^ n16271 ;
  assign n16267 = n14947 ^ n14920 ;
  assign n16268 = n16267 ^ n15678 ;
  assign n16612 = n16580 ^ n16268 ;
  assign n16613 = n16612 ^ n14084 ;
  assign n16659 = n16645 ^ n16613 ;
  assign n16713 = n16672 ^ n16659 ;
  assign n16714 = n16713 ^ n1463 ;
  assign n16717 = n16671 ^ n16660 ;
  assign n16718 = n16717 ^ n2304 ;
  assign n16719 = n16670 ^ n16669 ;
  assign n16720 = n16719 ^ n2191 ;
  assign n16721 = n16668 ^ n16667 ;
  assign n16722 = n16721 ^ n2171 ;
  assign n16725 = n16666 ^ n16661 ;
  assign n16726 = n16725 ^ n2175 ;
  assign n1873 = n1791 ^ x256 ;
  assign n1874 = n1873 ^ x448 ;
  assign n1875 = n1874 ^ x192 ;
  assign n16730 = n1875 & ~n16662 ;
  assign n16727 = n14844 ^ x287 ;
  assign n16728 = n16727 ^ x479 ;
  assign n16729 = n16728 ^ x223 ;
  assign n16731 = n16730 ^ n16729 ;
  assign n16732 = n16663 ^ n16662 ;
  assign n16733 = n16732 ^ n16729 ;
  assign n16734 = n16731 & ~n16733 ;
  assign n16735 = n16734 ^ n16730 ;
  assign n1929 = n1898 ^ x286 ;
  assign n1930 = n1929 ^ x478 ;
  assign n1931 = n1930 ^ x222 ;
  assign n16736 = n16735 ^ n1931 ;
  assign n16737 = n16665 ^ n16664 ;
  assign n16738 = n16737 ^ n1931 ;
  assign n16739 = n16736 & n16738 ;
  assign n16740 = n16739 ^ n1931 ;
  assign n16741 = n16740 ^ n16725 ;
  assign n16742 = n16726 & ~n16741 ;
  assign n16743 = n16742 ^ n2175 ;
  assign n16723 = n16719 ^ n2171 ;
  assign n16724 = n16723 ^ n16719 ;
  assign n16744 = n16743 ^ n16724 ;
  assign n16745 = ~n16722 & n16744 ;
  assign n16746 = n16745 ^ n16723 ;
  assign n16747 = ~n16720 & n16746 ;
  assign n16748 = n16747 ^ n2191 ;
  assign n16749 = n16748 ^ n2304 ;
  assign n16750 = ~n16718 & ~n16749 ;
  assign n16751 = n16750 ^ n16717 ;
  assign n16646 = n16645 ^ n16612 ;
  assign n16647 = n16613 & ~n16646 ;
  assign n16648 = n16647 ^ n14084 ;
  assign n16269 = n16268 ^ n16266 ;
  assign n16581 = n16269 & n16580 ;
  assign n16582 = n16581 ^ n16268 ;
  assign n16260 = n14942 ^ n14911 ;
  assign n16261 = n16260 ^ n15682 ;
  assign n16259 = n16179 ^ n16168 ;
  assign n16262 = n16261 ^ n16259 ;
  assign n16610 = n16582 ^ n16262 ;
  assign n16611 = n16610 ^ n14097 ;
  assign n16674 = n16648 ^ n16611 ;
  assign n16673 = n16659 & ~n16672 ;
  assign n16708 = n16674 ^ n16673 ;
  assign n16715 = n16708 ^ n1463 ;
  assign n16716 = n16715 ^ n16708 ;
  assign n16752 = n16751 ^ n16716 ;
  assign n16753 = n16714 & ~n16752 ;
  assign n16754 = n16753 ^ n16715 ;
  assign n16810 = n16754 ^ n16711 ;
  assign n16808 = n16210 ^ n16143 ;
  assign n16807 = n16304 ^ n15526 ;
  assign n16809 = n16808 ^ n16807 ;
  assign n16811 = n16810 ^ n16809 ;
  assign n16815 = n16751 ^ n16714 ;
  assign n16813 = n16207 ^ n16147 ;
  assign n16812 = n16310 ^ n15419 ;
  assign n16814 = n16813 ^ n16812 ;
  assign n16816 = n16815 ^ n16814 ;
  assign n16821 = n16748 ^ n16718 ;
  assign n16818 = n16203 ^ n1498 ;
  assign n16819 = n16818 ^ n16202 ;
  assign n16817 = n16246 ^ n14898 ;
  assign n16820 = n16819 ^ n16817 ;
  assign n16822 = n16821 ^ n16820 ;
  assign n17251 = n16746 ^ n2191 ;
  assign n17254 = n17251 ^ n16821 ;
  assign n16826 = n16743 ^ n16722 ;
  assign n16824 = n16196 ^ n16151 ;
  assign n16823 = n16126 ^ n14909 ;
  assign n16825 = n16824 ^ n16823 ;
  assign n16827 = n16826 ^ n16825 ;
  assign n16835 = n16740 ^ n16726 ;
  assign n16833 = n16111 ^ n14911 ;
  assign n16770 = n16194 ^ n16155 ;
  assign n16834 = n16833 ^ n16770 ;
  assign n16836 = n16835 ^ n16834 ;
  assign n16838 = n16070 ^ n14920 ;
  assign n16685 = n16191 ^ n16158 ;
  assign n16839 = n16838 ^ n16685 ;
  assign n16837 = n16738 ^ n16735 ;
  assign n16840 = n16839 ^ n16837 ;
  assign n16842 = n15678 ^ n14932 ;
  assign n16586 = n16186 ^ n2209 ;
  assign n16843 = n16842 ^ n16586 ;
  assign n16841 = n16662 ^ n1875 ;
  assign n16844 = n16843 ^ n16841 ;
  assign n16863 = n15260 ^ n14667 ;
  assign n16864 = n16863 ^ n16422 ;
  assign n16862 = n16484 ^ n16482 ;
  assign n16865 = n16864 ^ n16862 ;
  assign n16868 = n15870 ^ n15357 ;
  assign n16869 = n16868 ^ n16353 ;
  assign n16787 = n16480 ^ n1102 ;
  assign n16870 = n16869 ^ n16787 ;
  assign n16931 = n15836 ^ n15318 ;
  assign n16932 = n16931 ^ n16347 ;
  assign n16871 = n15821 ^ n15295 ;
  assign n16872 = n16871 ^ n16339 ;
  assign n16792 = n16236 ^ n1110 ;
  assign n16793 = n16792 ^ n16221 ;
  assign n16873 = n16872 ^ n16793 ;
  assign n16876 = n16218 ^ n16137 ;
  assign n16874 = n15770 ^ n15278 ;
  assign n16875 = n16874 ^ n16284 ;
  assign n16877 = n16876 ^ n16875 ;
  assign n16878 = n15762 ^ n15247 ;
  assign n16879 = n16878 ^ n15675 ;
  assign n16803 = n16215 ^ n16139 ;
  assign n16880 = n16879 ^ n16803 ;
  assign n16798 = n16213 ^ n688 ;
  assign n16914 = n16808 ^ n16798 ;
  assign n16881 = n15676 ^ n15144 ;
  assign n16882 = n16881 ^ n16293 ;
  assign n16883 = n16882 ^ n16808 ;
  assign n16884 = n15738 ^ n15099 ;
  assign n16885 = n16884 ^ n16295 ;
  assign n16886 = n16885 ^ n16813 ;
  assign n16908 = n16819 ^ n16813 ;
  assign n16829 = n16200 ^ n1492 ;
  assign n16895 = n16829 ^ n16824 ;
  assign n16887 = n15724 ^ n14907 ;
  assign n16888 = n16887 ^ n16310 ;
  assign n16889 = n16888 ^ n16824 ;
  assign n16892 = n16824 ^ n16770 ;
  assign n16263 = n16182 ^ n16166 ;
  assign n16264 = n16263 ^ n16259 ;
  assign n16265 = n16264 ^ n16263 ;
  assign n16583 = n16582 ^ n16265 ;
  assign n16584 = ~n16262 & n16583 ;
  assign n16585 = n16584 ^ n16264 ;
  assign n16590 = n16586 ^ n16263 ;
  assign n16587 = n14935 ^ n14909 ;
  assign n16588 = n16587 ^ n16070 ;
  assign n16589 = n16588 ^ n16586 ;
  assign n16591 = n16590 ^ n16589 ;
  assign n16592 = ~n16585 & n16591 ;
  assign n16593 = n16592 ^ n16590 ;
  assign n16594 = n16188 ^ n16162 ;
  assign n16598 = n16594 ^ n16586 ;
  assign n16595 = n14930 ^ n14900 ;
  assign n16596 = n16595 ^ n16111 ;
  assign n16597 = n16596 ^ n16594 ;
  assign n16599 = n16598 ^ n16597 ;
  assign n16600 = ~n16593 & ~n16599 ;
  assign n16601 = n16600 ^ n16598 ;
  assign n16687 = n16685 ^ n16594 ;
  assign n16602 = n14925 ^ n14898 ;
  assign n16603 = n16602 ^ n16126 ;
  assign n16686 = n16685 ^ n16603 ;
  assign n16688 = n16687 ^ n16686 ;
  assign n16689 = ~n16601 & ~n16688 ;
  assign n16690 = n16689 ^ n16687 ;
  assign n16772 = n16770 ^ n16685 ;
  assign n16691 = n15419 ^ n14917 ;
  assign n16692 = n16691 ^ n16231 ;
  assign n16771 = n16770 ^ n16692 ;
  assign n16773 = n16772 ^ n16771 ;
  assign n16774 = ~n16690 & n16773 ;
  assign n16775 = n16774 ^ n16772 ;
  assign n16776 = n15526 ^ n14914 ;
  assign n16777 = n16776 ^ n16246 ;
  assign n16890 = n16777 ^ n16770 ;
  assign n16891 = ~n16775 & n16890 ;
  assign n16893 = n16892 ^ n16891 ;
  assign n16894 = n16889 & n16893 ;
  assign n16896 = n16895 ^ n16894 ;
  assign n16898 = n16304 ^ n15717 ;
  assign n16899 = n16898 ^ n14903 ;
  assign n16897 = n16829 ^ n16819 ;
  assign n16900 = n16899 ^ n16897 ;
  assign n16901 = n16900 ^ n16819 ;
  assign n16902 = ~n16896 & n16901 ;
  assign n16903 = n16902 ^ n16897 ;
  assign n16904 = n15719 ^ n14351 ;
  assign n16905 = n16904 ^ n16300 ;
  assign n16906 = n16905 ^ n16819 ;
  assign n16907 = ~n16903 & ~n16906 ;
  assign n16909 = n16908 ^ n16907 ;
  assign n16910 = n16886 & ~n16909 ;
  assign n16911 = n16910 ^ n16885 ;
  assign n16912 = n16911 ^ n16808 ;
  assign n16913 = n16883 & n16912 ;
  assign n16915 = n16914 ^ n16913 ;
  assign n16918 = n15752 ^ n15228 ;
  assign n16919 = n16918 ^ n16287 ;
  assign n16916 = n16803 ^ n16798 ;
  assign n16917 = n16916 ^ n16803 ;
  assign n16920 = n16919 ^ n16917 ;
  assign n16921 = n16915 & n16920 ;
  assign n16922 = n16921 ^ n16916 ;
  assign n16923 = n16880 & ~n16922 ;
  assign n16924 = n16923 ^ n16803 ;
  assign n16925 = n16924 ^ n16875 ;
  assign n16926 = ~n16877 & n16925 ;
  assign n16927 = n16926 ^ n16876 ;
  assign n16928 = n16927 ^ n16872 ;
  assign n16929 = ~n16873 & n16928 ;
  assign n16930 = n16929 ^ n16793 ;
  assign n16933 = n16932 ^ n16930 ;
  assign n16257 = n16256 ^ n16240 ;
  assign n16934 = n16787 ^ n16257 ;
  assign n16935 = n16934 ^ n16787 ;
  assign n16936 = n16935 ^ n16930 ;
  assign n16937 = ~n16933 & n16936 ;
  assign n16938 = n16937 ^ n16934 ;
  assign n16939 = n16870 & n16938 ;
  assign n16940 = n16939 ^ n16787 ;
  assign n16866 = n15312 ^ n14669 ;
  assign n16867 = n16866 ^ n16528 ;
  assign n16941 = n16940 ^ n16867 ;
  assign n16942 = n16941 ^ n16862 ;
  assign n16943 = n16942 ^ n16867 ;
  assign n16944 = n16865 & n16943 ;
  assign n16945 = n16944 ^ n16941 ;
  assign n16949 = n16487 ^ n1276 ;
  assign n16946 = n15309 ^ n14662 ;
  assign n16947 = n16946 ^ n15956 ;
  assign n16950 = n16949 ^ n16947 ;
  assign n16948 = n16947 ^ n16867 ;
  assign n16951 = n16950 ^ n16948 ;
  assign n16952 = n16945 & n16951 ;
  assign n16953 = n16952 ^ n16948 ;
  assign n16955 = n16470 ^ n2788 ;
  assign n16956 = n16955 ^ n16489 ;
  assign n16859 = n15339 ^ n14682 ;
  assign n16860 = n16859 ^ n15961 ;
  assign n16957 = n16956 ^ n16860 ;
  assign n16954 = n16947 ^ n16860 ;
  assign n16958 = n16957 ^ n16954 ;
  assign n16959 = n16953 & n16958 ;
  assign n16960 = n16959 ^ n16954 ;
  assign n16858 = n16495 ^ n2544 ;
  assign n17048 = n16960 ^ n16858 ;
  assign n16970 = n16949 ^ n16945 ;
  assign n16971 = n16970 ^ n14020 ;
  assign n16973 = n16938 ^ n16869 ;
  assign n16974 = n16973 ^ n14572 ;
  assign n17025 = n16932 ^ n16257 ;
  assign n17026 = n17025 ^ n16930 ;
  assign n16976 = n16924 ^ n16877 ;
  assign n16977 = n16976 ^ n14465 ;
  assign n16979 = n16919 ^ n16915 ;
  assign n16980 = n16979 ^ n14389 ;
  assign n16982 = n16905 ^ n16903 ;
  assign n16983 = n16982 ^ n14402 ;
  assign n16984 = n16899 ^ n16896 ;
  assign n16985 = n16984 ^ n14408 ;
  assign n16986 = n16893 ^ n16888 ;
  assign n16987 = n16986 ^ n14416 ;
  assign n16778 = n16777 ^ n16775 ;
  assign n16779 = n16778 ^ n14418 ;
  assign n16693 = n16692 ^ n16690 ;
  assign n16694 = n16693 ^ n14426 ;
  assign n16606 = n16596 ^ n16593 ;
  assign n16607 = n16606 ^ n14190 ;
  assign n16608 = n16588 ^ n16585 ;
  assign n16609 = n16608 ^ n14176 ;
  assign n16649 = n16648 ^ n16610 ;
  assign n16650 = ~n16611 & ~n16649 ;
  assign n16651 = n16650 ^ n14097 ;
  assign n16652 = n16651 ^ n16608 ;
  assign n16653 = ~n16609 & ~n16652 ;
  assign n16654 = n16653 ^ n14176 ;
  assign n16655 = n16654 ^ n16606 ;
  assign n16656 = n16607 & n16655 ;
  assign n16657 = n16656 ^ n14190 ;
  assign n16604 = n16603 ^ n16601 ;
  assign n16681 = n16657 ^ n16604 ;
  assign n16682 = n16657 ^ n14333 ;
  assign n16683 = n16681 & n16682 ;
  assign n16684 = n16683 ^ n14333 ;
  assign n16767 = n16693 ^ n16684 ;
  assign n16768 = n16694 & n16767 ;
  assign n16769 = n16768 ^ n14426 ;
  assign n16988 = n16778 ^ n16769 ;
  assign n16989 = n16779 & n16988 ;
  assign n16990 = n16989 ^ n14418 ;
  assign n16991 = n16990 ^ n16986 ;
  assign n16992 = ~n16987 & n16991 ;
  assign n16993 = n16992 ^ n14416 ;
  assign n16994 = n16993 ^ n16984 ;
  assign n16995 = ~n16985 & n16994 ;
  assign n16996 = n16995 ^ n14408 ;
  assign n16997 = n16996 ^ n16982 ;
  assign n16998 = n16983 & n16997 ;
  assign n16999 = n16998 ^ n14402 ;
  assign n16981 = n16909 ^ n16885 ;
  assign n17000 = n16999 ^ n16981 ;
  assign n17001 = n16911 ^ n16883 ;
  assign n17002 = n17001 ^ n14447 ;
  assign n17003 = n17002 ^ n16981 ;
  assign n17004 = n17003 ^ n17001 ;
  assign n17005 = ~n17000 & ~n17004 ;
  assign n17006 = n17005 ^ n17002 ;
  assign n17008 = n16979 ^ n13725 ;
  assign n17007 = n17001 ^ n16979 ;
  assign n17009 = n17008 ^ n17007 ;
  assign n17010 = n17006 & n17009 ;
  assign n17011 = n17010 ^ n17008 ;
  assign n17012 = ~n16980 & ~n17011 ;
  assign n17013 = n17012 ^ n14389 ;
  assign n16978 = n16922 ^ n16879 ;
  assign n17014 = n17013 ^ n16978 ;
  assign n17015 = n17013 ^ n14383 ;
  assign n17016 = n17014 & n17015 ;
  assign n17017 = n17016 ^ n14383 ;
  assign n17018 = n17017 ^ n16976 ;
  assign n17019 = ~n16977 & n17018 ;
  assign n17020 = n17019 ^ n14465 ;
  assign n16975 = n16927 ^ n16873 ;
  assign n17021 = n17020 ^ n16975 ;
  assign n17022 = n17020 ^ n14468 ;
  assign n17023 = n17021 & ~n17022 ;
  assign n17024 = n17023 ^ n14468 ;
  assign n17027 = n17026 ^ n17024 ;
  assign n17028 = n16973 ^ n14472 ;
  assign n17029 = n17028 ^ n16973 ;
  assign n17030 = n17029 ^ n17024 ;
  assign n17031 = n17027 & n17030 ;
  assign n17032 = n17031 ^ n17028 ;
  assign n17033 = ~n16974 & n17032 ;
  assign n17034 = n17033 ^ n14572 ;
  assign n16972 = n16940 ^ n16865 ;
  assign n17035 = n17034 ^ n16972 ;
  assign n17036 = n16970 ^ n14025 ;
  assign n17037 = n17036 ^ n16972 ;
  assign n17038 = n17037 ^ n16970 ;
  assign n17039 = ~n17035 & n17038 ;
  assign n17040 = n17039 ^ n17036 ;
  assign n17041 = ~n16971 & n17040 ;
  assign n17042 = n17041 ^ n14020 ;
  assign n17043 = n17042 ^ n14018 ;
  assign n17044 = n16956 ^ n16953 ;
  assign n17045 = n17044 ^ n17042 ;
  assign n17046 = n17043 & n17045 ;
  assign n17047 = n17046 ^ n14018 ;
  assign n17049 = n17048 ^ n17047 ;
  assign n16861 = n16860 ^ n16858 ;
  assign n16961 = ~n16861 & n16960 ;
  assign n16962 = n16961 ^ n16860 ;
  assign n16856 = n16497 ^ n16467 ;
  assign n16854 = n15367 ^ n14651 ;
  assign n16855 = n16854 ^ n15952 ;
  assign n16857 = n16856 ^ n16855 ;
  assign n16968 = n16962 ^ n16857 ;
  assign n17050 = n16968 ^ n14009 ;
  assign n17051 = n17050 ^ n17047 ;
  assign n17052 = n17051 ^ n16968 ;
  assign n17053 = ~n17049 & n17052 ;
  assign n17054 = n17053 ^ n17050 ;
  assign n17098 = n17054 ^ n14004 ;
  assign n17060 = n17034 ^ n14025 ;
  assign n17061 = n17060 ^ n16972 ;
  assign n17062 = n17032 ^ n14572 ;
  assign n17063 = n16975 ^ n14468 ;
  assign n17064 = n17063 ^ n17020 ;
  assign n17065 = n17017 ^ n16977 ;
  assign n17066 = n16978 ^ n14383 ;
  assign n17067 = n17066 ^ n17013 ;
  assign n17068 = n17006 ^ n13725 ;
  assign n17069 = n16981 ^ n14447 ;
  assign n17070 = n17069 ^ n16999 ;
  assign n16780 = n16779 ^ n16769 ;
  assign n16605 = n16604 ^ n14333 ;
  assign n16658 = n16657 ^ n16605 ;
  assign n16675 = n16673 & ~n16674 ;
  assign n16676 = n16651 ^ n16609 ;
  assign n16677 = n16675 & n16676 ;
  assign n16678 = n16654 ^ n16607 ;
  assign n16679 = ~n16677 & ~n16678 ;
  assign n16680 = n16658 & ~n16679 ;
  assign n16695 = n16694 ^ n16684 ;
  assign n16781 = ~n16680 & n16695 ;
  assign n17071 = n16780 & ~n16781 ;
  assign n17072 = n16990 ^ n16987 ;
  assign n17073 = n17071 & n17072 ;
  assign n17074 = n16993 ^ n14408 ;
  assign n17075 = n17074 ^ n16984 ;
  assign n17076 = n17073 & n17075 ;
  assign n17077 = n16996 ^ n16983 ;
  assign n17078 = n17076 & ~n17077 ;
  assign n17079 = n17070 & ~n17078 ;
  assign n17080 = n17068 & n17079 ;
  assign n17081 = n17011 ^ n14389 ;
  assign n17082 = ~n17080 & ~n17081 ;
  assign n17083 = n17067 & n17082 ;
  assign n17084 = ~n17065 & ~n17083 ;
  assign n17085 = ~n17064 & ~n17084 ;
  assign n17086 = n17026 ^ n14472 ;
  assign n17087 = n17086 ^ n17024 ;
  assign n17088 = n17085 & ~n17087 ;
  assign n17089 = n17062 & ~n17088 ;
  assign n17090 = n17061 & ~n17089 ;
  assign n17091 = n17040 ^ n14020 ;
  assign n17092 = n17090 & ~n17091 ;
  assign n17093 = n17044 ^ n17043 ;
  assign n17094 = n17092 & ~n17093 ;
  assign n17095 = n17048 ^ n14009 ;
  assign n17096 = n17095 ^ n17047 ;
  assign n17097 = ~n17094 & ~n17096 ;
  assign n17112 = n17098 ^ n17097 ;
  assign n17113 = n17112 ^ n2694 ;
  assign n17114 = n17096 ^ n17094 ;
  assign n17115 = n17114 ^ n2450 ;
  assign n17116 = n17093 ^ n17092 ;
  assign n17117 = n17116 ^ n2496 ;
  assign n17177 = n17089 ^ n17061 ;
  assign n17119 = n17088 ^ n17062 ;
  assign n2864 = n2821 ^ x264 ;
  assign n2865 = n2864 ^ x456 ;
  assign n2866 = n2865 ^ x200 ;
  assign n17120 = n17119 ^ n2866 ;
  assign n17121 = n17087 ^ n17085 ;
  assign n17122 = n17121 ^ n2810 ;
  assign n17123 = n17082 ^ n17067 ;
  assign n17124 = n17123 ^ n1148 ;
  assign n17125 = n17081 ^ n17080 ;
  assign n966 = n896 ^ x269 ;
  assign n967 = n966 ^ x461 ;
  assign n968 = n967 ^ x205 ;
  assign n17126 = n17125 ^ n968 ;
  assign n17127 = n17079 ^ n17068 ;
  assign n17128 = n17127 ^ n971 ;
  assign n17151 = n17127 ^ n851 ;
  assign n17129 = n17078 ^ n17070 ;
  assign n17130 = n17129 ^ n851 ;
  assign n17131 = n17077 ^ n17076 ;
  assign n17132 = n17131 ^ n768 ;
  assign n17133 = n17075 ^ n17073 ;
  assign n17134 = n17133 ^ n756 ;
  assign n17135 = n17072 ^ n17071 ;
  assign n17136 = n17135 ^ n750 ;
  assign n16782 = n16781 ^ n16780 ;
  assign n16783 = n16782 ^ n1547 ;
  assign n16696 = n16695 ^ n16680 ;
  assign n16697 = n16696 ^ n1541 ;
  assign n16698 = n16679 ^ n16658 ;
  assign n16699 = n16698 ^ n521 ;
  assign n16702 = n16678 ^ n16677 ;
  assign n16703 = n16702 ^ n2929 ;
  assign n16704 = n16676 ^ n16675 ;
  assign n16705 = n16704 ^ n572 ;
  assign n16712 = n16711 ^ n16708 ;
  assign n16755 = n16712 & ~n16754 ;
  assign n16756 = n16755 ^ n16711 ;
  assign n16706 = n16702 ^ n572 ;
  assign n16707 = n16706 ^ n16702 ;
  assign n16757 = n16756 ^ n16707 ;
  assign n16758 = ~n16705 & n16757 ;
  assign n16759 = n16758 ^ n16706 ;
  assign n16760 = n16703 & ~n16759 ;
  assign n16761 = n16760 ^ n2929 ;
  assign n16700 = n16696 ^ n521 ;
  assign n16701 = n16700 ^ n16696 ;
  assign n16762 = n16761 ^ n16701 ;
  assign n16763 = n16699 & n16762 ;
  assign n16764 = n16763 ^ n16700 ;
  assign n16765 = ~n16697 & n16764 ;
  assign n16766 = n16765 ^ n1541 ;
  assign n17137 = n16766 ^ n1547 ;
  assign n17138 = n16783 & ~n17137 ;
  assign n17139 = n17138 ^ n16782 ;
  assign n17140 = n17139 ^ n750 ;
  assign n17141 = ~n17136 & ~n17140 ;
  assign n17142 = n17141 ^ n17135 ;
  assign n17143 = n17142 ^ n756 ;
  assign n17144 = ~n17134 & ~n17143 ;
  assign n17145 = n17144 ^ n756 ;
  assign n17146 = n17145 ^ n768 ;
  assign n17147 = n17132 & ~n17146 ;
  assign n17148 = n17147 ^ n17131 ;
  assign n17149 = n17148 ^ n851 ;
  assign n17150 = ~n17130 & n17149 ;
  assign n17152 = n17151 ^ n17150 ;
  assign n17153 = n17128 & ~n17152 ;
  assign n17154 = n17153 ^ n971 ;
  assign n17155 = n17154 ^ n17125 ;
  assign n17156 = ~n17126 & n17155 ;
  assign n17157 = n17156 ^ n968 ;
  assign n17158 = n17157 ^ n17123 ;
  assign n17159 = ~n17124 & n17158 ;
  assign n17160 = n17159 ^ n1148 ;
  assign n17161 = n17160 ^ n1409 ;
  assign n17162 = n17083 ^ n17065 ;
  assign n17163 = n17162 ^ n17160 ;
  assign n17164 = n17161 & ~n17163 ;
  assign n17165 = n17164 ^ n1409 ;
  assign n17166 = n17165 ^ n1382 ;
  assign n17167 = n17084 ^ n17064 ;
  assign n17168 = n17167 ^ n17165 ;
  assign n17169 = n17166 & n17168 ;
  assign n17170 = n17169 ^ n1382 ;
  assign n17171 = n17170 ^ n17121 ;
  assign n17172 = n17122 & ~n17171 ;
  assign n17173 = n17172 ^ n2810 ;
  assign n17174 = n17173 ^ n17119 ;
  assign n17175 = ~n17120 & n17174 ;
  assign n17176 = n17175 ^ n2866 ;
  assign n17178 = n17177 ^ n17176 ;
  assign n2573 = n2563 ^ x263 ;
  assign n2574 = n2573 ^ x455 ;
  assign n2575 = n2574 ^ x199 ;
  assign n17179 = n17177 ^ n2575 ;
  assign n17180 = ~n17178 & n17179 ;
  assign n17181 = n17180 ^ n2575 ;
  assign n17118 = n17091 ^ n17090 ;
  assign n17182 = n17181 ^ n17118 ;
  assign n17802 = n17118 ^ n2581 ;
  assign n17186 = ~n17182 & n17802 ;
  assign n17183 = n2581 ^ n2496 ;
  assign n17187 = n17186 ^ n17183 ;
  assign n17188 = n17117 & n17187 ;
  assign n17189 = n17188 ^ n2496 ;
  assign n17190 = n17189 ^ n17114 ;
  assign n17191 = n17115 & ~n17190 ;
  assign n17192 = n17191 ^ n2450 ;
  assign n17193 = n17192 ^ n17112 ;
  assign n17194 = n17113 & ~n17193 ;
  assign n17195 = n17194 ^ n2694 ;
  assign n17099 = ~n17097 & n17098 ;
  assign n16963 = n16962 ^ n16856 ;
  assign n16964 = ~n16857 & n16963 ;
  assign n16965 = n16964 ^ n16962 ;
  assign n16851 = n16465 ^ n2480 ;
  assign n16852 = n16851 ^ n16500 ;
  assign n16849 = n15948 ^ n14377 ;
  assign n16850 = n16849 ^ n14962 ;
  assign n16853 = n16852 ^ n16850 ;
  assign n17057 = n16965 ^ n16853 ;
  assign n17058 = n17057 ^ n13760 ;
  assign n16969 = n16968 ^ n14004 ;
  assign n17055 = n16969 & n17054 ;
  assign n17056 = n17055 ^ n14004 ;
  assign n17059 = n17058 ^ n17056 ;
  assign n17110 = n17099 ^ n17059 ;
  assign n17111 = n17110 ^ n1811 ;
  assign n17205 = n17195 ^ n17111 ;
  assign n17203 = n15689 ^ n14939 ;
  assign n17204 = n17203 ^ n16259 ;
  assign n17206 = n17205 ^ n17204 ;
  assign n17208 = n16266 ^ n15693 ;
  assign n17209 = n17208 ^ n14945 ;
  assign n17224 = n17209 ^ n17204 ;
  assign n17207 = n17192 ^ n17113 ;
  assign n17210 = n17209 ^ n17207 ;
  assign n17213 = n16275 ^ n15701 ;
  assign n17214 = n17213 ^ n14954 ;
  assign n17215 = n17187 ^ n17116 ;
  assign n17216 = n17214 & n17215 ;
  assign n17211 = n15699 ^ n14952 ;
  assign n17212 = n17211 ^ n16270 ;
  assign n17217 = n17216 ^ n17212 ;
  assign n17218 = n17189 ^ n17115 ;
  assign n17219 = n17218 ^ n17212 ;
  assign n17220 = n17217 & ~n17219 ;
  assign n17221 = n17220 ^ n17216 ;
  assign n17222 = n17221 ^ n17207 ;
  assign n17223 = n17210 & ~n17222 ;
  assign n17225 = n17224 ^ n17223 ;
  assign n17226 = ~n17206 & n17225 ;
  assign n17227 = n17226 ^ n17205 ;
  assign n17199 = n17057 ^ n17056 ;
  assign n17200 = n17058 & n17199 ;
  assign n17196 = n17195 ^ n17110 ;
  assign n17197 = n17111 & ~n17196 ;
  assign n17102 = n16525 ^ n1802 ;
  assign n17103 = n17102 ^ n15944 ;
  assign n17104 = n17103 ^ n14958 ;
  assign n17101 = n16506 ^ n3133 ;
  assign n17105 = n17104 ^ n17101 ;
  assign n17106 = n17105 ^ n1811 ;
  assign n17107 = n17106 ^ n13760 ;
  assign n17108 = n17107 ^ n16850 ;
  assign n17100 = ~n17059 & n17099 ;
  assign n17109 = n17108 ^ n17100 ;
  assign n17198 = n17197 ^ n17109 ;
  assign n17201 = n17200 ^ n17198 ;
  assign n16966 = n16965 ^ n16850 ;
  assign n16967 = ~n16853 & n16966 ;
  assign n17202 = n17201 ^ n16967 ;
  assign n17228 = n17227 ^ n17202 ;
  assign n17229 = n15685 ^ n14937 ;
  assign n17230 = n17229 ^ n16263 ;
  assign n17231 = n17230 ^ n17227 ;
  assign n17232 = ~n17228 & n17231 ;
  assign n17233 = n17232 ^ n17230 ;
  assign n16845 = n15682 ^ n14927 ;
  assign n16846 = n16845 ^ n16594 ;
  assign n16847 = n16846 ^ n16841 ;
  assign n16848 = n16847 ^ n16846 ;
  assign n17234 = n17233 ^ n16848 ;
  assign n17235 = n16844 & ~n17234 ;
  assign n17236 = n17235 ^ n16847 ;
  assign n17238 = n16732 ^ n16731 ;
  assign n17239 = n17238 ^ n16839 ;
  assign n17237 = n16846 ^ n16839 ;
  assign n17240 = n17239 ^ n17237 ;
  assign n17241 = ~n17236 & n17240 ;
  assign n17242 = n17241 ^ n17237 ;
  assign n17243 = ~n16840 & ~n17242 ;
  assign n17244 = n17243 ^ n16839 ;
  assign n17245 = n17244 ^ n16834 ;
  assign n17246 = n16836 & n17245 ;
  assign n17247 = n17246 ^ n16835 ;
  assign n16828 = n16231 ^ n14900 ;
  assign n16830 = n16829 ^ n16828 ;
  assign n16831 = n16830 ^ n16826 ;
  assign n16832 = n16831 ^ n16830 ;
  assign n17248 = n17247 ^ n16832 ;
  assign n17249 = n16827 & ~n17248 ;
  assign n17250 = n17249 ^ n16831 ;
  assign n17252 = n17251 ^ n16830 ;
  assign n17253 = n17250 & ~n17252 ;
  assign n17255 = n17254 ^ n17253 ;
  assign n17256 = ~n16822 & n17255 ;
  assign n17257 = n17256 ^ n16821 ;
  assign n17258 = n17257 ^ n16814 ;
  assign n17259 = ~n16816 & n17258 ;
  assign n17260 = n17259 ^ n16815 ;
  assign n17261 = n17260 ^ n16809 ;
  assign n17262 = ~n16811 & ~n17261 ;
  assign n17263 = n17262 ^ n16810 ;
  assign n16800 = n16756 ^ n16705 ;
  assign n16797 = n16300 ^ n15724 ;
  assign n16799 = n16798 ^ n16797 ;
  assign n16801 = n16800 ^ n16799 ;
  assign n17294 = n17263 ^ n16801 ;
  assign n17295 = n17294 ^ n14907 ;
  assign n17296 = n17260 ^ n16811 ;
  assign n17297 = n17296 ^ n14914 ;
  assign n17358 = n17257 ^ n16816 ;
  assign n17298 = n17255 ^ n16820 ;
  assign n17299 = n17298 ^ n14925 ;
  assign n17300 = n17251 ^ n17250 ;
  assign n17301 = n17300 ^ n14930 ;
  assign n17303 = n17244 ^ n16836 ;
  assign n17304 = n17303 ^ n14942 ;
  assign n17306 = n17230 ^ n17202 ;
  assign n17307 = n17306 ^ n17227 ;
  assign n17308 = n17307 ^ n14356 ;
  assign n17317 = n17221 ^ n17210 ;
  assign n17310 = n17215 ^ n17214 ;
  assign n17311 = ~n14696 & n17310 ;
  assign n17312 = n17311 ^ n14700 ;
  assign n17313 = n17218 ^ n17217 ;
  assign n17314 = n17313 ^ n17311 ;
  assign n17315 = n17312 & ~n17314 ;
  assign n17316 = n17315 ^ n14700 ;
  assign n17318 = n17317 ^ n17316 ;
  assign n17319 = n17317 ^ n14364 ;
  assign n17320 = ~n17318 & ~n17319 ;
  assign n17321 = n17320 ^ n14364 ;
  assign n17309 = n17225 ^ n17205 ;
  assign n17322 = n17321 ^ n17309 ;
  assign n17323 = n17307 ^ n14358 ;
  assign n17324 = n17323 ^ n17307 ;
  assign n17325 = n17324 ^ n17309 ;
  assign n17326 = ~n17322 & ~n17325 ;
  assign n17327 = n17326 ^ n17323 ;
  assign n17328 = n17308 & ~n17327 ;
  assign n17329 = n17328 ^ n14356 ;
  assign n17330 = n17329 ^ n14718 ;
  assign n17331 = n17233 ^ n16844 ;
  assign n17332 = n17331 ^ n17329 ;
  assign n17333 = ~n17330 & ~n17332 ;
  assign n17334 = n17333 ^ n14718 ;
  assign n17335 = n17334 ^ n14891 ;
  assign n17336 = n17238 ^ n17236 ;
  assign n17337 = n17336 ^ n17334 ;
  assign n17338 = n17335 & ~n17337 ;
  assign n17339 = n17338 ^ n14891 ;
  assign n17305 = n17242 ^ n16837 ;
  assign n17340 = n17339 ^ n17305 ;
  assign n17341 = n17339 ^ n14947 ;
  assign n17342 = ~n17340 & ~n17341 ;
  assign n17343 = n17342 ^ n14947 ;
  assign n17344 = n17343 ^ n17303 ;
  assign n17345 = n17304 & n17344 ;
  assign n17346 = n17345 ^ n14942 ;
  assign n17302 = n17247 ^ n16827 ;
  assign n17347 = n17346 ^ n17302 ;
  assign n17348 = n17300 ^ n14935 ;
  assign n17349 = n17348 ^ n17300 ;
  assign n17350 = n17349 ^ n17302 ;
  assign n17351 = n17347 & ~n17350 ;
  assign n17352 = n17351 ^ n17348 ;
  assign n17353 = n17301 & n17352 ;
  assign n17354 = n17353 ^ n14930 ;
  assign n17355 = n17354 ^ n17298 ;
  assign n17356 = ~n17299 & ~n17355 ;
  assign n17357 = n17356 ^ n14925 ;
  assign n17359 = n17358 ^ n17357 ;
  assign n17360 = n17358 ^ n14917 ;
  assign n17361 = n17359 & ~n17360 ;
  assign n17362 = n17361 ^ n14917 ;
  assign n17363 = n17362 ^ n17296 ;
  assign n17364 = n17297 & n17363 ;
  assign n17365 = n17364 ^ n14914 ;
  assign n17366 = n17365 ^ n17294 ;
  assign n17367 = ~n17295 & ~n17366 ;
  assign n17368 = n17367 ^ n14907 ;
  assign n17415 = n17368 ^ n14903 ;
  assign n17270 = n16759 ^ n2929 ;
  assign n16802 = n16295 ^ n15717 ;
  assign n16804 = n16803 ^ n16802 ;
  assign n16805 = n16804 ^ n16800 ;
  assign n16806 = n16805 ^ n16804 ;
  assign n17264 = n17263 ^ n16806 ;
  assign n17265 = n16801 & ~n17264 ;
  assign n17266 = n17265 ^ n16805 ;
  assign n17369 = n17270 ^ n17266 ;
  assign n17416 = n17415 ^ n17369 ;
  assign n17417 = n17362 ^ n17297 ;
  assign n17418 = n17354 ^ n17299 ;
  assign n17419 = n17305 ^ n14947 ;
  assign n17420 = n17419 ^ n17339 ;
  assign n17421 = n17336 ^ n17335 ;
  assign n17422 = n17331 ^ n17330 ;
  assign n17423 = n17310 ^ n14696 ;
  assign n17424 = n17313 ^ n17312 ;
  assign n17425 = ~n17423 & n17424 ;
  assign n17426 = n17319 ^ n17316 ;
  assign n17427 = n17425 & ~n17426 ;
  assign n17428 = n17309 ^ n14358 ;
  assign n17429 = n17428 ^ n17321 ;
  assign n17430 = n17427 & n17429 ;
  assign n17431 = n17327 ^ n14356 ;
  assign n17432 = n17430 & n17431 ;
  assign n17433 = n17422 & ~n17432 ;
  assign n17434 = ~n17421 & ~n17433 ;
  assign n17435 = ~n17420 & ~n17434 ;
  assign n17436 = n17343 ^ n17304 ;
  assign n17437 = n17435 & ~n17436 ;
  assign n17438 = n17302 ^ n14935 ;
  assign n17439 = n17438 ^ n17346 ;
  assign n17440 = n17437 & ~n17439 ;
  assign n17441 = n17352 ^ n14930 ;
  assign n17442 = ~n17440 & ~n17441 ;
  assign n17443 = n17418 & ~n17442 ;
  assign n17444 = n17360 ^ n17357 ;
  assign n17445 = ~n17443 & n17444 ;
  assign n17446 = n17417 & ~n17445 ;
  assign n17447 = n17365 ^ n17295 ;
  assign n17448 = n17446 & n17447 ;
  assign n17449 = ~n17416 & n17448 ;
  assign n17370 = n17369 ^ n17368 ;
  assign n17371 = n17369 ^ n14903 ;
  assign n17372 = ~n17370 & ~n17371 ;
  assign n17373 = n17372 ^ n14903 ;
  assign n17413 = n17373 ^ n14351 ;
  assign n17276 = n16761 ^ n16699 ;
  assign n17267 = n16293 ^ n15719 ;
  assign n17268 = n17267 ^ n16876 ;
  assign n17271 = n17270 ^ n17268 ;
  assign n17269 = n17268 ^ n16804 ;
  assign n17272 = n17271 ^ n17269 ;
  assign n17273 = n17266 & n17272 ;
  assign n17274 = n17273 ^ n17271 ;
  assign n17292 = n17276 ^ n17274 ;
  assign n17414 = n17413 ^ n17292 ;
  assign n17466 = n17449 ^ n17414 ;
  assign n17550 = n17466 ^ n937 ;
  assign n17467 = n17448 ^ n17416 ;
  assign n17468 = n17467 ^ n683 ;
  assign n17470 = n17445 ^ n17417 ;
  assign n17471 = n17470 ^ n540 ;
  assign n17472 = n17444 ^ n17443 ;
  assign n17473 = n17472 ^ n551 ;
  assign n17475 = n17442 ^ n17418 ;
  assign n17476 = n17475 ^ n604 ;
  assign n17477 = n17441 ^ n17440 ;
  assign n17481 = n17480 ^ n17477 ;
  assign n17484 = n17439 ^ n17437 ;
  assign n17529 = n17484 ^ n17477 ;
  assign n17482 = n17436 ^ n17435 ;
  assign n17483 = n17482 ^ n2436 ;
  assign n17488 = n17433 ^ n17421 ;
  assign n2202 = n2135 ^ x314 ;
  assign n2203 = n2202 ^ x506 ;
  assign n2204 = n2203 ^ x250 ;
  assign n17489 = n17488 ^ n2204 ;
  assign n17511 = n17432 ^ n17422 ;
  assign n17490 = n17431 ^ n17430 ;
  assign n2077 = n2019 ^ x316 ;
  assign n2078 = n2077 ^ x508 ;
  assign n2079 = n2078 ^ x252 ;
  assign n17491 = n17490 ^ n2079 ;
  assign n17492 = n17429 ^ n17427 ;
  assign n1985 = n1942 ^ x317 ;
  assign n1986 = n1985 ^ x509 ;
  assign n1987 = n1986 ^ x253 ;
  assign n17493 = n17492 ^ n1987 ;
  assign n17494 = n17426 ^ n17425 ;
  assign n1979 = n1936 ^ x318 ;
  assign n1980 = n1979 ^ x510 ;
  assign n1981 = n1980 ^ x254 ;
  assign n17495 = n17494 ^ n1981 ;
  assign n17497 = n17424 ^ n17423 ;
  assign n17501 = n17497 ^ n1981 ;
  assign n17496 = n1916 & n17423 ;
  assign n17498 = n17497 ^ n17496 ;
  assign n1920 = n1889 ^ x319 ;
  assign n1921 = n1920 ^ x511 ;
  assign n1922 = n1921 ^ x255 ;
  assign n17499 = n17496 ^ n1922 ;
  assign n17500 = ~n17498 & ~n17499 ;
  assign n17502 = n17501 ^ n17500 ;
  assign n17503 = ~n17495 & n17502 ;
  assign n17504 = n17503 ^ n17494 ;
  assign n17505 = n17504 ^ n1987 ;
  assign n17506 = n17493 & n17505 ;
  assign n17507 = n17506 ^ n17492 ;
  assign n17508 = n17507 ^ n2079 ;
  assign n17509 = n17491 & n17508 ;
  assign n17510 = n17509 ^ n2079 ;
  assign n17512 = n17511 ^ n17510 ;
  assign n17515 = n17510 ^ n2406 ;
  assign n17516 = ~n17512 & n17515 ;
  assign n17513 = n2406 ^ n2204 ;
  assign n17517 = n17516 ^ n17513 ;
  assign n17518 = n17489 & n17517 ;
  assign n17519 = n17518 ^ n2204 ;
  assign n17487 = n17434 ^ n17420 ;
  assign n17520 = n17519 ^ n17487 ;
  assign n17521 = n17519 ^ n2420 ;
  assign n17522 = n17520 & n17521 ;
  assign n17523 = n17522 ^ n2420 ;
  assign n17485 = n17484 ^ n2436 ;
  assign n17486 = n17485 ^ n17484 ;
  assign n17524 = n17523 ^ n17486 ;
  assign n17525 = n17483 & n17524 ;
  assign n17526 = n17525 ^ n17485 ;
  assign n17527 = n17484 ^ n1473 ;
  assign n17528 = n17526 & n17527 ;
  assign n17530 = n17529 ^ n17528 ;
  assign n17531 = n17481 & ~n17530 ;
  assign n17532 = n17531 ^ n17480 ;
  assign n17533 = n17532 ^ n17475 ;
  assign n17534 = n17476 & ~n17533 ;
  assign n17535 = n17534 ^ n604 ;
  assign n17474 = n551 ^ n540 ;
  assign n17536 = n17535 ^ n17474 ;
  assign n17537 = n17536 ^ n540 ;
  assign n17538 = ~n17473 & n17537 ;
  assign n17539 = n17538 ^ n17474 ;
  assign n17540 = n17471 & n17539 ;
  assign n17541 = n17540 ^ n540 ;
  assign n17545 = n17541 ^ n17467 ;
  assign n17469 = n17447 ^ n17446 ;
  assign n17542 = n17541 ^ n17469 ;
  assign n17543 = n17469 ^ n1602 ;
  assign n17544 = ~n17542 & n17543 ;
  assign n17546 = n17545 ^ n17544 ;
  assign n17547 = n17468 & ~n17546 ;
  assign n17548 = n17547 ^ n683 ;
  assign n18237 = n17550 ^ n17548 ;
  assign n17612 = n17507 ^ n17491 ;
  assign n17605 = n16813 ^ n16231 ;
  assign n17606 = n17605 ^ n17270 ;
  assign n17857 = n17612 ^ n17606 ;
  assign n17610 = n16819 ^ n16126 ;
  assign n17611 = n17610 ^ n16800 ;
  assign n17613 = n17612 ^ n17611 ;
  assign n17616 = n17504 ^ n17493 ;
  assign n17614 = n16829 ^ n16111 ;
  assign n17615 = n17614 ^ n16810 ;
  assign n17617 = n17616 ^ n17615 ;
  assign n17620 = n17502 ^ n17494 ;
  assign n17618 = n16824 ^ n16070 ;
  assign n17619 = n17618 ^ n16815 ;
  assign n17621 = n17620 ^ n17619 ;
  assign n17624 = n17499 ^ n17497 ;
  assign n17622 = n16770 ^ n15682 ;
  assign n17623 = n17622 ^ n16821 ;
  assign n17625 = n17624 ^ n17623 ;
  assign n17628 = n17423 ^ n1916 ;
  assign n17626 = n16685 ^ n15678 ;
  assign n17627 = n17626 ^ n17251 ;
  assign n17629 = n17628 ^ n17627 ;
  assign n17812 = n16594 ^ n15685 ;
  assign n17813 = n17812 ^ n16826 ;
  assign n17842 = n17813 ^ n17627 ;
  assign n17809 = n3028 ^ n2736 ;
  assign n17806 = n14377 ^ n14375 ;
  assign n17803 = n17802 ^ n17181 ;
  assign n17799 = n15707 ^ n14958 ;
  assign n17721 = n15711 ^ n14962 ;
  assign n17722 = n17721 ^ n16547 ;
  assign n17800 = n17799 ^ n17722 ;
  assign n17801 = n17800 ^ n16543 ;
  assign n17804 = n17803 ^ n17801 ;
  assign n17725 = n17179 ^ n17176 ;
  assign n17588 = n17173 ^ n2866 ;
  assign n17589 = n17588 ^ n17119 ;
  assign n17726 = n17725 ^ n17589 ;
  assign n17677 = n15944 ^ n15367 ;
  assign n17678 = n17677 ^ n16550 ;
  assign n17632 = n17170 ^ n17122 ;
  assign n17630 = n15948 ^ n15339 ;
  assign n17631 = n17630 ^ n16563 ;
  assign n17633 = n17632 ^ n17631 ;
  assign n17636 = n17167 ^ n17166 ;
  assign n17634 = n15952 ^ n15309 ;
  assign n17635 = n17634 ^ n16560 ;
  assign n17637 = n17636 ^ n17635 ;
  assign n17640 = n17162 ^ n17161 ;
  assign n17670 = n17640 ^ n17636 ;
  assign n17638 = n15961 ^ n15312 ;
  assign n17639 = n17638 ^ n17101 ;
  assign n17641 = n17640 ^ n17639 ;
  assign n17644 = n17157 ^ n1148 ;
  assign n17645 = n17644 ^ n17123 ;
  assign n17642 = n16852 ^ n15956 ;
  assign n17643 = n17642 ^ n15260 ;
  assign n17646 = n17645 ^ n17643 ;
  assign n17649 = n16528 ^ n15870 ;
  assign n17650 = n17649 ^ n16856 ;
  assign n17647 = n17154 ^ n17126 ;
  assign n17651 = n17650 ^ n17647 ;
  assign n17653 = n16422 ^ n15836 ;
  assign n17654 = n17653 ^ n16858 ;
  assign n17652 = n17152 ^ n971 ;
  assign n17655 = n17654 ^ n17652 ;
  assign n17579 = n16353 ^ n15821 ;
  assign n17580 = n17579 ^ n16956 ;
  assign n17578 = n17148 ^ n17130 ;
  assign n17581 = n17580 ^ n17578 ;
  assign n17403 = n16347 ^ n15770 ;
  assign n17404 = n17403 ^ n16949 ;
  assign n17388 = n16339 ^ n15762 ;
  assign n17389 = n17388 ^ n16862 ;
  assign n17405 = n17404 ^ n17389 ;
  assign n16784 = n16783 ^ n16766 ;
  assign n15677 = n15676 ^ n15675 ;
  assign n16258 = n16257 ^ n15677 ;
  assign n16785 = n16784 ^ n16258 ;
  assign n16795 = n16764 ^ n1541 ;
  assign n16791 = n16287 ^ n15738 ;
  assign n16794 = n16793 ^ n16791 ;
  assign n16796 = n16795 ^ n16794 ;
  assign n17277 = n17276 ^ n16794 ;
  assign n17275 = n17268 ^ n16794 ;
  assign n17278 = n17277 ^ n17275 ;
  assign n17279 = ~n17274 & n17278 ;
  assign n17280 = n17279 ^ n17277 ;
  assign n17281 = n16796 & n17280 ;
  assign n17282 = n17281 ^ n16795 ;
  assign n16786 = n16284 ^ n15752 ;
  assign n16788 = n16787 ^ n16786 ;
  assign n16789 = n16788 ^ n16784 ;
  assign n16790 = n16789 ^ n16788 ;
  assign n17283 = n17282 ^ n16790 ;
  assign n17284 = ~n16785 & ~n17283 ;
  assign n17285 = n17284 ^ n16789 ;
  assign n17286 = n17139 ^ n17136 ;
  assign n17391 = n17389 ^ n17286 ;
  assign n17390 = n17389 ^ n16788 ;
  assign n17392 = n17391 ^ n17390 ;
  assign n17393 = n17285 & ~n17392 ;
  assign n17394 = n17393 ^ n17390 ;
  assign n17395 = n17142 ^ n17134 ;
  assign n17401 = n17395 ^ n17389 ;
  assign n17402 = ~n17394 & ~n17401 ;
  assign n17406 = n17405 ^ n17402 ;
  assign n17407 = n17145 ^ n17132 ;
  assign n17575 = n17407 ^ n17404 ;
  assign n17576 = n17406 & ~n17575 ;
  assign n17577 = n17576 ^ n17404 ;
  assign n17658 = n17578 ^ n17577 ;
  assign n17659 = ~n17581 & ~n17658 ;
  assign n17660 = n17659 ^ n17580 ;
  assign n17661 = n17660 ^ n17652 ;
  assign n17662 = n17655 & n17661 ;
  assign n17656 = n17652 ^ n17647 ;
  assign n17663 = n17662 ^ n17656 ;
  assign n17664 = ~n17651 & ~n17663 ;
  assign n17648 = n17647 ^ n17643 ;
  assign n17665 = n17664 ^ n17648 ;
  assign n17666 = n17646 & ~n17665 ;
  assign n17667 = n17666 ^ n17645 ;
  assign n17668 = n17667 ^ n17640 ;
  assign n17669 = n17641 & ~n17668 ;
  assign n17671 = n17670 ^ n17669 ;
  assign n17672 = ~n17637 & ~n17671 ;
  assign n17673 = n17672 ^ n17636 ;
  assign n17674 = n17673 ^ n17631 ;
  assign n17675 = ~n17633 & ~n17674 ;
  assign n17676 = n17675 ^ n17632 ;
  assign n17679 = n17678 ^ n17676 ;
  assign n17723 = n17676 ^ n17589 ;
  assign n17724 = ~n17679 & ~n17723 ;
  assign n17727 = n17726 ^ n17724 ;
  assign n17797 = n17725 ^ n17722 ;
  assign n17798 = n17727 & n17797 ;
  assign n17805 = n17804 ^ n17798 ;
  assign n17807 = n17806 ^ n17805 ;
  assign n17680 = n17679 ^ n17589 ;
  assign n17731 = n17680 ^ n14651 ;
  assign n17681 = n17671 ^ n17635 ;
  assign n17682 = n17681 ^ n14662 ;
  assign n17684 = n17663 ^ n17650 ;
  assign n17685 = n17684 ^ n15357 ;
  assign n17686 = n17660 ^ n17655 ;
  assign n17687 = n17686 ^ n15318 ;
  assign n17582 = n17581 ^ n17577 ;
  assign n17688 = n17582 ^ n15295 ;
  assign n17408 = n17407 ^ n17406 ;
  assign n17409 = n17408 ^ n15278 ;
  assign n17396 = n17395 ^ n17394 ;
  assign n17287 = n17286 ^ n17285 ;
  assign n17288 = n17287 ^ n15228 ;
  assign n17290 = n17280 ^ n16795 ;
  assign n17291 = n17290 ^ n15099 ;
  assign n17293 = n17292 ^ n14351 ;
  assign n17374 = n17373 ^ n17292 ;
  assign n17375 = ~n17293 & ~n17374 ;
  assign n17376 = n17375 ^ n14351 ;
  assign n17377 = n17376 ^ n17290 ;
  assign n17378 = ~n17291 & n17377 ;
  assign n17379 = n17378 ^ n15099 ;
  assign n17289 = n17282 ^ n16785 ;
  assign n17380 = n17379 ^ n17289 ;
  assign n17381 = n17287 ^ n15144 ;
  assign n17382 = n17381 ^ n17287 ;
  assign n17383 = n17382 ^ n17289 ;
  assign n17384 = n17380 & ~n17383 ;
  assign n17385 = n17384 ^ n17381 ;
  assign n17386 = ~n17288 & ~n17385 ;
  assign n17387 = n17386 ^ n15228 ;
  assign n17397 = n17396 ^ n17387 ;
  assign n17398 = n17396 ^ n15247 ;
  assign n17399 = n17397 & ~n17398 ;
  assign n17400 = n17399 ^ n15247 ;
  assign n17571 = n17408 ^ n17400 ;
  assign n17572 = ~n17409 & ~n17571 ;
  assign n17573 = n17572 ^ n15278 ;
  assign n17689 = n17582 ^ n17573 ;
  assign n17690 = ~n17688 & n17689 ;
  assign n17691 = n17690 ^ n15295 ;
  assign n17692 = n17691 ^ n17686 ;
  assign n17693 = ~n17687 & n17692 ;
  assign n17694 = n17693 ^ n15318 ;
  assign n17695 = n17694 ^ n17684 ;
  assign n17696 = n17685 & ~n17695 ;
  assign n17697 = n17696 ^ n15357 ;
  assign n17683 = n17665 ^ n17645 ;
  assign n17698 = n17697 ^ n17683 ;
  assign n17699 = n17667 ^ n17641 ;
  assign n17700 = n17699 ^ n14667 ;
  assign n17701 = n17700 ^ n17683 ;
  assign n17702 = n17701 ^ n17699 ;
  assign n17703 = ~n17698 & n17702 ;
  assign n17704 = n17703 ^ n17700 ;
  assign n17706 = n17681 ^ n14669 ;
  assign n17705 = n17699 ^ n17681 ;
  assign n17707 = n17706 ^ n17705 ;
  assign n17708 = ~n17704 & n17707 ;
  assign n17709 = n17708 ^ n17706 ;
  assign n17710 = ~n17682 & ~n17709 ;
  assign n17711 = n17710 ^ n14662 ;
  assign n17712 = n17711 ^ n14682 ;
  assign n17713 = n17673 ^ n17633 ;
  assign n17714 = n17713 ^ n17711 ;
  assign n17715 = n17712 & ~n17714 ;
  assign n17716 = n17715 ^ n14682 ;
  assign n17732 = n17731 ^ n17716 ;
  assign n17733 = n17713 ^ n17712 ;
  assign n17734 = n17709 ^ n14662 ;
  assign n17574 = n17573 ^ n15295 ;
  assign n17583 = n17582 ^ n17574 ;
  assign n17410 = n17409 ^ n17400 ;
  assign n17411 = n17398 ^ n17387 ;
  assign n17412 = n17385 ^ n15228 ;
  assign n17450 = n17414 & n17449 ;
  assign n17451 = n17376 ^ n17291 ;
  assign n17452 = ~n17450 & n17451 ;
  assign n17453 = n17379 ^ n15144 ;
  assign n17454 = n17453 ^ n17289 ;
  assign n17455 = n17452 & n17454 ;
  assign n17456 = ~n17412 & ~n17455 ;
  assign n17457 = n17411 & n17456 ;
  assign n17584 = ~n17410 & ~n17457 ;
  assign n17735 = ~n17583 & ~n17584 ;
  assign n17736 = n17691 ^ n15318 ;
  assign n17737 = n17736 ^ n17686 ;
  assign n17738 = n17735 & ~n17737 ;
  assign n17739 = n17694 ^ n17685 ;
  assign n17740 = ~n17738 & ~n17739 ;
  assign n17741 = n17683 ^ n14667 ;
  assign n17742 = n17741 ^ n17697 ;
  assign n17743 = ~n17740 & n17742 ;
  assign n17744 = n17704 ^ n14669 ;
  assign n17745 = n17743 & n17744 ;
  assign n17746 = ~n17734 & n17745 ;
  assign n17747 = n17733 & ~n17746 ;
  assign n17748 = ~n17732 & ~n17747 ;
  assign n17728 = n17727 ^ n17722 ;
  assign n17791 = n17748 ^ n17728 ;
  assign n17717 = n17716 ^ n17680 ;
  assign n17718 = n17716 ^ n14651 ;
  assign n17719 = n17717 & ~n17718 ;
  assign n17720 = n17719 ^ n14651 ;
  assign n17794 = n17748 ^ n17720 ;
  assign n17795 = ~n17791 & ~n17794 ;
  assign n17792 = n17791 ^ n17720 ;
  assign n17793 = n14377 & ~n17792 ;
  assign n17796 = n17795 ^ n17793 ;
  assign n17808 = n17807 ^ n17796 ;
  assign n17810 = n17809 ^ n17808 ;
  assign n17729 = n17728 ^ n14377 ;
  assign n17730 = n17729 ^ n17720 ;
  assign n17749 = n17748 ^ n17730 ;
  assign n17750 = n17749 ^ n2736 ;
  assign n17751 = n17747 ^ n17732 ;
  assign n17752 = n17751 ^ n2680 ;
  assign n17753 = n17746 ^ n17733 ;
  assign n17754 = n17753 ^ n2665 ;
  assign n17755 = n17745 ^ n17734 ;
  assign n17756 = n17755 ^ n1835 ;
  assign n17757 = n17744 ^ n17743 ;
  assign n3119 = n3115 ^ x294 ;
  assign n3120 = n3119 ^ x486 ;
  assign n3121 = n3120 ^ x230 ;
  assign n17758 = n17757 ^ n3121 ;
  assign n17759 = n17742 ^ n17740 ;
  assign n17760 = n17759 ^ n3092 ;
  assign n17761 = n17739 ^ n17738 ;
  assign n17762 = n17761 ^ n2507 ;
  assign n17763 = n17737 ^ n17735 ;
  assign n17764 = n17763 ^ n3203 ;
  assign n17585 = n17584 ^ n17583 ;
  assign n17586 = n17585 ^ n2537 ;
  assign n17458 = n17457 ^ n17410 ;
  assign n17459 = n17458 ^ n1235 ;
  assign n17561 = n17456 ^ n17411 ;
  assign n17562 = n17561 ^ n1077 ;
  assign n17460 = n17455 ^ n17412 ;
  assign n17461 = n17460 ^ n1077 ;
  assign n17462 = n17454 ^ n17452 ;
  assign n17463 = n17462 ^ n955 ;
  assign n17464 = n17451 ^ n17450 ;
  assign n17465 = n17464 ^ n943 ;
  assign n17552 = n17548 ^ n943 ;
  assign n17549 = n17548 ^ n17466 ;
  assign n17551 = ~n17549 & n17550 ;
  assign n17553 = n17552 ^ n17551 ;
  assign n17554 = ~n17465 & ~n17553 ;
  assign n17555 = n17554 ^ n17464 ;
  assign n17556 = n17555 ^ n955 ;
  assign n17557 = n17463 & n17556 ;
  assign n17558 = n17557 ^ n17462 ;
  assign n17559 = n17558 ^ n1077 ;
  assign n17560 = ~n17461 & n17559 ;
  assign n17563 = n17562 ^ n17560 ;
  assign n17565 = n1235 ^ n1089 ;
  assign n17564 = n17561 ^ n1235 ;
  assign n17566 = n17565 ^ n17564 ;
  assign n17567 = n17563 & ~n17566 ;
  assign n17568 = n17567 ^ n17565 ;
  assign n17569 = n17459 & n17568 ;
  assign n17570 = n17569 ^ n1235 ;
  assign n17765 = n17585 ^ n17570 ;
  assign n17766 = ~n17586 & n17765 ;
  assign n17767 = n17766 ^ n2537 ;
  assign n17768 = n17767 ^ n17763 ;
  assign n17769 = n17764 & ~n17768 ;
  assign n17770 = n17769 ^ n3203 ;
  assign n17771 = n17770 ^ n17761 ;
  assign n17772 = n17762 & ~n17771 ;
  assign n17773 = n17772 ^ n2507 ;
  assign n17774 = n17773 ^ n17759 ;
  assign n17775 = n17760 & ~n17774 ;
  assign n17776 = n17775 ^ n3092 ;
  assign n17777 = n17776 ^ n17757 ;
  assign n17778 = ~n17758 & n17777 ;
  assign n17779 = n17778 ^ n3121 ;
  assign n17780 = n17779 ^ n17755 ;
  assign n17781 = n17756 & ~n17780 ;
  assign n17782 = n17781 ^ n1835 ;
  assign n17783 = n17782 ^ n17753 ;
  assign n17784 = ~n17754 & n17783 ;
  assign n17785 = n17784 ^ n2665 ;
  assign n17786 = n17785 ^ n17751 ;
  assign n17787 = ~n17752 & n17786 ;
  assign n17788 = n17787 ^ n2680 ;
  assign n17789 = n17788 ^ n2736 ;
  assign n17790 = n17750 & n17789 ;
  assign n17811 = n17810 ^ n17790 ;
  assign n17814 = n17813 ^ n17811 ;
  assign n17817 = n17788 ^ n17750 ;
  assign n17815 = n16586 ^ n15689 ;
  assign n17816 = n17815 ^ n16835 ;
  assign n17818 = n17817 ^ n17816 ;
  assign n17821 = n17785 ^ n17752 ;
  assign n17819 = n16263 ^ n15693 ;
  assign n17820 = n17819 ^ n16837 ;
  assign n17822 = n17821 ^ n17820 ;
  assign n17826 = n17779 ^ n17756 ;
  assign n17827 = n16266 ^ n15701 ;
  assign n17828 = n17827 ^ n16841 ;
  assign n17829 = n17826 & n17828 ;
  assign n17823 = n16259 ^ n15699 ;
  assign n17824 = n17823 ^ n17238 ;
  assign n17830 = n17829 ^ n17824 ;
  assign n17831 = n17782 ^ n17754 ;
  assign n17832 = n17831 ^ n17824 ;
  assign n17833 = n17830 & ~n17832 ;
  assign n17825 = n17824 ^ n17821 ;
  assign n17834 = n17833 ^ n17825 ;
  assign n17835 = ~n17822 & ~n17834 ;
  assign n17836 = n17835 ^ n17821 ;
  assign n17837 = n17836 ^ n17816 ;
  assign n17838 = ~n17818 & ~n17837 ;
  assign n17839 = n17838 ^ n17817 ;
  assign n17840 = n17839 ^ n17811 ;
  assign n17841 = n17814 & ~n17840 ;
  assign n17843 = n17842 ^ n17841 ;
  assign n17844 = n17629 & ~n17843 ;
  assign n17845 = n17844 ^ n17628 ;
  assign n17846 = n17845 ^ n17623 ;
  assign n17847 = ~n17625 & ~n17846 ;
  assign n17848 = n17847 ^ n17624 ;
  assign n17849 = n17848 ^ n17619 ;
  assign n17850 = n17621 & n17849 ;
  assign n17851 = n17850 ^ n17620 ;
  assign n17852 = n17851 ^ n17615 ;
  assign n17853 = n17617 & n17852 ;
  assign n17854 = n17853 ^ n17616 ;
  assign n17855 = n17854 ^ n17612 ;
  assign n17856 = n17613 & ~n17855 ;
  assign n17858 = n17857 ^ n17856 ;
  assign n17607 = n17511 ^ n2406 ;
  assign n17608 = n17607 ^ n17510 ;
  assign n17940 = n17858 ^ n17608 ;
  assign n17942 = n17940 ^ n14900 ;
  assign n17891 = n17854 ^ n17613 ;
  assign n17892 = n17891 ^ n14909 ;
  assign n17894 = n17848 ^ n17621 ;
  assign n17895 = n17894 ^ n14920 ;
  assign n17896 = n17845 ^ n17625 ;
  assign n17897 = n17896 ^ n14927 ;
  assign n17898 = n17839 ^ n17814 ;
  assign n17899 = n17898 ^ n14937 ;
  assign n17901 = n17834 ^ n17820 ;
  assign n17902 = n17901 ^ n14945 ;
  assign n17905 = n17831 ^ n17830 ;
  assign n17903 = n17828 ^ n17826 ;
  assign n17904 = ~n14954 & n17903 ;
  assign n17906 = n17905 ^ n17904 ;
  assign n17907 = n17905 ^ n14952 ;
  assign n17908 = n17906 & n17907 ;
  assign n17909 = n17908 ^ n14952 ;
  assign n17910 = n17909 ^ n17901 ;
  assign n17911 = n17902 & ~n17910 ;
  assign n17912 = n17911 ^ n14945 ;
  assign n17900 = n17836 ^ n17818 ;
  assign n17913 = n17912 ^ n17900 ;
  assign n17914 = n17898 ^ n14939 ;
  assign n17915 = n17914 ^ n17898 ;
  assign n17916 = n17915 ^ n17900 ;
  assign n17917 = n17913 & n17916 ;
  assign n17918 = n17917 ^ n17914 ;
  assign n17919 = ~n17899 & ~n17918 ;
  assign n17920 = n17919 ^ n14937 ;
  assign n17921 = n17920 ^ n14932 ;
  assign n17922 = n17843 ^ n17628 ;
  assign n17923 = n17922 ^ n17920 ;
  assign n17924 = ~n17921 & n17923 ;
  assign n17925 = n17924 ^ n14932 ;
  assign n17926 = n17925 ^ n17896 ;
  assign n17927 = n17897 & n17926 ;
  assign n17928 = n17927 ^ n14927 ;
  assign n17929 = n17928 ^ n17894 ;
  assign n17930 = n17895 & ~n17929 ;
  assign n17931 = n17930 ^ n14920 ;
  assign n17893 = n17851 ^ n17617 ;
  assign n17932 = n17931 ^ n17893 ;
  assign n17933 = n17891 ^ n14911 ;
  assign n17934 = n17933 ^ n17891 ;
  assign n17935 = n17934 ^ n17893 ;
  assign n17936 = n17932 & n17935 ;
  assign n17937 = n17936 ^ n17933 ;
  assign n17938 = ~n17892 & n17937 ;
  assign n17939 = n17938 ^ n14909 ;
  assign n17964 = n17942 ^ n17939 ;
  assign n17965 = n17900 ^ n14939 ;
  assign n17966 = n17965 ^ n17912 ;
  assign n17967 = n17909 ^ n17902 ;
  assign n17968 = n17903 ^ n14954 ;
  assign n17969 = n17904 ^ n14952 ;
  assign n17970 = n17969 ^ n17905 ;
  assign n17971 = ~n17968 & n17970 ;
  assign n17972 = ~n17967 & n17971 ;
  assign n17973 = ~n17966 & n17972 ;
  assign n17974 = n17918 ^ n14937 ;
  assign n17975 = n17973 & ~n17974 ;
  assign n17976 = n17922 ^ n17921 ;
  assign n17977 = ~n17975 & n17976 ;
  assign n17978 = n17925 ^ n17897 ;
  assign n17979 = ~n17977 & n17978 ;
  assign n17980 = n17928 ^ n17895 ;
  assign n17981 = ~n17979 & n17980 ;
  assign n17982 = n17893 ^ n14911 ;
  assign n17983 = n17982 ^ n17931 ;
  assign n17984 = n17981 & n17983 ;
  assign n17985 = n17937 ^ n14909 ;
  assign n17986 = n17984 & n17985 ;
  assign n17987 = ~n17964 & ~n17986 ;
  assign n17941 = n17940 ^ n17939 ;
  assign n17943 = n17941 & ~n17942 ;
  assign n17944 = n17943 ^ n14900 ;
  assign n17609 = n17608 ^ n17606 ;
  assign n17859 = ~n17609 & n17858 ;
  assign n17860 = n17859 ^ n17608 ;
  assign n17602 = n16808 ^ n16246 ;
  assign n17603 = n17602 ^ n17276 ;
  assign n17601 = n17517 ^ n17488 ;
  assign n17604 = n17603 ^ n17601 ;
  assign n17889 = n17860 ^ n17604 ;
  assign n17890 = n17889 ^ n14898 ;
  assign n17988 = n17944 ^ n17890 ;
  assign n17989 = ~n17987 & ~n17988 ;
  assign n17945 = n17944 ^ n17889 ;
  assign n17946 = n17890 & n17945 ;
  assign n17947 = n17946 ^ n14898 ;
  assign n17990 = n17947 ^ n15419 ;
  assign n17861 = n17860 ^ n17601 ;
  assign n17862 = ~n17604 & ~n17861 ;
  assign n17863 = n17862 ^ n17603 ;
  assign n17594 = n16798 ^ n16310 ;
  assign n17595 = n17594 ^ n16795 ;
  assign n17592 = n17487 ^ n2420 ;
  assign n17593 = n17592 ^ n17519 ;
  assign n17596 = n17595 ^ n17593 ;
  assign n17888 = n17863 ^ n17596 ;
  assign n17991 = n17990 ^ n17888 ;
  assign n17992 = ~n17989 & n17991 ;
  assign n17948 = n17947 ^ n17888 ;
  assign n17869 = n17523 ^ n17483 ;
  assign n17597 = n16803 ^ n16304 ;
  assign n17598 = n17597 ^ n16784 ;
  assign n17599 = n17598 ^ n17593 ;
  assign n17600 = n17599 ^ n17598 ;
  assign n17864 = n17863 ^ n17600 ;
  assign n17865 = ~n17596 & n17864 ;
  assign n17866 = n17865 ^ n17599 ;
  assign n17886 = n17869 ^ n17866 ;
  assign n17949 = n17886 ^ n15419 ;
  assign n17950 = n17949 ^ n17886 ;
  assign n17951 = n17950 ^ n17888 ;
  assign n17952 = n17948 & ~n17951 ;
  assign n17953 = n17952 ^ n17949 ;
  assign n17963 = n17953 ^ n15526 ;
  assign n18018 = n17992 ^ n17963 ;
  assign n18087 = n18018 ^ n671 ;
  assign n18016 = n17991 ^ n17989 ;
  assign n18017 = n18016 ^ n1516 ;
  assign n18021 = n17988 ^ n17987 ;
  assign n18022 = n18021 ^ n1507 ;
  assign n18024 = n17985 ^ n17984 ;
  assign n18028 = n18027 ^ n18024 ;
  assign n18029 = n17983 ^ n17981 ;
  assign n18030 = n18029 ^ n587 ;
  assign n18031 = n17980 ^ n17979 ;
  assign n18032 = n18031 ^ n2296 ;
  assign n18065 = n18031 ^ n2286 ;
  assign n18033 = n17976 ^ n17975 ;
  assign n18034 = n18033 ^ n2159 ;
  assign n18037 = n17974 ^ n17973 ;
  assign n18038 = n18037 ^ n2070 ;
  assign n18039 = n17972 ^ n17966 ;
  assign n18040 = n18039 ^ n2055 ;
  assign n3085 = n3051 ^ x351 ;
  assign n3086 = n3085 ^ n1871 ;
  assign n3087 = n3086 ^ x287 ;
  assign n2043 = n1994 ^ x350 ;
  assign n2047 = n2046 ^ n2043 ;
  assign n2048 = n2047 ^ x286 ;
  assign n18046 = n3087 ^ n2048 ;
  assign n18041 = n17970 ^ n17968 ;
  assign n18042 = n18041 ^ n3087 ;
  assign n3065 = n3037 ^ x320 ;
  assign n3069 = n3068 ^ n3065 ;
  assign n3070 = n3069 ^ x256 ;
  assign n18043 = n3070 & n17968 ;
  assign n18044 = n18043 ^ n18041 ;
  assign n18045 = ~n18042 & n18044 ;
  assign n18047 = n18046 ^ n18045 ;
  assign n18050 = n2055 ^ n2048 ;
  assign n18048 = n17971 ^ n17967 ;
  assign n18049 = n18048 ^ n2055 ;
  assign n18051 = n18050 ^ n18049 ;
  assign n18052 = n18047 & ~n18051 ;
  assign n18053 = n18052 ^ n18050 ;
  assign n18054 = ~n18040 & ~n18053 ;
  assign n18055 = n18054 ^ n18039 ;
  assign n18056 = n18055 ^ n18037 ;
  assign n18057 = ~n18038 & ~n18056 ;
  assign n18058 = n18057 ^ n2070 ;
  assign n18035 = n2286 ^ n2159 ;
  assign n18036 = n18035 ^ n2286 ;
  assign n18059 = n18058 ^ n18036 ;
  assign n18060 = n18034 & n18059 ;
  assign n18061 = n18060 ^ n18035 ;
  assign n18062 = n17978 ^ n17977 ;
  assign n18063 = n18062 ^ n2286 ;
  assign n18064 = n18061 & ~n18063 ;
  assign n18066 = n18065 ^ n18064 ;
  assign n18067 = n18032 & ~n18066 ;
  assign n18068 = n18067 ^ n2296 ;
  assign n18069 = n18068 ^ n18029 ;
  assign n18070 = ~n18030 & n18069 ;
  assign n18071 = n18070 ^ n587 ;
  assign n18072 = n18071 ^ n18027 ;
  assign n18073 = ~n18028 & n18072 ;
  assign n18074 = n18073 ^ n18027 ;
  assign n18078 = n18074 ^ n1507 ;
  assign n18023 = n17986 ^ n17964 ;
  assign n18075 = n18074 ^ n18023 ;
  assign n18076 = n18023 ^ n2924 ;
  assign n18077 = n18075 & ~n18076 ;
  assign n18079 = n18078 ^ n18077 ;
  assign n18080 = ~n18022 & n18079 ;
  assign n18081 = n18080 ^ n1507 ;
  assign n18019 = n18018 ^ n1516 ;
  assign n18020 = n18019 ^ n18018 ;
  assign n18082 = n18081 ^ n18020 ;
  assign n18083 = ~n18017 & n18082 ;
  assign n18084 = n18083 ^ n18019 ;
  assign n18085 = n18018 ^ n662 ;
  assign n18086 = ~n18084 & ~n18085 ;
  assign n18088 = n18087 ^ n18086 ;
  assign n17993 = ~n17963 & ~n17992 ;
  assign n17877 = n17526 ^ n1473 ;
  assign n17867 = n17286 ^ n16876 ;
  assign n17868 = n17867 ^ n16300 ;
  assign n17871 = n17868 ^ n17598 ;
  assign n17870 = n17869 ^ n17868 ;
  assign n17872 = n17871 ^ n17870 ;
  assign n17873 = n17866 & ~n17872 ;
  assign n17874 = n17873 ^ n17871 ;
  assign n17957 = n17877 ^ n17874 ;
  assign n17887 = n17886 ^ n15526 ;
  assign n17954 = ~n17887 & n17953 ;
  assign n17955 = n17954 ^ n15526 ;
  assign n17956 = n17955 ^ n15724 ;
  assign n17962 = n17957 ^ n17956 ;
  assign n18014 = n17993 ^ n17962 ;
  assign n18133 = n18088 ^ n18014 ;
  assign n19210 = n18237 ^ n18133 ;
  assign n19211 = n19210 ^ n17407 ;
  assign n18145 = n17546 ^ n683 ;
  assign n18138 = n18084 ^ n662 ;
  assign n19118 = n18145 ^ n18138 ;
  assign n19119 = n19118 ^ n17395 ;
  assign n18187 = n17608 ^ n16815 ;
  assign n18188 = n18187 ^ n16685 ;
  assign n18181 = n17601 ^ n16810 ;
  assign n18182 = n18181 ^ n16770 ;
  assign n18493 = n18188 ^ n18182 ;
  assign n18186 = n17968 ^ n3070 ;
  assign n18189 = n18188 ^ n18186 ;
  assign n18452 = n17799 ^ n16270 ;
  assign n18453 = n18452 ^ n17202 ;
  assign n18451 = n17776 ^ n17758 ;
  assign n18454 = n18453 ^ n18451 ;
  assign n18322 = n17770 ^ n2507 ;
  assign n18323 = n18322 ^ n17761 ;
  assign n18320 = n17207 ^ n15944 ;
  assign n18321 = n18320 ^ n16543 ;
  assign n18324 = n18323 ^ n18321 ;
  assign n18359 = n17773 ^ n17760 ;
  assign n18360 = n18359 ^ n18323 ;
  assign n18361 = n18360 ^ n18359 ;
  assign n18258 = n16547 ^ n15948 ;
  assign n18259 = n18258 ^ n17218 ;
  assign n18115 = n17767 ^ n17764 ;
  assign n18260 = n18259 ^ n18115 ;
  assign n18192 = n17215 ^ n16550 ;
  assign n18193 = n18192 ^ n15952 ;
  assign n17587 = n17586 ^ n17570 ;
  assign n18194 = n18193 ^ n17587 ;
  assign n18195 = n17803 ^ n16563 ;
  assign n18196 = n18195 ^ n15961 ;
  assign n18121 = n17568 ^ n17458 ;
  assign n18197 = n18196 ^ n18121 ;
  assign n18198 = n17725 ^ n15956 ;
  assign n18199 = n18198 ^ n16560 ;
  assign n18126 = n17563 ^ n1089 ;
  assign n18200 = n18199 ^ n18126 ;
  assign n18201 = n17589 ^ n16528 ;
  assign n18202 = n18201 ^ n17101 ;
  assign n18131 = n17558 ^ n17461 ;
  assign n18203 = n18202 ^ n18131 ;
  assign n18205 = n17632 ^ n16422 ;
  assign n18206 = n18205 ^ n16852 ;
  assign n18136 = n17555 ^ n17463 ;
  assign n18207 = n18206 ^ n18136 ;
  assign n18208 = n17636 ^ n16353 ;
  assign n18209 = n18208 ^ n16856 ;
  assign n18140 = n17553 ^ n17464 ;
  assign n18210 = n18209 ^ n18140 ;
  assign n18214 = n17640 ^ n16347 ;
  assign n18215 = n18214 ^ n16858 ;
  assign n18240 = n18215 ^ n18209 ;
  assign n18211 = n16956 ^ n16339 ;
  assign n18212 = n18211 ^ n17645 ;
  assign n18213 = n18212 ^ n18145 ;
  assign n18218 = n16949 ^ n16284 ;
  assign n18219 = n18218 ^ n17647 ;
  assign n18153 = n17543 ^ n17541 ;
  assign n18220 = n18219 ^ n18153 ;
  assign n18223 = n17539 ^ n17470 ;
  assign n18221 = n17652 ^ n16862 ;
  assign n18222 = n18221 ^ n15675 ;
  assign n18224 = n18223 ^ n18222 ;
  assign n18102 = n17535 ^ n17473 ;
  assign n18100 = n17578 ^ n16787 ;
  assign n18101 = n18100 ^ n16287 ;
  assign n18103 = n18102 ^ n18101 ;
  assign n18002 = n17532 ^ n17476 ;
  assign n18000 = n17407 ^ n16293 ;
  assign n18001 = n18000 ^ n16257 ;
  assign n18003 = n18002 ^ n18001 ;
  assign n17875 = n16793 ^ n16295 ;
  assign n17876 = n17875 ^ n17395 ;
  assign n17879 = n17876 ^ n17868 ;
  assign n17878 = n17877 ^ n17876 ;
  assign n17880 = n17879 ^ n17878 ;
  assign n17881 = n17874 & ~n17880 ;
  assign n17882 = n17881 ^ n17879 ;
  assign n17883 = n17530 ^ n17480 ;
  assign n18004 = n17883 ^ n17876 ;
  assign n18005 = n17882 & ~n18004 ;
  assign n18006 = n18005 ^ n17876 ;
  assign n18097 = n18006 ^ n18002 ;
  assign n18098 = n18003 & ~n18097 ;
  assign n18099 = n18098 ^ n18006 ;
  assign n18225 = n18101 ^ n18099 ;
  assign n18226 = n18103 & ~n18225 ;
  assign n18227 = n18226 ^ n18102 ;
  assign n18228 = n18227 ^ n18222 ;
  assign n18229 = n18224 & n18228 ;
  assign n18230 = n18229 ^ n18223 ;
  assign n18231 = n18230 ^ n18219 ;
  assign n18232 = ~n18220 & ~n18231 ;
  assign n18233 = n18232 ^ n18153 ;
  assign n18216 = n18215 ^ n18145 ;
  assign n18217 = n18216 ^ n18215 ;
  assign n18234 = n18233 ^ n18217 ;
  assign n18235 = n18213 & ~n18234 ;
  assign n18236 = n18235 ^ n18216 ;
  assign n18238 = n18237 ^ n18215 ;
  assign n18239 = ~n18236 & n18238 ;
  assign n18241 = n18240 ^ n18239 ;
  assign n18242 = ~n18210 & ~n18241 ;
  assign n18243 = n18242 ^ n18209 ;
  assign n18244 = n18243 ^ n18136 ;
  assign n18245 = n18207 & ~n18244 ;
  assign n18204 = n18202 ^ n18136 ;
  assign n18246 = n18245 ^ n18204 ;
  assign n18247 = n18203 & ~n18246 ;
  assign n18248 = n18247 ^ n18131 ;
  assign n18249 = n18248 ^ n18126 ;
  assign n18250 = n18200 & n18249 ;
  assign n18251 = n18250 ^ n18126 ;
  assign n18252 = n18251 ^ n18196 ;
  assign n18253 = ~n18197 & ~n18252 ;
  assign n18254 = n18253 ^ n18121 ;
  assign n18255 = n18254 ^ n17587 ;
  assign n18256 = n18194 & n18255 ;
  assign n18257 = n18256 ^ n18193 ;
  assign n18317 = n18259 ^ n18257 ;
  assign n18318 = ~n18260 & ~n18317 ;
  assign n18319 = n18318 ^ n18115 ;
  assign n18362 = n18361 ^ n18319 ;
  assign n18363 = ~n18324 & n18362 ;
  assign n18364 = n18363 ^ n18360 ;
  assign n18455 = n18454 ^ n18364 ;
  assign n3174 = n2763 ^ x322 ;
  assign n3175 = n3174 ^ n1796 ;
  assign n3176 = n3175 ^ x258 ;
  assign n18450 = n3176 ^ n1787 ;
  assign n18456 = n18455 ^ n18450 ;
  assign n18365 = n17205 ^ n16275 ;
  assign n18366 = n18365 ^ n15711 ;
  assign n18367 = n18366 ^ n18364 ;
  assign n18447 = n18367 ^ n14962 ;
  assign n18311 = n18254 ^ n18194 ;
  assign n18262 = n18251 ^ n18197 ;
  assign n18263 = n18262 ^ n15312 ;
  assign n18265 = n18246 ^ n18131 ;
  assign n18266 = n18265 ^ n15870 ;
  assign n18292 = n18241 ^ n18140 ;
  assign n18268 = n18237 ^ n18236 ;
  assign n18269 = n18268 ^ n15770 ;
  assign n18270 = n18233 ^ n18213 ;
  assign n18271 = n18270 ^ n15762 ;
  assign n18273 = n18227 ^ n18224 ;
  assign n18274 = n18273 ^ n15676 ;
  assign n18007 = n18006 ^ n18003 ;
  assign n18008 = n18007 ^ n15719 ;
  assign n17958 = n17957 ^ n17955 ;
  assign n17959 = ~n17956 & n17958 ;
  assign n17960 = n17959 ^ n15724 ;
  assign n17884 = n17883 ^ n17882 ;
  assign n17996 = n17960 ^ n17884 ;
  assign n17997 = n17960 ^ n15717 ;
  assign n17998 = ~n17996 & ~n17997 ;
  assign n17999 = n17998 ^ n15717 ;
  assign n18105 = n18007 ^ n17999 ;
  assign n18106 = ~n18008 & n18105 ;
  assign n18107 = n18106 ^ n15719 ;
  assign n18108 = n18107 ^ n15738 ;
  assign n18104 = n18103 ^ n18099 ;
  assign n18275 = n18107 ^ n18104 ;
  assign n18276 = n18108 & ~n18275 ;
  assign n18277 = n18276 ^ n15738 ;
  assign n18278 = n18277 ^ n18273 ;
  assign n18279 = n18274 & ~n18278 ;
  assign n18280 = n18279 ^ n15676 ;
  assign n18272 = n18230 ^ n18220 ;
  assign n18281 = n18280 ^ n18272 ;
  assign n18282 = n18270 ^ n15752 ;
  assign n18283 = n18282 ^ n18270 ;
  assign n18284 = n18283 ^ n18272 ;
  assign n18285 = ~n18281 & n18284 ;
  assign n18286 = n18285 ^ n18282 ;
  assign n18287 = ~n18271 & ~n18286 ;
  assign n18288 = n18287 ^ n15762 ;
  assign n18289 = n18288 ^ n18268 ;
  assign n18290 = ~n18269 & ~n18289 ;
  assign n18291 = n18290 ^ n15770 ;
  assign n18293 = n18292 ^ n18291 ;
  assign n18294 = n18292 ^ n15821 ;
  assign n18295 = n18293 & ~n18294 ;
  assign n18296 = n18295 ^ n15821 ;
  assign n18267 = n18243 ^ n18207 ;
  assign n18297 = n18296 ^ n18267 ;
  assign n18298 = n18296 ^ n15836 ;
  assign n18299 = n18297 & n18298 ;
  assign n18300 = n18299 ^ n15836 ;
  assign n18301 = n18300 ^ n18265 ;
  assign n18302 = ~n18266 & ~n18301 ;
  assign n18303 = n18302 ^ n15870 ;
  assign n18264 = n18248 ^ n18200 ;
  assign n18304 = n18303 ^ n18264 ;
  assign n18305 = n18303 ^ n15260 ;
  assign n18306 = n18304 & n18305 ;
  assign n18307 = n18306 ^ n15260 ;
  assign n18308 = n18307 ^ n18262 ;
  assign n18309 = ~n18263 & ~n18308 ;
  assign n18310 = n18309 ^ n15312 ;
  assign n18312 = n18311 ^ n18310 ;
  assign n18313 = n18311 ^ n15309 ;
  assign n18314 = n18312 & n18313 ;
  assign n18315 = n18314 ^ n15309 ;
  assign n18261 = n18260 ^ n18257 ;
  assign n18316 = n18315 ^ n18261 ;
  assign n18325 = n18324 ^ n18319 ;
  assign n18326 = n18325 ^ n15339 ;
  assign n18327 = n18326 ^ n18325 ;
  assign n18328 = n18327 ^ n18261 ;
  assign n18329 = ~n18316 & ~n18328 ;
  assign n18330 = n18329 ^ n18326 ;
  assign n18368 = n18325 ^ n15367 ;
  assign n18369 = ~n18330 & ~n18368 ;
  assign n18370 = n18369 ^ n15367 ;
  assign n18448 = n18370 ^ n18367 ;
  assign n18449 = ~n18447 & ~n18448 ;
  assign n18457 = n18456 ^ n18449 ;
  assign n18445 = n18366 ^ n18359 ;
  assign n18446 = ~n18364 & ~n18445 ;
  assign n18458 = n18457 ^ n18446 ;
  assign n18331 = n18330 ^ n15367 ;
  assign n18332 = n18261 ^ n15339 ;
  assign n18333 = n18332 ^ n18315 ;
  assign n18334 = n18313 ^ n18310 ;
  assign n18335 = n18307 ^ n18263 ;
  assign n18336 = n18264 ^ n15260 ;
  assign n18337 = n18336 ^ n18303 ;
  assign n18338 = n18300 ^ n18266 ;
  assign n18339 = n18298 ^ n18267 ;
  assign n18340 = n18294 ^ n18291 ;
  assign n18341 = n18286 ^ n15762 ;
  assign n17885 = n17884 ^ n15717 ;
  assign n17961 = n17960 ^ n17885 ;
  assign n17994 = n17962 & n17993 ;
  assign n17995 = n17961 & n17994 ;
  assign n18009 = n18008 ^ n17999 ;
  assign n18096 = n17995 & ~n18009 ;
  assign n18109 = n18108 ^ n18104 ;
  assign n18342 = ~n18096 & ~n18109 ;
  assign n18343 = n18277 ^ n18274 ;
  assign n18344 = n18342 & ~n18343 ;
  assign n18345 = n18272 ^ n15752 ;
  assign n18346 = n18345 ^ n18280 ;
  assign n18347 = ~n18344 & n18346 ;
  assign n18348 = ~n18341 & n18347 ;
  assign n18349 = n18288 ^ n18269 ;
  assign n18350 = ~n18348 & ~n18349 ;
  assign n18351 = ~n18340 & ~n18350 ;
  assign n18352 = ~n18339 & n18351 ;
  assign n18353 = n18338 & ~n18352 ;
  assign n18354 = n18337 & ~n18353 ;
  assign n18355 = n18335 & n18354 ;
  assign n18356 = n18334 & n18355 ;
  assign n18357 = ~n18333 & ~n18356 ;
  assign n18358 = ~n18331 & ~n18357 ;
  assign n18371 = n18370 ^ n14962 ;
  assign n18372 = n18371 ^ n18367 ;
  assign n18444 = n18358 & n18372 ;
  assign n18459 = n18458 ^ n18444 ;
  assign n18373 = n18372 ^ n18358 ;
  assign n18374 = n18373 ^ n3176 ;
  assign n18375 = n18357 ^ n18331 ;
  assign n18376 = n18375 ^ n1820 ;
  assign n18378 = n18355 ^ n18334 ;
  assign n18379 = n18378 ^ n3148 ;
  assign n18425 = n18354 ^ n18335 ;
  assign n18420 = n18353 ^ n18337 ;
  assign n18415 = n18352 ^ n18338 ;
  assign n18380 = n18351 ^ n18339 ;
  assign n18381 = n18380 ^ n2803 ;
  assign n18406 = n18350 ^ n18340 ;
  assign n18383 = n18347 ^ n18341 ;
  assign n18384 = n18383 ^ n1211 ;
  assign n18110 = n18109 ^ n18096 ;
  assign n18111 = n18110 ^ n742 ;
  assign n18010 = n18009 ^ n17995 ;
  assign n18011 = n18010 ^ n742 ;
  assign n18012 = n17994 ^ n17961 ;
  assign n18013 = n18012 ^ n733 ;
  assign n18090 = n733 ^ n671 ;
  assign n18015 = n18014 ^ n671 ;
  assign n18089 = ~n18015 & ~n18088 ;
  assign n18091 = n18090 ^ n18089 ;
  assign n18092 = ~n18013 & ~n18091 ;
  assign n18093 = n18092 ^ n18012 ;
  assign n18094 = n18093 ^ n742 ;
  assign n18095 = n18011 & ~n18094 ;
  assign n18112 = n18111 ^ n18095 ;
  assign n18386 = n18110 ^ n836 ;
  assign n18387 = ~n18112 & n18386 ;
  assign n18388 = n18387 ^ n836 ;
  assign n978 = n925 ^ x333 ;
  assign n979 = n978 ^ n974 ;
  assign n980 = n979 ^ x269 ;
  assign n18392 = n18388 ^ n980 ;
  assign n18385 = n18343 ^ n18342 ;
  assign n18389 = n18388 ^ n18385 ;
  assign n1191 = n1110 ^ x334 ;
  assign n1192 = n1191 ^ n830 ;
  assign n1193 = n1192 ^ x270 ;
  assign n18390 = n18385 ^ n1193 ;
  assign n18391 = ~n18389 & n18390 ;
  assign n18393 = n18392 ^ n18391 ;
  assign n18396 = n18383 ^ n980 ;
  assign n18394 = n18346 ^ n18344 ;
  assign n18395 = n18394 ^ n18383 ;
  assign n18397 = n18396 ^ n18395 ;
  assign n18398 = n18393 & n18397 ;
  assign n18399 = n18398 ^ n18396 ;
  assign n18400 = n18384 & ~n18399 ;
  assign n18401 = n18400 ^ n1211 ;
  assign n18382 = n18349 ^ n18348 ;
  assign n18402 = n18401 ^ n18382 ;
  assign n18403 = n18382 ^ n1229 ;
  assign n18404 = n18402 & ~n18403 ;
  assign n18405 = n18404 ^ n18401 ;
  assign n18407 = n18406 ^ n18405 ;
  assign n18408 = n18380 ^ n1368 ;
  assign n18409 = n18408 ^ n18380 ;
  assign n18410 = n18409 ^ n18405 ;
  assign n18411 = n18407 & n18410 ;
  assign n18412 = n18411 ^ n18408 ;
  assign n18413 = n18381 & ~n18412 ;
  assign n18414 = n18413 ^ n2803 ;
  assign n18416 = n18415 ^ n18414 ;
  assign n2548 = n2544 ^ x328 ;
  assign n2552 = n2551 ^ n2548 ;
  assign n2553 = n2552 ^ x264 ;
  assign n18417 = n18415 ^ n2553 ;
  assign n18418 = n18416 & ~n18417 ;
  assign n18419 = n18418 ^ n2553 ;
  assign n18421 = n18420 ^ n18419 ;
  assign n18422 = n18420 ^ n2624 ;
  assign n18423 = ~n18421 & n18422 ;
  assign n18424 = n18423 ^ n2624 ;
  assign n18426 = n18425 ^ n18424 ;
  assign n18427 = n18378 ^ n2486 ;
  assign n18428 = n18427 ^ n18378 ;
  assign n18429 = n18428 ^ n18424 ;
  assign n18430 = n18426 & n18429 ;
  assign n18431 = n18430 ^ n18427 ;
  assign n18432 = ~n18379 & n18431 ;
  assign n18433 = n18432 ^ n3148 ;
  assign n18377 = n18356 ^ n18333 ;
  assign n18434 = n18433 ^ n18377 ;
  assign n18477 = n18377 ^ n2468 ;
  assign n18438 = ~n18434 & n18477 ;
  assign n18435 = n2468 ^ n1820 ;
  assign n18439 = n18438 ^ n18435 ;
  assign n18440 = ~n18376 & n18439 ;
  assign n18441 = n18440 ^ n1820 ;
  assign n18442 = n18441 ^ n18373 ;
  assign n18443 = ~n18374 & n18442 ;
  assign n18460 = n18459 ^ n18443 ;
  assign n18190 = n16821 ^ n16594 ;
  assign n18191 = n18190 ^ n17612 ;
  assign n18461 = n18460 ^ n18191 ;
  assign n18464 = n18441 ^ n18374 ;
  assign n18462 = n17251 ^ n16586 ;
  assign n18463 = n18462 ^ n17616 ;
  assign n18465 = n18464 ^ n18463 ;
  assign n18467 = n16826 ^ n16263 ;
  assign n18468 = n18467 ^ n17620 ;
  assign n18484 = n18468 ^ n18463 ;
  assign n18466 = n18439 ^ n18375 ;
  assign n18469 = n18468 ^ n18466 ;
  assign n18474 = n17624 ^ n16835 ;
  assign n18475 = n18474 ^ n16259 ;
  assign n18481 = n18475 ^ n18468 ;
  assign n18470 = n18431 ^ n3148 ;
  assign n18471 = n17628 ^ n16837 ;
  assign n18472 = n18471 ^ n16266 ;
  assign n18473 = ~n18470 & n18472 ;
  assign n18476 = n18475 ^ n18473 ;
  assign n18478 = n18477 ^ n18433 ;
  assign n18479 = n18478 ^ n18475 ;
  assign n18480 = ~n18476 & ~n18479 ;
  assign n18482 = n18481 ^ n18480 ;
  assign n18483 = ~n18469 & ~n18482 ;
  assign n18485 = n18484 ^ n18483 ;
  assign n18486 = ~n18465 & ~n18485 ;
  assign n18487 = n18486 ^ n18464 ;
  assign n18488 = n18487 ^ n18191 ;
  assign n18489 = ~n18461 & n18488 ;
  assign n18490 = n18489 ^ n18460 ;
  assign n18491 = n18490 ^ n18186 ;
  assign n18492 = ~n18189 & n18491 ;
  assign n18494 = n18493 ^ n18492 ;
  assign n18183 = n18043 ^ n3087 ;
  assign n18184 = n18183 ^ n18041 ;
  assign n18581 = n18494 ^ n18184 ;
  assign n18582 = n18581 ^ n15682 ;
  assign n18583 = n18490 ^ n18189 ;
  assign n18584 = n18583 ^ n15678 ;
  assign n18585 = n18487 ^ n18461 ;
  assign n18586 = n18585 ^ n15685 ;
  assign n18590 = n18472 ^ n18470 ;
  assign n18591 = ~n15701 & ~n18590 ;
  assign n18589 = n18478 ^ n18476 ;
  assign n18592 = n18591 ^ n18589 ;
  assign n18593 = n18591 ^ n15699 ;
  assign n18594 = n18592 & n18593 ;
  assign n18595 = n18594 ^ n15699 ;
  assign n18588 = n18482 ^ n18466 ;
  assign n18596 = n18595 ^ n18588 ;
  assign n18597 = n18595 ^ n15693 ;
  assign n18598 = ~n18596 & ~n18597 ;
  assign n18599 = n18598 ^ n15693 ;
  assign n18587 = n18485 ^ n18464 ;
  assign n18600 = n18599 ^ n18587 ;
  assign n18601 = n18599 ^ n15689 ;
  assign n18602 = ~n18600 & n18601 ;
  assign n18603 = n18602 ^ n15689 ;
  assign n18604 = n18603 ^ n18585 ;
  assign n18605 = n18586 & n18604 ;
  assign n18606 = n18605 ^ n15685 ;
  assign n18607 = n18606 ^ n18583 ;
  assign n18608 = ~n18584 & ~n18607 ;
  assign n18609 = n18608 ^ n15678 ;
  assign n18610 = n18609 ^ n18581 ;
  assign n18611 = ~n18582 & ~n18610 ;
  assign n18612 = n18611 ^ n15682 ;
  assign n18185 = n18184 ^ n18182 ;
  assign n18495 = n18185 & ~n18494 ;
  assign n18496 = n18495 ^ n18184 ;
  assign n18179 = n18048 ^ n18047 ;
  assign n18177 = n17593 ^ n16824 ;
  assign n18178 = n18177 ^ n16800 ;
  assign n18180 = n18179 ^ n18178 ;
  assign n18579 = n18496 ^ n18180 ;
  assign n18580 = n18579 ^ n16070 ;
  assign n18738 = n18612 ^ n18580 ;
  assign n18723 = n18597 ^ n18588 ;
  assign n18724 = n18590 ^ n15701 ;
  assign n18725 = n18593 ^ n18589 ;
  assign n18726 = n18724 & ~n18725 ;
  assign n18727 = ~n18723 & n18726 ;
  assign n18728 = n18587 ^ n15689 ;
  assign n18729 = n18728 ^ n18599 ;
  assign n18730 = n18727 & ~n18729 ;
  assign n18731 = n18603 ^ n18586 ;
  assign n18732 = n18730 & ~n18731 ;
  assign n18733 = n18606 ^ n18584 ;
  assign n18734 = ~n18732 & n18733 ;
  assign n18735 = n18609 ^ n15682 ;
  assign n18736 = n18735 ^ n18581 ;
  assign n18737 = ~n18734 & n18736 ;
  assign n18816 = n18738 ^ n18737 ;
  assign n18817 = n18816 ^ n2385 ;
  assign n18818 = n18736 ^ n18734 ;
  assign n18819 = n18818 ^ n2266 ;
  assign n18822 = n18733 ^ n18732 ;
  assign n18823 = n18822 ^ n2240 ;
  assign n18843 = n18731 ^ n18730 ;
  assign n18824 = n18729 ^ n18727 ;
  assign n1971 = n1931 ^ x381 ;
  assign n1975 = n1974 ^ n1971 ;
  assign n1976 = n1975 ^ x317 ;
  assign n18825 = n18824 ^ n1976 ;
  assign n18829 = n18726 ^ n18723 ;
  assign n18826 = n16729 ^ x382 ;
  assign n18827 = n18826 ^ n1909 ;
  assign n18828 = n18827 ^ x318 ;
  assign n18830 = n18829 ^ n18828 ;
  assign n18832 = n18725 ^ n18724 ;
  assign n18836 = n18832 ^ n18828 ;
  assign n18831 = n1867 & ~n18724 ;
  assign n18833 = n18832 ^ n18831 ;
  assign n1900 = n1875 ^ x383 ;
  assign n1904 = n1903 ^ n1900 ;
  assign n1905 = n1904 ^ x319 ;
  assign n18834 = n18831 ^ n1905 ;
  assign n18835 = ~n18833 & ~n18834 ;
  assign n18837 = n18836 ^ n18835 ;
  assign n18838 = ~n18830 & n18837 ;
  assign n18839 = n18838 ^ n18829 ;
  assign n18840 = n18839 ^ n1976 ;
  assign n18841 = ~n18825 & n18840 ;
  assign n18842 = n18841 ^ n18824 ;
  assign n18844 = n18843 ^ n18842 ;
  assign n18847 = n18842 ^ n2247 ;
  assign n18848 = ~n18844 & ~n18847 ;
  assign n18845 = n2247 ^ n2240 ;
  assign n18849 = n18848 ^ n18845 ;
  assign n18850 = n18823 & n18849 ;
  assign n18851 = n18850 ^ n2240 ;
  assign n18820 = n18816 ^ n2266 ;
  assign n18821 = n18820 ^ n18816 ;
  assign n18852 = n18851 ^ n18821 ;
  assign n18853 = ~n18819 & n18852 ;
  assign n18854 = n18853 ^ n18820 ;
  assign n18855 = n18817 & n18854 ;
  assign n18856 = n18855 ^ n18816 ;
  assign n18613 = n18612 ^ n18579 ;
  assign n18614 = ~n18580 & n18613 ;
  assign n18615 = n18614 ^ n16070 ;
  assign n18740 = n18615 ^ n16111 ;
  assign n18175 = n18053 ^ n18039 ;
  assign n18499 = n18179 ^ n18175 ;
  assign n18497 = n18496 ^ n18179 ;
  assign n18498 = n18180 & n18497 ;
  assign n18500 = n18499 ^ n18498 ;
  assign n18173 = n17869 ^ n16829 ;
  assign n18174 = n18173 ^ n17270 ;
  assign n18578 = n18500 ^ n18174 ;
  assign n18741 = n18740 ^ n18578 ;
  assign n18739 = ~n18737 & n18738 ;
  assign n18814 = n18741 ^ n18739 ;
  assign n18815 = n18814 ^ n1466 ;
  assign n19058 = n18856 ^ n18815 ;
  assign n19120 = n19119 ^ n19058 ;
  assign n19123 = n18153 ^ n17286 ;
  assign n18143 = n18081 ^ n18017 ;
  assign n19124 = n19123 ^ n18143 ;
  assign n19065 = n18854 ^ n2385 ;
  assign n19125 = n19124 ^ n19065 ;
  assign n19070 = n18851 ^ n18819 ;
  assign n19203 = n19124 ^ n19070 ;
  assign n18156 = n18071 ^ n18028 ;
  assign n19129 = n18156 ^ n17276 ;
  assign n19130 = n19129 ^ n18002 ;
  assign n19126 = n18843 ^ n2247 ;
  assign n19127 = n19126 ^ n18842 ;
  assign n19131 = n19130 ^ n19127 ;
  assign n19134 = n18840 ^ n18824 ;
  assign n19132 = n17883 ^ n17270 ;
  assign n18512 = n18068 ^ n18030 ;
  assign n19133 = n19132 ^ n18512 ;
  assign n19135 = n19134 ^ n19133 ;
  assign n19136 = n18837 ^ n18829 ;
  assign n19185 = n19136 ^ n19134 ;
  assign n18162 = n18066 ^ n2296 ;
  assign n19137 = n18162 ^ n17877 ;
  assign n19138 = n19137 ^ n16800 ;
  assign n19139 = n19138 ^ n19136 ;
  assign n18160 = n18062 ^ n18061 ;
  assign n19140 = n18160 ^ n16810 ;
  assign n19141 = n19140 ^ n17869 ;
  assign n19081 = n18834 ^ n18832 ;
  assign n19142 = n19141 ^ n19081 ;
  assign n19145 = n18724 ^ n1867 ;
  assign n19179 = n19145 ^ n19081 ;
  assign n18167 = n18058 ^ n18034 ;
  assign n19143 = n18167 ^ n16815 ;
  assign n19144 = n19143 ^ n17593 ;
  assign n19146 = n19145 ^ n19144 ;
  assign n19168 = n17601 ^ n16821 ;
  assign n18171 = n18055 ^ n18038 ;
  assign n19169 = n19168 ^ n18171 ;
  assign n19176 = n19169 ^ n19144 ;
  assign n18778 = n2866 ^ x359 ;
  assign n18779 = n18778 ^ n3109 ;
  assign n18780 = n18779 ^ x295 ;
  assign n18682 = n18323 ^ n17101 ;
  assign n18683 = n18682 ^ n17803 ;
  assign n18681 = n18394 ^ n18393 ;
  assign n18684 = n18683 ^ n18681 ;
  assign n18113 = n18112 ^ n836 ;
  assign n17590 = n17589 ^ n17587 ;
  assign n17591 = n17590 ^ n16856 ;
  assign n18114 = n18113 ^ n17591 ;
  assign n18123 = n18093 ^ n18011 ;
  assign n18120 = n17632 ^ n16858 ;
  assign n18122 = n18121 ^ n18120 ;
  assign n18124 = n18123 ^ n18122 ;
  assign n18128 = n18091 ^ n18012 ;
  assign n18125 = n17636 ^ n16956 ;
  assign n18127 = n18126 ^ n18125 ;
  assign n18129 = n18128 ^ n18127 ;
  assign n18130 = n17640 ^ n16949 ;
  assign n18132 = n18131 ^ n18130 ;
  assign n18134 = n18133 ^ n18132 ;
  assign n18135 = n17645 ^ n16862 ;
  assign n18137 = n18136 ^ n18135 ;
  assign n18139 = n18138 ^ n18137 ;
  assign n18141 = n18140 ^ n16787 ;
  assign n18142 = n18141 ^ n17647 ;
  assign n18144 = n18143 ^ n18142 ;
  assign n18150 = n18079 ^ n18021 ;
  assign n18536 = n18150 ^ n18143 ;
  assign n18148 = n18076 ^ n18074 ;
  assign n18146 = n18145 ^ n16793 ;
  assign n18147 = n18146 ^ n17578 ;
  assign n18149 = n18148 ^ n18147 ;
  assign n18154 = n18153 ^ n17407 ;
  assign n18155 = n18154 ^ n16876 ;
  assign n18157 = n18156 ^ n18155 ;
  assign n18158 = n18002 ^ n16808 ;
  assign n18159 = n18158 ^ n16784 ;
  assign n18161 = n18160 ^ n18159 ;
  assign n18165 = n17883 ^ n16795 ;
  assign n18166 = n18165 ^ n16813 ;
  assign n18168 = n18167 ^ n18166 ;
  assign n18169 = n17877 ^ n17276 ;
  assign n18170 = n18169 ^ n16819 ;
  assign n18172 = n18171 ^ n18170 ;
  assign n18176 = n18175 ^ n18174 ;
  assign n18501 = ~n18176 & n18500 ;
  assign n18502 = n18501 ^ n18175 ;
  assign n18503 = n18502 ^ n18170 ;
  assign n18504 = ~n18172 & ~n18503 ;
  assign n18505 = n18504 ^ n18171 ;
  assign n18506 = n18505 ^ n18166 ;
  assign n18507 = n18168 & ~n18506 ;
  assign n18508 = n18507 ^ n18167 ;
  assign n18163 = n18162 ^ n18160 ;
  assign n18164 = n18163 ^ n18162 ;
  assign n18509 = n18508 ^ n18164 ;
  assign n18510 = n18161 & ~n18509 ;
  assign n18511 = n18510 ^ n18163 ;
  assign n18516 = n18512 ^ n18162 ;
  assign n18513 = n18102 ^ n16798 ;
  assign n18514 = n18513 ^ n17286 ;
  assign n18515 = n18514 ^ n18512 ;
  assign n18517 = n18516 ^ n18515 ;
  assign n18518 = ~n18511 & ~n18517 ;
  assign n18519 = n18518 ^ n18516 ;
  assign n18523 = n18512 ^ n18155 ;
  assign n18520 = n18223 ^ n17395 ;
  assign n18521 = n18520 ^ n16803 ;
  assign n18522 = n18521 ^ n18155 ;
  assign n18524 = n18523 ^ n18522 ;
  assign n18525 = ~n18519 & ~n18524 ;
  assign n18526 = n18525 ^ n18523 ;
  assign n18527 = n18157 & ~n18526 ;
  assign n18528 = n18527 ^ n18156 ;
  assign n18151 = n18150 ^ n18148 ;
  assign n18152 = n18151 ^ n18150 ;
  assign n18529 = n18528 ^ n18152 ;
  assign n18530 = ~n18149 & ~n18529 ;
  assign n18531 = n18530 ^ n18151 ;
  assign n18532 = n17652 ^ n16257 ;
  assign n18533 = n18532 ^ n18237 ;
  assign n18534 = n18533 ^ n18150 ;
  assign n18535 = ~n18531 & n18534 ;
  assign n18537 = n18536 ^ n18535 ;
  assign n18538 = ~n18144 & n18537 ;
  assign n18539 = n18538 ^ n18143 ;
  assign n18540 = n18539 ^ n18138 ;
  assign n18541 = ~n18139 & n18540 ;
  assign n18542 = n18541 ^ n18138 ;
  assign n18543 = n18542 ^ n18132 ;
  assign n18544 = ~n18134 & ~n18543 ;
  assign n18545 = n18544 ^ n18133 ;
  assign n18546 = n18545 ^ n18127 ;
  assign n18547 = ~n18129 & ~n18546 ;
  assign n18548 = n18547 ^ n18128 ;
  assign n18549 = n18548 ^ n18122 ;
  assign n18550 = n18124 & ~n18549 ;
  assign n18551 = n18550 ^ n18123 ;
  assign n18116 = n18115 ^ n17725 ;
  assign n18117 = n18116 ^ n16852 ;
  assign n18118 = n18117 ^ n18113 ;
  assign n18119 = n18118 ^ n18117 ;
  assign n18552 = n18551 ^ n18119 ;
  assign n18553 = n18114 & ~n18552 ;
  assign n18554 = n18553 ^ n18118 ;
  assign n18555 = n18390 ^ n18388 ;
  assign n18678 = n18555 ^ n18117 ;
  assign n18679 = ~n18554 & n18678 ;
  assign n18680 = n18679 ^ n18117 ;
  assign n18685 = n18684 ^ n18680 ;
  assign n18556 = n18555 ^ n18554 ;
  assign n18557 = n18556 ^ n16422 ;
  assign n18560 = n18545 ^ n18129 ;
  assign n18561 = n18560 ^ n16339 ;
  assign n18562 = n18542 ^ n18134 ;
  assign n18563 = n18562 ^ n16284 ;
  assign n18565 = n18533 ^ n18531 ;
  assign n18566 = n18565 ^ n16293 ;
  assign n18568 = n18526 ^ n18156 ;
  assign n18569 = n18568 ^ n16300 ;
  assign n18570 = n18521 ^ n18519 ;
  assign n18571 = n18570 ^ n16304 ;
  assign n18572 = n18514 ^ n18511 ;
  assign n18573 = n18572 ^ n16310 ;
  assign n18627 = n18508 ^ n18161 ;
  assign n18574 = n18505 ^ n18168 ;
  assign n18575 = n18574 ^ n16231 ;
  assign n18576 = n18502 ^ n18172 ;
  assign n18577 = n18576 ^ n16126 ;
  assign n18616 = n18615 ^ n18578 ;
  assign n18617 = n18576 ^ n16111 ;
  assign n18618 = n18617 ^ n18576 ;
  assign n18619 = n18618 ^ n18578 ;
  assign n18620 = ~n18616 & ~n18619 ;
  assign n18621 = n18620 ^ n18617 ;
  assign n18622 = n18577 & n18621 ;
  assign n18623 = n18622 ^ n16126 ;
  assign n18624 = n18623 ^ n18574 ;
  assign n18625 = n18575 & ~n18624 ;
  assign n18626 = n18625 ^ n16231 ;
  assign n18628 = n18627 ^ n18626 ;
  assign n18629 = n18572 ^ n16246 ;
  assign n18630 = n18629 ^ n18626 ;
  assign n18631 = n18630 ^ n18572 ;
  assign n18632 = ~n18628 & n18631 ;
  assign n18633 = n18632 ^ n18629 ;
  assign n18634 = n18573 & ~n18633 ;
  assign n18635 = n18634 ^ n16310 ;
  assign n18636 = n18635 ^ n18570 ;
  assign n18637 = n18571 & n18636 ;
  assign n18638 = n18637 ^ n16304 ;
  assign n18639 = n18638 ^ n18568 ;
  assign n18640 = ~n18569 & ~n18639 ;
  assign n18641 = n18640 ^ n16300 ;
  assign n18567 = n18528 ^ n18149 ;
  assign n18642 = n18641 ^ n18567 ;
  assign n18643 = n18565 ^ n16295 ;
  assign n18644 = n18643 ^ n18565 ;
  assign n18645 = n18644 ^ n18567 ;
  assign n18646 = ~n18642 & ~n18645 ;
  assign n18647 = n18646 ^ n18643 ;
  assign n18648 = ~n18566 & n18647 ;
  assign n18649 = n18648 ^ n16293 ;
  assign n18564 = n18537 ^ n18142 ;
  assign n18650 = n18649 ^ n18564 ;
  assign n18651 = n18539 ^ n18139 ;
  assign n18652 = n18651 ^ n16287 ;
  assign n18653 = n18652 ^ n18564 ;
  assign n18654 = n18653 ^ n18651 ;
  assign n18655 = n18650 & n18654 ;
  assign n18656 = n18655 ^ n18652 ;
  assign n18658 = n18562 ^ n15675 ;
  assign n18657 = n18651 ^ n18562 ;
  assign n18659 = n18658 ^ n18657 ;
  assign n18660 = ~n18656 & n18659 ;
  assign n18661 = n18660 ^ n18658 ;
  assign n18662 = ~n18563 & ~n18661 ;
  assign n18663 = n18662 ^ n16284 ;
  assign n18664 = n18663 ^ n18560 ;
  assign n18665 = n18561 & ~n18664 ;
  assign n18666 = n18665 ^ n16339 ;
  assign n18559 = n18548 ^ n18124 ;
  assign n18667 = n18666 ^ n18559 ;
  assign n18668 = n18666 ^ n16347 ;
  assign n18669 = ~n18667 & ~n18668 ;
  assign n18670 = n18669 ^ n16347 ;
  assign n18558 = n18551 ^ n18114 ;
  assign n18671 = n18670 ^ n18558 ;
  assign n18672 = n18670 ^ n16353 ;
  assign n18673 = n18671 & ~n18672 ;
  assign n18674 = n18673 ^ n16353 ;
  assign n18675 = n18674 ^ n18556 ;
  assign n18676 = n18557 & n18675 ;
  assign n18677 = n18676 ^ n16422 ;
  assign n18686 = n18685 ^ n18677 ;
  assign n18692 = n18359 ^ n17215 ;
  assign n18693 = n18692 ^ n16560 ;
  assign n18689 = n18681 ^ n18680 ;
  assign n18690 = n18684 & ~n18689 ;
  assign n18687 = n18399 ^ n1211 ;
  assign n18688 = n18687 ^ n18681 ;
  assign n18691 = n18690 ^ n18688 ;
  assign n18694 = n18693 ^ n18691 ;
  assign n18695 = n18694 ^ n16528 ;
  assign n18696 = n18695 ^ n18677 ;
  assign n18697 = n18696 ^ n18694 ;
  assign n18698 = n18686 & n18697 ;
  assign n18699 = n18698 ^ n18695 ;
  assign n18774 = n18699 ^ n15956 ;
  assign n18715 = n18663 ^ n18561 ;
  assign n18716 = n18656 ^ n15675 ;
  assign n18717 = n18564 ^ n16287 ;
  assign n18718 = n18717 ^ n18649 ;
  assign n18719 = n18641 ^ n16295 ;
  assign n18720 = n18719 ^ n18567 ;
  assign n18721 = n18633 ^ n16310 ;
  assign n18722 = n18623 ^ n18575 ;
  assign n18742 = n18739 & n18741 ;
  assign n18743 = n18621 ^ n16126 ;
  assign n18744 = n18742 & n18743 ;
  assign n18745 = n18722 & ~n18744 ;
  assign n18746 = n18627 ^ n16246 ;
  assign n18747 = n18746 ^ n18626 ;
  assign n18748 = ~n18745 & ~n18747 ;
  assign n18749 = n18721 & ~n18748 ;
  assign n18750 = n18635 ^ n16304 ;
  assign n18751 = n18750 ^ n18570 ;
  assign n18752 = ~n18749 & ~n18751 ;
  assign n18753 = n18638 ^ n16300 ;
  assign n18754 = n18753 ^ n18568 ;
  assign n18755 = n18752 & ~n18754 ;
  assign n18756 = n18720 & n18755 ;
  assign n18757 = n18647 ^ n16293 ;
  assign n18758 = n18756 & ~n18757 ;
  assign n18759 = ~n18718 & ~n18758 ;
  assign n18760 = n18716 & n18759 ;
  assign n18761 = n18661 ^ n16284 ;
  assign n18762 = ~n18760 & n18761 ;
  assign n18763 = n18715 & n18762 ;
  assign n18764 = n18668 ^ n18559 ;
  assign n18765 = ~n18763 & n18764 ;
  assign n18766 = n18558 ^ n16353 ;
  assign n18767 = n18766 ^ n18670 ;
  assign n18768 = ~n18765 & ~n18767 ;
  assign n18769 = n18674 ^ n18557 ;
  assign n18770 = n18768 & n18769 ;
  assign n18771 = n18685 ^ n16528 ;
  assign n18772 = n18771 ^ n18677 ;
  assign n18773 = ~n18770 & ~n18772 ;
  assign n18777 = n18774 ^ n18773 ;
  assign n18781 = n18780 ^ n18777 ;
  assign n18782 = n18772 ^ n18770 ;
  assign n18783 = n18782 ^ n2856 ;
  assign n18784 = n18769 ^ n18768 ;
  assign n18785 = n18784 ^ n2841 ;
  assign n18786 = n18767 ^ n18765 ;
  assign n18787 = n18786 ^ n2834 ;
  assign n18789 = n18761 ^ n18760 ;
  assign n18790 = n18789 ^ n1058 ;
  assign n18791 = n18759 ^ n18716 ;
  assign n18792 = n18791 ^ n903 ;
  assign n18886 = n18791 ^ n825 ;
  assign n18793 = n18758 ^ n18718 ;
  assign n18794 = n18793 ^ n825 ;
  assign n18795 = n18757 ^ n18756 ;
  assign n18796 = n18795 ^ n810 ;
  assign n18797 = n18755 ^ n18720 ;
  assign n18798 = n18797 ^ n801 ;
  assign n18799 = n18754 ^ n18752 ;
  assign n18800 = n18799 ^ n1557 ;
  assign n18801 = n18751 ^ n18749 ;
  assign n18802 = n18801 ^ n1567 ;
  assign n18804 = n18747 ^ n18745 ;
  assign n18805 = n18804 ^ n2938 ;
  assign n18806 = n18744 ^ n18722 ;
  assign n18807 = n18806 ^ n575 ;
  assign n18808 = n18743 ^ n18742 ;
  assign n18812 = n18811 ^ n18808 ;
  assign n18857 = n18856 ^ n18814 ;
  assign n18858 = ~n18815 & n18857 ;
  assign n18813 = n18811 ^ n1466 ;
  assign n18859 = n18858 ^ n18813 ;
  assign n18860 = ~n18812 & n18859 ;
  assign n18861 = n18860 ^ n18811 ;
  assign n18862 = n18861 ^ n18806 ;
  assign n18863 = ~n18807 & n18862 ;
  assign n18864 = n18863 ^ n575 ;
  assign n18865 = n18864 ^ n18804 ;
  assign n18866 = ~n18805 & n18865 ;
  assign n18867 = n18866 ^ n2938 ;
  assign n18803 = n18748 ^ n18721 ;
  assign n18868 = n18867 ^ n18803 ;
  assign n18869 = n18867 ^ n527 ;
  assign n18870 = n18868 & n18869 ;
  assign n18871 = n18870 ^ n527 ;
  assign n18872 = n18871 ^ n1567 ;
  assign n18873 = ~n18802 & ~n18872 ;
  assign n18874 = n18873 ^ n18801 ;
  assign n18875 = n18874 ^ n1557 ;
  assign n18876 = n18800 & n18875 ;
  assign n18877 = n18876 ^ n18799 ;
  assign n18878 = n18877 ^ n801 ;
  assign n18879 = ~n18798 & ~n18878 ;
  assign n18880 = n18879 ^ n18797 ;
  assign n18881 = n18880 ^ n810 ;
  assign n18882 = n18796 & n18881 ;
  assign n18883 = n18882 ^ n18795 ;
  assign n18884 = n18883 ^ n825 ;
  assign n18885 = n18794 & n18884 ;
  assign n18887 = n18886 ^ n18885 ;
  assign n18888 = n18792 & n18887 ;
  assign n18889 = n18888 ^ n18791 ;
  assign n18890 = n18889 ^ n18789 ;
  assign n18891 = n18790 & ~n18890 ;
  assign n18892 = n18891 ^ n1058 ;
  assign n1050 = n968 ^ x364 ;
  assign n1054 = n1053 ^ n1050 ;
  assign n1055 = n1054 ^ x300 ;
  assign n18893 = n18892 ^ n1055 ;
  assign n18894 = n18762 ^ n18715 ;
  assign n18895 = n18894 ^ n18892 ;
  assign n18896 = n18893 & n18895 ;
  assign n18897 = n18896 ^ n1055 ;
  assign n18788 = n18764 ^ n18763 ;
  assign n18898 = n18897 ^ n18788 ;
  assign n18899 = n18786 ^ n1250 ;
  assign n18900 = n18899 ^ n18786 ;
  assign n18901 = n18900 ^ n18788 ;
  assign n18902 = n18898 & ~n18901 ;
  assign n18903 = n18902 ^ n18899 ;
  assign n18904 = ~n18787 & n18903 ;
  assign n18905 = n18904 ^ n2834 ;
  assign n18906 = n18905 ^ n18784 ;
  assign n18907 = ~n18785 & n18906 ;
  assign n18908 = n18907 ^ n2841 ;
  assign n18909 = n18908 ^ n18782 ;
  assign n18910 = n18783 & ~n18909 ;
  assign n18911 = n18910 ^ n2856 ;
  assign n18912 = n18911 ^ n18777 ;
  assign n18913 = n18781 & ~n18912 ;
  assign n18914 = n18913 ^ n18780 ;
  assign n18775 = ~n18773 & n18774 ;
  assign n18705 = n17218 ^ n16563 ;
  assign n18706 = n18705 ^ n18451 ;
  assign n18703 = n18401 ^ n1229 ;
  assign n18704 = n18703 ^ n18382 ;
  assign n18707 = n18706 ^ n18704 ;
  assign n18700 = n18693 ^ n18687 ;
  assign n18701 = n18691 & ~n18700 ;
  assign n18702 = n18701 ^ n18687 ;
  assign n18708 = n18707 ^ n18702 ;
  assign n18710 = n18708 ^ n15956 ;
  assign n18709 = n18708 ^ n18694 ;
  assign n18711 = n18710 ^ n18709 ;
  assign n18712 = n18699 & ~n18711 ;
  assign n18713 = n18712 ^ n18710 ;
  assign n18714 = n18713 ^ n15961 ;
  assign n18776 = n18775 ^ n18714 ;
  assign n18915 = n18914 ^ n18776 ;
  assign n18930 = ~n18714 & n18775 ;
  assign n18926 = n18708 ^ n15961 ;
  assign n18927 = n18713 & n18926 ;
  assign n18928 = n18927 ^ n15961 ;
  assign n18922 = n18406 ^ n1368 ;
  assign n18923 = n18922 ^ n18405 ;
  assign n18918 = n17207 ^ n16550 ;
  assign n18919 = n18918 ^ n17826 ;
  assign n18920 = n18919 ^ n18704 ;
  assign n18916 = n18704 ^ n18702 ;
  assign n18917 = ~n18707 & n18916 ;
  assign n18921 = n18920 ^ n18917 ;
  assign n18924 = n18923 ^ n18921 ;
  assign n18925 = n18924 ^ n15952 ;
  assign n18929 = n18928 ^ n18925 ;
  assign n18931 = n18930 ^ n18929 ;
  assign n2588 = n2575 ^ x358 ;
  assign n2589 = n2588 ^ n1829 ;
  assign n2590 = n2589 ^ x294 ;
  assign n18932 = n18931 ^ n2590 ;
  assign n18933 = n18932 ^ n18776 ;
  assign n18934 = n18933 ^ n18931 ;
  assign n18935 = ~n18915 & n18934 ;
  assign n18936 = n18935 ^ n18932 ;
  assign n18951 = n18412 ^ n2803 ;
  assign n18949 = n17831 ^ n17205 ;
  assign n18950 = n18949 ^ n16547 ;
  assign n18952 = n18951 ^ n18950 ;
  assign n18946 = n18923 ^ n18919 ;
  assign n18947 = ~n18921 & ~n18946 ;
  assign n18948 = n18947 ^ n18923 ;
  assign n18953 = n18952 ^ n18948 ;
  assign n18954 = n18953 ^ n15948 ;
  assign n18942 = n18928 ^ n18924 ;
  assign n18943 = n18928 ^ n15952 ;
  assign n18944 = ~n18942 & n18943 ;
  assign n18945 = n18944 ^ n15952 ;
  assign n18955 = n18954 ^ n18945 ;
  assign n18941 = n18929 & n18930 ;
  assign n18956 = n18955 ^ n18941 ;
  assign n18958 = n18956 ^ n2596 ;
  assign n18957 = n18956 ^ n18931 ;
  assign n18959 = n18958 ^ n18957 ;
  assign n18960 = n18936 & ~n18959 ;
  assign n18961 = n18960 ^ n18958 ;
  assign n18979 = n17821 ^ n17202 ;
  assign n18980 = n18979 ^ n16543 ;
  assign n18972 = n18414 ^ n2553 ;
  assign n18973 = n18972 ^ n18415 ;
  assign n18974 = n18973 ^ n18951 ;
  assign n18975 = n18974 ^ n18973 ;
  assign n18976 = n18975 ^ n18948 ;
  assign n18977 = n18952 & ~n18976 ;
  assign n18978 = n18977 ^ n18974 ;
  assign n18981 = n18980 ^ n18978 ;
  assign n18982 = n18981 ^ n15944 ;
  assign n18969 = n18953 ^ n18945 ;
  assign n18970 = ~n18954 & ~n18969 ;
  assign n18971 = n18970 ^ n15948 ;
  assign n18983 = n18982 ^ n18971 ;
  assign n18968 = ~n18941 & n18955 ;
  assign n18984 = n18983 ^ n18968 ;
  assign n18986 = n18984 ^ n2530 ;
  assign n18985 = n18984 ^ n18956 ;
  assign n18987 = n18986 ^ n18985 ;
  assign n18988 = n18961 & ~n18987 ;
  assign n18989 = n18988 ^ n18986 ;
  assign n19032 = n18422 ^ n18419 ;
  assign n19030 = n17817 ^ n16275 ;
  assign n19031 = n19030 ^ n16841 ;
  assign n19033 = n19032 ^ n19031 ;
  assign n19027 = n18980 ^ n18973 ;
  assign n19028 = ~n18978 & ~n19027 ;
  assign n19029 = n19028 ^ n18973 ;
  assign n19034 = n19033 ^ n19029 ;
  assign n19035 = n19034 ^ n15944 ;
  assign n19036 = n19035 ^ n19034 ;
  assign n19037 = n19036 ^ n18971 ;
  assign n19038 = ~n18982 & n19037 ;
  assign n19039 = n19038 ^ n19035 ;
  assign n19040 = n19039 ^ n15711 ;
  assign n19026 = ~n18968 & n18983 ;
  assign n19041 = n19040 ^ n19026 ;
  assign n19043 = n19041 ^ n18984 ;
  assign n19042 = n19041 ^ n2456 ;
  assign n19044 = n19043 ^ n19042 ;
  assign n19045 = ~n18989 & n19044 ;
  assign n19046 = n19045 ^ n19042 ;
  assign n19165 = n19041 ^ n2744 ;
  assign n19166 = n19046 & ~n19165 ;
  assign n19161 = n19039 ^ n19026 ;
  assign n19162 = ~n15711 & n19161 ;
  assign n19157 = n19031 ^ n15707 ;
  assign n19154 = n18425 ^ n2486 ;
  assign n19155 = n19154 ^ n18424 ;
  assign n19152 = n17811 ^ n17238 ;
  assign n19153 = n19152 ^ n16270 ;
  assign n19156 = n19155 ^ n19153 ;
  assign n19158 = n19157 ^ n19156 ;
  assign n19151 = n2744 ^ n1858 ;
  assign n19159 = n19158 ^ n19151 ;
  assign n19149 = n19031 ^ n19029 ;
  assign n19150 = ~n19033 & n19149 ;
  assign n19160 = n19159 ^ n19150 ;
  assign n19163 = n19162 ^ n19160 ;
  assign n19147 = n19034 ^ n19026 ;
  assign n19148 = ~n19039 & n19147 ;
  assign n19164 = n19163 ^ n19148 ;
  assign n19167 = n19166 ^ n19164 ;
  assign n19170 = n19169 ^ n19167 ;
  assign n19047 = n19046 ^ n2744 ;
  assign n19173 = n19167 ^ n19047 ;
  assign n19048 = n18175 ^ n17608 ;
  assign n19049 = n19048 ^ n17251 ;
  assign n19050 = n19049 ^ n19047 ;
  assign n18990 = n18989 ^ n2456 ;
  assign n18962 = n18961 ^ n2530 ;
  assign n18991 = n18990 ^ n18962 ;
  assign n18937 = n18936 ^ n2596 ;
  assign n18938 = n18186 ^ n17620 ;
  assign n18939 = n18938 ^ n16837 ;
  assign n18940 = ~n18937 & n18939 ;
  assign n18963 = n18962 ^ n18940 ;
  assign n18964 = n18184 ^ n16835 ;
  assign n18965 = n18964 ^ n17616 ;
  assign n18966 = n18965 ^ n18940 ;
  assign n18967 = ~n18963 & ~n18966 ;
  assign n18992 = n18991 ^ n18967 ;
  assign n18993 = n17612 ^ n16826 ;
  assign n18994 = n18993 ^ n18179 ;
  assign n19023 = n18994 ^ n18990 ;
  assign n19024 = ~n18992 & n19023 ;
  assign n19025 = n19024 ^ n18990 ;
  assign n19171 = n19047 ^ n19025 ;
  assign n19172 = ~n19050 & ~n19171 ;
  assign n19174 = n19173 ^ n19172 ;
  assign n19175 = n19170 & ~n19174 ;
  assign n19177 = n19176 ^ n19175 ;
  assign n19178 = ~n19146 & n19177 ;
  assign n19180 = n19179 ^ n19178 ;
  assign n19181 = n19142 & n19180 ;
  assign n19182 = n19181 ^ n19081 ;
  assign n19183 = n19182 ^ n19136 ;
  assign n19184 = ~n19139 & ~n19183 ;
  assign n19186 = n19185 ^ n19184 ;
  assign n19187 = ~n19135 & n19186 ;
  assign n19188 = n19187 ^ n19134 ;
  assign n19189 = n19188 ^ n19127 ;
  assign n19190 = ~n19131 & n19189 ;
  assign n19076 = n18849 ^ n18822 ;
  assign n19128 = n19127 ^ n19076 ;
  assign n19191 = n19190 ^ n19128 ;
  assign n19193 = n18148 ^ n16795 ;
  assign n19194 = n19193 ^ n18102 ;
  assign n19192 = n19076 ^ n19070 ;
  assign n19195 = n19194 ^ n19192 ;
  assign n19196 = n19195 ^ n19070 ;
  assign n19197 = n19191 & n19196 ;
  assign n19198 = n19197 ^ n19192 ;
  assign n19199 = n18223 ^ n16784 ;
  assign n19200 = n19199 ^ n18150 ;
  assign n19201 = n19200 ^ n19070 ;
  assign n19202 = ~n19198 & n19201 ;
  assign n19204 = n19203 ^ n19202 ;
  assign n19205 = ~n19125 & ~n19204 ;
  assign n19206 = n19205 ^ n19065 ;
  assign n19062 = n18859 ^ n18808 ;
  assign n19121 = n19062 ^ n19058 ;
  assign n19122 = n19121 ^ n19062 ;
  assign n19207 = n19206 ^ n19122 ;
  assign n19208 = n19120 & ~n19207 ;
  assign n19209 = n19208 ^ n19121 ;
  assign n19257 = n19211 ^ n19209 ;
  assign n19258 = n19257 ^ n16876 ;
  assign n19309 = n19206 ^ n19120 ;
  assign n19259 = n19204 ^ n19065 ;
  assign n19260 = n19259 ^ n16798 ;
  assign n19261 = n19200 ^ n19198 ;
  assign n19262 = n19261 ^ n16808 ;
  assign n19263 = n19194 ^ n19191 ;
  assign n19264 = n19263 ^ n16813 ;
  assign n19266 = n19186 ^ n19133 ;
  assign n19267 = n19266 ^ n16829 ;
  assign n19268 = n19182 ^ n19139 ;
  assign n19269 = n19268 ^ n16824 ;
  assign n19270 = n19180 ^ n19141 ;
  assign n19271 = n19270 ^ n16770 ;
  assign n19272 = n19177 ^ n19145 ;
  assign n19273 = n19272 ^ n16685 ;
  assign n19051 = n19050 ^ n19025 ;
  assign n19052 = n19051 ^ n16586 ;
  assign n18995 = n18994 ^ n18992 ;
  assign n18996 = n18995 ^ n16263 ;
  assign n18997 = n18939 ^ n18937 ;
  assign n18998 = n16266 & ~n18997 ;
  assign n18999 = n18998 ^ n16259 ;
  assign n19000 = n18966 ^ n18962 ;
  assign n19001 = n19000 ^ n18998 ;
  assign n19002 = n18999 & n19001 ;
  assign n19003 = n19002 ^ n16259 ;
  assign n19020 = n19003 ^ n18995 ;
  assign n19021 = n18996 & n19020 ;
  assign n19022 = n19021 ^ n16263 ;
  assign n19275 = n19051 ^ n19022 ;
  assign n19276 = ~n19052 & ~n19275 ;
  assign n19277 = n19276 ^ n16586 ;
  assign n19274 = n19174 ^ n19169 ;
  assign n19278 = n19277 ^ n19274 ;
  assign n19279 = n19272 ^ n16594 ;
  assign n19280 = n19279 ^ n19272 ;
  assign n19281 = n19280 ^ n19274 ;
  assign n19282 = n19278 & n19281 ;
  assign n19283 = n19282 ^ n19279 ;
  assign n19284 = n19273 & n19283 ;
  assign n19285 = n19284 ^ n16685 ;
  assign n19286 = n19285 ^ n19270 ;
  assign n19287 = n19271 & n19286 ;
  assign n19288 = n19287 ^ n16770 ;
  assign n19289 = n19288 ^ n19268 ;
  assign n19290 = ~n19269 & n19289 ;
  assign n19291 = n19290 ^ n16824 ;
  assign n19292 = n19291 ^ n19266 ;
  assign n19293 = ~n19267 & ~n19292 ;
  assign n19294 = n19293 ^ n16829 ;
  assign n19265 = n19188 ^ n19131 ;
  assign n19295 = n19294 ^ n19265 ;
  assign n19296 = n19263 ^ n16819 ;
  assign n19297 = n19296 ^ n19263 ;
  assign n19298 = n19297 ^ n19265 ;
  assign n19299 = n19295 & n19298 ;
  assign n19300 = n19299 ^ n19296 ;
  assign n19301 = ~n19264 & n19300 ;
  assign n19302 = n19301 ^ n16813 ;
  assign n19303 = n19302 ^ n19261 ;
  assign n19304 = ~n19262 & n19303 ;
  assign n19305 = n19304 ^ n16808 ;
  assign n19306 = n19305 ^ n19259 ;
  assign n19307 = ~n19260 & n19306 ;
  assign n19308 = n19307 ^ n16798 ;
  assign n19310 = n19309 ^ n19308 ;
  assign n19311 = n19309 ^ n16803 ;
  assign n19312 = n19310 & n19311 ;
  assign n19313 = n19312 ^ n16803 ;
  assign n19314 = n19313 ^ n19257 ;
  assign n19315 = ~n19258 & n19314 ;
  assign n19316 = n19315 ^ n16876 ;
  assign n19114 = n18861 ^ n18807 ;
  assign n19214 = n19114 ^ n19062 ;
  assign n19212 = n19211 ^ n19062 ;
  assign n19213 = n19209 & n19212 ;
  assign n19215 = n19214 ^ n19213 ;
  assign n19115 = n18128 ^ n17578 ;
  assign n19116 = n19115 ^ n18140 ;
  assign n19255 = n19215 ^ n19116 ;
  assign n19256 = n19255 ^ n16793 ;
  assign n19356 = n19316 ^ n19256 ;
  assign n19357 = n19311 ^ n19308 ;
  assign n19053 = n19052 ^ n19022 ;
  assign n19004 = n19003 ^ n18996 ;
  assign n19005 = n18997 ^ n16266 ;
  assign n19006 = n19000 ^ n18999 ;
  assign n19007 = ~n19005 & ~n19006 ;
  assign n19054 = n19004 & n19007 ;
  assign n19358 = n19053 & n19054 ;
  assign n19359 = n19274 ^ n16594 ;
  assign n19360 = n19359 ^ n19277 ;
  assign n19361 = n19358 & n19360 ;
  assign n19362 = n19283 ^ n16685 ;
  assign n19363 = ~n19361 & n19362 ;
  assign n19364 = n19285 ^ n19271 ;
  assign n19365 = ~n19363 & n19364 ;
  assign n19366 = n19288 ^ n19269 ;
  assign n19367 = ~n19365 & ~n19366 ;
  assign n19368 = n19291 ^ n19267 ;
  assign n19369 = n19367 & ~n19368 ;
  assign n19370 = n19265 ^ n16819 ;
  assign n19371 = n19370 ^ n19294 ;
  assign n19372 = n19369 & ~n19371 ;
  assign n19373 = n19300 ^ n16813 ;
  assign n19374 = ~n19372 & n19373 ;
  assign n19375 = n19302 ^ n19262 ;
  assign n19376 = ~n19374 & ~n19375 ;
  assign n19377 = n19305 ^ n19260 ;
  assign n19378 = ~n19376 & n19377 ;
  assign n19379 = n19357 & ~n19378 ;
  assign n19380 = n19313 ^ n19258 ;
  assign n19381 = n19379 & n19380 ;
  assign n19382 = n19356 & n19381 ;
  assign n19317 = n19316 ^ n19255 ;
  assign n19318 = ~n19256 & n19317 ;
  assign n19319 = n19318 ^ n16793 ;
  assign n19117 = n19116 ^ n19114 ;
  assign n19216 = n19117 & ~n19215 ;
  assign n19217 = n19216 ^ n19116 ;
  assign n19111 = n18123 ^ n17652 ;
  assign n19112 = n19111 ^ n18136 ;
  assign n19110 = n18864 ^ n18805 ;
  assign n19113 = n19112 ^ n19110 ;
  assign n19253 = n19217 ^ n19113 ;
  assign n19254 = n19253 ^ n16257 ;
  assign n19383 = n19319 ^ n19254 ;
  assign n19384 = n19382 & ~n19383 ;
  assign n19320 = n19319 ^ n19253 ;
  assign n19321 = n19254 & ~n19320 ;
  assign n19322 = n19321 ^ n16257 ;
  assign n19218 = n19217 ^ n19110 ;
  assign n19219 = ~n19113 & ~n19218 ;
  assign n19220 = n19219 ^ n19112 ;
  assign n19104 = n18131 ^ n18113 ;
  assign n19105 = n19104 ^ n17647 ;
  assign n19102 = n18803 ^ n527 ;
  assign n19103 = n19102 ^ n18867 ;
  assign n19106 = n19105 ^ n19103 ;
  assign n19251 = n19220 ^ n19106 ;
  assign n19252 = n19251 ^ n16787 ;
  assign n19385 = n19322 ^ n19252 ;
  assign n19386 = ~n19384 & ~n19385 ;
  assign n19323 = n19322 ^ n19251 ;
  assign n19324 = ~n19252 & n19323 ;
  assign n19325 = n19324 ^ n16787 ;
  assign n19354 = n19325 ^ n16862 ;
  assign n19225 = n18126 ^ n17645 ;
  assign n19226 = n19225 ^ n18555 ;
  assign n19107 = n18871 ^ n18802 ;
  assign n19108 = n19107 ^ n19103 ;
  assign n19109 = n19108 ^ n19107 ;
  assign n19221 = n19220 ^ n19109 ;
  assign n19222 = ~n19106 & ~n19221 ;
  assign n19223 = n19222 ^ n19108 ;
  assign n19250 = n19226 ^ n19223 ;
  assign n19355 = n19354 ^ n19250 ;
  assign n19467 = n19386 ^ n19355 ;
  assign n19468 = n19467 ^ n1021 ;
  assign n19469 = n19385 ^ n19384 ;
  assign n19470 = n19469 ^ n1015 ;
  assign n19548 = n19383 ^ n19382 ;
  assign n19471 = n19381 ^ n19356 ;
  assign n19472 = n19471 ^ n1623 ;
  assign n19473 = n19380 ^ n19379 ;
  assign n19474 = n19473 ^ n648 ;
  assign n19475 = n19378 ^ n19357 ;
  assign n19476 = n19475 ^ n557 ;
  assign n19477 = n19377 ^ n19376 ;
  assign n19478 = n19477 ^ n616 ;
  assign n19535 = n19482 ^ n616 ;
  assign n19479 = n19375 ^ n19374 ;
  assign n19483 = n19482 ^ n19479 ;
  assign n19484 = n19373 ^ n19372 ;
  assign n19485 = n19484 ^ n1482 ;
  assign n2280 = n2204 ^ x409 ;
  assign n2281 = n2280 ^ n581 ;
  assign n2282 = n2281 ^ x345 ;
  assign n19514 = n19513 ^ n2282 ;
  assign n19507 = n19366 ^ n19365 ;
  assign n19486 = n19364 ^ n19363 ;
  assign n19490 = n19489 ^ n19486 ;
  assign n19491 = n19362 ^ n19361 ;
  assign n2137 = n2079 ^ x411 ;
  assign n2141 = n2140 ^ n2137 ;
  assign n2142 = n2141 ^ x347 ;
  assign n19492 = n19491 ^ n2142 ;
  assign n19493 = n19360 ^ n19358 ;
  assign n2033 = n1987 ^ x412 ;
  assign n2034 = n2033 ^ n2030 ;
  assign n2035 = n2034 ^ x348 ;
  assign n19494 = n19493 ^ n2035 ;
  assign n2024 = n1981 ^ x413 ;
  assign n2025 = n2024 ^ n1968 ;
  assign n2026 = n2025 ^ x349 ;
  assign n19497 = n19493 ^ n2026 ;
  assign n19055 = n19054 ^ n19053 ;
  assign n19056 = n19055 ^ n2026 ;
  assign n19008 = n19007 ^ n19004 ;
  assign n1959 = n1922 ^ x414 ;
  assign n1960 = n1959 ^ n1956 ;
  assign n1961 = n1960 ^ x350 ;
  assign n19009 = n19008 ^ n1961 ;
  assign n19011 = n19006 ^ n19005 ;
  assign n3056 = n3028 ^ x384 ;
  assign n3057 = n3056 ^ n3021 ;
  assign n3058 = n3057 ^ x320 ;
  assign n19010 = n3058 & n19005 ;
  assign n19012 = n19011 ^ n19010 ;
  assign n1950 = n1916 ^ x415 ;
  assign n1951 = n1950 ^ n1949 ;
  assign n1952 = n1951 ^ x351 ;
  assign n19073 = n19010 ^ n1952 ;
  assign n19016 = ~n19012 & n19073 ;
  assign n19013 = n1961 ^ n1952 ;
  assign n19017 = n19016 ^ n19013 ;
  assign n19018 = n19009 & ~n19017 ;
  assign n19019 = n19018 ^ n19008 ;
  assign n19495 = n19019 ^ n2026 ;
  assign n19496 = n19056 & n19495 ;
  assign n19498 = n19497 ^ n19496 ;
  assign n19499 = n19494 & n19498 ;
  assign n19500 = n19499 ^ n19493 ;
  assign n19501 = n19500 ^ n2142 ;
  assign n19502 = n19492 & ~n19501 ;
  assign n19503 = n19502 ^ n19491 ;
  assign n19504 = n19503 ^ n19486 ;
  assign n19505 = ~n19490 & n19504 ;
  assign n19506 = n19505 ^ n19489 ;
  assign n19508 = n19507 ^ n19506 ;
  assign n19509 = n19507 ^ n2282 ;
  assign n19510 = n19508 & ~n19509 ;
  assign n19515 = n19514 ^ n19510 ;
  assign n19519 = n19368 ^ n19367 ;
  assign n19516 = n19371 ^ n19369 ;
  assign n19517 = n19516 ^ n19513 ;
  assign n19518 = n19517 ^ n19516 ;
  assign n19520 = n19519 ^ n19518 ;
  assign n19521 = n19515 & n19520 ;
  assign n19522 = n19521 ^ n19517 ;
  assign n19527 = n19526 ^ n19484 ;
  assign n19523 = n19516 ^ n19484 ;
  assign n19528 = n19527 ^ n19523 ;
  assign n19529 = ~n19522 & n19528 ;
  assign n19530 = n19529 ^ n19527 ;
  assign n19531 = ~n19485 & ~n19530 ;
  assign n19532 = n19531 ^ n19484 ;
  assign n19533 = n19532 ^ n19482 ;
  assign n19534 = ~n19483 & ~n19533 ;
  assign n19536 = n19535 ^ n19534 ;
  assign n19537 = ~n19478 & n19536 ;
  assign n19538 = n19537 ^ n616 ;
  assign n19539 = n19538 ^ n19475 ;
  assign n19540 = n19476 & ~n19539 ;
  assign n19541 = n19540 ^ n557 ;
  assign n19542 = n19541 ^ n648 ;
  assign n19543 = ~n19474 & ~n19542 ;
  assign n19544 = n19543 ^ n19473 ;
  assign n19545 = n19544 ^ n1623 ;
  assign n19546 = ~n19472 & n19545 ;
  assign n19547 = n19546 ^ n19471 ;
  assign n19549 = n19548 ^ n19547 ;
  assign n19550 = n19469 ^ n728 ;
  assign n19551 = n19550 ^ n19469 ;
  assign n19552 = n19551 ^ n19547 ;
  assign n19553 = n19549 & ~n19552 ;
  assign n19554 = n19553 ^ n19550 ;
  assign n19555 = n19470 & n19554 ;
  assign n19556 = n19555 ^ n19469 ;
  assign n19557 = n19556 ^ n1021 ;
  assign n19558 = ~n19468 & n19557 ;
  assign n19560 = n19559 ^ n19558 ;
  assign n19326 = n19325 ^ n19250 ;
  assign n19232 = n18121 ^ n17640 ;
  assign n19233 = n19232 ^ n18681 ;
  assign n19224 = n18874 ^ n18800 ;
  assign n19228 = n19224 ^ n19107 ;
  assign n19227 = n19226 ^ n19224 ;
  assign n19229 = n19228 ^ n19227 ;
  assign n19230 = n19223 & n19229 ;
  assign n19231 = n19230 ^ n19228 ;
  assign n19327 = n19233 ^ n19231 ;
  assign n19328 = n19327 ^ n16862 ;
  assign n19329 = n19328 ^ n19250 ;
  assign n19330 = n19329 ^ n19327 ;
  assign n19331 = n19326 & ~n19330 ;
  assign n19332 = n19331 ^ n19328 ;
  assign n19388 = n19332 ^ n16949 ;
  assign n19387 = ~n19355 & n19386 ;
  assign n19561 = n19388 ^ n19387 ;
  assign n19562 = n19561 ^ n1167 ;
  assign n19563 = n19562 ^ n1036 ;
  assign n19564 = n19563 ^ n1167 ;
  assign n19565 = ~n19560 & ~n19564 ;
  assign n19566 = n19565 ^ n19562 ;
  assign n19389 = ~n19387 & ~n19388 ;
  assign n19099 = n18687 ^ n17587 ;
  assign n19100 = n19099 ^ n17636 ;
  assign n19235 = n19224 ^ n19100 ;
  assign n19234 = n19233 ^ n19100 ;
  assign n19236 = n19235 ^ n19234 ;
  assign n19237 = n19231 & ~n19236 ;
  assign n19238 = n19237 ^ n19235 ;
  assign n19098 = n18877 ^ n18798 ;
  assign n19248 = n19238 ^ n19098 ;
  assign n19334 = n19248 ^ n16949 ;
  assign n19333 = n19327 ^ n19248 ;
  assign n19335 = n19334 ^ n19333 ;
  assign n19336 = ~n19332 & n19335 ;
  assign n19337 = n19336 ^ n19334 ;
  assign n19353 = n19337 ^ n16956 ;
  assign n19465 = n19389 ^ n19353 ;
  assign n19914 = n19566 ^ n19465 ;
  assign n19409 = n18894 ^ n18893 ;
  assign n21309 = n19914 ^ n19409 ;
  assign n19778 = n18143 ^ n18102 ;
  assign n19779 = n19778 ^ n19114 ;
  assign n19059 = n19058 ^ n18148 ;
  assign n19060 = n19059 ^ n17883 ;
  assign n19057 = n19056 ^ n19019 ;
  assign n19061 = n19060 ^ n19057 ;
  assign n19068 = n19017 ^ n19008 ;
  assign n19066 = n19065 ^ n17877 ;
  assign n19067 = n19066 ^ n18156 ;
  assign n19069 = n19068 ^ n19067 ;
  assign n19074 = n19073 ^ n19011 ;
  assign n19071 = n19070 ^ n17869 ;
  assign n19072 = n19071 ^ n18512 ;
  assign n19075 = n19074 ^ n19072 ;
  assign n19079 = n19005 ^ n3058 ;
  assign n19077 = n19076 ^ n18162 ;
  assign n19078 = n19077 ^ n17593 ;
  assign n19080 = n19079 ^ n19078 ;
  assign n19402 = n18973 ^ n18451 ;
  assign n19403 = n19402 ^ n17803 ;
  assign n19401 = n18889 ^ n18790 ;
  assign n19404 = n19403 ^ n19401 ;
  assign n19410 = n19409 ^ n19401 ;
  assign n19411 = n19410 ^ n19409 ;
  assign n19085 = n18951 ^ n17725 ;
  assign n19086 = n19085 ^ n18359 ;
  assign n19084 = n18887 ^ n903 ;
  assign n19087 = n19086 ^ n19084 ;
  assign n19090 = n18883 ^ n18794 ;
  assign n19088 = n18323 ^ n17589 ;
  assign n19089 = n19088 ^ n18923 ;
  assign n19091 = n19090 ^ n19089 ;
  assign n19093 = n18704 ^ n17632 ;
  assign n19094 = n19093 ^ n18115 ;
  assign n19092 = n18880 ^ n18796 ;
  assign n19095 = n19094 ^ n19092 ;
  assign n19101 = n19100 ^ n19098 ;
  assign n19239 = ~n19101 & ~n19238 ;
  assign n19240 = n19239 ^ n19100 ;
  assign n19241 = n19240 ^ n19092 ;
  assign n19242 = ~n19095 & ~n19241 ;
  assign n19096 = n19092 ^ n19090 ;
  assign n19243 = n19242 ^ n19096 ;
  assign n19244 = n19091 & ~n19243 ;
  assign n19245 = n19244 ^ n19090 ;
  assign n19398 = n19245 ^ n19086 ;
  assign n19399 = ~n19087 & n19398 ;
  assign n19400 = n19399 ^ n19245 ;
  assign n19412 = n19411 ^ n19400 ;
  assign n19413 = n19404 & n19412 ;
  assign n19414 = n19413 ^ n19410 ;
  assign n19415 = n19032 ^ n17215 ;
  assign n19416 = n19415 ^ n17826 ;
  assign n19433 = n19416 ^ n19409 ;
  assign n19434 = ~n19414 & ~n19433 ;
  assign n19435 = n19434 ^ n19409 ;
  assign n19430 = n18788 ^ n1250 ;
  assign n19431 = n19430 ^ n18897 ;
  assign n19428 = n19155 ^ n17218 ;
  assign n19429 = n19428 ^ n17831 ;
  assign n19432 = n19431 ^ n19429 ;
  assign n19436 = n19435 ^ n19432 ;
  assign n19437 = n19436 ^ n16563 ;
  assign n19405 = n19404 ^ n19400 ;
  assign n19406 = n19405 ^ n17101 ;
  assign n19249 = n19248 ^ n16956 ;
  assign n19338 = n19249 & ~n19337 ;
  assign n19339 = n19338 ^ n16956 ;
  assign n19340 = n19339 ^ n16858 ;
  assign n19341 = n19240 ^ n19095 ;
  assign n19342 = n19341 ^ n19339 ;
  assign n19343 = ~n19340 & n19342 ;
  assign n19344 = n19343 ^ n16858 ;
  assign n19345 = n19344 ^ n16856 ;
  assign n19346 = n19243 ^ n19089 ;
  assign n19347 = n19346 ^ n19344 ;
  assign n19348 = ~n19345 & ~n19347 ;
  assign n19349 = n19348 ^ n16856 ;
  assign n19246 = n19245 ^ n19087 ;
  assign n19394 = n19349 ^ n19246 ;
  assign n19395 = n19349 ^ n16852 ;
  assign n19396 = ~n19394 & ~n19395 ;
  assign n19397 = n19396 ^ n16852 ;
  assign n19419 = n19405 ^ n19397 ;
  assign n19420 = n19406 & n19419 ;
  assign n19421 = n19420 ^ n17101 ;
  assign n19417 = n19416 ^ n19414 ;
  assign n19424 = n19421 ^ n19417 ;
  assign n19425 = n19421 ^ n16560 ;
  assign n19426 = n19424 & ~n19425 ;
  assign n19427 = n19426 ^ n16560 ;
  assign n19450 = n19436 ^ n19427 ;
  assign n19451 = n19437 & n19450 ;
  assign n19452 = n19451 ^ n16563 ;
  assign n19446 = n18470 ^ n17207 ;
  assign n19447 = n19446 ^ n17821 ;
  assign n19440 = n18903 ^ n2834 ;
  assign n19441 = n19440 ^ n19435 ;
  assign n19442 = n19441 ^ n19431 ;
  assign n19443 = n19442 ^ n19440 ;
  assign n19444 = n19432 & n19443 ;
  assign n19445 = n19444 ^ n19441 ;
  assign n19448 = n19447 ^ n19445 ;
  assign n19597 = n19452 ^ n19448 ;
  assign n19603 = n18905 ^ n18785 ;
  assign n19601 = n18478 ^ n17205 ;
  assign n19602 = n19601 ^ n17817 ;
  assign n19604 = n19603 ^ n19602 ;
  assign n19598 = n19447 ^ n19440 ;
  assign n19599 = n19445 & ~n19598 ;
  assign n19600 = n19599 ^ n19440 ;
  assign n19605 = n19604 ^ n19600 ;
  assign n19606 = n19605 ^ n16550 ;
  assign n19607 = n19606 ^ n19448 ;
  assign n19608 = n19607 ^ n19605 ;
  assign n19609 = ~n19597 & n19608 ;
  assign n19610 = n19609 ^ n19606 ;
  assign n19611 = n19610 ^ n16547 ;
  assign n19247 = n19246 ^ n16852 ;
  assign n19350 = n19349 ^ n19247 ;
  assign n19351 = n19346 ^ n19345 ;
  assign n19352 = n19341 ^ n19340 ;
  assign n19390 = ~n19353 & n19389 ;
  assign n19391 = n19352 & ~n19390 ;
  assign n19392 = ~n19351 & ~n19391 ;
  assign n19393 = n19350 & n19392 ;
  assign n19407 = n19406 ^ n19397 ;
  assign n19408 = ~n19393 & ~n19407 ;
  assign n19418 = n19417 ^ n16560 ;
  assign n19422 = n19421 ^ n19418 ;
  assign n19423 = ~n19408 & ~n19422 ;
  assign n19438 = n19437 ^ n19427 ;
  assign n19439 = n19423 & n19438 ;
  assign n19449 = n19448 ^ n16550 ;
  assign n19453 = n19452 ^ n19449 ;
  assign n19596 = n19439 & ~n19453 ;
  assign n19612 = n19611 ^ n19596 ;
  assign n19454 = n19453 ^ n19439 ;
  assign n3125 = n3121 ^ x389 ;
  assign n3126 = n3125 ^ n2462 ;
  assign n3127 = n3126 ^ x325 ;
  assign n19455 = n19454 ^ n3127 ;
  assign n19592 = n3127 ^ n1838 ;
  assign n19456 = n19438 ^ n19423 ;
  assign n19457 = n19456 ^ n3098 ;
  assign n19459 = n19407 ^ n19393 ;
  assign n19460 = n19459 ^ n3206 ;
  assign n19461 = n19392 ^ n19350 ;
  assign n19462 = n19461 ^ n2540 ;
  assign n19463 = n19391 ^ n19351 ;
  assign n19464 = n19463 ^ n1340 ;
  assign n19569 = n19390 ^ n19352 ;
  assign n19466 = n19465 ^ n1167 ;
  assign n19567 = n19466 & n19566 ;
  assign n19568 = n19567 ^ n19465 ;
  assign n19570 = n19569 ^ n19568 ;
  assign n19571 = n19569 ^ n1182 ;
  assign n19572 = n19570 & ~n19571 ;
  assign n19573 = n19572 ^ n1182 ;
  assign n19574 = n19573 ^ n19463 ;
  assign n19575 = ~n19464 & n19574 ;
  assign n19576 = n19575 ^ n1340 ;
  assign n19577 = n19576 ^ n19461 ;
  assign n19578 = ~n19462 & n19577 ;
  assign n19579 = n19578 ^ n2540 ;
  assign n19580 = n19579 ^ n19459 ;
  assign n19581 = n19460 & ~n19580 ;
  assign n19582 = n19581 ^ n3206 ;
  assign n19458 = n19422 ^ n19408 ;
  assign n19583 = n19582 ^ n19458 ;
  assign n19586 = n19458 ^ n2510 ;
  assign n19587 = n19583 & ~n19586 ;
  assign n19584 = n3098 ^ n2510 ;
  assign n19588 = n19587 ^ n19584 ;
  assign n19589 = ~n19457 & n19588 ;
  assign n19590 = n19589 ^ n3098 ;
  assign n19591 = n19590 ^ n1838 ;
  assign n19593 = n19592 ^ n19591 ;
  assign n19594 = n19455 & n19593 ;
  assign n19595 = n19594 ^ n19592 ;
  assign n19613 = n19612 ^ n19595 ;
  assign n19082 = n19081 ^ n18175 ;
  assign n19083 = n19082 ^ n17616 ;
  assign n19614 = n19613 ^ n19083 ;
  assign n19638 = n19590 ^ n19455 ;
  assign n19639 = n19145 ^ n17620 ;
  assign n19640 = n19639 ^ n18179 ;
  assign n19641 = n19638 & n19640 ;
  assign n19625 = n18908 ^ n18783 ;
  assign n19622 = n17811 ^ n17202 ;
  assign n19623 = n19622 ^ n18466 ;
  assign n19619 = n19602 ^ n19600 ;
  assign n19620 = ~n19604 & n19619 ;
  assign n19621 = n19620 ^ n19603 ;
  assign n19624 = n19623 ^ n19621 ;
  assign n19626 = n19625 ^ n19624 ;
  assign n19627 = n19626 ^ n16543 ;
  assign n19616 = n19605 ^ n16547 ;
  assign n19617 = ~n19610 & ~n19616 ;
  assign n19618 = n19617 ^ n16547 ;
  assign n19628 = n19627 ^ n19618 ;
  assign n19615 = ~n19596 & ~n19611 ;
  assign n19629 = n19628 ^ n19615 ;
  assign n19631 = n19629 ^ n1838 ;
  assign n19630 = n19629 ^ n19612 ;
  assign n19632 = n19631 ^ n19630 ;
  assign n19633 = n19595 & n19632 ;
  assign n19634 = n19633 ^ n19631 ;
  assign n19635 = n19634 ^ n2713 ;
  assign n19636 = n19635 ^ n19613 ;
  assign n19637 = n19636 ^ n19635 ;
  assign n19642 = n19641 ^ n19637 ;
  assign n19643 = ~n19614 & n19642 ;
  assign n19644 = n19643 ^ n19636 ;
  assign n19658 = n19626 ^ n19618 ;
  assign n19659 = ~n19627 & n19658 ;
  assign n19660 = n19659 ^ n16543 ;
  assign n19654 = n18464 ^ n17628 ;
  assign n19655 = n19654 ^ n16841 ;
  assign n19648 = n18911 ^ n18781 ;
  assign n19649 = n19648 ^ n19625 ;
  assign n19650 = n19649 ^ n19648 ;
  assign n19651 = n19650 ^ n19621 ;
  assign n19652 = ~n19624 & ~n19651 ;
  assign n19653 = n19652 ^ n19649 ;
  assign n19656 = n19655 ^ n19653 ;
  assign n19657 = n19656 ^ n16275 ;
  assign n19661 = n19660 ^ n19657 ;
  assign n19647 = ~n19615 & ~n19628 ;
  assign n19662 = n19661 ^ n19647 ;
  assign n19664 = n19662 ^ n19629 ;
  assign n19663 = n19662 ^ n2713 ;
  assign n19665 = n19664 ^ n19663 ;
  assign n19666 = n19634 & ~n19665 ;
  assign n19667 = n19666 ^ n19663 ;
  assign n19668 = n19667 ^ n2730 ;
  assign n19670 = n19668 ^ n19635 ;
  assign n19645 = n19136 ^ n17612 ;
  assign n19646 = n19645 ^ n18171 ;
  assign n19669 = n19668 ^ n19646 ;
  assign n19671 = n19670 ^ n19669 ;
  assign n19672 = ~n19644 & ~n19671 ;
  assign n19673 = n19672 ^ n19670 ;
  assign n19693 = n19647 & n19661 ;
  assign n19690 = n19655 ^ n19648 ;
  assign n19691 = ~n19653 & n19690 ;
  assign n19682 = n18776 ^ n2590 ;
  assign n19683 = n19682 ^ n18914 ;
  assign n19680 = n18460 ^ n17624 ;
  assign n19681 = n19680 ^ n17238 ;
  assign n19684 = n19683 ^ n19681 ;
  assign n19685 = n19684 ^ n19655 ;
  assign n19679 = n16275 ^ n16270 ;
  assign n19686 = n19685 ^ n19679 ;
  assign n19687 = n19686 ^ n3014 ;
  assign n19688 = n19687 ^ n2730 ;
  assign n19676 = n19660 ^ n19656 ;
  assign n19677 = n19660 ^ n16275 ;
  assign n19678 = n19676 & ~n19677 ;
  assign n19689 = n19688 ^ n19678 ;
  assign n19692 = n19691 ^ n19689 ;
  assign n19694 = n19693 ^ n19692 ;
  assign n19674 = n19662 ^ n2730 ;
  assign n19675 = n19667 & ~n19674 ;
  assign n19695 = n19694 ^ n19675 ;
  assign n19699 = n19695 ^ n19668 ;
  assign n19696 = n19134 ^ n17608 ;
  assign n19697 = n19696 ^ n18167 ;
  assign n19698 = n19697 ^ n19695 ;
  assign n19700 = n19699 ^ n19698 ;
  assign n19701 = n19673 & ~n19700 ;
  assign n19702 = n19701 ^ n19699 ;
  assign n19706 = n19695 ^ n19079 ;
  assign n19703 = n18160 ^ n17601 ;
  assign n19704 = n19703 ^ n19127 ;
  assign n19705 = n19704 ^ n19079 ;
  assign n19707 = n19706 ^ n19705 ;
  assign n19708 = ~n19702 & ~n19707 ;
  assign n19709 = n19708 ^ n19706 ;
  assign n19710 = ~n19080 & n19709 ;
  assign n19711 = n19710 ^ n19079 ;
  assign n19712 = n19711 ^ n19072 ;
  assign n19713 = n19075 & ~n19712 ;
  assign n19714 = n19713 ^ n19074 ;
  assign n19715 = n19714 ^ n19067 ;
  assign n19716 = ~n19069 & n19715 ;
  assign n19717 = n19716 ^ n19068 ;
  assign n19063 = n19062 ^ n18150 ;
  assign n19064 = n19063 ^ n18002 ;
  assign n19718 = n19717 ^ n19064 ;
  assign n19719 = n19718 ^ n19057 ;
  assign n19720 = n19719 ^ n19064 ;
  assign n19721 = n19061 & n19720 ;
  assign n19722 = n19721 ^ n19718 ;
  assign n19772 = n19501 ^ n19491 ;
  assign n19774 = n19772 ^ n19064 ;
  assign n19723 = n19498 ^ n2035 ;
  assign n19773 = n19772 ^ n19723 ;
  assign n19775 = n19774 ^ n19773 ;
  assign n19776 = n19722 & n19775 ;
  assign n19777 = n19776 ^ n19774 ;
  assign n19780 = n19779 ^ n19777 ;
  assign n19725 = n19714 ^ n19069 ;
  assign n19726 = n19725 ^ n16800 ;
  assign n19754 = n19711 ^ n19075 ;
  assign n19727 = n19709 ^ n19078 ;
  assign n19728 = n19727 ^ n16815 ;
  assign n19742 = n19697 ^ n19673 ;
  assign n19730 = n19640 ^ n19638 ;
  assign n19731 = n16837 & n19730 ;
  assign n19732 = n19731 ^ n16835 ;
  assign n19733 = n19641 ^ n19614 ;
  assign n19734 = n19733 ^ n19731 ;
  assign n19735 = n19732 & n19734 ;
  assign n19736 = n19735 ^ n16835 ;
  assign n19737 = n19736 ^ n16826 ;
  assign n19738 = n19646 ^ n19644 ;
  assign n19739 = n19738 ^ n19736 ;
  assign n19740 = ~n19737 & n19739 ;
  assign n19741 = n19740 ^ n16826 ;
  assign n19743 = n19742 ^ n19741 ;
  assign n19744 = n19742 ^ n17251 ;
  assign n19745 = n19743 & ~n19744 ;
  assign n19746 = n19745 ^ n17251 ;
  assign n19729 = n19704 ^ n19702 ;
  assign n19747 = n19746 ^ n19729 ;
  assign n19748 = n19746 ^ n16821 ;
  assign n19749 = n19747 & n19748 ;
  assign n19750 = n19749 ^ n16821 ;
  assign n19751 = n19750 ^ n19727 ;
  assign n19752 = n19728 & ~n19751 ;
  assign n19753 = n19752 ^ n16815 ;
  assign n19755 = n19754 ^ n19753 ;
  assign n19756 = n19725 ^ n16810 ;
  assign n19757 = n19756 ^ n19753 ;
  assign n19758 = n19757 ^ n19725 ;
  assign n19759 = n19755 & ~n19758 ;
  assign n19760 = n19759 ^ n19756 ;
  assign n19761 = n19726 & n19760 ;
  assign n19762 = n19761 ^ n16800 ;
  assign n19763 = n19762 ^ n17270 ;
  assign n19764 = n19717 ^ n19061 ;
  assign n19765 = n19764 ^ n19762 ;
  assign n19766 = ~n19763 & ~n19765 ;
  assign n19767 = n19766 ^ n17270 ;
  assign n19724 = n19723 ^ n19722 ;
  assign n19768 = n19767 ^ n19724 ;
  assign n19769 = n19767 ^ n17276 ;
  assign n19770 = ~n19768 & n19769 ;
  assign n19771 = n19770 ^ n17276 ;
  assign n19781 = n19780 ^ n19771 ;
  assign n19789 = n19503 ^ n19490 ;
  assign n19782 = n19110 ^ n18223 ;
  assign n19783 = n19782 ^ n18138 ;
  assign n19785 = n19783 ^ n19779 ;
  assign n19784 = n19783 ^ n19772 ;
  assign n19786 = n19785 ^ n19784 ;
  assign n19787 = n19777 & ~n19786 ;
  assign n19788 = n19787 ^ n19784 ;
  assign n19790 = n19789 ^ n19788 ;
  assign n19791 = n19790 ^ n16795 ;
  assign n19792 = n19791 ^ n19790 ;
  assign n19793 = n19792 ^ n19771 ;
  assign n19794 = n19781 & ~n19793 ;
  assign n19795 = n19794 ^ n19791 ;
  assign n19898 = n19790 ^ n16784 ;
  assign n19899 = ~n19795 & ~n19898 ;
  assign n19900 = n19899 ^ n16784 ;
  assign n19901 = n19900 ^ n17286 ;
  assign n19895 = n19103 ^ n18133 ;
  assign n19896 = n19895 ^ n18153 ;
  assign n19889 = n19509 ^ n19506 ;
  assign n19891 = n19889 ^ n19783 ;
  assign n19890 = n19889 ^ n19789 ;
  assign n19892 = n19891 ^ n19890 ;
  assign n19893 = n19788 & ~n19892 ;
  assign n19894 = n19893 ^ n19891 ;
  assign n19897 = n19896 ^ n19894 ;
  assign n19902 = n19901 ^ n19897 ;
  assign n19796 = n19795 ^ n16784 ;
  assign n19797 = n19750 ^ n19728 ;
  assign n19798 = n19729 ^ n16821 ;
  assign n19799 = n19798 ^ n19746 ;
  assign n19800 = n19744 ^ n19741 ;
  assign n19801 = n19730 ^ n16837 ;
  assign n19802 = n19733 ^ n19732 ;
  assign n19803 = n19801 & ~n19802 ;
  assign n19804 = n19738 ^ n19737 ;
  assign n19805 = n19803 & n19804 ;
  assign n19806 = n19800 & n19805 ;
  assign n19807 = n19799 & n19806 ;
  assign n19808 = n19797 & ~n19807 ;
  assign n19809 = n19754 ^ n16810 ;
  assign n19810 = n19809 ^ n19753 ;
  assign n19811 = ~n19808 & ~n19810 ;
  assign n19812 = n19760 ^ n16800 ;
  assign n19813 = ~n19811 & ~n19812 ;
  assign n19814 = n19764 ^ n19763 ;
  assign n19815 = n19813 & ~n19814 ;
  assign n19816 = n19724 ^ n17276 ;
  assign n19817 = n19816 ^ n19767 ;
  assign n19818 = n19815 & ~n19817 ;
  assign n19819 = n19780 ^ n16795 ;
  assign n19820 = n19819 ^ n19771 ;
  assign n19821 = ~n19818 & n19820 ;
  assign n19903 = ~n19796 & ~n19821 ;
  assign n20114 = n19902 & ~n19903 ;
  assign n19962 = n19896 ^ n19889 ;
  assign n19963 = ~n19894 & ~n19962 ;
  assign n19964 = n19963 ^ n19889 ;
  assign n19960 = n19519 ^ n19515 ;
  assign n19958 = n19107 ^ n18128 ;
  assign n19959 = n19958 ^ n18145 ;
  assign n19961 = n19960 ^ n19959 ;
  assign n20050 = n19964 ^ n19961 ;
  assign n20115 = n20050 ^ n17395 ;
  assign n20051 = n19900 ^ n19897 ;
  assign n20052 = ~n19901 & n20051 ;
  assign n20053 = n20052 ^ n17286 ;
  assign n20116 = n20115 ^ n20053 ;
  assign n20117 = ~n20114 & ~n20116 ;
  assign n20054 = n20053 ^ n20050 ;
  assign n20055 = n20053 ^ n17395 ;
  assign n20056 = ~n20054 & ~n20055 ;
  assign n20057 = n20056 ^ n17395 ;
  assign n19965 = n19964 ^ n19959 ;
  assign n19966 = n19961 & n19965 ;
  assign n19967 = n19966 ^ n19960 ;
  assign n19956 = n19526 ^ n19522 ;
  assign n19954 = n18237 ^ n18123 ;
  assign n19955 = n19954 ^ n19224 ;
  assign n19957 = n19956 ^ n19955 ;
  assign n20048 = n19967 ^ n19957 ;
  assign n20049 = n20048 ^ n17407 ;
  assign n20118 = n20057 ^ n20049 ;
  assign n20119 = n20117 & n20118 ;
  assign n19968 = n19967 ^ n19955 ;
  assign n19969 = ~n19957 & n19968 ;
  assign n19970 = n19969 ^ n19956 ;
  assign n19949 = n19098 ^ n18140 ;
  assign n19950 = n19949 ^ n18113 ;
  assign n19948 = n19530 ^ n1482 ;
  assign n19951 = n19950 ^ n19948 ;
  assign n20047 = n19970 ^ n19951 ;
  assign n20120 = n20047 ^ n17578 ;
  assign n20058 = n20057 ^ n20048 ;
  assign n20059 = ~n20049 & n20058 ;
  assign n20060 = n20059 ^ n17407 ;
  assign n20121 = n20120 ^ n20060 ;
  assign n20122 = n20119 & ~n20121 ;
  assign n20061 = n20060 ^ n20047 ;
  assign n20062 = n20060 ^ n17578 ;
  assign n20063 = n20061 & ~n20062 ;
  assign n20064 = n20063 ^ n17578 ;
  assign n19971 = n19970 ^ n19948 ;
  assign n19972 = ~n19951 & ~n19971 ;
  assign n19945 = n19092 ^ n18555 ;
  assign n19946 = n19945 ^ n18136 ;
  assign n19952 = n19948 ^ n19946 ;
  assign n19973 = n19972 ^ n19952 ;
  assign n19944 = n19532 ^ n19483 ;
  assign n20045 = n19973 ^ n19944 ;
  assign n20046 = n20045 ^ n17652 ;
  assign n20123 = n20064 ^ n20046 ;
  assign n20124 = n20122 & n20123 ;
  assign n19947 = n19946 ^ n19944 ;
  assign n19974 = ~n19947 & n19973 ;
  assign n19975 = n19974 ^ n19946 ;
  assign n19942 = n19536 ^ n19477 ;
  assign n19940 = n19090 ^ n18131 ;
  assign n19941 = n19940 ^ n18681 ;
  assign n19943 = n19942 ^ n19941 ;
  assign n20044 = n19975 ^ n19943 ;
  assign n20112 = n20044 ^ n17647 ;
  assign n20065 = n20064 ^ n20045 ;
  assign n20066 = n20046 & n20065 ;
  assign n20067 = n20066 ^ n17652 ;
  assign n20113 = n20112 ^ n20067 ;
  assign n20163 = n20124 ^ n20113 ;
  assign n20164 = n20163 ^ n790 ;
  assign n20168 = n20123 ^ n20122 ;
  assign n20169 = n20168 ^ n781 ;
  assign n20170 = n20121 ^ n20119 ;
  assign n20171 = n20170 ^ n713 ;
  assign n20172 = n20118 ^ n20117 ;
  assign n20173 = n20172 ^ n704 ;
  assign n20183 = n1534 ^ n704 ;
  assign n19904 = n19903 ^ n19902 ;
  assign n19822 = n19821 ^ n19796 ;
  assign n19823 = n19822 ^ n2933 ;
  assign n19824 = n19820 ^ n19818 ;
  assign n19828 = n19827 ^ n19824 ;
  assign n19829 = n19817 ^ n19815 ;
  assign n19830 = n19829 ^ n590 ;
  assign n19831 = n19812 ^ n19811 ;
  assign n19873 = n19831 ^ n2377 ;
  assign n19832 = n19831 ^ n2368 ;
  assign n19833 = n19810 ^ n19808 ;
  assign n19834 = n19833 ^ n2228 ;
  assign n19864 = n19807 ^ n19797 ;
  assign n19837 = n19806 ^ n19799 ;
  assign n19838 = n19837 ^ n2115 ;
  assign n19839 = n19805 ^ n19800 ;
  assign n2103 = n2048 ^ x445 ;
  assign n2107 = n2106 ^ n2103 ;
  assign n2108 = n2107 ^ x381 ;
  assign n19840 = n19839 ^ n2108 ;
  assign n19842 = n3087 ^ x446 ;
  assign n19843 = n19842 ^ n1898 ;
  assign n19844 = n19843 ^ x382 ;
  assign n19857 = n19844 ^ n2108 ;
  assign n19841 = n19804 ^ n19803 ;
  assign n19845 = n19844 ^ n19841 ;
  assign n19847 = n19802 ^ n19801 ;
  assign n19854 = n19847 ^ n19844 ;
  assign n19846 = n1793 & ~n19801 ;
  assign n19848 = n19847 ^ n19846 ;
  assign n19849 = n3070 ^ x447 ;
  assign n19850 = n19849 ^ n14844 ;
  assign n19851 = n19850 ^ x383 ;
  assign n19852 = n19851 ^ n19846 ;
  assign n19853 = ~n19848 & ~n19852 ;
  assign n19855 = n19854 ^ n19853 ;
  assign n19856 = n19845 & ~n19855 ;
  assign n19858 = n19857 ^ n19856 ;
  assign n19859 = n19840 & n19858 ;
  assign n19860 = n19859 ^ n2108 ;
  assign n19861 = n19860 ^ n2115 ;
  assign n19862 = n19838 & ~n19861 ;
  assign n19863 = n19862 ^ n19837 ;
  assign n19865 = n19864 ^ n19863 ;
  assign n19866 = n19864 ^ n2130 ;
  assign n19867 = ~n19865 & n19866 ;
  assign n19868 = n19867 ^ n2130 ;
  assign n19835 = n19831 ^ n2228 ;
  assign n19836 = n19835 ^ n19831 ;
  assign n19869 = n19868 ^ n19836 ;
  assign n19870 = n19834 & n19869 ;
  assign n19871 = n19870 ^ n19835 ;
  assign n19872 = ~n19832 & ~n19871 ;
  assign n19874 = n19873 ^ n19872 ;
  assign n19877 = n2377 ^ n590 ;
  assign n19875 = n19814 ^ n19813 ;
  assign n19876 = n19875 ^ n590 ;
  assign n19878 = n19877 ^ n19876 ;
  assign n19879 = ~n19874 & n19878 ;
  assign n19880 = n19879 ^ n19877 ;
  assign n19881 = n19830 & n19880 ;
  assign n19882 = n19881 ^ n590 ;
  assign n19883 = n19882 ^ n19824 ;
  assign n19884 = ~n19828 & n19883 ;
  assign n19885 = n19884 ^ n19827 ;
  assign n19886 = n19885 ^ n2933 ;
  assign n19887 = ~n19823 & ~n19886 ;
  assign n19888 = n19887 ^ n19822 ;
  assign n20174 = n19904 ^ n19888 ;
  assign n20177 = n19888 ^ n1525 ;
  assign n20178 = ~n20174 & ~n20177 ;
  assign n20175 = n1534 ^ n1525 ;
  assign n20179 = n20178 ^ n20175 ;
  assign n20180 = n20116 ^ n20114 ;
  assign n20181 = n20180 ^ n1534 ;
  assign n20182 = n20179 & ~n20181 ;
  assign n20184 = n20183 ^ n20182 ;
  assign n20185 = ~n20173 & ~n20184 ;
  assign n20186 = n20185 ^ n20172 ;
  assign n20187 = n20186 ^ n713 ;
  assign n20188 = n20171 & n20187 ;
  assign n20189 = n20188 ^ n20170 ;
  assign n20190 = n20189 ^ n781 ;
  assign n20191 = ~n20169 & ~n20190 ;
  assign n20192 = n20191 ^ n20168 ;
  assign n20068 = n20067 ^ n20044 ;
  assign n20069 = n20067 ^ n17647 ;
  assign n20070 = n20068 & ~n20069 ;
  assign n20071 = n20070 ^ n17647 ;
  assign n20126 = n20071 ^ n17645 ;
  assign n19938 = n19538 ^ n19476 ;
  assign n19976 = n19975 ^ n19938 ;
  assign n19977 = n19976 ^ n19941 ;
  assign n19978 = n19977 ^ n19938 ;
  assign n19979 = ~n19943 & n19978 ;
  assign n19980 = n19979 ^ n19976 ;
  assign n19936 = n18687 ^ n18126 ;
  assign n19937 = n19936 ^ n19084 ;
  assign n20072 = n19980 ^ n19937 ;
  assign n20127 = n20126 ^ n20072 ;
  assign n20125 = n20113 & ~n20124 ;
  assign n20165 = n20127 ^ n20125 ;
  assign n20166 = n20165 ^ n790 ;
  assign n20167 = n20166 ^ n20165 ;
  assign n20193 = n20192 ^ n20167 ;
  assign n20194 = ~n20164 & ~n20193 ;
  assign n20195 = n20194 ^ n20166 ;
  assign n20479 = n20195 ^ n915 ;
  assign n21310 = n21309 ^ n20479 ;
  assign n20540 = n19107 ^ n18138 ;
  assign n20541 = n20540 ^ n19944 ;
  assign n20514 = n19960 ^ n19114 ;
  assign n20515 = n20514 ^ n18148 ;
  assign n20472 = n19858 ^ n19839 ;
  assign n20516 = n20515 ^ n20472 ;
  assign n20423 = n19855 ^ n19841 ;
  assign n20374 = n19852 ^ n19847 ;
  assign n20424 = n20423 ^ n20374 ;
  assign n20372 = n19789 ^ n19058 ;
  assign n20373 = n20372 ^ n18512 ;
  assign n20375 = n20374 ^ n20373 ;
  assign n20357 = n19801 ^ n1793 ;
  assign n20021 = n18466 ^ n17821 ;
  assign n20022 = n20021 ^ n18937 ;
  assign n20015 = n19573 ^ n19464 ;
  assign n20008 = n19571 ^ n19568 ;
  assign n20016 = n20015 ^ n20008 ;
  assign n20009 = n20008 ^ n19914 ;
  assign n19912 = n19648 ^ n17826 ;
  assign n19913 = n19912 ^ n18470 ;
  assign n19915 = n19914 ^ n19913 ;
  assign n19918 = n19561 ^ n19560 ;
  assign n19916 = n19625 ^ n19155 ;
  assign n19917 = n19916 ^ n18451 ;
  assign n19919 = n19918 ^ n19917 ;
  assign n19922 = n19556 ^ n19468 ;
  assign n19920 = n19603 ^ n18359 ;
  assign n19921 = n19920 ^ n19032 ;
  assign n19923 = n19922 ^ n19921 ;
  assign n19926 = n19554 ^ n1015 ;
  assign n19999 = n19926 ^ n19922 ;
  assign n19924 = n19440 ^ n18973 ;
  assign n19925 = n19924 ^ n18323 ;
  assign n19927 = n19926 ^ n19925 ;
  assign n19930 = n19548 ^ n728 ;
  assign n19931 = n19930 ^ n19547 ;
  assign n19928 = n19431 ^ n18951 ;
  assign n19929 = n19928 ^ n18115 ;
  assign n19932 = n19931 ^ n19929 ;
  assign n19985 = n19544 ^ n19472 ;
  assign n19908 = n19541 ^ n19474 ;
  assign n19986 = n19985 ^ n19908 ;
  assign n19933 = n19401 ^ n18704 ;
  assign n19934 = n19933 ^ n18121 ;
  assign n19935 = n19934 ^ n19908 ;
  assign n19939 = n19938 ^ n19937 ;
  assign n19981 = ~n19939 & ~n19980 ;
  assign n19982 = n19981 ^ n19938 ;
  assign n19983 = n19982 ^ n19908 ;
  assign n19984 = ~n19935 & ~n19983 ;
  assign n19987 = n19986 ^ n19984 ;
  assign n19990 = n18923 ^ n17587 ;
  assign n19991 = n19990 ^ n19409 ;
  assign n19992 = n19991 ^ n19985 ;
  assign n19993 = ~n19987 & ~n19992 ;
  assign n19988 = n19985 ^ n19929 ;
  assign n19994 = n19993 ^ n19988 ;
  assign n19995 = n19932 & n19994 ;
  assign n19996 = n19995 ^ n19931 ;
  assign n19997 = n19996 ^ n19926 ;
  assign n19998 = n19927 & ~n19997 ;
  assign n20000 = n19999 ^ n19998 ;
  assign n20001 = n19923 & ~n20000 ;
  assign n20002 = n20001 ^ n19922 ;
  assign n20003 = n20002 ^ n19917 ;
  assign n20004 = ~n19919 & n20003 ;
  assign n20005 = n20004 ^ n19918 ;
  assign n20006 = n20005 ^ n19914 ;
  assign n20007 = n19915 & n20006 ;
  assign n20010 = n20009 ^ n20007 ;
  assign n20011 = n19683 ^ n18478 ;
  assign n20012 = n20011 ^ n17831 ;
  assign n20013 = n20012 ^ n20008 ;
  assign n20014 = n20010 & n20013 ;
  assign n20017 = n20016 ^ n20014 ;
  assign n20030 = n20022 ^ n20017 ;
  assign n20031 = n20030 ^ n17207 ;
  assign n20032 = n20012 ^ n20010 ;
  assign n20033 = n20032 ^ n17218 ;
  assign n20098 = n20005 ^ n19915 ;
  assign n20034 = n20002 ^ n19919 ;
  assign n20035 = n20034 ^ n17803 ;
  assign n20036 = n20000 ^ n19921 ;
  assign n20037 = n20036 ^ n17725 ;
  assign n20087 = n19996 ^ n19927 ;
  assign n20038 = n19994 ^ n19931 ;
  assign n20039 = n20038 ^ n17632 ;
  assign n20040 = n19991 ^ n19987 ;
  assign n20041 = n20040 ^ n17636 ;
  assign n20042 = n19982 ^ n19935 ;
  assign n20043 = n20042 ^ n17640 ;
  assign n20073 = n20072 ^ n20071 ;
  assign n20074 = n20042 ^ n17645 ;
  assign n20075 = n20074 ^ n20042 ;
  assign n20076 = n20075 ^ n20071 ;
  assign n20077 = n20073 & n20076 ;
  assign n20078 = n20077 ^ n20074 ;
  assign n20079 = ~n20043 & ~n20078 ;
  assign n20080 = n20079 ^ n17640 ;
  assign n20081 = n20080 ^ n20040 ;
  assign n20082 = ~n20041 & ~n20081 ;
  assign n20083 = n20082 ^ n17636 ;
  assign n20084 = n20083 ^ n20038 ;
  assign n20085 = n20039 & n20084 ;
  assign n20086 = n20085 ^ n17632 ;
  assign n20088 = n20087 ^ n20086 ;
  assign n20089 = n20087 ^ n17589 ;
  assign n20090 = n20088 & n20089 ;
  assign n20091 = n20090 ^ n17589 ;
  assign n20092 = n20091 ^ n20036 ;
  assign n20093 = n20037 & n20092 ;
  assign n20094 = n20093 ^ n17725 ;
  assign n20095 = n20094 ^ n20034 ;
  assign n20096 = n20035 & ~n20095 ;
  assign n20097 = n20096 ^ n17803 ;
  assign n20099 = n20098 ^ n20097 ;
  assign n20100 = n20098 ^ n17215 ;
  assign n20101 = n20099 & ~n20100 ;
  assign n20102 = n20101 ^ n17215 ;
  assign n20103 = n20102 ^ n20032 ;
  assign n20104 = ~n20033 & n20103 ;
  assign n20105 = n20104 ^ n17218 ;
  assign n20106 = n20105 ^ n20030 ;
  assign n20107 = ~n20031 & n20106 ;
  assign n20108 = n20107 ^ n17207 ;
  assign n20026 = n18464 ^ n17817 ;
  assign n20027 = n20026 ^ n18962 ;
  assign n20018 = n19576 ^ n19462 ;
  assign n20019 = n20018 ^ n20015 ;
  assign n20020 = n20019 ^ n20018 ;
  assign n20023 = n20022 ^ n20020 ;
  assign n20024 = n20017 & n20023 ;
  assign n20025 = n20024 ^ n20019 ;
  assign n20028 = n20027 ^ n20025 ;
  assign n20029 = n20028 ^ n17205 ;
  assign n20109 = n20108 ^ n20029 ;
  assign n20110 = n20091 ^ n20037 ;
  assign n20111 = n20089 ^ n20086 ;
  assign n20128 = n20125 & n20127 ;
  assign n20129 = n20078 ^ n17640 ;
  assign n20130 = ~n20128 & ~n20129 ;
  assign n20131 = n20080 ^ n17636 ;
  assign n20132 = n20131 ^ n20040 ;
  assign n20133 = n20130 & n20132 ;
  assign n20134 = n20083 ^ n20039 ;
  assign n20135 = ~n20133 & ~n20134 ;
  assign n20136 = ~n20111 & ~n20135 ;
  assign n20137 = n20110 & n20136 ;
  assign n20138 = n20094 ^ n20035 ;
  assign n20139 = ~n20137 & n20138 ;
  assign n20140 = n20100 ^ n20097 ;
  assign n20141 = ~n20139 & n20140 ;
  assign n20142 = n20102 ^ n20033 ;
  assign n20143 = n20141 & n20142 ;
  assign n20144 = n20105 ^ n20031 ;
  assign n20145 = n20143 & n20144 ;
  assign n20250 = n20109 & ~n20145 ;
  assign n20245 = n18460 ^ n17811 ;
  assign n20246 = n20245 ^ n18990 ;
  assign n20239 = n19579 ^ n19460 ;
  assign n20241 = n20239 ^ n20018 ;
  assign n20240 = n20239 ^ n20027 ;
  assign n20242 = n20241 ^ n20240 ;
  assign n20243 = n20025 & ~n20242 ;
  assign n20244 = n20243 ^ n20241 ;
  assign n20247 = n20246 ^ n20244 ;
  assign n20248 = n20247 ^ n17202 ;
  assign n20236 = n20108 ^ n20028 ;
  assign n20237 = n20029 & ~n20236 ;
  assign n20238 = n20237 ^ n17205 ;
  assign n20249 = n20248 ^ n20238 ;
  assign n20251 = n20250 ^ n20249 ;
  assign n20252 = n20251 ^ n2474 ;
  assign n20280 = n20238 ^ n17202 ;
  assign n20281 = n20247 ^ n20238 ;
  assign n20282 = ~n20280 & n20281 ;
  assign n20283 = n20282 ^ n20247 ;
  assign n20284 = n20283 ^ n16841 ;
  assign n20277 = n18186 ^ n17628 ;
  assign n20278 = n20277 ^ n19047 ;
  assign n20270 = n19582 ^ n2510 ;
  assign n20271 = n20270 ^ n19458 ;
  assign n20273 = n20271 ^ n20239 ;
  assign n20272 = n20271 ^ n20246 ;
  assign n20274 = n20273 ^ n20272 ;
  assign n20275 = ~n20244 & ~n20274 ;
  assign n20276 = n20275 ^ n20273 ;
  assign n20279 = n20278 ^ n20276 ;
  assign n20285 = n20284 ^ n20279 ;
  assign n20269 = ~n20249 & ~n20250 ;
  assign n20286 = n20285 ^ n20269 ;
  assign n20287 = n20286 ^ n2474 ;
  assign n20288 = n20287 ^ n20286 ;
  assign n20146 = n20145 ^ n20109 ;
  assign n20147 = n20146 ^ n3166 ;
  assign n20227 = n20144 ^ n20143 ;
  assign n20148 = n20142 ^ n20141 ;
  assign n20149 = n20148 ^ n2627 ;
  assign n20218 = n20140 ^ n20139 ;
  assign n20150 = n20138 ^ n20137 ;
  assign n20151 = n20150 ^ n2827 ;
  assign n20152 = n20136 ^ n20110 ;
  assign n20153 = n20152 ^ n2816 ;
  assign n20155 = n20134 ^ n20133 ;
  assign n20156 = n20155 ^ n1313 ;
  assign n20157 = n20132 ^ n20130 ;
  assign n1065 = n980 ^ x428 ;
  assign n1066 = n1065 ^ n1061 ;
  assign n1067 = n1066 ^ x364 ;
  assign n20158 = n20157 ^ n1067 ;
  assign n20161 = n20129 ^ n20128 ;
  assign n1293 = n1193 ^ x429 ;
  assign n1294 = n1293 ^ n896 ;
  assign n1295 = n1294 ^ x365 ;
  assign n20162 = n20161 ^ n1295 ;
  assign n20197 = n20161 ^ n915 ;
  assign n20196 = n20165 ^ n20161 ;
  assign n20198 = n20197 ^ n20196 ;
  assign n20199 = ~n20195 & n20198 ;
  assign n20200 = n20199 ^ n20197 ;
  assign n20201 = ~n20162 & ~n20200 ;
  assign n20202 = n20201 ^ n20161 ;
  assign n20159 = n20155 ^ n1067 ;
  assign n20160 = n20159 ^ n20155 ;
  assign n20203 = n20202 ^ n20160 ;
  assign n20204 = ~n20158 & ~n20203 ;
  assign n20205 = n20204 ^ n20159 ;
  assign n20206 = n20156 & ~n20205 ;
  assign n20207 = n20206 ^ n1313 ;
  assign n20211 = n20207 ^ n20152 ;
  assign n20154 = n20135 ^ n20111 ;
  assign n20208 = n20207 ^ n20154 ;
  assign n20209 = n20154 ^ n1331 ;
  assign n20210 = ~n20208 & n20209 ;
  assign n20212 = n20211 ^ n20210 ;
  assign n20213 = ~n20153 & n20212 ;
  assign n20214 = n20213 ^ n2816 ;
  assign n20215 = n20214 ^ n20150 ;
  assign n20216 = ~n20151 & n20215 ;
  assign n20217 = n20216 ^ n2827 ;
  assign n20219 = n20218 ^ n20217 ;
  assign n2560 = n2553 ^ x423 ;
  assign n2564 = n2563 ^ n2560 ;
  assign n2565 = n2564 ^ x359 ;
  assign n20220 = n20148 ^ n2565 ;
  assign n20221 = n20220 ^ n20148 ;
  assign n20222 = n20221 ^ n20217 ;
  assign n20223 = ~n20219 & n20222 ;
  assign n20224 = n20223 ^ n20220 ;
  assign n20225 = ~n20149 & n20224 ;
  assign n20226 = n20225 ^ n2627 ;
  assign n20228 = n20227 ^ n20226 ;
  assign n20229 = n20146 ^ n2492 ;
  assign n20230 = n20229 ^ n20146 ;
  assign n20231 = n20230 ^ n20226 ;
  assign n20232 = n20228 & n20231 ;
  assign n20233 = n20232 ^ n20229 ;
  assign n20234 = ~n20147 & n20233 ;
  assign n20235 = n20234 ^ n3166 ;
  assign n20289 = n20288 ^ n20235 ;
  assign n20290 = ~n20252 & n20289 ;
  assign n20291 = n20290 ^ n20287 ;
  assign n20340 = n20286 ^ n1823 ;
  assign n20341 = n20291 & ~n20340 ;
  assign n20336 = n20278 ^ n20271 ;
  assign n20337 = n20276 & n20336 ;
  assign n20330 = n3176 ^ x417 ;
  assign n20331 = n20330 ^ n1799 ;
  assign n20332 = n20331 ^ x353 ;
  assign n20333 = n20332 ^ n1823 ;
  assign n20328 = n17238 ^ n16841 ;
  assign n20324 = n19167 ^ n18184 ;
  assign n20325 = n20324 ^ n17624 ;
  assign n20326 = n20325 ^ n20278 ;
  assign n20323 = n19588 ^ n19456 ;
  assign n20327 = n20326 ^ n20323 ;
  assign n20329 = n20328 ^ n20327 ;
  assign n20334 = n20333 ^ n20329 ;
  assign n20320 = n20279 ^ n16841 ;
  assign n20321 = n20283 ^ n20279 ;
  assign n20322 = ~n20320 & ~n20321 ;
  assign n20335 = n20334 ^ n20322 ;
  assign n20338 = n20337 ^ n20335 ;
  assign n20319 = n20269 & n20285 ;
  assign n20339 = n20338 ^ n20319 ;
  assign n20342 = n20341 ^ n20339 ;
  assign n20358 = n20357 ^ n20342 ;
  assign n20317 = n19723 ^ n19070 ;
  assign n20318 = n20317 ^ n18160 ;
  assign n20343 = n20342 ^ n20318 ;
  assign n20292 = n20291 ^ n1823 ;
  assign n20253 = n20252 ^ n20235 ;
  assign n20293 = n20292 ^ n20253 ;
  assign n19910 = n19127 ^ n19068 ;
  assign n19911 = n19910 ^ n18171 ;
  assign n20254 = n20253 ^ n19911 ;
  assign n20257 = n20227 ^ n2492 ;
  assign n20258 = n20257 ^ n20226 ;
  assign n20259 = n19079 ^ n18179 ;
  assign n20260 = n20259 ^ n19136 ;
  assign n20261 = ~n20258 & ~n20260 ;
  assign n20255 = n19134 ^ n18175 ;
  assign n20256 = n20255 ^ n19074 ;
  assign n20262 = n20261 ^ n20256 ;
  assign n20263 = n20233 ^ n3166 ;
  assign n20264 = n20263 ^ n20256 ;
  assign n20265 = ~n20262 & n20264 ;
  assign n20266 = n20265 ^ n20256 ;
  assign n20267 = n20266 ^ n20253 ;
  assign n20268 = ~n20254 & n20267 ;
  assign n20294 = n20293 ^ n20268 ;
  assign n20295 = n19076 ^ n19057 ;
  assign n20296 = n20295 ^ n18167 ;
  assign n20314 = n20296 ^ n20292 ;
  assign n20315 = ~n20294 & ~n20314 ;
  assign n20316 = n20315 ^ n20296 ;
  assign n20355 = n20342 ^ n20316 ;
  assign n20356 = ~n20343 & ~n20355 ;
  assign n20359 = n20358 ^ n20356 ;
  assign n20360 = n19772 ^ n18162 ;
  assign n20361 = n20360 ^ n19065 ;
  assign n20369 = n20361 ^ n20357 ;
  assign n20370 = n20359 & ~n20369 ;
  assign n20371 = n20370 ^ n20357 ;
  assign n20421 = n20374 ^ n20371 ;
  assign n20422 = n20375 & n20421 ;
  assign n20425 = n20424 ^ n20422 ;
  assign n20426 = n19889 ^ n19062 ;
  assign n20427 = n20426 ^ n18156 ;
  assign n20520 = n20427 ^ n20423 ;
  assign n20521 = ~n20425 & n20520 ;
  assign n20522 = n20521 ^ n20427 ;
  assign n20517 = n19860 ^ n19838 ;
  assign n20518 = n20517 ^ n20472 ;
  assign n20519 = n20518 ^ n20517 ;
  assign n20523 = n20522 ^ n20519 ;
  assign n20524 = ~n20516 & ~n20523 ;
  assign n20525 = n20524 ^ n20518 ;
  assign n20468 = n19866 ^ n19863 ;
  assign n20529 = n20517 ^ n20468 ;
  assign n20526 = n19110 ^ n18150 ;
  assign n20527 = n20526 ^ n19956 ;
  assign n20528 = n20527 ^ n20468 ;
  assign n20530 = n20529 ^ n20528 ;
  assign n20531 = n20525 & n20530 ;
  assign n20532 = n20531 ^ n20529 ;
  assign n20462 = n19868 ^ n19834 ;
  assign n20536 = n20468 ^ n20462 ;
  assign n20533 = n19103 ^ n18143 ;
  assign n20534 = n20533 ^ n19948 ;
  assign n20535 = n20534 ^ n20462 ;
  assign n20537 = n20536 ^ n20535 ;
  assign n20538 = n20532 & ~n20537 ;
  assign n20539 = n20538 ^ n20536 ;
  assign n20602 = n20541 ^ n20539 ;
  assign n20603 = n20602 ^ n18223 ;
  assign n20604 = n20534 ^ n20532 ;
  assign n20605 = n20604 ^ n18102 ;
  assign n20606 = n20527 ^ n20525 ;
  assign n20607 = n20606 ^ n18002 ;
  assign n20428 = n20427 ^ n20425 ;
  assign n20429 = n20428 ^ n17877 ;
  assign n20362 = n20361 ^ n20359 ;
  assign n20363 = n20362 ^ n17593 ;
  assign n20344 = n20343 ^ n20316 ;
  assign n20345 = n20344 ^ n17601 ;
  assign n20297 = n20296 ^ n20294 ;
  assign n20298 = n20297 ^ n17608 ;
  assign n20299 = n20266 ^ n20254 ;
  assign n20300 = n20299 ^ n17612 ;
  assign n20302 = n20260 ^ n20258 ;
  assign n20303 = n17620 & n20302 ;
  assign n20301 = n20263 ^ n20262 ;
  assign n20304 = n20303 ^ n20301 ;
  assign n20305 = n20303 ^ n17616 ;
  assign n20306 = ~n20304 & ~n20305 ;
  assign n20307 = n20306 ^ n17616 ;
  assign n20308 = n20307 ^ n20299 ;
  assign n20309 = n20300 & n20308 ;
  assign n20310 = n20309 ^ n17612 ;
  assign n20311 = n20310 ^ n20297 ;
  assign n20312 = n20298 & ~n20311 ;
  assign n20313 = n20312 ^ n17608 ;
  assign n20364 = n20344 ^ n20313 ;
  assign n20365 = ~n20345 & n20364 ;
  assign n20366 = n20365 ^ n17601 ;
  assign n20378 = n20366 ^ n20362 ;
  assign n20379 = ~n20363 & ~n20378 ;
  assign n20380 = n20379 ^ n17593 ;
  assign n20376 = n20375 ^ n20371 ;
  assign n20417 = n20380 ^ n20376 ;
  assign n20418 = n20380 ^ n17869 ;
  assign n20419 = ~n20417 & ~n20418 ;
  assign n20420 = n20419 ^ n17869 ;
  assign n20609 = n20428 ^ n20420 ;
  assign n20610 = ~n20429 & n20609 ;
  assign n20611 = n20610 ^ n17877 ;
  assign n20608 = n20522 ^ n20516 ;
  assign n20612 = n20611 ^ n20608 ;
  assign n20613 = n20611 ^ n17883 ;
  assign n20614 = ~n20612 & n20613 ;
  assign n20615 = n20614 ^ n17883 ;
  assign n20616 = n20615 ^ n20606 ;
  assign n20617 = n20607 & ~n20616 ;
  assign n20618 = n20617 ^ n18002 ;
  assign n20619 = n20618 ^ n20604 ;
  assign n20620 = n20605 & n20619 ;
  assign n20621 = n20620 ^ n18102 ;
  assign n20622 = n20621 ^ n20602 ;
  assign n20623 = n20603 & n20622 ;
  assign n20624 = n20623 ^ n18223 ;
  assign n20547 = n19942 ^ n18133 ;
  assign n20548 = n20547 ^ n19224 ;
  assign n20458 = n19871 ^ n2368 ;
  assign n20543 = n20462 ^ n20458 ;
  assign n20542 = n20541 ^ n20458 ;
  assign n20544 = n20543 ^ n20542 ;
  assign n20545 = n20539 & n20544 ;
  assign n20546 = n20545 ^ n20543 ;
  assign n20600 = n20548 ^ n20546 ;
  assign n20601 = n20600 ^ n18153 ;
  assign n20692 = n20624 ^ n20601 ;
  assign n20682 = n20608 ^ n17883 ;
  assign n20683 = n20682 ^ n20611 ;
  assign n20346 = n20345 ^ n20313 ;
  assign n20347 = n20307 ^ n20300 ;
  assign n20348 = n20302 ^ n17620 ;
  assign n20349 = n20305 ^ n20301 ;
  assign n20350 = n20348 & ~n20349 ;
  assign n20351 = ~n20347 & n20350 ;
  assign n20352 = n20310 ^ n20298 ;
  assign n20353 = n20351 & n20352 ;
  assign n20354 = ~n20346 & n20353 ;
  assign n20367 = n20366 ^ n20363 ;
  assign n20368 = ~n20354 & n20367 ;
  assign n20377 = n20376 ^ n17869 ;
  assign n20381 = n20380 ^ n20377 ;
  assign n20416 = ~n20368 & n20381 ;
  assign n20430 = n20429 ^ n20420 ;
  assign n20684 = ~n20416 & n20430 ;
  assign n20685 = ~n20683 & n20684 ;
  assign n20686 = n20615 ^ n20607 ;
  assign n20687 = n20685 & ~n20686 ;
  assign n20688 = n20618 ^ n20605 ;
  assign n20689 = ~n20687 & n20688 ;
  assign n20690 = n20621 ^ n20603 ;
  assign n20691 = ~n20689 & n20690 ;
  assign n20753 = n20692 ^ n20691 ;
  assign n20754 = n20753 ^ n2947 ;
  assign n20755 = n20690 ^ n20689 ;
  assign n20756 = n20755 ^ n578 ;
  assign n20757 = n20688 ^ n20687 ;
  assign n20761 = n20760 ^ n20757 ;
  assign n20762 = n20686 ^ n20685 ;
  assign n20763 = n20762 ^ n1469 ;
  assign n20769 = n20684 ^ n20683 ;
  assign n20770 = n20769 ^ n20768 ;
  assign n20431 = n20430 ^ n20416 ;
  assign n20432 = n20431 ^ n2347 ;
  assign n20771 = n20769 ^ n2347 ;
  assign n20772 = n20771 ^ n20769 ;
  assign n20382 = n20381 ^ n20368 ;
  assign n20383 = n20382 ^ n2321 ;
  assign n20384 = n20367 ^ n20354 ;
  assign n20385 = n20384 ^ n2328 ;
  assign n2016 = n1976 ^ x476 ;
  assign n2020 = n2019 ^ n2016 ;
  assign n2021 = n2020 ^ x412 ;
  assign n20409 = n20384 ^ n2021 ;
  assign n20386 = n20353 ^ n20346 ;
  assign n20387 = n20386 ^ n2021 ;
  assign n20391 = n20352 ^ n20351 ;
  assign n20388 = n18828 ^ x477 ;
  assign n20389 = n20388 ^ n1942 ;
  assign n20390 = n20389 ^ x413 ;
  assign n20392 = n20391 ^ n20390 ;
  assign n1880 = n1858 ^ x448 ;
  assign n1884 = n1883 ^ n1880 ;
  assign n1885 = n1884 ^ x384 ;
  assign n20393 = n1885 & ~n20348 ;
  assign n1892 = n1867 ^ x479 ;
  assign n1893 = n1892 ^ n1889 ;
  assign n1894 = n1893 ^ x415 ;
  assign n20394 = n20393 ^ n1894 ;
  assign n20395 = n20349 ^ n20348 ;
  assign n20396 = n20395 ^ n1894 ;
  assign n20397 = n20394 & n20396 ;
  assign n20398 = n20397 ^ n20393 ;
  assign n1933 = n1905 ^ x478 ;
  assign n1937 = n1936 ^ n1933 ;
  assign n1938 = n1937 ^ x414 ;
  assign n20399 = n20398 ^ n1938 ;
  assign n20400 = n20350 ^ n20347 ;
  assign n20401 = n20400 ^ n1938 ;
  assign n20402 = n20399 & ~n20401 ;
  assign n20403 = n20402 ^ n1938 ;
  assign n20404 = n20403 ^ n20390 ;
  assign n20405 = n20392 & ~n20404 ;
  assign n20406 = n20405 ^ n20391 ;
  assign n20407 = n20406 ^ n2021 ;
  assign n20408 = ~n20387 & n20407 ;
  assign n20410 = n20409 ^ n20408 ;
  assign n20411 = n20385 & ~n20410 ;
  assign n20412 = n20411 ^ n2328 ;
  assign n20413 = n20412 ^ n20382 ;
  assign n20414 = ~n20383 & n20413 ;
  assign n20415 = n20414 ^ n2321 ;
  assign n20773 = n20772 ^ n20415 ;
  assign n20774 = n20432 & n20773 ;
  assign n20775 = n20774 ^ n20771 ;
  assign n20776 = n20770 & n20775 ;
  assign n20777 = n20776 ^ n20769 ;
  assign n20764 = n20757 ^ n1469 ;
  assign n20765 = n20764 ^ n20757 ;
  assign n20778 = n20777 ^ n20765 ;
  assign n20779 = n20763 & n20778 ;
  assign n20780 = n20779 ^ n20764 ;
  assign n20781 = ~n20761 & n20780 ;
  assign n20782 = n20781 ^ n20760 ;
  assign n20783 = n20782 ^ n20755 ;
  assign n20784 = n20756 & ~n20783 ;
  assign n20785 = n20784 ^ n578 ;
  assign n20786 = n20785 ^ n20753 ;
  assign n20787 = ~n20754 & n20786 ;
  assign n20788 = n20787 ^ n2947 ;
  assign n20625 = n20624 ^ n20600 ;
  assign n20626 = n20601 & n20625 ;
  assign n20627 = n20626 ^ n18153 ;
  assign n20453 = n19875 ^ n19874 ;
  assign n20550 = n20458 ^ n20453 ;
  assign n20549 = n20548 ^ n20453 ;
  assign n20551 = n20550 ^ n20549 ;
  assign n20552 = ~n20546 & ~n20551 ;
  assign n20553 = n20552 ^ n20550 ;
  assign n20511 = n19938 ^ n19098 ;
  assign n20512 = n20511 ^ n18128 ;
  assign n20598 = n20553 ^ n20512 ;
  assign n20599 = n20598 ^ n18145 ;
  assign n20694 = n20627 ^ n20599 ;
  assign n20693 = ~n20691 & n20692 ;
  assign n20749 = n20694 ^ n20693 ;
  assign n20750 = n20749 ^ n533 ;
  assign n21308 = n20788 ^ n20750 ;
  assign n21311 = n21310 ^ n21308 ;
  assign n21314 = n20785 ^ n20754 ;
  assign n21321 = n21314 ^ n21308 ;
  assign n21312 = n19918 ^ n19401 ;
  assign n20475 = n20192 ^ n20164 ;
  assign n21313 = n21312 ^ n20475 ;
  assign n21315 = n21314 ^ n21313 ;
  assign n21248 = n20782 ^ n20756 ;
  assign n21246 = n19922 ^ n19084 ;
  assign n20482 = n20189 ^ n20169 ;
  assign n21247 = n21246 ^ n20482 ;
  assign n21249 = n21248 ^ n21247 ;
  assign n21133 = n20780 ^ n20760 ;
  assign n21125 = n20777 ^ n20763 ;
  assign n21134 = n21133 ^ n21125 ;
  assign n20492 = n20184 ^ n20172 ;
  assign n21123 = n20492 ^ n19092 ;
  assign n21124 = n21123 ^ n19931 ;
  assign n21126 = n21125 ^ n21124 ;
  assign n21015 = n20775 ^ n20768 ;
  assign n20433 = n20432 ^ n20415 ;
  assign n21016 = n21015 ^ n20433 ;
  assign n19905 = n19904 ^ n1525 ;
  assign n19906 = n19905 ^ n19888 ;
  assign n19907 = n19906 ^ n19224 ;
  assign n19909 = n19908 ^ n19907 ;
  assign n20434 = n20433 ^ n19909 ;
  assign n20438 = n20412 ^ n20383 ;
  assign n20435 = n19885 ^ n19823 ;
  assign n20436 = n20435 ^ n19107 ;
  assign n20437 = n20436 ^ n19938 ;
  assign n20439 = n20438 ^ n20437 ;
  assign n20443 = n20410 ^ n2328 ;
  assign n20441 = n19882 ^ n19828 ;
  assign n20440 = n19942 ^ n19103 ;
  assign n20442 = n20441 ^ n20440 ;
  assign n20444 = n20443 ^ n20442 ;
  assign n20450 = n20406 ^ n20387 ;
  assign n20448 = n19880 ^ n19829 ;
  assign n20447 = n19944 ^ n19110 ;
  assign n20449 = n20448 ^ n20447 ;
  assign n20451 = n20450 ^ n20449 ;
  assign n20452 = n20403 ^ n20392 ;
  assign n21004 = n20452 ^ n20450 ;
  assign n20454 = n20453 ^ n19114 ;
  assign n20455 = n20454 ^ n19948 ;
  assign n20456 = n20455 ^ n20452 ;
  assign n20459 = n20458 ^ n19956 ;
  assign n20460 = n20459 ^ n19062 ;
  assign n20457 = n20401 ^ n20398 ;
  assign n20461 = n20460 ^ n20457 ;
  assign n20465 = n20395 ^ n20394 ;
  assign n20998 = n20465 ^ n20457 ;
  assign n20463 = n20462 ^ n19058 ;
  assign n20464 = n20463 ^ n19960 ;
  assign n20466 = n20465 ^ n20464 ;
  assign n20469 = n20468 ^ n19065 ;
  assign n20470 = n20469 ^ n19889 ;
  assign n20467 = n20348 ^ n1885 ;
  assign n20471 = n20470 ^ n20467 ;
  assign n20966 = n19789 ^ n19070 ;
  assign n20967 = n20966 ^ n20517 ;
  assign n20486 = n20186 ^ n20171 ;
  assign n20572 = n20492 ^ n20486 ;
  assign n20490 = n19918 ^ n19431 ;
  assign n20491 = n20490 ^ n18704 ;
  assign n20493 = n20492 ^ n20491 ;
  assign n20495 = n19922 ^ n18687 ;
  assign n20496 = n20495 ^ n19409 ;
  assign n20494 = n20180 ^ n20179 ;
  assign n20497 = n20496 ^ n20494 ;
  assign n20566 = n20494 ^ n19906 ;
  assign n20498 = n19926 ^ n18681 ;
  assign n20499 = n20498 ^ n19401 ;
  assign n20500 = n20499 ^ n19906 ;
  assign n20501 = n19931 ^ n18555 ;
  assign n20502 = n20501 ^ n19084 ;
  assign n20503 = n20502 ^ n20435 ;
  assign n20560 = n20441 ^ n20435 ;
  assign n20504 = n19985 ^ n18113 ;
  assign n20505 = n20504 ^ n19090 ;
  assign n20506 = n20505 ^ n20441 ;
  assign n20507 = n19092 ^ n18123 ;
  assign n20508 = n20507 ^ n19908 ;
  assign n20557 = n20508 ^ n20441 ;
  assign n20509 = n20508 ^ n20448 ;
  assign n20513 = n20512 ^ n20453 ;
  assign n20554 = ~n20513 & n20553 ;
  assign n20510 = n20453 ^ n20448 ;
  assign n20555 = n20554 ^ n20510 ;
  assign n20556 = ~n20509 & n20555 ;
  assign n20558 = n20557 ^ n20556 ;
  assign n20559 = ~n20506 & n20558 ;
  assign n20561 = n20560 ^ n20559 ;
  assign n20562 = ~n20503 & n20561 ;
  assign n20563 = n20562 ^ n20435 ;
  assign n20564 = n20563 ^ n20499 ;
  assign n20565 = n20500 & n20564 ;
  assign n20567 = n20566 ^ n20565 ;
  assign n20568 = ~n20497 & n20567 ;
  assign n20569 = n20568 ^ n20496 ;
  assign n20570 = n20569 ^ n20492 ;
  assign n20571 = ~n20493 & ~n20570 ;
  assign n20573 = n20572 ^ n20571 ;
  assign n20487 = n19440 ^ n18923 ;
  assign n20488 = n20487 ^ n19914 ;
  assign n20651 = n20573 ^ n20488 ;
  assign n20588 = n20569 ^ n20493 ;
  assign n20589 = n20588 ^ n18121 ;
  assign n20643 = n20567 ^ n20496 ;
  assign n20590 = n20563 ^ n20500 ;
  assign n20591 = n20590 ^ n18131 ;
  assign n20592 = n20561 ^ n20502 ;
  assign n20593 = n20592 ^ n18136 ;
  assign n20594 = n20558 ^ n20505 ;
  assign n20595 = n20594 ^ n18140 ;
  assign n20596 = n20555 ^ n20508 ;
  assign n20597 = n20596 ^ n18237 ;
  assign n20628 = n20627 ^ n20598 ;
  assign n20629 = n20599 & n20628 ;
  assign n20630 = n20629 ^ n18145 ;
  assign n20631 = n20630 ^ n20596 ;
  assign n20632 = ~n20597 & ~n20631 ;
  assign n20633 = n20632 ^ n18237 ;
  assign n20634 = n20633 ^ n20594 ;
  assign n20635 = ~n20595 & n20634 ;
  assign n20636 = n20635 ^ n18140 ;
  assign n20637 = n20636 ^ n20592 ;
  assign n20638 = ~n20593 & n20637 ;
  assign n20639 = n20638 ^ n18136 ;
  assign n20640 = n20639 ^ n20590 ;
  assign n20641 = n20591 & ~n20640 ;
  assign n20642 = n20641 ^ n18131 ;
  assign n20644 = n20643 ^ n20642 ;
  assign n20645 = n20643 ^ n18126 ;
  assign n20646 = ~n20644 & n20645 ;
  assign n20647 = n20646 ^ n18126 ;
  assign n20648 = n20647 ^ n20588 ;
  assign n20649 = ~n20589 & ~n20648 ;
  assign n20650 = n20649 ^ n18121 ;
  assign n20652 = n20651 ^ n20650 ;
  assign n20653 = n20651 ^ n17587 ;
  assign n20654 = n20652 & n20653 ;
  assign n20655 = n20654 ^ n17587 ;
  assign n20489 = n20488 ^ n20486 ;
  assign n20574 = n20489 & ~n20573 ;
  assign n20575 = n20574 ^ n20488 ;
  assign n20483 = n20008 ^ n18951 ;
  assign n20484 = n20483 ^ n19603 ;
  assign n20485 = n20484 ^ n20482 ;
  assign n20586 = n20575 ^ n20485 ;
  assign n20587 = n20586 ^ n18115 ;
  assign n20678 = n20655 ^ n20587 ;
  assign n20679 = n20653 ^ n20650 ;
  assign n20680 = n20647 ^ n20589 ;
  assign n20681 = n20645 ^ n20642 ;
  assign n20695 = ~n20693 & n20694 ;
  assign n20696 = n20630 ^ n18237 ;
  assign n20697 = n20696 ^ n20596 ;
  assign n20698 = n20695 & n20697 ;
  assign n20699 = n20633 ^ n18140 ;
  assign n20700 = n20699 ^ n20594 ;
  assign n20701 = n20698 & ~n20700 ;
  assign n20702 = n20636 ^ n20593 ;
  assign n20703 = n20701 & ~n20702 ;
  assign n20704 = n20639 ^ n20591 ;
  assign n20705 = ~n20703 & ~n20704 ;
  assign n20706 = ~n20681 & n20705 ;
  assign n20707 = ~n20680 & ~n20706 ;
  assign n20708 = ~n20679 & n20707 ;
  assign n20709 = ~n20678 & ~n20708 ;
  assign n20576 = n20575 ^ n20482 ;
  assign n20577 = ~n20485 & n20576 ;
  assign n20578 = n20577 ^ n20482 ;
  assign n20476 = n20015 ^ n19625 ;
  assign n20477 = n20476 ^ n18973 ;
  assign n20478 = n20477 ^ n20475 ;
  assign n20659 = n20578 ^ n20478 ;
  assign n20661 = n20659 ^ n18323 ;
  assign n20656 = n20655 ^ n20586 ;
  assign n20657 = n20587 & n20656 ;
  assign n20658 = n20657 ^ n18115 ;
  assign n20710 = n20661 ^ n20658 ;
  assign n20711 = ~n20709 & n20710 ;
  assign n20660 = n20659 ^ n20658 ;
  assign n20662 = n20660 & ~n20661 ;
  assign n20663 = n20662 ^ n18323 ;
  assign n20582 = n20018 ^ n19032 ;
  assign n20583 = n20582 ^ n19648 ;
  assign n20480 = n20479 ^ n20475 ;
  assign n20481 = n20480 ^ n20479 ;
  assign n20579 = n20578 ^ n20481 ;
  assign n20580 = n20478 & ~n20579 ;
  assign n20581 = n20580 ^ n20480 ;
  assign n20584 = n20583 ^ n20581 ;
  assign n20585 = n20584 ^ n18359 ;
  assign n20712 = n20663 ^ n20585 ;
  assign n20713 = n20711 & n20712 ;
  assign n20673 = n19683 ^ n19155 ;
  assign n20674 = n20673 ^ n20239 ;
  assign n20667 = n20200 ^ n1295 ;
  assign n20669 = n20667 ^ n20479 ;
  assign n20668 = n20667 ^ n20583 ;
  assign n20670 = n20669 ^ n20668 ;
  assign n20671 = n20581 & ~n20670 ;
  assign n20672 = n20671 ^ n20669 ;
  assign n20675 = n20674 ^ n20672 ;
  assign n20676 = n20675 ^ n18451 ;
  assign n20664 = n20663 ^ n20584 ;
  assign n20665 = ~n20585 & n20664 ;
  assign n20666 = n20665 ^ n18359 ;
  assign n20677 = n20676 ^ n20666 ;
  assign n20730 = n20713 ^ n20677 ;
  assign n2884 = n2841 ^ x456 ;
  assign n2885 = n2884 ^ n2504 ;
  assign n2886 = n2885 ^ x392 ;
  assign n20731 = n20730 ^ n2886 ;
  assign n20732 = n20712 ^ n20711 ;
  assign n20733 = n20732 ^ n2879 ;
  assign n20735 = n20708 ^ n20678 ;
  assign n1137 = n1055 ^ x459 ;
  assign n1141 = n1140 ^ n1137 ;
  assign n1142 = n1141 ^ x395 ;
  assign n20736 = n20735 ^ n1142 ;
  assign n20809 = n20707 ^ n20679 ;
  assign n20737 = n20706 ^ n20680 ;
  assign n20738 = n20737 ^ n995 ;
  assign n20805 = n20737 ^ n891 ;
  assign n20739 = n20705 ^ n20681 ;
  assign n20740 = n20739 ^ n891 ;
  assign n20741 = n20704 ^ n20703 ;
  assign n20742 = n20741 ^ n876 ;
  assign n20743 = n20702 ^ n20701 ;
  assign n20744 = n20743 ^ n867 ;
  assign n20745 = n20700 ^ n20698 ;
  assign n20746 = n20745 ^ n1589 ;
  assign n20747 = n20697 ^ n20695 ;
  assign n20748 = n20747 ^ n1583 ;
  assign n20751 = n20747 ^ n533 ;
  assign n20752 = n20751 ^ n20747 ;
  assign n20789 = n20788 ^ n20752 ;
  assign n20790 = n20750 & n20789 ;
  assign n20791 = n20790 ^ n20751 ;
  assign n20792 = ~n20748 & ~n20791 ;
  assign n20793 = n20792 ^ n20747 ;
  assign n20794 = n20793 ^ n1589 ;
  assign n20795 = n20746 & n20794 ;
  assign n20796 = n20795 ^ n20745 ;
  assign n20797 = n20796 ^ n867 ;
  assign n20798 = n20744 & ~n20797 ;
  assign n20799 = n20798 ^ n20743 ;
  assign n20800 = n20799 ^ n876 ;
  assign n20801 = n20742 & ~n20800 ;
  assign n20802 = n20801 ^ n20741 ;
  assign n20803 = n20802 ^ n891 ;
  assign n20804 = ~n20740 & n20803 ;
  assign n20806 = n20805 ^ n20804 ;
  assign n20807 = ~n20738 & ~n20806 ;
  assign n20808 = n20807 ^ n20737 ;
  assign n20810 = n20809 ^ n20808 ;
  assign n20811 = n20735 ^ n1145 ;
  assign n20812 = n20811 ^ n20735 ;
  assign n20813 = n20812 ^ n20808 ;
  assign n20814 = n20810 & ~n20813 ;
  assign n20815 = n20814 ^ n20811 ;
  assign n20816 = n20736 & ~n20815 ;
  assign n20817 = n20816 ^ n1142 ;
  assign n20734 = n20710 ^ n20709 ;
  assign n20818 = n20817 ^ n20734 ;
  assign n20819 = n20732 ^ n1349 ;
  assign n20820 = n20819 ^ n20732 ;
  assign n20821 = n20820 ^ n20734 ;
  assign n20822 = ~n20818 & n20821 ;
  assign n20823 = n20822 ^ n20819 ;
  assign n20824 = ~n20733 & n20823 ;
  assign n20825 = n20824 ^ n2879 ;
  assign n20826 = n20825 ^ n20730 ;
  assign n20827 = n20731 & ~n20826 ;
  assign n20828 = n20827 ^ n2886 ;
  assign n20725 = n20675 ^ n20666 ;
  assign n20726 = ~n20676 & ~n20725 ;
  assign n20727 = n20726 ^ n18451 ;
  assign n20721 = n20271 ^ n18470 ;
  assign n20722 = n20721 ^ n18937 ;
  assign n20715 = n20202 ^ n20158 ;
  assign n20717 = n20715 ^ n20667 ;
  assign n20716 = n20715 ^ n20674 ;
  assign n20718 = n20717 ^ n20716 ;
  assign n20719 = ~n20672 & n20718 ;
  assign n20720 = n20719 ^ n20717 ;
  assign n20723 = n20722 ^ n20720 ;
  assign n20724 = n20723 ^ n17826 ;
  assign n20728 = n20727 ^ n20724 ;
  assign n20714 = ~n20677 & ~n20713 ;
  assign n20729 = n20728 ^ n20714 ;
  assign n20829 = n20828 ^ n20729 ;
  assign n20841 = n20323 ^ n18962 ;
  assign n20842 = n20841 ^ n18478 ;
  assign n20835 = n20205 ^ n1313 ;
  assign n20837 = n20835 ^ n20715 ;
  assign n20836 = n20835 ^ n20722 ;
  assign n20838 = n20837 ^ n20836 ;
  assign n20839 = ~n20720 & ~n20838 ;
  assign n20840 = n20839 ^ n20837 ;
  assign n20843 = n20842 ^ n20840 ;
  assign n20844 = n20843 ^ n17831 ;
  assign n20831 = n20727 ^ n20723 ;
  assign n20832 = n20727 ^ n17826 ;
  assign n20833 = n20831 & ~n20832 ;
  assign n20834 = n20833 ^ n17826 ;
  assign n20845 = n20844 ^ n20834 ;
  assign n20830 = ~n20714 & n20728 ;
  assign n20846 = n20845 ^ n20830 ;
  assign n20847 = n20846 ^ n2901 ;
  assign n20848 = n20847 ^ n20729 ;
  assign n20849 = n20848 ^ n20846 ;
  assign n20850 = ~n20829 & n20849 ;
  assign n20851 = n20850 ^ n20847 ;
  assign n20869 = n18780 ^ x454 ;
  assign n20870 = n20869 ^ n3115 ;
  assign n20871 = n20870 ^ x390 ;
  assign n20862 = n19638 ^ n18466 ;
  assign n20863 = n20862 ^ n18990 ;
  assign n20856 = n20209 ^ n20207 ;
  assign n20858 = n20856 ^ n20835 ;
  assign n20857 = n20856 ^ n20842 ;
  assign n20859 = n20858 ^ n20857 ;
  assign n20860 = n20840 & n20859 ;
  assign n20861 = n20860 ^ n20858 ;
  assign n20864 = n20863 ^ n20861 ;
  assign n20865 = n20864 ^ n17821 ;
  assign n20853 = n20843 ^ n20834 ;
  assign n20854 = ~n20844 & ~n20853 ;
  assign n20855 = n20854 ^ n17831 ;
  assign n20866 = n20865 ^ n20855 ;
  assign n20852 = n20830 & n20845 ;
  assign n20867 = n20866 ^ n20852 ;
  assign n20872 = n20871 ^ n20867 ;
  assign n20868 = n20867 ^ n20846 ;
  assign n20873 = n20872 ^ n20868 ;
  assign n20874 = n20851 & ~n20873 ;
  assign n20875 = n20874 ^ n20872 ;
  assign n20887 = n20864 ^ n20855 ;
  assign n20888 = ~n20865 & n20887 ;
  assign n20889 = n20888 ^ n17821 ;
  assign n20883 = n19613 ^ n19047 ;
  assign n20884 = n20883 ^ n18464 ;
  assign n20877 = n20212 ^ n2816 ;
  assign n20879 = n20877 ^ n20856 ;
  assign n20878 = n20877 ^ n20863 ;
  assign n20880 = n20879 ^ n20878 ;
  assign n20881 = ~n20861 & n20880 ;
  assign n20882 = n20881 ^ n20879 ;
  assign n20885 = n20884 ^ n20882 ;
  assign n20886 = n20885 ^ n17817 ;
  assign n20890 = n20889 ^ n20886 ;
  assign n20876 = n20852 & ~n20866 ;
  assign n20891 = n20890 ^ n20876 ;
  assign n2603 = n2590 ^ x453 ;
  assign n2604 = n2603 ^ n1832 ;
  assign n2605 = n2604 ^ x389 ;
  assign n20893 = n20891 ^ n2605 ;
  assign n20892 = n20891 ^ n20867 ;
  assign n20894 = n20893 ^ n20892 ;
  assign n20895 = ~n20875 & n20894 ;
  assign n20896 = n20895 ^ n20893 ;
  assign n20912 = ~n20876 & ~n20890 ;
  assign n20907 = n19635 ^ n18460 ;
  assign n20908 = n20907 ^ n19167 ;
  assign n20901 = n20214 ^ n20151 ;
  assign n20903 = n20901 ^ n20877 ;
  assign n20902 = n20901 ^ n20884 ;
  assign n20904 = n20903 ^ n20902 ;
  assign n20905 = n20882 & ~n20904 ;
  assign n20906 = n20905 ^ n20903 ;
  assign n20909 = n20908 ^ n20906 ;
  assign n20910 = n20909 ^ n17811 ;
  assign n20897 = n20889 ^ n20885 ;
  assign n20898 = n20889 ^ n17817 ;
  assign n20899 = n20897 & ~n20898 ;
  assign n20900 = n20899 ^ n17817 ;
  assign n20911 = n20910 ^ n20900 ;
  assign n20913 = n20912 ^ n20911 ;
  assign n20915 = n20913 ^ n2611 ;
  assign n20914 = n20913 ^ n20891 ;
  assign n20916 = n20915 ^ n20914 ;
  assign n20917 = ~n20896 & n20916 ;
  assign n20918 = n20917 ^ n20915 ;
  assign n20930 = n20909 ^ n20900 ;
  assign n20931 = ~n20910 & n20930 ;
  assign n20932 = n20931 ^ n17811 ;
  assign n20933 = n20932 ^ n17628 ;
  assign n20927 = n19668 ^ n19145 ;
  assign n20928 = n20927 ^ n18186 ;
  assign n20920 = n20218 ^ n2565 ;
  assign n20921 = n20920 ^ n20217 ;
  assign n20923 = n20921 ^ n20901 ;
  assign n20922 = n20921 ^ n20908 ;
  assign n20924 = n20923 ^ n20922 ;
  assign n20925 = n20906 & n20924 ;
  assign n20926 = n20925 ^ n20923 ;
  assign n20929 = n20928 ^ n20926 ;
  assign n20934 = n20933 ^ n20929 ;
  assign n20919 = n20911 & ~n20912 ;
  assign n20935 = n20934 ^ n20919 ;
  assign n20937 = n20935 ^ n20913 ;
  assign n20936 = n20935 ^ n2701 ;
  assign n20938 = n20937 ^ n20936 ;
  assign n20939 = ~n20918 & n20938 ;
  assign n20940 = n20939 ^ n20936 ;
  assign n20941 = n20940 ^ n2690 ;
  assign n20473 = n20472 ^ n19772 ;
  assign n20474 = n20473 ^ n19076 ;
  assign n20942 = n20941 ^ n20474 ;
  assign n20945 = n20357 ^ n19068 ;
  assign n20946 = n20945 ^ n19136 ;
  assign n20947 = n20875 ^ n2605 ;
  assign n20948 = ~n20946 & n20947 ;
  assign n20943 = n20374 ^ n19134 ;
  assign n20944 = n20943 ^ n19057 ;
  assign n20949 = n20948 ^ n20944 ;
  assign n20952 = n20896 ^ n2611 ;
  assign n20950 = n20918 ^ n2701 ;
  assign n20951 = n20950 ^ n20944 ;
  assign n20953 = n20952 ^ n20951 ;
  assign n20954 = n20953 ^ n20950 ;
  assign n20955 = ~n20949 & ~n20954 ;
  assign n20956 = n20955 ^ n20951 ;
  assign n20960 = n20950 ^ n20941 ;
  assign n20957 = n19723 ^ n19127 ;
  assign n20958 = n20957 ^ n20423 ;
  assign n20959 = n20958 ^ n20941 ;
  assign n20961 = n20960 ^ n20959 ;
  assign n20962 = ~n20956 & ~n20961 ;
  assign n20963 = n20962 ^ n20960 ;
  assign n20964 = ~n20942 & ~n20963 ;
  assign n20965 = n20964 ^ n20941 ;
  assign n20968 = n20967 ^ n20965 ;
  assign n20986 = n20935 ^ n2690 ;
  assign n20987 = n20940 & ~n20986 ;
  assign n20981 = n3000 ^ n2690 ;
  assign n20979 = n17628 ^ n17624 ;
  assign n20977 = n20224 ^ n2627 ;
  assign n20974 = n19695 ^ n19081 ;
  assign n20975 = n20974 ^ n18184 ;
  assign n20976 = n20975 ^ n20928 ;
  assign n20978 = n20977 ^ n20976 ;
  assign n20980 = n20979 ^ n20978 ;
  assign n20982 = n20981 ^ n20980 ;
  assign n20972 = n20932 ^ n20929 ;
  assign n20973 = n20933 & n20972 ;
  assign n20983 = n20982 ^ n20973 ;
  assign n20970 = n20928 ^ n20921 ;
  assign n20971 = n20926 & n20970 ;
  assign n20984 = n20983 ^ n20971 ;
  assign n20969 = n20919 & n20934 ;
  assign n20985 = n20984 ^ n20969 ;
  assign n20988 = n20987 ^ n20985 ;
  assign n20991 = n20988 ^ n20965 ;
  assign n20992 = n20968 & n20991 ;
  assign n20989 = n20988 ^ n20467 ;
  assign n20993 = n20992 ^ n20989 ;
  assign n20994 = n20471 & ~n20993 ;
  assign n20995 = n20994 ^ n20470 ;
  assign n20996 = n20995 ^ n20465 ;
  assign n20997 = n20466 & n20996 ;
  assign n20999 = n20998 ^ n20997 ;
  assign n21000 = ~n20461 & ~n20999 ;
  assign n21001 = n21000 ^ n20460 ;
  assign n21002 = n21001 ^ n20452 ;
  assign n21003 = ~n20456 & n21002 ;
  assign n21005 = n21004 ^ n21003 ;
  assign n21006 = n20451 & ~n21005 ;
  assign n21007 = n21006 ^ n20450 ;
  assign n21008 = n21007 ^ n20443 ;
  assign n21009 = ~n20444 & ~n21008 ;
  assign n20445 = n20443 ^ n20438 ;
  assign n21010 = n21009 ^ n20445 ;
  assign n21011 = ~n20439 & ~n21010 ;
  assign n21012 = n21011 ^ n20438 ;
  assign n21013 = n21012 ^ n19909 ;
  assign n21014 = n20434 & n21013 ;
  assign n21017 = n21016 ^ n21014 ;
  assign n21018 = n19985 ^ n19098 ;
  assign n21019 = n21018 ^ n20494 ;
  assign n21120 = n21019 ^ n21015 ;
  assign n21121 = n21017 & n21120 ;
  assign n21122 = n21121 ^ n21015 ;
  assign n21131 = n21125 ^ n21122 ;
  assign n21132 = ~n21126 & n21131 ;
  assign n21135 = n21134 ^ n21132 ;
  assign n21136 = n19926 ^ n19090 ;
  assign n21137 = n21136 ^ n20486 ;
  assign n21243 = n21137 ^ n21133 ;
  assign n21244 = n21135 & n21243 ;
  assign n21245 = n21244 ^ n21137 ;
  assign n21316 = n21247 ^ n21245 ;
  assign n21317 = n21249 & n21316 ;
  assign n21318 = n21317 ^ n21248 ;
  assign n21319 = n21318 ^ n21313 ;
  assign n21320 = n21315 & n21319 ;
  assign n21322 = n21321 ^ n21320 ;
  assign n21323 = n21311 & n21322 ;
  assign n21324 = n21323 ^ n21310 ;
  assign n21306 = n20791 ^ n1583 ;
  assign n21304 = n20008 ^ n19431 ;
  assign n21305 = n21304 ^ n20667 ;
  assign n21307 = n21306 ^ n21305 ;
  assign n21399 = n21324 ^ n21307 ;
  assign n21400 = n21399 ^ n18704 ;
  assign n21401 = n21322 ^ n21310 ;
  assign n21402 = n21401 ^ n18687 ;
  assign n21406 = n21318 ^ n21315 ;
  assign n21250 = n21249 ^ n21245 ;
  assign n21251 = n21250 ^ n18555 ;
  assign n21138 = n21137 ^ n21135 ;
  assign n21139 = n21138 ^ n18113 ;
  assign n21127 = n21126 ^ n21122 ;
  assign n21128 = n21127 ^ n18123 ;
  assign n21022 = n21012 ^ n20434 ;
  assign n21023 = n21022 ^ n18133 ;
  assign n21025 = n21007 ^ n20444 ;
  assign n21026 = n21025 ^ n18143 ;
  assign n21027 = n21005 ^ n20449 ;
  assign n21028 = n21027 ^ n18150 ;
  assign n21029 = n21001 ^ n20456 ;
  assign n21030 = n21029 ^ n18148 ;
  assign n21032 = n20995 ^ n20466 ;
  assign n21033 = n21032 ^ n18512 ;
  assign n21057 = n20993 ^ n20470 ;
  assign n21034 = n20988 ^ n20967 ;
  assign n21035 = n21034 ^ n20965 ;
  assign n21036 = n21035 ^ n18160 ;
  assign n21038 = n20958 ^ n20956 ;
  assign n21039 = n21038 ^ n18171 ;
  assign n21042 = n20952 ^ n20949 ;
  assign n21040 = n20947 ^ n20946 ;
  assign n21041 = ~n18179 & ~n21040 ;
  assign n21043 = n21042 ^ n21041 ;
  assign n21044 = n21042 ^ n18175 ;
  assign n21045 = n21043 & n21044 ;
  assign n21046 = n21045 ^ n18175 ;
  assign n21047 = n21046 ^ n21038 ;
  assign n21048 = n21039 & n21047 ;
  assign n21049 = n21048 ^ n18171 ;
  assign n21037 = n20963 ^ n20474 ;
  assign n21050 = n21049 ^ n21037 ;
  assign n21051 = n21049 ^ n18167 ;
  assign n21052 = n21050 & n21051 ;
  assign n21053 = n21052 ^ n18167 ;
  assign n21054 = n21053 ^ n21035 ;
  assign n21055 = ~n21036 & ~n21054 ;
  assign n21056 = n21055 ^ n18160 ;
  assign n21058 = n21057 ^ n21056 ;
  assign n21059 = n21057 ^ n18162 ;
  assign n21060 = ~n21058 & ~n21059 ;
  assign n21061 = n21060 ^ n18162 ;
  assign n21062 = n21061 ^ n21032 ;
  assign n21063 = n21033 & n21062 ;
  assign n21064 = n21063 ^ n18512 ;
  assign n21031 = n20999 ^ n20460 ;
  assign n21065 = n21064 ^ n21031 ;
  assign n21066 = n21064 ^ n18156 ;
  assign n21067 = n21065 & n21066 ;
  assign n21068 = n21067 ^ n18156 ;
  assign n21069 = n21068 ^ n21029 ;
  assign n21070 = ~n21030 & ~n21069 ;
  assign n21071 = n21070 ^ n18148 ;
  assign n21072 = n21071 ^ n21027 ;
  assign n21073 = ~n21028 & ~n21072 ;
  assign n21074 = n21073 ^ n18150 ;
  assign n21075 = n21074 ^ n21025 ;
  assign n21076 = ~n21026 & n21075 ;
  assign n21077 = n21076 ^ n18143 ;
  assign n21024 = n21010 ^ n20437 ;
  assign n21078 = n21077 ^ n21024 ;
  assign n21079 = n21077 ^ n18138 ;
  assign n21080 = ~n21078 & n21079 ;
  assign n21081 = n21080 ^ n18138 ;
  assign n21082 = n21081 ^ n21022 ;
  assign n21083 = ~n21023 & ~n21082 ;
  assign n21084 = n21083 ^ n18133 ;
  assign n21020 = n21019 ^ n21017 ;
  assign n21116 = n21084 ^ n21020 ;
  assign n21117 = n21084 ^ n18128 ;
  assign n21118 = ~n21116 & ~n21117 ;
  assign n21119 = n21118 ^ n18128 ;
  assign n21140 = n21127 ^ n21119 ;
  assign n21141 = n21128 & ~n21140 ;
  assign n21142 = n21141 ^ n18123 ;
  assign n21240 = n21142 ^ n21138 ;
  assign n21241 = n21139 & n21240 ;
  assign n21242 = n21241 ^ n18113 ;
  assign n21403 = n21250 ^ n21242 ;
  assign n21404 = n21251 & n21403 ;
  assign n21405 = n21404 ^ n18555 ;
  assign n21407 = n21406 ^ n21405 ;
  assign n21408 = n21406 ^ n18681 ;
  assign n21409 = n21407 & n21408 ;
  assign n21410 = n21409 ^ n18681 ;
  assign n21411 = n21410 ^ n21401 ;
  assign n21412 = ~n21402 & n21411 ;
  assign n21413 = n21412 ^ n18687 ;
  assign n21414 = n21413 ^ n21399 ;
  assign n21415 = n21400 & ~n21414 ;
  assign n21416 = n21415 ^ n18704 ;
  assign n21300 = n20793 ^ n20746 ;
  assign n21327 = n21306 ^ n21300 ;
  assign n21325 = n21324 ^ n21305 ;
  assign n21326 = n21307 & n21325 ;
  assign n21328 = n21327 ^ n21326 ;
  assign n21301 = n20015 ^ n19440 ;
  assign n21302 = n21301 ^ n20715 ;
  assign n21397 = n21328 ^ n21302 ;
  assign n21398 = n21397 ^ n18923 ;
  assign n21462 = n21416 ^ n21398 ;
  assign n21455 = n21410 ^ n21402 ;
  assign n21456 = n21408 ^ n21405 ;
  assign n21021 = n21020 ^ n18128 ;
  assign n21085 = n21084 ^ n21021 ;
  assign n21086 = n21081 ^ n21023 ;
  assign n21087 = n21024 ^ n18138 ;
  assign n21088 = n21087 ^ n21077 ;
  assign n21089 = n21068 ^ n21030 ;
  assign n21090 = n21031 ^ n18156 ;
  assign n21091 = n21090 ^ n21064 ;
  assign n21092 = n21061 ^ n21033 ;
  assign n21093 = n21059 ^ n21056 ;
  assign n21094 = n21053 ^ n21036 ;
  assign n21095 = n21037 ^ n18167 ;
  assign n21096 = n21095 ^ n21049 ;
  assign n21097 = n21041 ^ n18175 ;
  assign n21098 = n21097 ^ n21042 ;
  assign n21099 = n21040 ^ n18179 ;
  assign n21100 = n21098 & n21099 ;
  assign n21101 = n21046 ^ n21039 ;
  assign n21102 = n21100 & ~n21101 ;
  assign n21103 = ~n21096 & n21102 ;
  assign n21104 = ~n21094 & n21103 ;
  assign n21105 = ~n21093 & ~n21104 ;
  assign n21106 = n21092 & ~n21105 ;
  assign n21107 = ~n21091 & ~n21106 ;
  assign n21108 = ~n21089 & n21107 ;
  assign n21109 = n21071 ^ n21028 ;
  assign n21110 = n21108 & n21109 ;
  assign n21111 = n21074 ^ n21026 ;
  assign n21112 = ~n21110 & n21111 ;
  assign n21113 = n21088 & ~n21112 ;
  assign n21114 = n21086 & ~n21113 ;
  assign n21115 = n21085 & ~n21114 ;
  assign n21129 = n21128 ^ n21119 ;
  assign n21130 = n21115 & n21129 ;
  assign n21143 = n21142 ^ n21139 ;
  assign n21239 = n21130 & n21143 ;
  assign n21252 = n21251 ^ n21242 ;
  assign n21457 = n21239 & ~n21252 ;
  assign n21458 = ~n21456 & ~n21457 ;
  assign n21459 = ~n21455 & n21458 ;
  assign n21460 = n21413 ^ n21400 ;
  assign n21461 = ~n21459 & ~n21460 ;
  assign n21539 = n21462 ^ n21461 ;
  assign n21417 = n21416 ^ n21397 ;
  assign n21418 = ~n21398 & ~n21417 ;
  assign n21419 = n21418 ^ n18923 ;
  assign n21303 = n21302 ^ n21300 ;
  assign n21329 = ~n21303 & ~n21328 ;
  assign n21330 = n21329 ^ n21302 ;
  assign n21297 = n20018 ^ n19603 ;
  assign n21298 = n21297 ^ n20835 ;
  assign n21256 = n20796 ^ n20744 ;
  assign n21299 = n21298 ^ n21256 ;
  assign n21395 = n21330 ^ n21299 ;
  assign n21396 = n21395 ^ n18951 ;
  assign n21464 = n21419 ^ n21396 ;
  assign n21463 = n21461 & n21462 ;
  assign n21518 = n21464 ^ n21463 ;
  assign n21542 = n21539 ^ n21518 ;
  assign n21520 = n21460 ^ n21459 ;
  assign n1096 = n1021 ^ x493 ;
  assign n1097 = n1096 ^ n925 ;
  assign n1098 = n1097 ^ x429 ;
  assign n21521 = n21520 ^ n1098 ;
  assign n21534 = n21520 ^ n1112 ;
  assign n21522 = n21458 ^ n21455 ;
  assign n21523 = n21522 ^ n1112 ;
  assign n21527 = n21457 ^ n21456 ;
  assign n21253 = n21252 ^ n21239 ;
  assign n21254 = n21253 ^ n1644 ;
  assign n21144 = n21143 ^ n21130 ;
  assign n21145 = n21144 ^ n690 ;
  assign n21146 = n21129 ^ n21115 ;
  assign n21147 = n21146 ^ n637 ;
  assign n21232 = n21146 ^ n628 ;
  assign n21148 = n21114 ^ n21085 ;
  assign n21149 = n21148 ^ n628 ;
  assign n21153 = n21113 ^ n21086 ;
  assign n21154 = n21153 ^ n21152 ;
  assign n21155 = n21112 ^ n21088 ;
  assign n21156 = n21155 ^ n1494 ;
  assign n21160 = n21111 ^ n21110 ;
  assign n21161 = n21160 ^ n21159 ;
  assign n21162 = n21109 ^ n21108 ;
  assign n21166 = n21165 ^ n21162 ;
  assign n21169 = n21107 ^ n21089 ;
  assign n2361 = n2282 ^ x504 ;
  assign n2362 = n2361 ^ n584 ;
  assign n2363 = n2362 ^ x440 ;
  assign n21170 = n21169 ^ n2363 ;
  assign n21171 = n21106 ^ n21091 ;
  assign n21175 = n21174 ^ n21171 ;
  assign n21178 = n21105 ^ n21092 ;
  assign n2206 = n2142 ^ x506 ;
  assign n2210 = n2209 ^ n2206 ;
  assign n2211 = n2210 ^ x442 ;
  assign n21179 = n21178 ^ n2211 ;
  assign n21180 = n21104 ^ n21093 ;
  assign n2093 = n2035 ^ x507 ;
  assign n2094 = n2093 ^ n2090 ;
  assign n2095 = n2094 ^ x443 ;
  assign n21181 = n21180 ^ n2095 ;
  assign n21182 = n21103 ^ n21094 ;
  assign n2084 = n2026 ^ x508 ;
  assign n2085 = n2084 ^ n2013 ;
  assign n2086 = n2085 ^ x444 ;
  assign n21183 = n21182 ^ n2086 ;
  assign n21186 = n21102 ^ n21096 ;
  assign n2004 = n1961 ^ x509 ;
  assign n2005 = n2004 ^ n2001 ;
  assign n2006 = n2005 ^ x445 ;
  assign n21187 = n21186 ^ n2006 ;
  assign n21188 = n21101 ^ n21100 ;
  assign n1995 = n1952 ^ x510 ;
  assign n1996 = n1995 ^ n1994 ;
  assign n1997 = n1996 ^ x446 ;
  assign n21189 = n21188 ^ n1997 ;
  assign n21193 = n3058 ^ x511 ;
  assign n21194 = n21193 ^ n3051 ;
  assign n21195 = n21194 ^ x447 ;
  assign n3042 = n3014 ^ x480 ;
  assign n3043 = n3042 ^ n3037 ;
  assign n3044 = n3043 ^ x416 ;
  assign n21192 = n3044 & ~n21099 ;
  assign n21196 = n21195 ^ n21192 ;
  assign n21197 = n21099 ^ n21098 ;
  assign n21198 = n21197 ^ n21192 ;
  assign n21199 = n21196 & ~n21198 ;
  assign n21200 = n21199 ^ n21195 ;
  assign n21190 = n21186 ^ n1997 ;
  assign n21191 = n21190 ^ n21186 ;
  assign n21201 = n21200 ^ n21191 ;
  assign n21202 = ~n21189 & n21201 ;
  assign n21203 = n21202 ^ n21190 ;
  assign n21204 = ~n21187 & ~n21203 ;
  assign n21205 = n21204 ^ n21186 ;
  assign n21184 = n21180 ^ n2086 ;
  assign n21185 = n21184 ^ n21180 ;
  assign n21206 = n21205 ^ n21185 ;
  assign n21207 = ~n21183 & ~n21206 ;
  assign n21208 = n21207 ^ n21184 ;
  assign n21209 = ~n21181 & ~n21208 ;
  assign n21210 = n21209 ^ n21180 ;
  assign n21211 = n21210 ^ n2211 ;
  assign n21212 = ~n21179 & n21211 ;
  assign n21213 = n21212 ^ n21178 ;
  assign n21176 = n21174 ^ n21169 ;
  assign n21177 = n21176 ^ n21169 ;
  assign n21214 = n21213 ^ n21177 ;
  assign n21215 = ~n21175 & ~n21214 ;
  assign n21216 = n21215 ^ n21176 ;
  assign n21217 = n21170 & ~n21216 ;
  assign n21218 = n21217 ^ n2363 ;
  assign n21219 = n21218 ^ n21165 ;
  assign n21220 = ~n21166 & n21219 ;
  assign n21167 = n21165 ^ n21160 ;
  assign n21221 = n21220 ^ n21167 ;
  assign n21222 = ~n21161 & ~n21221 ;
  assign n21223 = n21222 ^ n21160 ;
  assign n21224 = n21223 ^ n1494 ;
  assign n21225 = n21156 & n21224 ;
  assign n21226 = n21225 ^ n21155 ;
  assign n21227 = n21226 ^ n21152 ;
  assign n21228 = ~n21154 & ~n21227 ;
  assign n21229 = n21228 ^ n21153 ;
  assign n21230 = n21229 ^ n628 ;
  assign n21231 = n21149 & ~n21230 ;
  assign n21233 = n21232 ^ n21231 ;
  assign n21234 = ~n21147 & ~n21233 ;
  assign n21235 = n21234 ^ n21146 ;
  assign n21236 = n21235 ^ n690 ;
  assign n21237 = ~n21145 & n21236 ;
  assign n21238 = n21237 ^ n21144 ;
  assign n21524 = n21238 ^ n1644 ;
  assign n21525 = n21254 & n21524 ;
  assign n21526 = n21525 ^ n21253 ;
  assign n21528 = n21527 ^ n21526 ;
  assign n21529 = n21527 ^ n776 ;
  assign n21530 = ~n21528 & n21529 ;
  assign n21531 = n21530 ^ n776 ;
  assign n21532 = n21531 ^ n1112 ;
  assign n21533 = ~n21523 & n21532 ;
  assign n21535 = n21534 ^ n21533 ;
  assign n21536 = ~n21521 & ~n21535 ;
  assign n21537 = n21536 ^ n21520 ;
  assign n21538 = n21537 ^ n1123 ;
  assign n21540 = n21539 ^ n1123 ;
  assign n21541 = n21538 & ~n21540 ;
  assign n21543 = n21542 ^ n21541 ;
  assign n21940 = n21543 ^ n1269 ;
  assign n21282 = n20815 ^ n1142 ;
  assign n23200 = n21940 ^ n21282 ;
  assign n21759 = n20482 ^ n19931 ;
  assign n21760 = n21759 ^ n21306 ;
  assign n21260 = n21203 ^ n2006 ;
  assign n21258 = n20441 ^ n19948 ;
  assign n21259 = n21258 ^ n21015 ;
  assign n21261 = n21260 ^ n21259 ;
  assign n21266 = n20448 ^ n19956 ;
  assign n21267 = n21266 ^ n20433 ;
  assign n21265 = n21200 ^ n21189 ;
  assign n21268 = n21267 ^ n21265 ;
  assign n21272 = n20458 ^ n19889 ;
  assign n21273 = n21272 ^ n20443 ;
  assign n21271 = n21099 ^ n3044 ;
  assign n21274 = n21273 ^ n21271 ;
  assign n21355 = n19635 ^ n18990 ;
  assign n21356 = n21355 ^ n20258 ;
  assign n21279 = n19638 ^ n18937 ;
  assign n21280 = n21279 ^ n20921 ;
  assign n21277 = n20809 ^ n1145 ;
  assign n21278 = n21277 ^ n20808 ;
  assign n21281 = n21280 ^ n21278 ;
  assign n21286 = n20323 ^ n19683 ;
  assign n21287 = n21286 ^ n20901 ;
  assign n21285 = n20806 ^ n995 ;
  assign n21288 = n21287 ^ n21285 ;
  assign n21290 = n20271 ^ n19648 ;
  assign n21291 = n21290 ^ n20877 ;
  assign n21289 = n20802 ^ n20740 ;
  assign n21292 = n21291 ^ n21289 ;
  assign n21295 = n20799 ^ n20742 ;
  assign n21336 = n21295 ^ n21289 ;
  assign n21293 = n20239 ^ n19625 ;
  assign n21294 = n21293 ^ n20856 ;
  assign n21296 = n21295 ^ n21294 ;
  assign n21331 = n21330 ^ n21256 ;
  assign n21332 = n21299 & ~n21331 ;
  assign n21333 = n21332 ^ n21298 ;
  assign n21334 = n21333 ^ n21295 ;
  assign n21335 = ~n21296 & n21334 ;
  assign n21337 = n21336 ^ n21335 ;
  assign n21338 = ~n21292 & n21337 ;
  assign n21339 = n21338 ^ n21291 ;
  assign n21340 = n21339 ^ n21285 ;
  assign n21341 = ~n21288 & n21340 ;
  assign n21342 = n21341 ^ n21287 ;
  assign n21283 = n21282 ^ n21278 ;
  assign n21284 = n21283 ^ n21282 ;
  assign n21343 = n21342 ^ n21284 ;
  assign n21344 = n21281 & ~n21343 ;
  assign n21345 = n21344 ^ n21283 ;
  assign n21346 = n20734 ^ n1349 ;
  assign n21347 = n21346 ^ n20817 ;
  assign n21351 = n21347 ^ n21282 ;
  assign n21348 = n19613 ^ n18962 ;
  assign n21349 = n21348 ^ n20977 ;
  assign n21350 = n21349 ^ n21347 ;
  assign n21352 = n21351 ^ n21350 ;
  assign n21353 = ~n21345 & n21352 ;
  assign n21354 = n21353 ^ n21351 ;
  assign n21385 = n21356 ^ n21354 ;
  assign n21386 = n21385 ^ n18466 ;
  assign n21435 = n21349 ^ n21345 ;
  assign n21387 = n21342 ^ n21281 ;
  assign n21388 = n21387 ^ n18470 ;
  assign n21389 = n21339 ^ n21288 ;
  assign n21390 = n21389 ^ n19155 ;
  assign n21391 = n21337 ^ n21291 ;
  assign n21392 = n21391 ^ n19032 ;
  assign n21393 = n21333 ^ n21296 ;
  assign n21394 = n21393 ^ n18973 ;
  assign n21420 = n21419 ^ n21395 ;
  assign n21421 = n21396 & n21420 ;
  assign n21422 = n21421 ^ n18951 ;
  assign n21423 = n21422 ^ n21393 ;
  assign n21424 = n21394 & n21423 ;
  assign n21425 = n21424 ^ n18973 ;
  assign n21426 = n21425 ^ n21391 ;
  assign n21427 = ~n21392 & ~n21426 ;
  assign n21428 = n21427 ^ n19032 ;
  assign n21429 = n21428 ^ n21389 ;
  assign n21430 = n21390 & n21429 ;
  assign n21431 = n21430 ^ n19155 ;
  assign n21432 = n21431 ^ n21387 ;
  assign n21433 = ~n21388 & n21432 ;
  assign n21434 = n21433 ^ n18470 ;
  assign n21436 = n21435 ^ n21434 ;
  assign n21437 = n21435 ^ n18478 ;
  assign n21438 = ~n21436 & ~n21437 ;
  assign n21439 = n21438 ^ n18478 ;
  assign n21440 = n21439 ^ n21385 ;
  assign n21441 = ~n21386 & ~n21440 ;
  assign n21442 = n21441 ^ n18466 ;
  assign n21363 = n19668 ^ n19047 ;
  assign n21364 = n21363 ^ n20263 ;
  assign n21357 = n20823 ^ n2879 ;
  assign n21359 = n21357 ^ n21347 ;
  assign n21358 = n21357 ^ n21356 ;
  assign n21360 = n21359 ^ n21358 ;
  assign n21361 = n21354 & n21360 ;
  assign n21362 = n21361 ^ n21359 ;
  assign n21383 = n21364 ^ n21362 ;
  assign n21384 = n21383 ^ n18464 ;
  assign n21453 = n21442 ^ n21384 ;
  assign n21454 = n21437 ^ n21434 ;
  assign n21465 = ~n21463 & ~n21464 ;
  assign n21466 = n21422 ^ n21394 ;
  assign n21467 = ~n21465 & ~n21466 ;
  assign n21468 = n21425 ^ n21392 ;
  assign n21469 = n21467 & ~n21468 ;
  assign n21470 = n21428 ^ n21390 ;
  assign n21471 = ~n21469 & n21470 ;
  assign n21472 = n21431 ^ n21388 ;
  assign n21473 = ~n21471 & ~n21472 ;
  assign n21474 = ~n21454 & n21473 ;
  assign n21475 = n21439 ^ n21386 ;
  assign n21476 = n21474 & n21475 ;
  assign n21477 = n21453 & ~n21476 ;
  assign n21373 = n19695 ^ n19167 ;
  assign n21374 = n21373 ^ n20253 ;
  assign n21365 = n20825 ^ n20731 ;
  assign n21367 = n21365 ^ n21357 ;
  assign n21366 = n21365 ^ n21364 ;
  assign n21368 = n21367 ^ n21366 ;
  assign n21369 = ~n21362 & n21368 ;
  assign n21370 = n21369 ^ n21367 ;
  assign n21446 = n21374 ^ n21370 ;
  assign n21448 = n21446 ^ n18460 ;
  assign n21443 = n21442 ^ n21383 ;
  assign n21444 = ~n21384 & n21443 ;
  assign n21445 = n21444 ^ n18464 ;
  assign n21478 = n21448 ^ n21445 ;
  assign n21479 = ~n21477 & n21478 ;
  assign n21447 = n21446 ^ n21445 ;
  assign n21449 = ~n21447 & n21448 ;
  assign n21450 = n21449 ^ n18460 ;
  assign n21451 = n21450 ^ n18186 ;
  assign n21380 = n19145 ^ n19079 ;
  assign n21381 = n21380 ^ n20292 ;
  assign n21371 = n20729 ^ n2901 ;
  assign n21372 = n21371 ^ n20828 ;
  assign n21376 = n21372 ^ n21365 ;
  assign n21375 = n21374 ^ n21372 ;
  assign n21377 = n21376 ^ n21375 ;
  assign n21378 = ~n21370 & n21377 ;
  assign n21379 = n21378 ^ n21376 ;
  assign n21382 = n21381 ^ n21379 ;
  assign n21452 = n21451 ^ n21382 ;
  assign n21497 = n21479 ^ n21452 ;
  assign n21498 = n21497 ^ n2765 ;
  assign n21499 = n21478 ^ n21477 ;
  assign n21500 = n21499 ^ n1841 ;
  assign n21503 = n21476 ^ n21453 ;
  assign n3140 = n3127 ^ x484 ;
  assign n3141 = n3140 ^ n2465 ;
  assign n3142 = n3141 ^ x420 ;
  assign n21504 = n21503 ^ n3142 ;
  assign n21505 = n21475 ^ n21474 ;
  assign n21506 = n21505 ^ n3135 ;
  assign n21509 = n21473 ^ n21454 ;
  assign n21510 = n21509 ^ n2513 ;
  assign n21558 = n21472 ^ n21471 ;
  assign n21511 = n21470 ^ n21469 ;
  assign n21512 = n21511 ^ n2546 ;
  assign n21513 = n21468 ^ n21467 ;
  assign n21517 = n21516 ^ n21513 ;
  assign n21546 = n21466 ^ n21465 ;
  assign n21519 = n21518 ^ n1269 ;
  assign n21544 = n21519 & ~n21543 ;
  assign n21545 = n21544 ^ n21518 ;
  assign n21547 = n21546 ^ n21545 ;
  assign n21548 = n21513 ^ n1284 ;
  assign n21549 = n21548 ^ n21513 ;
  assign n21550 = n21549 ^ n21545 ;
  assign n21551 = n21547 & n21550 ;
  assign n21552 = n21551 ^ n21548 ;
  assign n21553 = n21517 & ~n21552 ;
  assign n21554 = n21553 ^ n21516 ;
  assign n21555 = n21554 ^ n21511 ;
  assign n21556 = ~n21512 & n21555 ;
  assign n21557 = n21556 ^ n2546 ;
  assign n21559 = n21558 ^ n21557 ;
  assign n21560 = n21509 ^ n3209 ;
  assign n21561 = n21560 ^ n21509 ;
  assign n21562 = n21561 ^ n21557 ;
  assign n21563 = n21559 & n21562 ;
  assign n21564 = n21563 ^ n21560 ;
  assign n21565 = n21510 & ~n21564 ;
  assign n21566 = n21565 ^ n2513 ;
  assign n21507 = n21503 ^ n3135 ;
  assign n21508 = n21507 ^ n21503 ;
  assign n21567 = n21566 ^ n21508 ;
  assign n21568 = ~n21506 & n21567 ;
  assign n21569 = n21568 ^ n21507 ;
  assign n21570 = ~n21504 & n21569 ;
  assign n21571 = n21570 ^ n3142 ;
  assign n21501 = n21497 ^ n1841 ;
  assign n21502 = n21501 ^ n21497 ;
  assign n21572 = n21571 ^ n21502 ;
  assign n21573 = n21500 & n21572 ;
  assign n21574 = n21573 ^ n21501 ;
  assign n21575 = ~n21498 & n21574 ;
  assign n21492 = n2781 ^ n2765 ;
  assign n21490 = n18186 ^ n18184 ;
  assign n21486 = n19081 ^ n19074 ;
  assign n21487 = n21486 ^ n20342 ;
  assign n21488 = n21487 ^ n21381 ;
  assign n21485 = n20871 ^ n20851 ;
  assign n21489 = n21488 ^ n21485 ;
  assign n21491 = n21490 ^ n21489 ;
  assign n21493 = n21492 ^ n21491 ;
  assign n21483 = n21450 ^ n21382 ;
  assign n21484 = ~n21451 & n21483 ;
  assign n21494 = n21493 ^ n21484 ;
  assign n21481 = n21381 ^ n21372 ;
  assign n21482 = ~n21379 & n21481 ;
  assign n21495 = n21494 ^ n21482 ;
  assign n21480 = n21452 & n21479 ;
  assign n21496 = n21495 ^ n21480 ;
  assign n21576 = n21575 ^ n21496 ;
  assign n21275 = n20462 ^ n19789 ;
  assign n21276 = n21275 ^ n20450 ;
  assign n21577 = n21576 ^ n21276 ;
  assign n21580 = n20468 ^ n19772 ;
  assign n21581 = n21580 ^ n20452 ;
  assign n21578 = n21574 ^ n2765 ;
  assign n21582 = n21581 ^ n21578 ;
  assign n21584 = n20517 ^ n19723 ;
  assign n21585 = n21584 ^ n20457 ;
  assign n21583 = n21571 ^ n21500 ;
  assign n21586 = n21585 ^ n21583 ;
  assign n21589 = n20423 ^ n19068 ;
  assign n21590 = n21589 ^ n20467 ;
  assign n21591 = n21566 ^ n21506 ;
  assign n21592 = n21590 & ~n21591 ;
  assign n21597 = n21592 ^ n21583 ;
  assign n21587 = n20472 ^ n19057 ;
  assign n21588 = n21587 ^ n20465 ;
  assign n21593 = n21592 ^ n21588 ;
  assign n21594 = n21569 ^ n3142 ;
  assign n21595 = n21594 ^ n21592 ;
  assign n21596 = ~n21593 & ~n21595 ;
  assign n21598 = n21597 ^ n21596 ;
  assign n21599 = ~n21586 & ~n21598 ;
  assign n21600 = n21599 ^ n21585 ;
  assign n21601 = n21600 ^ n21578 ;
  assign n21602 = ~n21582 & n21601 ;
  assign n21579 = n21578 ^ n21576 ;
  assign n21603 = n21602 ^ n21579 ;
  assign n21604 = ~n21577 & n21603 ;
  assign n21605 = n21604 ^ n21576 ;
  assign n21606 = n21605 ^ n21271 ;
  assign n21607 = ~n21274 & n21606 ;
  assign n21608 = n21607 ^ n21271 ;
  assign n21613 = n21608 ^ n21265 ;
  assign n21269 = n20453 ^ n19960 ;
  assign n21270 = n21269 ^ n20438 ;
  assign n21609 = n21608 ^ n21270 ;
  assign n21610 = n21197 ^ n21196 ;
  assign n21611 = n21610 ^ n21270 ;
  assign n21612 = ~n21609 & ~n21611 ;
  assign n21614 = n21613 ^ n21612 ;
  assign n21615 = ~n21268 & ~n21614 ;
  assign n21616 = n21615 ^ n21267 ;
  assign n21262 = n21205 ^ n21183 ;
  assign n21263 = n21262 ^ n21260 ;
  assign n21264 = n21263 ^ n21262 ;
  assign n21617 = n21616 ^ n21264 ;
  assign n21618 = ~n21261 & ~n21617 ;
  assign n21619 = n21618 ^ n21263 ;
  assign n21622 = n21208 ^ n2095 ;
  assign n21624 = n21622 ^ n21262 ;
  assign n21620 = n20435 ^ n19944 ;
  assign n21621 = n21620 ^ n21125 ;
  assign n21623 = n21622 ^ n21621 ;
  assign n21625 = n21624 ^ n21623 ;
  assign n21626 = ~n21619 & ~n21625 ;
  assign n21627 = n21626 ^ n21624 ;
  assign n21628 = n21210 ^ n21179 ;
  assign n21632 = n21628 ^ n21622 ;
  assign n21629 = n19942 ^ n19906 ;
  assign n21630 = n21629 ^ n21133 ;
  assign n21631 = n21630 ^ n21628 ;
  assign n21633 = n21632 ^ n21631 ;
  assign n21634 = ~n21627 & ~n21633 ;
  assign n21635 = n21634 ^ n21632 ;
  assign n21636 = n21213 ^ n21175 ;
  assign n21640 = n21636 ^ n21628 ;
  assign n21637 = n20494 ^ n19938 ;
  assign n21638 = n21637 ^ n21248 ;
  assign n21639 = n21638 ^ n21636 ;
  assign n21641 = n21640 ^ n21639 ;
  assign n21642 = ~n21635 & ~n21641 ;
  assign n21643 = n21642 ^ n21640 ;
  assign n21736 = n21216 ^ n2363 ;
  assign n21738 = n21736 ^ n21636 ;
  assign n21644 = n20492 ^ n19908 ;
  assign n21645 = n21644 ^ n21314 ;
  assign n21737 = n21736 ^ n21645 ;
  assign n21739 = n21738 ^ n21737 ;
  assign n21740 = n21643 & ~n21739 ;
  assign n21741 = n21740 ^ n21738 ;
  assign n21753 = n21218 ^ n21166 ;
  assign n21755 = n21753 ^ n21736 ;
  assign n21742 = n20486 ^ n19985 ;
  assign n21743 = n21742 ^ n21308 ;
  assign n21754 = n21753 ^ n21743 ;
  assign n21756 = n21755 ^ n21754 ;
  assign n21757 = n21741 & ~n21756 ;
  assign n21758 = n21757 ^ n21755 ;
  assign n21761 = n21760 ^ n21758 ;
  assign n21744 = n21743 ^ n21741 ;
  assign n21745 = n21744 ^ n19098 ;
  assign n21700 = n21638 ^ n21635 ;
  assign n21648 = n21630 ^ n21627 ;
  assign n21649 = n21648 ^ n19103 ;
  assign n21692 = n21621 ^ n21619 ;
  assign n21650 = n21616 ^ n21261 ;
  assign n21651 = n21650 ^ n19114 ;
  assign n21652 = n21614 ^ n21267 ;
  assign n21653 = n21652 ^ n19062 ;
  assign n21654 = n21611 ^ n21608 ;
  assign n21655 = n21654 ^ n19058 ;
  assign n21674 = n21603 ^ n21276 ;
  assign n21657 = n21600 ^ n21582 ;
  assign n21658 = n21657 ^ n19076 ;
  assign n21666 = n21598 ^ n21585 ;
  assign n21661 = n21594 ^ n21593 ;
  assign n21659 = n21591 ^ n21590 ;
  assign n21660 = n19136 & ~n21659 ;
  assign n21662 = n21661 ^ n21660 ;
  assign n21663 = n21661 ^ n19134 ;
  assign n21664 = ~n21662 & n21663 ;
  assign n21665 = n21664 ^ n19134 ;
  assign n21667 = n21666 ^ n21665 ;
  assign n21668 = n21666 ^ n19127 ;
  assign n21669 = n21667 & ~n21668 ;
  assign n21670 = n21669 ^ n19127 ;
  assign n21671 = n21670 ^ n21657 ;
  assign n21672 = n21658 & ~n21671 ;
  assign n21673 = n21672 ^ n19076 ;
  assign n21675 = n21674 ^ n21673 ;
  assign n21676 = n21674 ^ n19070 ;
  assign n21677 = ~n21675 & ~n21676 ;
  assign n21678 = n21677 ^ n19070 ;
  assign n21656 = n21605 ^ n21274 ;
  assign n21679 = n21678 ^ n21656 ;
  assign n21680 = n21678 ^ n19065 ;
  assign n21681 = n21679 & ~n21680 ;
  assign n21682 = n21681 ^ n19065 ;
  assign n21683 = n21682 ^ n21654 ;
  assign n21684 = n21655 & n21683 ;
  assign n21685 = n21684 ^ n19058 ;
  assign n21686 = n21685 ^ n21652 ;
  assign n21687 = ~n21653 & n21686 ;
  assign n21688 = n21687 ^ n19062 ;
  assign n21689 = n21688 ^ n21650 ;
  assign n21690 = n21651 & ~n21689 ;
  assign n21691 = n21690 ^ n19114 ;
  assign n21693 = n21692 ^ n21691 ;
  assign n21694 = n21692 ^ n19110 ;
  assign n21695 = n21693 & ~n21694 ;
  assign n21696 = n21695 ^ n19110 ;
  assign n21697 = n21696 ^ n21648 ;
  assign n21698 = n21649 & ~n21697 ;
  assign n21699 = n21698 ^ n19103 ;
  assign n21701 = n21700 ^ n21699 ;
  assign n21702 = n21700 ^ n19107 ;
  assign n21703 = n21701 & ~n21702 ;
  assign n21704 = n21703 ^ n19107 ;
  assign n21646 = n21645 ^ n21643 ;
  assign n21732 = n21704 ^ n21646 ;
  assign n21733 = n21704 ^ n19224 ;
  assign n21734 = ~n21732 & n21733 ;
  assign n21735 = n21734 ^ n19224 ;
  assign n21749 = n21744 ^ n21735 ;
  assign n21750 = n21745 & ~n21749 ;
  assign n21751 = n21750 ^ n19098 ;
  assign n21752 = n21751 ^ n19092 ;
  assign n21762 = n21761 ^ n21752 ;
  assign n21647 = n21646 ^ n19224 ;
  assign n21705 = n21704 ^ n21647 ;
  assign n21706 = n21682 ^ n21655 ;
  assign n21707 = n21656 ^ n19065 ;
  assign n21708 = n21707 ^ n21678 ;
  assign n21709 = n21676 ^ n21673 ;
  assign n21710 = n21670 ^ n21658 ;
  assign n21711 = n21668 ^ n21665 ;
  assign n21712 = n21659 ^ n19136 ;
  assign n21713 = n21660 ^ n19134 ;
  assign n21714 = n21713 ^ n21661 ;
  assign n21715 = ~n21712 & n21714 ;
  assign n21716 = ~n21711 & n21715 ;
  assign n21717 = n21710 & n21716 ;
  assign n21718 = ~n21709 & n21717 ;
  assign n21719 = n21708 & ~n21718 ;
  assign n21720 = n21706 & ~n21719 ;
  assign n21721 = n21685 ^ n21653 ;
  assign n21722 = ~n21720 & ~n21721 ;
  assign n21723 = n21688 ^ n21651 ;
  assign n21724 = n21722 & n21723 ;
  assign n21725 = n21694 ^ n21691 ;
  assign n21726 = n21724 & ~n21725 ;
  assign n21727 = n21696 ^ n21649 ;
  assign n21728 = ~n21726 & ~n21727 ;
  assign n21729 = n21702 ^ n21699 ;
  assign n21730 = ~n21728 & ~n21729 ;
  assign n21731 = ~n21705 & ~n21730 ;
  assign n21746 = n21745 ^ n21735 ;
  assign n21763 = ~n21731 & n21746 ;
  assign n22069 = ~n21762 & n21763 ;
  assign n21991 = n21761 ^ n21751 ;
  assign n21992 = n21752 & n21991 ;
  assign n21993 = n21992 ^ n19092 ;
  assign n21893 = n21221 ^ n21159 ;
  assign n21899 = n21893 ^ n21753 ;
  assign n21897 = n21760 ^ n21753 ;
  assign n21898 = ~n21758 & n21897 ;
  assign n21900 = n21899 ^ n21898 ;
  assign n21894 = n20475 ^ n19926 ;
  assign n21895 = n21894 ^ n21300 ;
  assign n21989 = n21900 ^ n21895 ;
  assign n21990 = n21989 ^ n19090 ;
  assign n22070 = n21993 ^ n21990 ;
  assign n22071 = n22069 & ~n22070 ;
  assign n21896 = n21895 ^ n21893 ;
  assign n21901 = n21896 & ~n21900 ;
  assign n21902 = n21901 ^ n21895 ;
  assign n21891 = n21223 ^ n21156 ;
  assign n21889 = n20479 ^ n19922 ;
  assign n21890 = n21889 ^ n21256 ;
  assign n21892 = n21891 ^ n21890 ;
  assign n21997 = n21902 ^ n21892 ;
  assign n21999 = n21997 ^ n19084 ;
  assign n21994 = n21993 ^ n21989 ;
  assign n21995 = ~n21990 & ~n21994 ;
  assign n21996 = n21995 ^ n19090 ;
  assign n22072 = n21999 ^ n21996 ;
  assign n22073 = n22071 & n22072 ;
  assign n21998 = n21997 ^ n21996 ;
  assign n22000 = n21998 & ~n21999 ;
  assign n22001 = n22000 ^ n19084 ;
  assign n21903 = n21902 ^ n21890 ;
  assign n21904 = n21892 & ~n21903 ;
  assign n21905 = n21904 ^ n21891 ;
  assign n21886 = n20667 ^ n19918 ;
  assign n21887 = n21886 ^ n21295 ;
  assign n21884 = n21226 ^ n21154 ;
  assign n21888 = n21887 ^ n21884 ;
  assign n21987 = n21905 ^ n21888 ;
  assign n21988 = n21987 ^ n19401 ;
  assign n22074 = n22001 ^ n21988 ;
  assign n22075 = ~n22073 & n22074 ;
  assign n21906 = n21905 ^ n21884 ;
  assign n21907 = ~n21888 & n21906 ;
  assign n21882 = n21229 ^ n21149 ;
  assign n21885 = n21884 ^ n21882 ;
  assign n21908 = n21907 ^ n21885 ;
  assign n21880 = n20715 ^ n19914 ;
  assign n21881 = n21880 ^ n21289 ;
  assign n22005 = n21908 ^ n21881 ;
  assign n22007 = n22005 ^ n19409 ;
  assign n22002 = n22001 ^ n21987 ;
  assign n22003 = n21988 & ~n22002 ;
  assign n22004 = n22003 ^ n19401 ;
  assign n22076 = n22007 ^ n22004 ;
  assign n22077 = n22075 & ~n22076 ;
  assign n21883 = n21882 ^ n21881 ;
  assign n21909 = ~n21883 & n21908 ;
  assign n21910 = n21909 ^ n21882 ;
  assign n21877 = n20835 ^ n20008 ;
  assign n21878 = n21877 ^ n21285 ;
  assign n21875 = n21233 ^ n637 ;
  assign n21879 = n21878 ^ n21875 ;
  assign n21986 = n21910 ^ n21879 ;
  assign n22067 = n21986 ^ n19431 ;
  assign n22006 = n22005 ^ n22004 ;
  assign n22008 = ~n22006 & ~n22007 ;
  assign n22009 = n22008 ^ n19409 ;
  assign n22068 = n22067 ^ n22009 ;
  assign n22115 = n22077 ^ n22068 ;
  assign n854 = n830 ^ n790 ;
  assign n855 = n854 ^ n851 ;
  assign n856 = n855 ^ x462 ;
  assign n22139 = n22115 ^ n856 ;
  assign n22117 = n22076 ^ n22075 ;
  assign n22118 = n22117 ^ n856 ;
  assign n22119 = n22074 ^ n22073 ;
  assign n22120 = n22119 ^ n847 ;
  assign n22121 = n22072 ^ n22071 ;
  assign n22122 = n22121 ^ n761 ;
  assign n22123 = n22070 ^ n22069 ;
  assign n22124 = n22123 ^ n752 ;
  assign n21747 = n21746 ^ n21731 ;
  assign n21748 = n21747 ^ n1543 ;
  assign n21767 = n21730 ^ n21705 ;
  assign n21768 = n21767 ^ n2942 ;
  assign n21769 = n21729 ^ n21728 ;
  assign n21773 = n21772 ^ n21769 ;
  assign n21774 = n21727 ^ n21726 ;
  assign n21775 = n21774 ^ n593 ;
  assign n21776 = n21725 ^ n21724 ;
  assign n21780 = n21779 ^ n21776 ;
  assign n21786 = n21723 ^ n21722 ;
  assign n21787 = n21786 ^ n21785 ;
  assign n21833 = n21786 ^ n2309 ;
  assign n21788 = n21721 ^ n21720 ;
  assign n21789 = n21788 ^ n2309 ;
  assign n21790 = n21719 ^ n21706 ;
  assign n21791 = n21790 ^ n2199 ;
  assign n21792 = n21718 ^ n21708 ;
  assign n21793 = n21792 ^ n2184 ;
  assign n21794 = n21717 ^ n21709 ;
  assign n2172 = n2108 ^ n2062 ;
  assign n2176 = n2175 ^ n2172 ;
  assign n2177 = n2176 ^ x476 ;
  assign n21795 = n21794 ^ n2177 ;
  assign n21799 = n19844 ^ n2042 ;
  assign n21800 = n21799 ^ n1931 ;
  assign n21801 = n21800 ^ x477 ;
  assign n21798 = n21716 ^ n21710 ;
  assign n21802 = n21801 ^ n21798 ;
  assign n21806 = n21715 ^ n21711 ;
  assign n21803 = n19851 ^ n2046 ;
  assign n21804 = n21803 ^ n16729 ;
  assign n21805 = n21804 ^ x478 ;
  assign n21807 = n21806 ^ n21805 ;
  assign n21808 = n20332 ^ n3068 ;
  assign n21809 = n21808 ^ n1802 ;
  assign n21810 = n21809 ^ x448 ;
  assign n21811 = n21712 & n21810 ;
  assign n1872 = n1871 ^ n1793 ;
  assign n1876 = n1875 ^ n1872 ;
  assign n1877 = n1876 ^ x479 ;
  assign n21812 = n21811 ^ n1877 ;
  assign n21813 = n21714 ^ n21712 ;
  assign n21814 = n21813 ^ n1877 ;
  assign n21815 = n21812 & n21814 ;
  assign n21816 = n21815 ^ n21811 ;
  assign n21817 = n21816 ^ n21805 ;
  assign n21818 = ~n21807 & n21817 ;
  assign n21819 = n21818 ^ n21805 ;
  assign n21820 = n21819 ^ n21798 ;
  assign n21821 = n21802 & ~n21820 ;
  assign n21822 = n21821 ^ n21801 ;
  assign n21796 = n21792 ^ n2177 ;
  assign n21797 = n21796 ^ n21792 ;
  assign n21823 = n21822 ^ n21797 ;
  assign n21824 = ~n21795 & n21823 ;
  assign n21825 = n21824 ^ n21796 ;
  assign n21826 = n21793 & n21825 ;
  assign n21827 = n21826 ^ n21792 ;
  assign n21828 = n21827 ^ n21790 ;
  assign n21829 = ~n21791 & n21828 ;
  assign n21830 = n21829 ^ n2199 ;
  assign n21831 = n21830 ^ n2309 ;
  assign n21832 = ~n21789 & n21831 ;
  assign n21834 = n21833 ^ n21832 ;
  assign n21835 = ~n21787 & ~n21834 ;
  assign n21836 = n21835 ^ n21786 ;
  assign n21781 = n21779 ^ n21774 ;
  assign n21782 = n21781 ^ n21774 ;
  assign n21837 = n21836 ^ n21782 ;
  assign n21838 = n21780 & ~n21837 ;
  assign n21839 = n21838 ^ n21781 ;
  assign n21840 = n21775 & ~n21839 ;
  assign n21841 = n21840 ^ n593 ;
  assign n21842 = n21841 ^ n21769 ;
  assign n21843 = ~n21773 & n21842 ;
  assign n21844 = n21843 ^ n21772 ;
  assign n21845 = n21844 ^ n2942 ;
  assign n21846 = n21768 & ~n21845 ;
  assign n21847 = n21846 ^ n21767 ;
  assign n21764 = n21763 ^ n21762 ;
  assign n21765 = n21764 ^ n1543 ;
  assign n21766 = n21765 ^ n21764 ;
  assign n21848 = n21847 ^ n21766 ;
  assign n21849 = n21748 & n21848 ;
  assign n21850 = n21849 ^ n21765 ;
  assign n22125 = n21764 ^ n1552 ;
  assign n22126 = n21850 & n22125 ;
  assign n22127 = n22126 ^ n21764 ;
  assign n22128 = n22127 ^ n752 ;
  assign n22129 = n22124 & ~n22128 ;
  assign n22130 = n22129 ^ n22123 ;
  assign n22131 = n22130 ^ n761 ;
  assign n22132 = ~n22122 & ~n22131 ;
  assign n22133 = n22132 ^ n22121 ;
  assign n22134 = n22133 ^ n847 ;
  assign n22135 = ~n22120 & n22134 ;
  assign n22136 = n22135 ^ n22119 ;
  assign n22137 = n22136 ^ n856 ;
  assign n22138 = ~n22118 & ~n22137 ;
  assign n22140 = n22139 ^ n22138 ;
  assign n22436 = n22140 ^ n977 ;
  assign n23201 = n23200 ^ n22436 ;
  assign n22408 = n21830 ^ n21789 ;
  assign n22404 = n21834 ^ n21785 ;
  assign n22499 = n22408 ^ n22404 ;
  assign n22477 = n21306 ^ n20492 ;
  assign n22478 = n22477 ^ n21884 ;
  assign n22479 = n22478 ^ n22408 ;
  assign n22482 = n21827 ^ n21791 ;
  assign n22480 = n21308 ^ n20494 ;
  assign n22481 = n22480 ^ n21891 ;
  assign n22483 = n22482 ^ n22481 ;
  assign n22484 = n21314 ^ n19906 ;
  assign n22485 = n22484 ^ n21893 ;
  assign n22413 = n21825 ^ n2184 ;
  assign n22486 = n22485 ^ n22413 ;
  assign n22301 = n21819 ^ n21802 ;
  assign n22273 = n21816 ^ n21807 ;
  assign n22302 = n22301 ^ n22273 ;
  assign n21855 = n21813 ^ n21812 ;
  assign n22274 = n22273 ^ n21855 ;
  assign n21858 = n20458 ^ n20433 ;
  assign n21859 = n21858 ^ n21622 ;
  assign n21856 = n21810 ^ n21712 ;
  assign n21860 = n21859 ^ n21856 ;
  assign n22203 = n20462 ^ n20438 ;
  assign n22204 = n22203 ^ n21262 ;
  assign n22235 = n22204 ^ n21856 ;
  assign n22196 = n21564 ^ n2513 ;
  assign n22193 = n20374 ^ n19074 ;
  assign n22059 = n20357 ^ n19079 ;
  assign n22060 = n22059 ^ n20941 ;
  assign n22194 = n22193 ^ n22060 ;
  assign n22195 = n22194 ^ n20988 ;
  assign n22197 = n22196 ^ n22195 ;
  assign n22198 = n22197 ^ n19179 ;
  assign n21863 = n21529 ^ n21526 ;
  assign n21861 = n20901 ^ n20239 ;
  assign n21862 = n21861 ^ n21347 ;
  assign n21864 = n21863 ^ n21862 ;
  assign n21868 = n20877 ^ n20018 ;
  assign n21869 = n21868 ^ n21282 ;
  assign n21255 = n21254 ^ n21238 ;
  assign n21870 = n21869 ^ n21255 ;
  assign n21873 = n21235 ^ n21145 ;
  assign n21871 = n20856 ^ n20015 ;
  assign n21872 = n21871 ^ n21278 ;
  assign n21874 = n21873 ^ n21872 ;
  assign n21911 = n21910 ^ n21875 ;
  assign n21912 = ~n21879 & n21911 ;
  assign n21876 = n21875 ^ n21873 ;
  assign n21913 = n21912 ^ n21876 ;
  assign n21914 = ~n21874 & ~n21913 ;
  assign n21915 = n21914 ^ n21873 ;
  assign n21916 = n21915 ^ n21869 ;
  assign n21917 = ~n21870 & ~n21916 ;
  assign n21918 = n21917 ^ n21255 ;
  assign n21865 = n21531 ^ n21523 ;
  assign n21866 = n21865 ^ n21863 ;
  assign n21867 = n21866 ^ n21865 ;
  assign n21919 = n21918 ^ n21867 ;
  assign n21920 = ~n21864 & ~n21919 ;
  assign n21921 = n21920 ^ n21866 ;
  assign n21922 = n21535 ^ n1098 ;
  assign n21926 = n21922 ^ n21865 ;
  assign n21923 = n20921 ^ n20271 ;
  assign n21924 = n21923 ^ n21357 ;
  assign n21925 = n21924 ^ n21922 ;
  assign n21927 = n21926 ^ n21925 ;
  assign n21928 = ~n21921 & ~n21927 ;
  assign n21929 = n21928 ^ n21926 ;
  assign n21932 = n21540 ^ n21537 ;
  assign n21934 = n21932 ^ n21922 ;
  assign n21930 = n20977 ^ n20323 ;
  assign n21931 = n21930 ^ n21365 ;
  assign n21933 = n21932 ^ n21931 ;
  assign n21935 = n21934 ^ n21933 ;
  assign n21936 = n21929 & ~n21935 ;
  assign n21937 = n21936 ^ n21934 ;
  assign n21942 = n21940 ^ n21932 ;
  assign n21938 = n20258 ^ n19638 ;
  assign n21939 = n21938 ^ n21372 ;
  assign n21941 = n21940 ^ n21939 ;
  assign n21943 = n21942 ^ n21941 ;
  assign n21944 = ~n21937 & ~n21943 ;
  assign n21945 = n21944 ^ n21942 ;
  assign n21948 = n21546 ^ n1284 ;
  assign n21949 = n21948 ^ n21545 ;
  assign n21951 = n21949 ^ n21940 ;
  assign n21946 = n20263 ^ n19613 ;
  assign n21947 = n21946 ^ n21485 ;
  assign n21950 = n21949 ^ n21947 ;
  assign n21952 = n21951 ^ n21950 ;
  assign n21953 = ~n21945 & ~n21952 ;
  assign n21954 = n21953 ^ n21951 ;
  assign n21957 = n21552 ^ n21516 ;
  assign n21959 = n21957 ^ n21949 ;
  assign n21955 = n20253 ^ n19635 ;
  assign n21956 = n21955 ^ n20947 ;
  assign n21958 = n21957 ^ n21956 ;
  assign n21960 = n21959 ^ n21958 ;
  assign n21961 = n21954 & ~n21960 ;
  assign n21962 = n21961 ^ n21959 ;
  assign n21965 = n21554 ^ n21512 ;
  assign n21967 = n21965 ^ n21957 ;
  assign n21963 = n20292 ^ n19668 ;
  assign n21964 = n21963 ^ n20952 ;
  assign n21966 = n21965 ^ n21964 ;
  assign n21968 = n21967 ^ n21966 ;
  assign n21969 = ~n21962 & n21968 ;
  assign n21970 = n21969 ^ n21967 ;
  assign n22052 = n21558 ^ n3209 ;
  assign n22053 = n22052 ^ n21557 ;
  assign n21971 = n20342 ^ n19695 ;
  assign n21972 = n21971 ^ n20950 ;
  assign n22055 = n22053 ^ n21972 ;
  assign n22054 = n22053 ^ n21965 ;
  assign n22056 = n22055 ^ n22054 ;
  assign n22057 = ~n21970 & n22056 ;
  assign n22058 = n22057 ^ n22054 ;
  assign n22191 = n22060 ^ n22053 ;
  assign n22192 = ~n22058 & ~n22191 ;
  assign n22199 = n22198 ^ n22192 ;
  assign n22061 = n22060 ^ n22058 ;
  assign n21973 = n21972 ^ n21970 ;
  assign n21974 = n21973 ^ n19167 ;
  assign n22043 = n21964 ^ n21962 ;
  assign n21975 = n21956 ^ n21954 ;
  assign n21976 = n21975 ^ n18990 ;
  assign n22035 = n21947 ^ n21945 ;
  assign n21977 = n21939 ^ n21937 ;
  assign n21978 = n21977 ^ n18937 ;
  assign n21979 = n21931 ^ n21929 ;
  assign n21980 = n21979 ^ n19683 ;
  assign n21981 = n21924 ^ n21921 ;
  assign n21982 = n21981 ^ n19648 ;
  assign n22021 = n21918 ^ n21864 ;
  assign n21984 = n21913 ^ n21872 ;
  assign n21985 = n21984 ^ n19440 ;
  assign n22010 = n22009 ^ n21986 ;
  assign n22011 = n22009 ^ n19431 ;
  assign n22012 = n22010 & n22011 ;
  assign n22013 = n22012 ^ n19431 ;
  assign n22014 = n22013 ^ n21984 ;
  assign n22015 = ~n21985 & n22014 ;
  assign n22016 = n22015 ^ n19440 ;
  assign n21983 = n21915 ^ n21870 ;
  assign n22017 = n22016 ^ n21983 ;
  assign n22018 = n22016 ^ n19603 ;
  assign n22019 = ~n22017 & n22018 ;
  assign n22020 = n22019 ^ n19603 ;
  assign n22022 = n22021 ^ n22020 ;
  assign n22023 = n22021 ^ n19625 ;
  assign n22024 = n22022 & n22023 ;
  assign n22025 = n22024 ^ n19625 ;
  assign n22026 = n22025 ^ n21981 ;
  assign n22027 = ~n21982 & n22026 ;
  assign n22028 = n22027 ^ n19648 ;
  assign n22029 = n22028 ^ n21979 ;
  assign n22030 = n21980 & ~n22029 ;
  assign n22031 = n22030 ^ n19683 ;
  assign n22032 = n22031 ^ n21977 ;
  assign n22033 = ~n21978 & ~n22032 ;
  assign n22034 = n22033 ^ n18937 ;
  assign n22036 = n22035 ^ n22034 ;
  assign n22037 = n22035 ^ n18962 ;
  assign n22038 = ~n22036 & n22037 ;
  assign n22039 = n22038 ^ n18962 ;
  assign n22040 = n22039 ^ n21975 ;
  assign n22041 = n21976 & n22040 ;
  assign n22042 = n22041 ^ n18990 ;
  assign n22044 = n22043 ^ n22042 ;
  assign n22045 = n22043 ^ n19047 ;
  assign n22046 = n22044 & n22045 ;
  assign n22047 = n22046 ^ n19047 ;
  assign n22048 = n22047 ^ n21973 ;
  assign n22049 = ~n21974 & n22048 ;
  assign n22050 = n22049 ^ n19167 ;
  assign n22185 = n22061 ^ n22050 ;
  assign n22063 = n22028 ^ n21980 ;
  assign n22064 = n21983 ^ n19603 ;
  assign n22065 = n22064 ^ n22016 ;
  assign n22066 = n22013 ^ n21985 ;
  assign n22078 = ~n22068 & ~n22077 ;
  assign n22079 = ~n22066 & n22078 ;
  assign n22080 = ~n22065 & ~n22079 ;
  assign n22081 = n22023 ^ n22020 ;
  assign n22082 = ~n22080 & n22081 ;
  assign n22083 = n22025 ^ n21982 ;
  assign n22084 = n22082 & n22083 ;
  assign n22085 = n22063 & ~n22084 ;
  assign n22086 = n22031 ^ n21978 ;
  assign n22087 = ~n22085 & n22086 ;
  assign n22088 = n22037 ^ n22034 ;
  assign n22089 = n22087 & n22088 ;
  assign n22090 = n22039 ^ n21976 ;
  assign n22091 = n22089 & n22090 ;
  assign n22092 = n22045 ^ n22042 ;
  assign n22093 = ~n22091 & n22092 ;
  assign n22094 = n22047 ^ n21974 ;
  assign n22095 = ~n22093 & ~n22094 ;
  assign n22188 = n22185 ^ n22095 ;
  assign n22189 = ~n19145 & n22188 ;
  assign n22186 = n22095 ^ n22050 ;
  assign n22187 = n22185 & ~n22186 ;
  assign n22190 = n22189 ^ n22187 ;
  assign n22200 = n22199 ^ n22190 ;
  assign n22184 = n2696 ^ n1826 ;
  assign n22201 = n22200 ^ n22184 ;
  assign n22051 = n22050 ^ n19145 ;
  assign n22062 = n22061 ^ n22051 ;
  assign n22096 = n22095 ^ n22062 ;
  assign n22097 = n22096 ^ n2696 ;
  assign n22098 = n22086 ^ n22085 ;
  assign n2870 = n2827 ^ n2557 ;
  assign n2871 = n2870 ^ n2866 ;
  assign n2872 = n2871 ^ x455 ;
  assign n22099 = n22098 ^ n2872 ;
  assign n22103 = n22084 ^ n22063 ;
  assign n22104 = n22103 ^ n2861 ;
  assign n22105 = n22083 ^ n22082 ;
  assign n22106 = n22105 ^ n1445 ;
  assign n22107 = n22081 ^ n22080 ;
  assign n22108 = n22107 ^ n1427 ;
  assign n22111 = n22079 ^ n22065 ;
  assign n1155 = n1154 ^ n1067 ;
  assign n1156 = n1155 ^ n1148 ;
  assign n1157 = n1156 ^ x459 ;
  assign n22112 = n22111 ^ n1157 ;
  assign n1414 = n1295 ^ n1203 ;
  assign n1415 = n1414 ^ n968 ;
  assign n1416 = n1415 ^ x460 ;
  assign n22145 = n22111 ^ n1416 ;
  assign n22113 = n22078 ^ n22066 ;
  assign n22114 = n22113 ^ n1416 ;
  assign n22116 = n22115 ^ n977 ;
  assign n22141 = ~n22116 & n22140 ;
  assign n22142 = n22141 ^ n977 ;
  assign n22143 = n22142 ^ n1416 ;
  assign n22144 = n22114 & n22143 ;
  assign n22146 = n22145 ^ n22144 ;
  assign n22147 = n22112 & ~n22146 ;
  assign n22148 = n22147 ^ n1157 ;
  assign n22109 = n22105 ^ n1427 ;
  assign n22110 = n22109 ^ n22105 ;
  assign n22149 = n22148 ^ n22110 ;
  assign n22150 = n22108 & n22149 ;
  assign n22151 = n22150 ^ n22109 ;
  assign n22152 = ~n22106 & ~n22151 ;
  assign n22153 = n22152 ^ n22105 ;
  assign n22154 = n22153 ^ n22103 ;
  assign n22155 = ~n22104 & ~n22154 ;
  assign n22156 = n22155 ^ n2861 ;
  assign n22100 = n22088 ^ n22087 ;
  assign n22101 = n22100 ^ n2872 ;
  assign n22102 = n22101 ^ n22100 ;
  assign n22157 = n22156 ^ n22102 ;
  assign n22158 = n22099 & n22157 ;
  assign n22159 = n22158 ^ n22101 ;
  assign n22160 = n22090 ^ n22089 ;
  assign n2572 = n2565 ^ n2484 ;
  assign n2576 = n2575 ^ n2572 ;
  assign n2577 = n2576 ^ x454 ;
  assign n22162 = n22160 ^ n2577 ;
  assign n22161 = n22160 ^ n22100 ;
  assign n22163 = n22162 ^ n22161 ;
  assign n22164 = n22159 & ~n22163 ;
  assign n22165 = n22164 ^ n22162 ;
  assign n22166 = n22092 ^ n22091 ;
  assign n22168 = n22166 ^ n2630 ;
  assign n22167 = n22166 ^ n22160 ;
  assign n22169 = n22168 ^ n22167 ;
  assign n22170 = n22165 & ~n22169 ;
  assign n22171 = n22170 ^ n22168 ;
  assign n22172 = n22094 ^ n22093 ;
  assign n22174 = n22172 ^ n2498 ;
  assign n22173 = n22172 ^ n22166 ;
  assign n22175 = n22174 ^ n22173 ;
  assign n22176 = n22171 & ~n22175 ;
  assign n22177 = n22176 ^ n22174 ;
  assign n22179 = n22172 ^ n22096 ;
  assign n22178 = n22096 ^ n3188 ;
  assign n22180 = n22179 ^ n22178 ;
  assign n22181 = n22177 & ~n22180 ;
  assign n22182 = n22181 ^ n22178 ;
  assign n22183 = n22097 & ~n22182 ;
  assign n22202 = n22201 ^ n22183 ;
  assign n22205 = n22204 ^ n22202 ;
  assign n22222 = n22182 ^ n2696 ;
  assign n22232 = n22222 ^ n22202 ;
  assign n22208 = n20457 ^ n20423 ;
  assign n22209 = n22208 ^ n21271 ;
  assign n22210 = n22165 ^ n2630 ;
  assign n22211 = ~n22209 & ~n22210 ;
  assign n22206 = n20472 ^ n20452 ;
  assign n22207 = n22206 ^ n21610 ;
  assign n22212 = n22211 ^ n22207 ;
  assign n22216 = n22171 ^ n2498 ;
  assign n22213 = n22177 ^ n3188 ;
  assign n22214 = n22213 ^ n22207 ;
  assign n22215 = n22214 ^ n22213 ;
  assign n22217 = n22216 ^ n22215 ;
  assign n22218 = n22212 & ~n22217 ;
  assign n22219 = n22218 ^ n22214 ;
  assign n22224 = n22222 ^ n22213 ;
  assign n22220 = n20517 ^ n20450 ;
  assign n22221 = n22220 ^ n21265 ;
  assign n22223 = n22222 ^ n22221 ;
  assign n22225 = n22224 ^ n22223 ;
  assign n22226 = ~n22219 & ~n22225 ;
  assign n22227 = n22226 ^ n22224 ;
  assign n22228 = n20468 ^ n20443 ;
  assign n22229 = n22228 ^ n21260 ;
  assign n22230 = n22229 ^ n22222 ;
  assign n22231 = ~n22227 & ~n22230 ;
  assign n22233 = n22232 ^ n22231 ;
  assign n22234 = n22205 & n22233 ;
  assign n22236 = n22235 ^ n22234 ;
  assign n22237 = n21860 & ~n22236 ;
  assign n21857 = n21856 ^ n21855 ;
  assign n22238 = n22237 ^ n21857 ;
  assign n21853 = n21015 ^ n20453 ;
  assign n21854 = n21853 ^ n21628 ;
  assign n22271 = n21855 ^ n21854 ;
  assign n22272 = ~n22238 & n22271 ;
  assign n22275 = n22274 ^ n22272 ;
  assign n22276 = n21125 ^ n20448 ;
  assign n22277 = n22276 ^ n21636 ;
  assign n22299 = n22277 ^ n22273 ;
  assign n22300 = n22275 & ~n22299 ;
  assign n22303 = n22302 ^ n22300 ;
  assign n22353 = n21822 ^ n21795 ;
  assign n22354 = n22353 ^ n22301 ;
  assign n22304 = n21133 ^ n20441 ;
  assign n22305 = n22304 ^ n21736 ;
  assign n22355 = n22354 ^ n22305 ;
  assign n22356 = n22355 ^ n22353 ;
  assign n22357 = ~n22303 & n22356 ;
  assign n22358 = n22357 ^ n22354 ;
  assign n22359 = n21248 ^ n20435 ;
  assign n22360 = n22359 ^ n21753 ;
  assign n22487 = n22360 ^ n22353 ;
  assign n22488 = ~n22358 & ~n22487 ;
  assign n22489 = n22488 ^ n22353 ;
  assign n22490 = n22489 ^ n22482 ;
  assign n22491 = n22490 ^ n22413 ;
  assign n22492 = n22491 ^ n22482 ;
  assign n22493 = ~n22486 & ~n22492 ;
  assign n22494 = n22493 ^ n22490 ;
  assign n22495 = ~n22483 & n22494 ;
  assign n22496 = n22495 ^ n22482 ;
  assign n22497 = n22496 ^ n22408 ;
  assign n22498 = n22479 & n22497 ;
  assign n22500 = n22499 ^ n22498 ;
  assign n22474 = n21300 ^ n20486 ;
  assign n22475 = n22474 ^ n21882 ;
  assign n22598 = n22500 ^ n22475 ;
  assign n22599 = n22598 ^ n19985 ;
  assign n22600 = n22496 ^ n22479 ;
  assign n22601 = n22600 ^ n19908 ;
  assign n22602 = n22494 ^ n22481 ;
  assign n22603 = n22602 ^ n19938 ;
  assign n22361 = n22360 ^ n22358 ;
  assign n22362 = n22361 ^ n19944 ;
  assign n22306 = n22305 ^ n22303 ;
  assign n22307 = n22306 ^ n19948 ;
  assign n22278 = n22277 ^ n22275 ;
  assign n22279 = n22278 ^ n19956 ;
  assign n22239 = n22238 ^ n21854 ;
  assign n22240 = n22239 ^ n19960 ;
  assign n22241 = n22236 ^ n21859 ;
  assign n22242 = n22241 ^ n19889 ;
  assign n22243 = n22233 ^ n22204 ;
  assign n22244 = n22243 ^ n19789 ;
  assign n22257 = n22229 ^ n22227 ;
  assign n22245 = n22221 ^ n22219 ;
  assign n22246 = n22245 ^ n19723 ;
  assign n22247 = n22210 ^ n22209 ;
  assign n22248 = n19068 & n22247 ;
  assign n22249 = n22248 ^ n19057 ;
  assign n22250 = n22216 ^ n22212 ;
  assign n22251 = n22250 ^ n22248 ;
  assign n22252 = n22249 & n22251 ;
  assign n22253 = n22252 ^ n19057 ;
  assign n22254 = n22253 ^ n22245 ;
  assign n22255 = ~n22246 & n22254 ;
  assign n22256 = n22255 ^ n19723 ;
  assign n22258 = n22257 ^ n22256 ;
  assign n22259 = n22257 ^ n19772 ;
  assign n22260 = ~n22258 & n22259 ;
  assign n22261 = n22260 ^ n19772 ;
  assign n22262 = n22261 ^ n22243 ;
  assign n22263 = ~n22244 & ~n22262 ;
  assign n22264 = n22263 ^ n19789 ;
  assign n22265 = n22264 ^ n22241 ;
  assign n22266 = n22242 & ~n22265 ;
  assign n22267 = n22266 ^ n19889 ;
  assign n22268 = n22267 ^ n22239 ;
  assign n22269 = n22240 & n22268 ;
  assign n22270 = n22269 ^ n19960 ;
  assign n22296 = n22278 ^ n22270 ;
  assign n22297 = n22279 & ~n22296 ;
  assign n22298 = n22297 ^ n19956 ;
  assign n22350 = n22306 ^ n22298 ;
  assign n22351 = n22307 & n22350 ;
  assign n22352 = n22351 ^ n19948 ;
  assign n22605 = n22361 ^ n22352 ;
  assign n22606 = ~n22362 & ~n22605 ;
  assign n22607 = n22606 ^ n19944 ;
  assign n22604 = n22489 ^ n22486 ;
  assign n22608 = n22607 ^ n22604 ;
  assign n22609 = n22607 ^ n19942 ;
  assign n22610 = n22608 & ~n22609 ;
  assign n22611 = n22610 ^ n19942 ;
  assign n22612 = n22611 ^ n22602 ;
  assign n22613 = n22603 & n22612 ;
  assign n22614 = n22613 ^ n19938 ;
  assign n22615 = n22614 ^ n22600 ;
  assign n22616 = n22601 & n22615 ;
  assign n22617 = n22616 ^ n19908 ;
  assign n22618 = n22617 ^ n22598 ;
  assign n22619 = ~n22599 & ~n22618 ;
  assign n22620 = n22619 ^ n19985 ;
  assign n22476 = n22475 ^ n22404 ;
  assign n22501 = n22476 & ~n22500 ;
  assign n22502 = n22501 ^ n22475 ;
  assign n22471 = n21256 ^ n20482 ;
  assign n22472 = n22471 ^ n21875 ;
  assign n22398 = n21836 ^ n21780 ;
  assign n22473 = n22472 ^ n22398 ;
  assign n22596 = n22502 ^ n22473 ;
  assign n22597 = n22596 ^ n19931 ;
  assign n22694 = n22620 ^ n22597 ;
  assign n22684 = n22611 ^ n22603 ;
  assign n22685 = n22604 ^ n19942 ;
  assign n22686 = n22685 ^ n22607 ;
  assign n22363 = n22362 ^ n22352 ;
  assign n22308 = n22307 ^ n22298 ;
  assign n22280 = n22279 ^ n22270 ;
  assign n22281 = n22259 ^ n22256 ;
  assign n22282 = n22253 ^ n22246 ;
  assign n22283 = n22247 ^ n19068 ;
  assign n22284 = n22250 ^ n22249 ;
  assign n22285 = n22283 & ~n22284 ;
  assign n22286 = ~n22282 & n22285 ;
  assign n22287 = n22281 & n22286 ;
  assign n22288 = n22261 ^ n22244 ;
  assign n22289 = n22287 & ~n22288 ;
  assign n22290 = n22264 ^ n22242 ;
  assign n22291 = ~n22289 & n22290 ;
  assign n22292 = n22267 ^ n22240 ;
  assign n22293 = ~n22291 & ~n22292 ;
  assign n22309 = ~n22280 & ~n22293 ;
  assign n22364 = ~n22308 & n22309 ;
  assign n22687 = ~n22363 & n22364 ;
  assign n22688 = n22686 & ~n22687 ;
  assign n22689 = n22684 & ~n22688 ;
  assign n22690 = n22614 ^ n22601 ;
  assign n22691 = ~n22689 & n22690 ;
  assign n22692 = n22617 ^ n22599 ;
  assign n22693 = ~n22691 & ~n22692 ;
  assign n22767 = n22694 ^ n22693 ;
  assign n22794 = n22767 ^ n2956 ;
  assign n22769 = n22692 ^ n22691 ;
  assign n22770 = n22769 ^ n2956 ;
  assign n22771 = n22690 ^ n22689 ;
  assign n22772 = n22771 ^ n606 ;
  assign n22773 = n22688 ^ n22684 ;
  assign n22777 = n22776 ^ n22773 ;
  assign n22778 = n22687 ^ n22686 ;
  assign n22779 = n22778 ^ n1475 ;
  assign n22365 = n22364 ^ n22363 ;
  assign n22782 = n22778 ^ n22365 ;
  assign n22294 = n22293 ^ n22280 ;
  assign n2400 = n2321 ^ n2274 ;
  assign n2401 = n2400 ^ n2204 ;
  assign n2402 = n2401 ^ x505 ;
  assign n22295 = n22294 ^ n2402 ;
  assign n22313 = n22292 ^ n22291 ;
  assign n22314 = n22313 ^ n2409 ;
  assign n22315 = n22290 ^ n22289 ;
  assign n2076 = n2075 ^ n2021 ;
  assign n2080 = n2079 ^ n2076 ;
  assign n2081 = n2080 ^ x507 ;
  assign n22316 = n22315 ^ n2081 ;
  assign n22317 = n20390 ^ n2244 ;
  assign n22318 = n22317 ^ n1987 ;
  assign n22319 = n22318 ^ x508 ;
  assign n22340 = n22319 ^ n22315 ;
  assign n22320 = n22288 ^ n22287 ;
  assign n22321 = n22320 ^ n22319 ;
  assign n22322 = n22286 ^ n22281 ;
  assign n1978 = n1974 ^ n1938 ;
  assign n1982 = n1981 ^ n1978 ;
  assign n1983 = n1982 ^ x509 ;
  assign n22323 = n22322 ^ n1983 ;
  assign n22324 = n22285 ^ n22282 ;
  assign n1925 = n1909 ^ n1894 ;
  assign n1926 = n1925 ^ n1922 ;
  assign n1927 = n1926 ^ x510 ;
  assign n22325 = n22324 ^ n1927 ;
  assign n22326 = n3030 & ~n22283 ;
  assign n1913 = n1885 ^ x511 ;
  assign n1917 = n1916 ^ n1913 ;
  assign n1918 = n1917 ^ n1903 ;
  assign n22327 = n22326 ^ n1918 ;
  assign n22328 = n22284 ^ n22283 ;
  assign n22329 = n22328 ^ n22326 ;
  assign n22330 = n22327 & n22329 ;
  assign n22331 = n22330 ^ n1918 ;
  assign n22332 = n22331 ^ n1927 ;
  assign n22333 = ~n22325 & ~n22332 ;
  assign n22334 = n22333 ^ n22324 ;
  assign n22335 = n22334 ^ n22322 ;
  assign n22336 = n22323 & n22335 ;
  assign n22337 = n22336 ^ n1983 ;
  assign n22338 = n22337 ^ n22319 ;
  assign n22339 = ~n22321 & n22338 ;
  assign n22341 = n22340 ^ n22339 ;
  assign n22342 = n22316 & n22341 ;
  assign n22343 = n22342 ^ n22315 ;
  assign n22344 = n22343 ^ n22313 ;
  assign n22345 = n22314 & ~n22344 ;
  assign n22346 = n22345 ^ n2409 ;
  assign n22310 = n22309 ^ n22308 ;
  assign n22311 = n22310 ^ n2402 ;
  assign n22312 = n22311 ^ n22310 ;
  assign n22347 = n22346 ^ n22312 ;
  assign n22348 = ~n22295 & n22347 ;
  assign n22349 = n22348 ^ n22311 ;
  assign n2426 = n2347 ^ n1451 ;
  assign n2427 = n2426 ^ n2420 ;
  assign n2428 = n2427 ^ x504 ;
  assign n22367 = n22365 ^ n2428 ;
  assign n22366 = n22365 ^ n22310 ;
  assign n22368 = n22367 ^ n22366 ;
  assign n22369 = ~n22349 & n22368 ;
  assign n22370 = n22369 ^ n22367 ;
  assign n22780 = n22373 ^ n22365 ;
  assign n22781 = n22370 & n22780 ;
  assign n22783 = n22782 ^ n22781 ;
  assign n22784 = ~n22779 & n22783 ;
  assign n22785 = n22784 ^ n1475 ;
  assign n22786 = n22785 ^ n22773 ;
  assign n22787 = n22777 & ~n22786 ;
  assign n22788 = n22787 ^ n22776 ;
  assign n22789 = n22788 ^ n22771 ;
  assign n22790 = ~n22772 & n22789 ;
  assign n22791 = n22790 ^ n606 ;
  assign n22792 = n22791 ^ n2956 ;
  assign n22793 = ~n22770 & n22792 ;
  assign n22795 = n22794 ^ n22793 ;
  assign n23197 = n22795 ^ n542 ;
  assign n23169 = n22791 ^ n22770 ;
  assign n23198 = n23197 ^ n23169 ;
  assign n23015 = n22788 ^ n22772 ;
  assign n23013 = n21922 ^ n21285 ;
  assign n22444 = n22133 ^ n22120 ;
  assign n23014 = n23013 ^ n22444 ;
  assign n23016 = n23015 ^ n23014 ;
  assign n23170 = n23169 ^ n23015 ;
  assign n23171 = n23170 ^ n23169 ;
  assign n23003 = n22785 ^ n22777 ;
  assign n22918 = n22783 ^ n1475 ;
  assign n23004 = n23003 ^ n22918 ;
  assign n22919 = n21863 ^ n21295 ;
  assign n22452 = n22127 ^ n22124 ;
  assign n22920 = n22919 ^ n22452 ;
  assign n22921 = n22920 ^ n22918 ;
  assign n22374 = n22373 ^ n22370 ;
  assign n21851 = n21850 ^ n1552 ;
  assign n21257 = n21256 ^ n21255 ;
  assign n21852 = n21851 ^ n21257 ;
  assign n22375 = n22374 ^ n21852 ;
  assign n22379 = n21847 ^ n21748 ;
  assign n22378 = n21873 ^ n21300 ;
  assign n22380 = n22379 ^ n22378 ;
  assign n22376 = n22349 ^ n2428 ;
  assign n22381 = n22380 ^ n22376 ;
  assign n22385 = n22346 ^ n22295 ;
  assign n22383 = n21844 ^ n21768 ;
  assign n22382 = n21875 ^ n21306 ;
  assign n22384 = n22383 ^ n22382 ;
  assign n22386 = n22385 ^ n22384 ;
  assign n22390 = n22343 ^ n22314 ;
  assign n22388 = n21841 ^ n21773 ;
  assign n22387 = n21882 ^ n21308 ;
  assign n22389 = n22388 ^ n22387 ;
  assign n22391 = n22390 ^ n22389 ;
  assign n22395 = n22341 ^ n2081 ;
  assign n22906 = n22395 ^ n22390 ;
  assign n22393 = n21839 ^ n593 ;
  assign n22392 = n21884 ^ n21314 ;
  assign n22394 = n22393 ^ n22392 ;
  assign n22396 = n22395 ^ n22394 ;
  assign n22399 = n22398 ^ n21891 ;
  assign n22400 = n22399 ^ n21248 ;
  assign n22397 = n22337 ^ n22321 ;
  assign n22401 = n22400 ^ n22397 ;
  assign n22402 = n22334 ^ n22323 ;
  assign n22900 = n22402 ^ n22397 ;
  assign n22403 = n21893 ^ n21133 ;
  assign n22405 = n22404 ^ n22403 ;
  assign n22406 = n22405 ^ n22402 ;
  assign n22410 = n22331 ^ n22325 ;
  assign n22407 = n21753 ^ n21125 ;
  assign n22409 = n22408 ^ n22407 ;
  assign n22411 = n22410 ^ n22409 ;
  assign n22887 = n22328 ^ n22327 ;
  assign n22414 = n22413 ^ n21636 ;
  assign n22415 = n22414 ^ n20433 ;
  assign n22412 = n22283 ^ n3030 ;
  assign n22416 = n22415 ^ n22412 ;
  assign n22431 = n22142 ^ n22114 ;
  assign n22429 = n20947 ^ n20258 ;
  assign n22430 = n22429 ^ n22053 ;
  assign n22432 = n22431 ^ n22430 ;
  assign n22437 = n21485 ^ n20977 ;
  assign n22438 = n22437 ^ n21965 ;
  assign n22439 = n22438 ^ n22436 ;
  assign n22441 = n21372 ^ n20921 ;
  assign n22442 = n22441 ^ n21957 ;
  assign n22440 = n22136 ^ n22118 ;
  assign n22443 = n22442 ^ n22440 ;
  assign n22529 = n22444 ^ n22440 ;
  assign n22445 = n21365 ^ n20901 ;
  assign n22446 = n22445 ^ n21949 ;
  assign n22447 = n22446 ^ n22444 ;
  assign n22449 = n21357 ^ n20877 ;
  assign n22450 = n22449 ^ n21940 ;
  assign n22448 = n22130 ^ n22122 ;
  assign n22451 = n22450 ^ n22448 ;
  assign n22453 = n21347 ^ n20856 ;
  assign n22454 = n22453 ^ n21932 ;
  assign n22455 = n22454 ^ n22452 ;
  assign n22520 = n22452 ^ n21851 ;
  assign n22456 = n21282 ^ n20835 ;
  assign n22457 = n22456 ^ n21922 ;
  assign n22458 = n22457 ^ n21851 ;
  assign n22459 = n21278 ^ n20715 ;
  assign n22460 = n22459 ^ n21865 ;
  assign n22461 = n22460 ^ n22379 ;
  assign n22514 = n22383 ^ n22379 ;
  assign n22462 = n21285 ^ n20667 ;
  assign n22463 = n22462 ^ n21863 ;
  assign n22464 = n22463 ^ n22383 ;
  assign n22465 = n21289 ^ n20479 ;
  assign n22466 = n22465 ^ n21255 ;
  assign n22467 = n22466 ^ n22388 ;
  assign n22468 = n21295 ^ n20475 ;
  assign n22469 = n22468 ^ n21873 ;
  assign n22470 = n22469 ^ n22393 ;
  assign n22505 = n22398 ^ n22393 ;
  assign n22503 = n22502 ^ n22472 ;
  assign n22504 = ~n22473 & n22503 ;
  assign n22506 = n22505 ^ n22504 ;
  assign n22507 = n22470 & ~n22506 ;
  assign n22508 = n22507 ^ n22393 ;
  assign n22509 = n22508 ^ n22466 ;
  assign n22510 = ~n22467 & ~n22509 ;
  assign n22511 = n22510 ^ n22388 ;
  assign n22512 = n22511 ^ n22463 ;
  assign n22513 = n22464 & n22512 ;
  assign n22515 = n22514 ^ n22513 ;
  assign n22516 = n22461 & n22515 ;
  assign n22517 = n22516 ^ n22379 ;
  assign n22518 = n22517 ^ n22457 ;
  assign n22519 = ~n22458 & n22518 ;
  assign n22521 = n22520 ^ n22519 ;
  assign n22522 = ~n22455 & ~n22521 ;
  assign n22523 = n22522 ^ n22454 ;
  assign n22524 = n22523 ^ n22448 ;
  assign n22525 = n22451 & ~n22524 ;
  assign n22526 = n22525 ^ n22450 ;
  assign n22527 = n22526 ^ n22444 ;
  assign n22528 = n22447 & ~n22527 ;
  assign n22530 = n22529 ^ n22528 ;
  assign n22531 = n22443 & ~n22530 ;
  assign n22532 = n22531 ^ n22442 ;
  assign n22533 = n22532 ^ n22436 ;
  assign n22534 = n22439 & n22533 ;
  assign n22535 = n22534 ^ n22438 ;
  assign n22433 = n22146 ^ n1157 ;
  assign n22434 = n22433 ^ n22431 ;
  assign n22435 = n22434 ^ n22433 ;
  assign n22536 = n22535 ^ n22435 ;
  assign n22537 = n22432 & ~n22536 ;
  assign n22538 = n22537 ^ n22434 ;
  assign n22539 = n22148 ^ n22108 ;
  assign n22543 = n22539 ^ n22433 ;
  assign n22540 = n20952 ^ n20263 ;
  assign n22541 = n22540 ^ n22196 ;
  assign n22542 = n22541 ^ n22539 ;
  assign n22544 = n22543 ^ n22542 ;
  assign n22545 = n22538 & ~n22544 ;
  assign n22546 = n22545 ^ n22543 ;
  assign n22547 = n22151 ^ n1445 ;
  assign n22551 = n22547 ^ n22539 ;
  assign n22548 = n20950 ^ n20253 ;
  assign n22549 = n22548 ^ n21591 ;
  assign n22550 = n22549 ^ n22547 ;
  assign n22552 = n22551 ^ n22550 ;
  assign n22553 = n22546 & n22552 ;
  assign n22554 = n22553 ^ n22551 ;
  assign n22555 = n22153 ^ n22104 ;
  assign n22559 = n22555 ^ n22547 ;
  assign n22556 = n20941 ^ n20292 ;
  assign n22557 = n22556 ^ n21594 ;
  assign n22558 = n22557 ^ n22555 ;
  assign n22560 = n22559 ^ n22558 ;
  assign n22561 = ~n22554 & n22560 ;
  assign n22562 = n22561 ^ n22559 ;
  assign n22563 = n22156 ^ n22099 ;
  assign n22567 = n22563 ^ n22555 ;
  assign n22564 = n20988 ^ n20342 ;
  assign n22565 = n22564 ^ n21583 ;
  assign n22566 = n22565 ^ n22563 ;
  assign n22568 = n22567 ^ n22566 ;
  assign n22569 = ~n22562 & n22568 ;
  assign n22570 = n22569 ^ n22567 ;
  assign n22426 = n20467 ^ n20357 ;
  assign n22427 = n22426 ^ n21578 ;
  assign n22850 = n22563 ^ n22427 ;
  assign n22851 = ~n22570 & ~n22850 ;
  assign n22572 = n22565 ^ n22562 ;
  assign n22573 = n22572 ^ n19695 ;
  assign n22575 = n22549 ^ n22546 ;
  assign n22576 = n22575 ^ n19635 ;
  assign n22578 = n22535 ^ n22432 ;
  assign n22579 = n22578 ^ n19638 ;
  assign n22580 = n22532 ^ n22439 ;
  assign n22581 = n22580 ^ n20323 ;
  assign n22582 = n22530 ^ n22442 ;
  assign n22583 = n22582 ^ n20271 ;
  assign n22647 = n22526 ^ n22447 ;
  assign n22584 = n22523 ^ n22451 ;
  assign n22585 = n22584 ^ n20018 ;
  assign n22639 = n22521 ^ n22454 ;
  assign n22586 = n22517 ^ n22458 ;
  assign n22587 = n22586 ^ n20008 ;
  assign n22588 = n22515 ^ n22460 ;
  assign n22589 = n22588 ^ n19914 ;
  assign n22590 = n22511 ^ n22464 ;
  assign n22591 = n22590 ^ n19918 ;
  assign n22592 = n22508 ^ n22467 ;
  assign n22593 = n22592 ^ n19922 ;
  assign n22594 = n22506 ^ n22469 ;
  assign n22595 = n22594 ^ n19926 ;
  assign n22621 = n22620 ^ n22596 ;
  assign n22622 = ~n22597 & ~n22621 ;
  assign n22623 = n22622 ^ n19931 ;
  assign n22624 = n22623 ^ n22594 ;
  assign n22625 = ~n22595 & ~n22624 ;
  assign n22626 = n22625 ^ n19926 ;
  assign n22627 = n22626 ^ n22592 ;
  assign n22628 = n22593 & n22627 ;
  assign n22629 = n22628 ^ n19922 ;
  assign n22630 = n22629 ^ n22590 ;
  assign n22631 = n22591 & ~n22630 ;
  assign n22632 = n22631 ^ n19918 ;
  assign n22633 = n22632 ^ n22588 ;
  assign n22634 = ~n22589 & n22633 ;
  assign n22635 = n22634 ^ n19914 ;
  assign n22636 = n22635 ^ n22586 ;
  assign n22637 = n22587 & ~n22636 ;
  assign n22638 = n22637 ^ n20008 ;
  assign n22640 = n22639 ^ n22638 ;
  assign n22641 = n22639 ^ n20015 ;
  assign n22642 = ~n22640 & n22641 ;
  assign n22643 = n22642 ^ n20015 ;
  assign n22644 = n22643 ^ n22584 ;
  assign n22645 = n22585 & ~n22644 ;
  assign n22646 = n22645 ^ n20018 ;
  assign n22648 = n22647 ^ n22646 ;
  assign n22649 = n22647 ^ n20239 ;
  assign n22650 = ~n22648 & ~n22649 ;
  assign n22651 = n22650 ^ n20239 ;
  assign n22652 = n22651 ^ n22582 ;
  assign n22653 = ~n22583 & ~n22652 ;
  assign n22654 = n22653 ^ n20271 ;
  assign n22655 = n22654 ^ n22580 ;
  assign n22656 = ~n22581 & n22655 ;
  assign n22657 = n22656 ^ n20323 ;
  assign n22658 = n22657 ^ n22578 ;
  assign n22659 = ~n22579 & ~n22658 ;
  assign n22660 = n22659 ^ n19638 ;
  assign n22577 = n22541 ^ n22538 ;
  assign n22661 = n22660 ^ n22577 ;
  assign n22662 = n22660 ^ n19613 ;
  assign n22663 = n22661 & n22662 ;
  assign n22664 = n22663 ^ n19613 ;
  assign n22665 = n22664 ^ n22575 ;
  assign n22666 = ~n22576 & ~n22665 ;
  assign n22667 = n22666 ^ n19635 ;
  assign n22574 = n22557 ^ n22554 ;
  assign n22668 = n22667 ^ n22574 ;
  assign n22669 = n22667 ^ n19668 ;
  assign n22670 = n22668 & n22669 ;
  assign n22671 = n22670 ^ n19668 ;
  assign n22672 = n22671 ^ n22572 ;
  assign n22673 = ~n22573 & ~n22672 ;
  assign n22674 = n22673 ^ n19695 ;
  assign n22675 = n22674 ^ n19079 ;
  assign n22571 = n22570 ^ n22427 ;
  assign n22847 = n22674 ^ n22571 ;
  assign n22848 = n22675 & n22847 ;
  assign n22677 = n22574 ^ n19668 ;
  assign n22678 = n22677 ^ n22667 ;
  assign n22679 = n22577 ^ n19613 ;
  assign n22680 = n22679 ^ n22660 ;
  assign n22681 = n22651 ^ n22583 ;
  assign n22682 = n22649 ^ n22646 ;
  assign n22683 = n22641 ^ n22638 ;
  assign n22695 = n22693 & n22694 ;
  assign n22696 = n22623 ^ n22595 ;
  assign n22697 = n22695 & ~n22696 ;
  assign n22698 = n22626 ^ n22593 ;
  assign n22699 = n22697 & ~n22698 ;
  assign n22700 = n22629 ^ n22591 ;
  assign n22701 = ~n22699 & ~n22700 ;
  assign n22702 = n22632 ^ n22589 ;
  assign n22703 = n22701 & n22702 ;
  assign n22704 = n22635 ^ n22587 ;
  assign n22705 = ~n22703 & n22704 ;
  assign n22706 = n22683 & n22705 ;
  assign n22707 = n22643 ^ n22585 ;
  assign n22708 = ~n22706 & ~n22707 ;
  assign n22709 = ~n22682 & ~n22708 ;
  assign n22710 = n22681 & n22709 ;
  assign n22711 = n22654 ^ n22581 ;
  assign n22712 = ~n22710 & n22711 ;
  assign n22713 = n22657 ^ n22579 ;
  assign n22714 = ~n22712 & ~n22713 ;
  assign n22715 = n22680 & n22714 ;
  assign n22716 = n22664 ^ n22576 ;
  assign n22717 = n22715 & n22716 ;
  assign n22718 = n22678 & ~n22717 ;
  assign n22719 = n22671 ^ n22573 ;
  assign n22720 = ~n22718 & ~n22719 ;
  assign n22676 = n22675 ^ n22571 ;
  assign n22723 = n22720 ^ n22676 ;
  assign n22724 = n22723 ^ n2748 ;
  assign n22725 = n22719 ^ n22718 ;
  assign n22726 = n22725 ^ n2675 ;
  assign n22728 = n22717 ^ n22678 ;
  assign n2667 = n2605 ^ n2528 ;
  assign n2668 = n2667 ^ n1835 ;
  assign n2669 = n2668 ^ x484 ;
  assign n22729 = n22728 ^ n2669 ;
  assign n22731 = n20871 ^ n2586 ;
  assign n22732 = n22731 ^ n3121 ;
  assign n22733 = n22732 ^ x485 ;
  assign n22730 = n22716 ^ n22715 ;
  assign n22734 = n22733 ^ n22730 ;
  assign n22736 = n22714 ^ n22680 ;
  assign n22737 = n22736 ^ n3101 ;
  assign n22739 = n3109 ^ n2886 ;
  assign n22740 = n22739 ^ n2507 ;
  assign n22741 = n22740 ^ x487 ;
  assign n22738 = n22713 ^ n22712 ;
  assign n22742 = n22741 ^ n22738 ;
  assign n22745 = n22711 ^ n22710 ;
  assign n22749 = n22748 ^ n22745 ;
  assign n22750 = n22709 ^ n22681 ;
  assign n22751 = n22750 ^ n2639 ;
  assign n22753 = n22707 ^ n22706 ;
  assign n22754 = n22753 ^ n1247 ;
  assign n22815 = n22753 ^ n1082 ;
  assign n22755 = n22705 ^ n22683 ;
  assign n22756 = n22755 ^ n1082 ;
  assign n22757 = n22704 ^ n22703 ;
  assign n22758 = n22757 ^ n963 ;
  assign n22809 = n22757 ^ n948 ;
  assign n22759 = n22702 ^ n22701 ;
  assign n22760 = n22759 ^ n948 ;
  assign n22761 = n22700 ^ n22699 ;
  assign n22762 = n22761 ^ n939 ;
  assign n22763 = n22698 ^ n22697 ;
  assign n22764 = n22763 ^ n1610 ;
  assign n22765 = n22696 ^ n22695 ;
  assign n22766 = n22765 ^ n1604 ;
  assign n22768 = n22767 ^ n542 ;
  assign n22796 = ~n22768 & ~n22795 ;
  assign n22797 = n22796 ^ n22767 ;
  assign n22798 = n22797 ^ n1604 ;
  assign n22799 = n22766 & n22798 ;
  assign n22800 = n22799 ^ n22765 ;
  assign n22801 = n22800 ^ n1610 ;
  assign n22802 = n22764 & ~n22801 ;
  assign n22803 = n22802 ^ n22763 ;
  assign n22804 = n22803 ^ n939 ;
  assign n22805 = n22762 & ~n22804 ;
  assign n22806 = n22805 ^ n22761 ;
  assign n22807 = n22806 ^ n948 ;
  assign n22808 = n22760 & n22807 ;
  assign n22810 = n22809 ^ n22808 ;
  assign n22811 = n22758 & n22810 ;
  assign n22812 = n22811 ^ n22757 ;
  assign n22813 = n22812 ^ n1082 ;
  assign n22814 = ~n22756 & n22813 ;
  assign n22816 = n22815 ^ n22814 ;
  assign n22817 = n22754 & ~n22816 ;
  assign n22818 = n22817 ^ n1247 ;
  assign n22752 = n22708 ^ n22682 ;
  assign n22819 = n22818 ^ n22752 ;
  assign n1239 = n1238 ^ n1235 ;
  assign n1240 = n1239 ^ n1142 ;
  assign n1241 = n1240 ^ x490 ;
  assign n22820 = n22750 ^ n1241 ;
  assign n22821 = n22820 ^ n22750 ;
  assign n22822 = n22821 ^ n22752 ;
  assign n22823 = n22819 & ~n22822 ;
  assign n22824 = n22823 ^ n22820 ;
  assign n22825 = ~n22751 & n22824 ;
  assign n22826 = n22825 ^ n2639 ;
  assign n22827 = n22826 ^ n22745 ;
  assign n22828 = ~n22749 & n22827 ;
  assign n22829 = n22828 ^ n22748 ;
  assign n22743 = n22741 ^ n22736 ;
  assign n22744 = n22743 ^ n22736 ;
  assign n22830 = n22829 ^ n22744 ;
  assign n22831 = ~n22742 & n22830 ;
  assign n22832 = n22831 ^ n22743 ;
  assign n22833 = ~n22737 & n22832 ;
  assign n22834 = n22833 ^ n3101 ;
  assign n22735 = n22733 ^ n22728 ;
  assign n22835 = n22834 ^ n22735 ;
  assign n22836 = n22835 ^ n22728 ;
  assign n22837 = ~n22734 & n22836 ;
  assign n22838 = n22837 ^ n22735 ;
  assign n22839 = ~n22729 & n22838 ;
  assign n22840 = n22839 ^ n2669 ;
  assign n22727 = n22723 ^ n2675 ;
  assign n22841 = n22840 ^ n22727 ;
  assign n22842 = n22841 ^ n22723 ;
  assign n22843 = ~n22726 & n22842 ;
  assign n22844 = n22843 ^ n22727 ;
  assign n22845 = ~n22724 & n22844 ;
  assign n22721 = n22676 & n22720 ;
  assign n22421 = n22159 ^ n2577 ;
  assign n22419 = n22193 ^ n20465 ;
  assign n22420 = n22419 ^ n21576 ;
  assign n22422 = n22421 ^ n22420 ;
  assign n22423 = n22422 ^ n2738 ;
  assign n22424 = n22423 ^ n2748 ;
  assign n22425 = n22424 ^ n19079 ;
  assign n22428 = n22427 ^ n22425 ;
  assign n22722 = n22721 ^ n22428 ;
  assign n22846 = n22845 ^ n22722 ;
  assign n22849 = n22848 ^ n22846 ;
  assign n22852 = n22851 ^ n22849 ;
  assign n22417 = n21628 ^ n20438 ;
  assign n22418 = n22417 ^ n22353 ;
  assign n22853 = n22852 ^ n22418 ;
  assign n22855 = n21622 ^ n20443 ;
  assign n22856 = n22855 ^ n22301 ;
  assign n22854 = n22844 ^ n2748 ;
  assign n22857 = n22856 ^ n22854 ;
  assign n22862 = n22840 ^ n22726 ;
  assign n22860 = n21262 ^ n20450 ;
  assign n22861 = n22860 ^ n22273 ;
  assign n22863 = n22862 ^ n22861 ;
  assign n22868 = n21260 ^ n20452 ;
  assign n22869 = n22868 ^ n21855 ;
  assign n22864 = n21265 ^ n20457 ;
  assign n22865 = n22864 ^ n21856 ;
  assign n22866 = n22834 ^ n22734 ;
  assign n22867 = n22865 & ~n22866 ;
  assign n22870 = n22869 ^ n22867 ;
  assign n22872 = n22838 ^ n2669 ;
  assign n22871 = n22867 ^ n22862 ;
  assign n22873 = n22872 ^ n22871 ;
  assign n22874 = n22873 ^ n22862 ;
  assign n22875 = n22870 & ~n22874 ;
  assign n22876 = n22875 ^ n22871 ;
  assign n22877 = ~n22863 & ~n22876 ;
  assign n22878 = n22877 ^ n22862 ;
  assign n22879 = n22878 ^ n22854 ;
  assign n22880 = n22857 & n22879 ;
  assign n22858 = n22854 ^ n22852 ;
  assign n22881 = n22880 ^ n22858 ;
  assign n22882 = n22853 & ~n22881 ;
  assign n22883 = n22882 ^ n22852 ;
  assign n22884 = n22883 ^ n22412 ;
  assign n22885 = ~n22416 & n22884 ;
  assign n22886 = n22885 ^ n22415 ;
  assign n22888 = n22887 ^ n22886 ;
  assign n22889 = n21736 ^ n21015 ;
  assign n22890 = n22889 ^ n22482 ;
  assign n22893 = n22890 ^ n22886 ;
  assign n22894 = n22888 & ~n22893 ;
  assign n22891 = n22890 ^ n22410 ;
  assign n22895 = n22894 ^ n22891 ;
  assign n22896 = ~n22411 & n22895 ;
  assign n22897 = n22896 ^ n22410 ;
  assign n22898 = n22897 ^ n22402 ;
  assign n22899 = n22406 & n22898 ;
  assign n22901 = n22900 ^ n22899 ;
  assign n22902 = ~n22401 & ~n22901 ;
  assign n22903 = n22902 ^ n22400 ;
  assign n22904 = n22903 ^ n22395 ;
  assign n22905 = n22396 & n22904 ;
  assign n22907 = n22906 ^ n22905 ;
  assign n22908 = n22391 & n22907 ;
  assign n22909 = n22908 ^ n22390 ;
  assign n22910 = n22909 ^ n22384 ;
  assign n22911 = ~n22386 & ~n22910 ;
  assign n22912 = n22911 ^ n22385 ;
  assign n22913 = n22912 ^ n22376 ;
  assign n22914 = ~n22381 & ~n22913 ;
  assign n22377 = n22376 ^ n22374 ;
  assign n22915 = n22914 ^ n22377 ;
  assign n22916 = ~n22375 & n22915 ;
  assign n22917 = n22916 ^ n22374 ;
  assign n23001 = n22918 ^ n22917 ;
  assign n23002 = ~n22921 & ~n23001 ;
  assign n23005 = n23004 ^ n23002 ;
  assign n23006 = n21865 ^ n21289 ;
  assign n23007 = n23006 ^ n22448 ;
  assign n23010 = n23007 ^ n23003 ;
  assign n23011 = ~n23005 & ~n23010 ;
  assign n23012 = n23011 ^ n23003 ;
  assign n23172 = n23171 ^ n23012 ;
  assign n23173 = ~n23016 & ~n23172 ;
  assign n23174 = n23173 ^ n23170 ;
  assign n23175 = n21932 ^ n21278 ;
  assign n23176 = n23175 ^ n22440 ;
  assign n23195 = n23176 ^ n23169 ;
  assign n23196 = n23174 & n23195 ;
  assign n23199 = n23198 ^ n23196 ;
  assign n23202 = n23201 ^ n23199 ;
  assign n23203 = n23202 ^ n20835 ;
  assign n23008 = n23007 ^ n23005 ;
  assign n22923 = n22915 ^ n21852 ;
  assign n22924 = n22923 ^ n20482 ;
  assign n22925 = n22912 ^ n22381 ;
  assign n22926 = n22925 ^ n20486 ;
  assign n22981 = n22907 ^ n22389 ;
  assign n22928 = n22903 ^ n22396 ;
  assign n22929 = n22928 ^ n19906 ;
  assign n22973 = n22901 ^ n22400 ;
  assign n22931 = n22895 ^ n22409 ;
  assign n22932 = n22931 ^ n20448 ;
  assign n22935 = n22883 ^ n22416 ;
  assign n22936 = n22935 ^ n20458 ;
  assign n22937 = n22881 ^ n22418 ;
  assign n22938 = n22937 ^ n20462 ;
  assign n22940 = n22876 ^ n22861 ;
  assign n22941 = n22940 ^ n20517 ;
  assign n22944 = n22872 ^ n22870 ;
  assign n22942 = n22866 ^ n22865 ;
  assign n22943 = ~n20423 & ~n22942 ;
  assign n22945 = n22944 ^ n22943 ;
  assign n22946 = n22944 ^ n20472 ;
  assign n22947 = n22945 & ~n22946 ;
  assign n22948 = n22947 ^ n20472 ;
  assign n22949 = n22948 ^ n22940 ;
  assign n22950 = ~n22941 & n22949 ;
  assign n22951 = n22950 ^ n20517 ;
  assign n22939 = n22878 ^ n22857 ;
  assign n22952 = n22951 ^ n22939 ;
  assign n22953 = n22951 ^ n20468 ;
  assign n22954 = n22952 & n22953 ;
  assign n22955 = n22954 ^ n20468 ;
  assign n22956 = n22955 ^ n22937 ;
  assign n22957 = ~n22938 & n22956 ;
  assign n22958 = n22957 ^ n20462 ;
  assign n22959 = n22958 ^ n22935 ;
  assign n22960 = n22936 & n22959 ;
  assign n22961 = n22960 ^ n20458 ;
  assign n22933 = n22890 ^ n22887 ;
  assign n22934 = n22933 ^ n22886 ;
  assign n22962 = n22961 ^ n22934 ;
  assign n22963 = n22961 ^ n20453 ;
  assign n22964 = n22962 & n22963 ;
  assign n22965 = n22964 ^ n20453 ;
  assign n22966 = n22965 ^ n22931 ;
  assign n22967 = n22932 & n22966 ;
  assign n22968 = n22967 ^ n20448 ;
  assign n22930 = n22897 ^ n22406 ;
  assign n22969 = n22968 ^ n22930 ;
  assign n22970 = n22968 ^ n20441 ;
  assign n22971 = n22969 & ~n22970 ;
  assign n22972 = n22971 ^ n20441 ;
  assign n22974 = n22973 ^ n22972 ;
  assign n22975 = n22973 ^ n20435 ;
  assign n22976 = n22974 & ~n22975 ;
  assign n22977 = n22976 ^ n20435 ;
  assign n22978 = n22977 ^ n22928 ;
  assign n22979 = n22929 & n22978 ;
  assign n22980 = n22979 ^ n19906 ;
  assign n22982 = n22981 ^ n22980 ;
  assign n22983 = n22981 ^ n20494 ;
  assign n22984 = ~n22982 & ~n22983 ;
  assign n22985 = n22984 ^ n20494 ;
  assign n22927 = n22909 ^ n22386 ;
  assign n22986 = n22985 ^ n22927 ;
  assign n22987 = n22925 ^ n20492 ;
  assign n22988 = n22987 ^ n22925 ;
  assign n22989 = n22988 ^ n22927 ;
  assign n22990 = ~n22986 & n22989 ;
  assign n22991 = n22990 ^ n22987 ;
  assign n22992 = ~n22926 & n22991 ;
  assign n22993 = n22992 ^ n20486 ;
  assign n22994 = n22993 ^ n22923 ;
  assign n22995 = n22924 & ~n22994 ;
  assign n22996 = n22995 ^ n20482 ;
  assign n22922 = n22921 ^ n22917 ;
  assign n22997 = n22996 ^ n22922 ;
  assign n22998 = n22996 ^ n20475 ;
  assign n22999 = ~n22997 & ~n22998 ;
  assign n23000 = n22999 ^ n20475 ;
  assign n23009 = n23008 ^ n23000 ;
  assign n23017 = n23016 ^ n23012 ;
  assign n23018 = n23017 ^ n20479 ;
  assign n23019 = n23018 ^ n23017 ;
  assign n23020 = n23019 ^ n23000 ;
  assign n23021 = ~n23009 & n23020 ;
  assign n23022 = n23021 ^ n23018 ;
  assign n23179 = n23017 ^ n20667 ;
  assign n23180 = n23022 & n23179 ;
  assign n23181 = n23180 ^ n20667 ;
  assign n23177 = n23176 ^ n23174 ;
  assign n23191 = n23181 ^ n23177 ;
  assign n23192 = n23181 ^ n20715 ;
  assign n23193 = ~n23191 & ~n23192 ;
  assign n23194 = n23193 ^ n20715 ;
  assign n23221 = n23202 ^ n23194 ;
  assign n23222 = n23203 & ~n23221 ;
  assign n23223 = n23222 ^ n20835 ;
  assign n23217 = n22797 ^ n22766 ;
  assign n23215 = n21949 ^ n21347 ;
  assign n23216 = n23215 ^ n22431 ;
  assign n23218 = n23217 ^ n23216 ;
  assign n23212 = n23201 ^ n23197 ;
  assign n23213 = n23199 & ~n23212 ;
  assign n23214 = n23213 ^ n23197 ;
  assign n23219 = n23218 ^ n23214 ;
  assign n23229 = n23223 ^ n23219 ;
  assign n23235 = n21957 ^ n21357 ;
  assign n23236 = n23235 ^ n22433 ;
  assign n23232 = n22800 ^ n22764 ;
  assign n23233 = n23232 ^ n23217 ;
  assign n23230 = n23217 ^ n23214 ;
  assign n23231 = n23218 & n23230 ;
  assign n23234 = n23233 ^ n23231 ;
  assign n23237 = n23236 ^ n23234 ;
  assign n23238 = n23237 ^ n20856 ;
  assign n23239 = n23238 ^ n23237 ;
  assign n23240 = n23239 ^ n23223 ;
  assign n23241 = n23229 & ~n23240 ;
  assign n23242 = n23241 ^ n23238 ;
  assign n23394 = n23237 ^ n20877 ;
  assign n23395 = n23242 & ~n23394 ;
  assign n23396 = n23395 ^ n20877 ;
  assign n23443 = n23396 ^ n20901 ;
  assign n23298 = n22803 ^ n22762 ;
  assign n23361 = n23298 ^ n23236 ;
  assign n23359 = n23236 ^ n23232 ;
  assign n23360 = n23234 & ~n23359 ;
  assign n23362 = n23361 ^ n23360 ;
  assign n23356 = n21965 ^ n21365 ;
  assign n23357 = n23356 ^ n22539 ;
  assign n23397 = n23362 ^ n23357 ;
  assign n23444 = n23443 ^ n23397 ;
  assign n23243 = n23242 ^ n20877 ;
  assign n23220 = n23219 ^ n20856 ;
  assign n23224 = n23223 ^ n23220 ;
  assign n23204 = n23203 ^ n23194 ;
  assign n23178 = n23177 ^ n20715 ;
  assign n23182 = n23181 ^ n23178 ;
  assign n23023 = n23022 ^ n20667 ;
  assign n23024 = n22983 ^ n22980 ;
  assign n23025 = n22975 ^ n22972 ;
  assign n23026 = n22930 ^ n20441 ;
  assign n23027 = n23026 ^ n22968 ;
  assign n23028 = n22965 ^ n22932 ;
  assign n23029 = n22934 ^ n20453 ;
  assign n23030 = n23029 ^ n22961 ;
  assign n23031 = n22942 ^ n20423 ;
  assign n23032 = n22943 ^ n20472 ;
  assign n23033 = n23032 ^ n22944 ;
  assign n23034 = n23031 & ~n23033 ;
  assign n23035 = n22948 ^ n22941 ;
  assign n23036 = n23034 & ~n23035 ;
  assign n23037 = n22939 ^ n20468 ;
  assign n23038 = n23037 ^ n22951 ;
  assign n23039 = n23036 & ~n23038 ;
  assign n23040 = n22955 ^ n22938 ;
  assign n23041 = n23039 & ~n23040 ;
  assign n23042 = n22958 ^ n22936 ;
  assign n23043 = ~n23041 & ~n23042 ;
  assign n23044 = n23030 & ~n23043 ;
  assign n23045 = n23028 & ~n23044 ;
  assign n23046 = ~n23027 & n23045 ;
  assign n23047 = ~n23025 & n23046 ;
  assign n23048 = n22977 ^ n22929 ;
  assign n23049 = ~n23047 & ~n23048 ;
  assign n23050 = n23024 & ~n23049 ;
  assign n23051 = n22927 ^ n20492 ;
  assign n23052 = n23051 ^ n22985 ;
  assign n23053 = ~n23050 & ~n23052 ;
  assign n23054 = n22991 ^ n20486 ;
  assign n23055 = ~n23053 & ~n23054 ;
  assign n23056 = n22993 ^ n22924 ;
  assign n23057 = n23055 & n23056 ;
  assign n23058 = n22922 ^ n20475 ;
  assign n23059 = n23058 ^ n22996 ;
  assign n23060 = n23057 & ~n23059 ;
  assign n23061 = n23008 ^ n20479 ;
  assign n23062 = n23061 ^ n23000 ;
  assign n23063 = n23060 & ~n23062 ;
  assign n23183 = n23023 & ~n23063 ;
  assign n23205 = n23182 & n23183 ;
  assign n23225 = ~n23204 & ~n23205 ;
  assign n23244 = ~n23224 & n23225 ;
  assign n23442 = n23243 & ~n23244 ;
  assign n23476 = n23444 ^ n23442 ;
  assign n23477 = n23476 ^ n1360 ;
  assign n23245 = n23244 ^ n23243 ;
  assign n1199 = n1098 ^ n1046 ;
  assign n1200 = n1199 ^ n980 ;
  assign n1204 = n1203 ^ n1200 ;
  assign n23246 = n23245 ^ n1204 ;
  assign n23184 = n23183 ^ n23182 ;
  assign n23064 = n23063 ^ n23023 ;
  assign n1662 = n1644 ^ n1013 ;
  assign n1663 = n1662 ^ n742 ;
  assign n1664 = n1663 ^ n833 ;
  assign n23065 = n23064 ^ n1664 ;
  assign n23066 = n23062 ^ n23060 ;
  assign n23067 = n23066 ^ n738 ;
  assign n23068 = n23059 ^ n23057 ;
  assign n23069 = n23068 ^ n679 ;
  assign n23148 = n23056 ^ n23055 ;
  assign n23159 = n23148 ^ n23068 ;
  assign n23145 = n23054 ^ n23053 ;
  assign n23146 = n23145 ^ n1512 ;
  assign n23141 = n23052 ^ n23050 ;
  assign n23073 = n23049 ^ n23024 ;
  assign n23074 = n23073 ^ n23072 ;
  assign n23129 = n23048 ^ n23047 ;
  assign n23075 = n23046 ^ n23025 ;
  assign n2910 = n2906 ^ n2363 ;
  assign n2911 = n2910 ^ n587 ;
  assign n2915 = n2914 ^ n2911 ;
  assign n23076 = n23075 ^ n2915 ;
  assign n23077 = n23045 ^ n23027 ;
  assign n23081 = n23080 ^ n23077 ;
  assign n23082 = n23044 ^ n23028 ;
  assign n2287 = n2286 ^ n2211 ;
  assign n2288 = n2287 ^ n581 ;
  assign n2292 = n2291 ^ n2288 ;
  assign n23083 = n23082 ^ n2292 ;
  assign n23084 = n23043 ^ n23030 ;
  assign n2162 = n2146 ^ n2095 ;
  assign n2163 = n2162 ^ n2159 ;
  assign n2164 = n2163 ^ n1457 ;
  assign n23085 = n23084 ^ n2164 ;
  assign n23086 = n23040 ^ n23039 ;
  assign n2058 = n2030 ^ n2006 ;
  assign n2059 = n2058 ^ n2055 ;
  assign n2063 = n2062 ^ n2059 ;
  assign n23087 = n23086 ^ n2063 ;
  assign n23091 = n23038 ^ n23036 ;
  assign n2049 = n1997 ^ n1968 ;
  assign n2050 = n2049 ^ n2048 ;
  assign n2051 = n2050 ^ n2042 ;
  assign n23092 = n23091 ^ n2051 ;
  assign n23094 = n21195 ^ n1956 ;
  assign n23095 = n23094 ^ n3087 ;
  assign n23096 = n23095 ^ n2046 ;
  assign n23093 = n23035 ^ n23034 ;
  assign n23097 = n23096 ^ n23093 ;
  assign n3072 = n3021 ^ n2781 ;
  assign n3073 = n3072 ^ n1787 ;
  assign n3074 = n3073 ^ n3068 ;
  assign n23098 = n3074 & ~n23031 ;
  assign n3078 = n3044 ^ n1949 ;
  assign n3079 = n3078 ^ n3070 ;
  assign n3080 = n3079 ^ n1871 ;
  assign n23099 = n23098 ^ n3080 ;
  assign n23100 = n23033 ^ n23031 ;
  assign n23101 = n23100 ^ n3080 ;
  assign n23102 = n23099 & n23101 ;
  assign n23103 = n23102 ^ n23098 ;
  assign n23104 = n23103 ^ n23093 ;
  assign n23105 = ~n23097 & n23104 ;
  assign n23106 = n23105 ^ n23096 ;
  assign n23107 = n23106 ^ n2051 ;
  assign n23108 = ~n23092 & n23107 ;
  assign n23109 = n23108 ^ n2051 ;
  assign n23088 = n23042 ^ n23041 ;
  assign n23089 = n23088 ^ n2063 ;
  assign n23090 = n23089 ^ n23088 ;
  assign n23110 = n23109 ^ n23090 ;
  assign n23111 = ~n23087 & n23110 ;
  assign n23112 = n23111 ^ n23089 ;
  assign n2150 = n2140 ^ n2086 ;
  assign n2151 = n2150 ^ n2070 ;
  assign n2155 = n2154 ^ n2151 ;
  assign n23114 = n23084 ^ n2155 ;
  assign n23113 = n23088 ^ n23084 ;
  assign n23115 = n23114 ^ n23113 ;
  assign n23116 = ~n23112 & ~n23115 ;
  assign n23117 = n23116 ^ n23113 ;
  assign n23118 = ~n23085 & n23117 ;
  assign n23119 = n23118 ^ n23084 ;
  assign n23120 = n23119 ^ n2292 ;
  assign n23121 = n23083 & ~n23120 ;
  assign n23122 = n23121 ^ n2292 ;
  assign n23123 = n23122 ^ n23077 ;
  assign n23124 = n23081 & ~n23123 ;
  assign n23125 = n23124 ^ n23080 ;
  assign n23126 = n23125 ^ n23075 ;
  assign n23127 = n23076 & ~n23126 ;
  assign n23128 = n23127 ^ n2915 ;
  assign n23130 = n23129 ^ n23128 ;
  assign n23136 = n23133 ^ n23128 ;
  assign n23137 = ~n23130 & n23136 ;
  assign n23134 = n23133 ^ n23072 ;
  assign n23138 = n23137 ^ n23134 ;
  assign n23139 = n23074 & ~n23138 ;
  assign n23140 = n23139 ^ n23073 ;
  assign n23142 = n23141 ^ n23140 ;
  assign n23143 = n23140 ^ n1512 ;
  assign n23144 = ~n23142 & n23143 ;
  assign n23147 = n23146 ^ n23144 ;
  assign n23149 = n23148 ^ n23145 ;
  assign n23150 = n23149 ^ n23148 ;
  assign n23154 = n23153 ^ n23150 ;
  assign n23155 = ~n23147 & ~n23154 ;
  assign n23156 = n23155 ^ n23149 ;
  assign n23157 = n23148 ^ n667 ;
  assign n23158 = n23156 & ~n23157 ;
  assign n23160 = n23159 ^ n23158 ;
  assign n23161 = n23069 & ~n23160 ;
  assign n23162 = n23161 ^ n23068 ;
  assign n23163 = n23162 ^ n738 ;
  assign n23164 = n23067 & ~n23163 ;
  assign n23165 = n23164 ^ n23066 ;
  assign n23166 = n23165 ^ n1664 ;
  assign n23167 = ~n23065 & ~n23166 ;
  assign n23168 = n23167 ^ n23064 ;
  assign n23185 = n23184 ^ n23168 ;
  assign n840 = n839 ^ n776 ;
  assign n841 = n840 ^ n836 ;
  assign n842 = n841 ^ n830 ;
  assign n23188 = n23168 ^ n842 ;
  assign n23189 = n23185 & ~n23188 ;
  assign n1190 = n1112 ^ n1028 ;
  assign n1194 = n1193 ^ n1190 ;
  assign n1195 = n1194 ^ n974 ;
  assign n23186 = n1195 ^ n842 ;
  assign n23190 = n23189 ^ n23186 ;
  assign n23208 = n1204 ^ n1195 ;
  assign n23206 = n23205 ^ n23204 ;
  assign n23207 = n23206 ^ n1204 ;
  assign n23209 = n23208 ^ n23207 ;
  assign n23210 = n23190 & ~n23209 ;
  assign n23211 = n23210 ^ n23208 ;
  assign n23226 = n23225 ^ n23224 ;
  assign n23227 = n23226 ^ n1204 ;
  assign n23228 = n23211 & n23227 ;
  assign n23247 = n23246 ^ n23228 ;
  assign n23478 = n23245 ^ n1219 ;
  assign n23479 = ~n23247 & ~n23478 ;
  assign n23480 = n23479 ^ n23245 ;
  assign n23481 = n23480 ^ n1360 ;
  assign n23482 = ~n23477 & n23481 ;
  assign n23483 = n23482 ^ n23476 ;
  assign n23398 = n23397 ^ n23396 ;
  assign n23399 = n23397 ^ n20901 ;
  assign n23400 = n23398 & ~n23399 ;
  assign n23401 = n23400 ^ n20901 ;
  assign n23358 = n23357 ^ n23298 ;
  assign n23363 = ~n23358 & ~n23362 ;
  assign n23364 = n23363 ^ n23298 ;
  assign n23353 = n22053 ^ n21372 ;
  assign n23354 = n23353 ^ n22547 ;
  assign n23294 = n22806 ^ n22760 ;
  assign n23355 = n23354 ^ n23294 ;
  assign n23392 = n23364 ^ n23355 ;
  assign n23393 = n23392 ^ n20921 ;
  assign n23446 = n23401 ^ n23393 ;
  assign n23445 = ~n23442 & ~n23444 ;
  assign n23474 = n23446 ^ n23445 ;
  assign n23475 = n23474 ^ n1396 ;
  assign n24022 = n23483 ^ n23475 ;
  assign n24020 = n22222 ^ n21578 ;
  assign n24021 = n24020 ^ n22872 ;
  assign n24023 = n24022 ^ n24021 ;
  assign n23648 = n22213 ^ n21583 ;
  assign n23649 = n23648 ^ n22866 ;
  assign n23647 = n23480 ^ n23477 ;
  assign n23650 = n23649 ^ n23647 ;
  assign n23250 = n22832 ^ n3101 ;
  assign n23249 = n22216 ^ n21594 ;
  assign n23251 = n23250 ^ n23249 ;
  assign n23248 = n23247 ^ n1219 ;
  assign n23252 = n23251 ^ n23248 ;
  assign n23256 = n23226 ^ n23211 ;
  assign n23643 = n23256 ^ n23251 ;
  assign n23254 = n22829 ^ n22742 ;
  assign n23253 = n22210 ^ n21591 ;
  assign n23255 = n23254 ^ n23253 ;
  assign n23257 = n23256 ^ n23255 ;
  assign n23261 = n23206 ^ n23190 ;
  assign n23640 = n23261 ^ n23256 ;
  assign n23259 = n22826 ^ n22749 ;
  assign n23258 = n22421 ^ n22196 ;
  assign n23260 = n23259 ^ n23258 ;
  assign n23262 = n23261 ^ n23260 ;
  assign n23266 = n23185 ^ n842 ;
  assign n23264 = n22824 ^ n2639 ;
  assign n23263 = n22563 ^ n22053 ;
  assign n23265 = n23264 ^ n23263 ;
  assign n23267 = n23266 ^ n23265 ;
  assign n23272 = n23165 ^ n23065 ;
  assign n23634 = n23272 ^ n23266 ;
  assign n23269 = n22752 ^ n1241 ;
  assign n23270 = n23269 ^ n22818 ;
  assign n23268 = n22555 ^ n21965 ;
  assign n23271 = n23270 ^ n23268 ;
  assign n23273 = n23272 ^ n23271 ;
  assign n23277 = n23162 ^ n23067 ;
  assign n23275 = n22816 ^ n1247 ;
  assign n23274 = n22547 ^ n21957 ;
  assign n23276 = n23275 ^ n23274 ;
  assign n23278 = n23277 ^ n23276 ;
  assign n23284 = n23160 ^ n679 ;
  assign n23282 = n22812 ^ n22756 ;
  assign n23281 = n22539 ^ n21949 ;
  assign n23283 = n23282 ^ n23281 ;
  assign n23285 = n23284 ^ n23283 ;
  assign n23289 = n23156 ^ n667 ;
  assign n23287 = n22810 ^ n963 ;
  assign n23286 = n22433 ^ n21940 ;
  assign n23288 = n23287 ^ n23286 ;
  assign n23290 = n23289 ^ n23288 ;
  assign n23293 = n22431 ^ n21932 ;
  assign n23295 = n23294 ^ n23293 ;
  assign n23291 = n23153 ^ n23147 ;
  assign n23296 = n23295 ^ n23291 ;
  assign n23300 = n23142 ^ n1512 ;
  assign n23297 = n22436 ^ n21922 ;
  assign n23299 = n23298 ^ n23297 ;
  assign n23301 = n23300 ^ n23299 ;
  assign n23304 = n23138 ^ n23073 ;
  assign n23302 = n22440 ^ n21865 ;
  assign n23303 = n23302 ^ n23232 ;
  assign n23305 = n23304 ^ n23303 ;
  assign n23607 = n22444 ^ n21863 ;
  assign n23608 = n23607 ^ n23217 ;
  assign n23308 = n23125 ^ n23076 ;
  assign n23306 = n22448 ^ n21255 ;
  assign n23307 = n23306 ^ n23197 ;
  assign n23309 = n23308 ^ n23307 ;
  assign n23312 = n23122 ^ n23081 ;
  assign n23310 = n22452 ^ n21873 ;
  assign n23311 = n23310 ^ n23169 ;
  assign n23313 = n23312 ^ n23311 ;
  assign n23576 = n23112 ^ n2155 ;
  assign n23314 = n23109 ^ n23087 ;
  assign n23577 = n23576 ^ n23314 ;
  assign n23315 = n22388 ^ n21891 ;
  assign n23316 = n23315 ^ n22374 ;
  assign n23317 = n23316 ^ n23314 ;
  assign n23320 = n23106 ^ n23092 ;
  assign n23318 = n22393 ^ n21893 ;
  assign n23319 = n23318 ^ n22376 ;
  assign n23321 = n23320 ^ n23319 ;
  assign n23323 = n22398 ^ n21753 ;
  assign n23324 = n23323 ^ n22385 ;
  assign n23322 = n23103 ^ n23097 ;
  assign n23325 = n23324 ^ n23322 ;
  assign n23328 = n23100 ^ n23099 ;
  assign n23326 = n22404 ^ n21736 ;
  assign n23327 = n23326 ^ n22390 ;
  assign n23329 = n23328 ^ n23327 ;
  assign n23332 = n23031 ^ n3074 ;
  assign n23564 = n23332 ^ n23327 ;
  assign n23330 = n22408 ^ n21636 ;
  assign n23331 = n23330 ^ n22395 ;
  assign n23333 = n23332 ^ n23331 ;
  assign n23526 = n3009 ^ n2765 ;
  assign n23527 = n23526 ^ n3176 ;
  assign n23528 = n23527 ^ n1785 ;
  assign n23529 = n23528 ^ n1844 ;
  assign n23522 = n20374 ^ n20357 ;
  assign n23518 = n21610 ^ n20465 ;
  assign n23432 = n21271 ^ n20467 ;
  assign n23433 = n23432 ^ n22222 ;
  assign n23519 = n23518 ^ n23433 ;
  assign n23520 = n23519 ^ n22202 ;
  assign n23521 = n23520 ^ n23250 ;
  assign n23523 = n23522 ^ n23521 ;
  assign n23434 = n23433 ^ n23254 ;
  assign n23336 = n21578 ^ n20941 ;
  assign n23337 = n23336 ^ n22216 ;
  assign n23338 = n23337 ^ n23264 ;
  assign n23341 = n21583 ^ n20950 ;
  assign n23342 = n23341 ^ n22210 ;
  assign n23343 = n23342 ^ n23270 ;
  assign n23344 = n21594 ^ n20952 ;
  assign n23345 = n23344 ^ n22421 ;
  assign n23346 = n23345 ^ n23275 ;
  assign n23347 = n21591 ^ n20947 ;
  assign n23348 = n23347 ^ n22563 ;
  assign n23349 = n23348 ^ n23282 ;
  assign n23350 = n22196 ^ n21485 ;
  assign n23351 = n23350 ^ n22555 ;
  assign n23352 = n23351 ^ n23287 ;
  assign n23365 = n23364 ^ n23294 ;
  assign n23366 = n23355 & n23365 ;
  assign n23367 = n23366 ^ n23294 ;
  assign n23368 = n23367 ^ n23351 ;
  assign n23369 = ~n23352 & n23368 ;
  assign n23370 = n23369 ^ n23287 ;
  assign n23371 = n23370 ^ n23348 ;
  assign n23372 = n23349 & n23371 ;
  assign n23373 = n23372 ^ n23282 ;
  assign n23374 = n23373 ^ n23345 ;
  assign n23375 = n23346 & n23374 ;
  assign n23376 = n23375 ^ n23275 ;
  assign n23377 = n23376 ^ n23342 ;
  assign n23378 = n23343 & n23377 ;
  assign n23379 = n23378 ^ n23270 ;
  assign n23380 = n23379 ^ n23264 ;
  assign n23381 = n23338 & n23380 ;
  assign n23339 = n23264 ^ n23259 ;
  assign n23382 = n23381 ^ n23339 ;
  assign n23383 = n21576 ^ n20988 ;
  assign n23384 = n23383 ^ n22213 ;
  assign n23429 = n23384 ^ n23259 ;
  assign n23430 = n23382 & n23429 ;
  assign n23431 = n23430 ^ n23259 ;
  assign n23516 = n23433 ^ n23431 ;
  assign n23517 = ~n23434 & ~n23516 ;
  assign n23524 = n23523 ^ n23517 ;
  assign n23385 = n23384 ^ n23382 ;
  assign n23438 = n23385 ^ n20342 ;
  assign n23386 = n23379 ^ n23338 ;
  assign n23387 = n23386 ^ n20292 ;
  assign n23416 = n23376 ^ n23343 ;
  assign n23388 = n23373 ^ n23346 ;
  assign n23389 = n23388 ^ n20263 ;
  assign n23390 = n23370 ^ n23349 ;
  assign n23391 = n23390 ^ n20258 ;
  assign n23402 = n23401 ^ n23392 ;
  assign n23403 = n23393 & n23402 ;
  assign n23404 = n23403 ^ n20921 ;
  assign n23405 = n23404 ^ n20977 ;
  assign n23406 = n23367 ^ n23352 ;
  assign n23407 = n23406 ^ n23404 ;
  assign n23408 = ~n23405 & n23407 ;
  assign n23409 = n23408 ^ n20977 ;
  assign n23410 = n23409 ^ n23390 ;
  assign n23411 = ~n23391 & n23410 ;
  assign n23412 = n23411 ^ n20258 ;
  assign n23413 = n23412 ^ n23388 ;
  assign n23414 = n23389 & ~n23413 ;
  assign n23415 = n23414 ^ n20263 ;
  assign n23417 = n23416 ^ n23415 ;
  assign n23418 = n23386 ^ n20253 ;
  assign n23419 = n23418 ^ n23386 ;
  assign n23420 = n23419 ^ n23415 ;
  assign n23421 = n23417 & n23420 ;
  assign n23422 = n23421 ^ n23418 ;
  assign n23423 = n23387 & ~n23422 ;
  assign n23424 = n23423 ^ n20292 ;
  assign n23439 = n23438 ^ n23424 ;
  assign n23440 = n23422 ^ n20292 ;
  assign n23441 = n23412 ^ n23389 ;
  assign n23447 = n23445 & n23446 ;
  assign n23448 = n23406 ^ n23405 ;
  assign n23449 = ~n23447 & n23448 ;
  assign n23450 = n23409 ^ n23391 ;
  assign n23451 = ~n23449 & ~n23450 ;
  assign n23452 = n23441 & n23451 ;
  assign n23453 = n23415 ^ n20253 ;
  assign n23454 = n23453 ^ n23416 ;
  assign n23455 = n23452 & ~n23454 ;
  assign n23456 = ~n23440 & ~n23455 ;
  assign n23457 = n23439 & ~n23456 ;
  assign n23435 = n23434 ^ n23431 ;
  assign n23509 = n23457 ^ n23435 ;
  assign n23425 = n23424 ^ n23385 ;
  assign n23426 = n23424 ^ n20342 ;
  assign n23427 = ~n23425 & n23426 ;
  assign n23428 = n23427 ^ n20342 ;
  assign n23511 = n23435 ^ n23428 ;
  assign n23514 = n23509 & n23511 ;
  assign n23512 = n23511 ^ n23457 ;
  assign n23513 = ~n20357 & n23512 ;
  assign n23515 = n23514 ^ n23513 ;
  assign n23525 = n23524 ^ n23515 ;
  assign n23530 = n23529 ^ n23525 ;
  assign n23436 = n23435 ^ n20357 ;
  assign n23437 = n23436 ^ n23428 ;
  assign n23458 = n23457 ^ n23437 ;
  assign n23459 = n23458 ^ n1844 ;
  assign n23460 = n23456 ^ n23439 ;
  assign n3155 = n3142 ^ n2711 ;
  assign n3156 = n3155 ^ n2468 ;
  assign n3157 = n3156 ^ n1805 ;
  assign n23461 = n23460 ^ n3157 ;
  assign n23462 = n23455 ^ n23440 ;
  assign n23463 = n23462 ^ n3150 ;
  assign n23465 = n23451 ^ n23441 ;
  assign n23466 = n23465 ^ n3212 ;
  assign n23467 = n23450 ^ n23449 ;
  assign n2547 = n2546 ^ n2478 ;
  assign n2554 = n2553 ^ n2547 ;
  assign n2558 = n2557 ^ n2554 ;
  assign n23468 = n23467 ^ n2558 ;
  assign n23469 = n23448 ^ n23447 ;
  assign n23473 = n23472 ^ n23469 ;
  assign n23484 = n23483 ^ n23474 ;
  assign n23485 = ~n23475 & ~n23484 ;
  assign n23486 = n23485 ^ n1396 ;
  assign n23487 = n23486 ^ n23469 ;
  assign n23488 = ~n23473 & n23487 ;
  assign n23489 = n23488 ^ n23472 ;
  assign n23490 = n23489 ^ n23467 ;
  assign n23491 = ~n23468 & n23490 ;
  assign n23492 = n23491 ^ n2558 ;
  assign n23493 = n23492 ^ n23465 ;
  assign n23494 = ~n23466 & n23493 ;
  assign n23495 = n23494 ^ n3212 ;
  assign n23464 = n23454 ^ n23452 ;
  assign n23496 = n23495 ^ n23464 ;
  assign n23497 = n23462 ^ n2516 ;
  assign n23498 = n23497 ^ n23462 ;
  assign n23499 = n23498 ^ n23464 ;
  assign n23500 = ~n23496 & n23499 ;
  assign n23501 = n23500 ^ n23497 ;
  assign n23502 = n23463 & ~n23501 ;
  assign n23503 = n23502 ^ n3150 ;
  assign n23504 = n23503 ^ n23460 ;
  assign n23505 = n23461 & ~n23504 ;
  assign n23506 = n23505 ^ n3157 ;
  assign n23507 = n23506 ^ n1844 ;
  assign n23508 = n23459 & n23507 ;
  assign n23531 = n23530 ^ n23508 ;
  assign n23334 = n22482 ^ n21628 ;
  assign n23335 = n23334 ^ n22397 ;
  assign n23532 = n23531 ^ n23335 ;
  assign n23533 = n23506 ^ n23459 ;
  assign n23558 = n23533 ^ n23335 ;
  assign n23534 = n22413 ^ n21622 ;
  assign n23535 = n23534 ^ n22402 ;
  assign n23536 = n23535 ^ n23533 ;
  assign n23538 = n22353 ^ n21262 ;
  assign n23539 = n23538 ^ n22410 ;
  assign n23537 = n23503 ^ n23461 ;
  assign n23540 = n23539 ^ n23537 ;
  assign n23544 = n22273 ^ n21265 ;
  assign n23545 = n23544 ^ n22412 ;
  assign n23546 = n23464 ^ n2516 ;
  assign n23547 = n23546 ^ n23495 ;
  assign n23548 = ~n23545 & n23547 ;
  assign n23541 = n22301 ^ n21260 ;
  assign n23542 = n23541 ^ n22887 ;
  assign n23549 = n23548 ^ n23542 ;
  assign n23550 = n23501 ^ n3150 ;
  assign n23551 = n23550 ^ n23542 ;
  assign n23552 = n23549 & n23551 ;
  assign n23543 = n23542 ^ n23539 ;
  assign n23553 = n23552 ^ n23543 ;
  assign n23554 = n23540 & n23553 ;
  assign n23555 = n23554 ^ n23539 ;
  assign n23556 = n23555 ^ n23533 ;
  assign n23557 = n23536 & n23556 ;
  assign n23559 = n23558 ^ n23557 ;
  assign n23560 = n23532 & ~n23559 ;
  assign n23561 = n23560 ^ n23531 ;
  assign n23562 = n23561 ^ n23332 ;
  assign n23563 = n23333 & ~n23562 ;
  assign n23565 = n23564 ^ n23563 ;
  assign n23566 = n23329 & ~n23565 ;
  assign n23567 = n23566 ^ n23328 ;
  assign n23568 = n23567 ^ n23322 ;
  assign n23569 = n23325 & ~n23568 ;
  assign n23570 = n23569 ^ n23324 ;
  assign n23571 = n23570 ^ n23319 ;
  assign n23572 = n23321 & ~n23571 ;
  assign n23573 = n23572 ^ n23320 ;
  assign n23574 = n23573 ^ n23314 ;
  assign n23575 = ~n23317 & n23574 ;
  assign n23578 = n23577 ^ n23575 ;
  assign n23582 = n22383 ^ n21884 ;
  assign n23583 = n23582 ^ n22918 ;
  assign n23579 = n23117 ^ n2164 ;
  assign n23580 = n23579 ^ n23576 ;
  assign n23581 = n23580 ^ n23579 ;
  assign n23584 = n23583 ^ n23581 ;
  assign n23585 = n23578 & ~n23584 ;
  assign n23586 = n23585 ^ n23580 ;
  assign n23587 = n21875 ^ n21851 ;
  assign n23588 = n23587 ^ n23015 ;
  assign n23592 = n23588 ^ n23579 ;
  assign n23589 = n22379 ^ n21882 ;
  assign n23590 = n23589 ^ n23003 ;
  assign n23591 = n23590 ^ n23588 ;
  assign n23593 = n23592 ^ n23591 ;
  assign n23594 = n23586 & ~n23593 ;
  assign n23595 = n23594 ^ n23591 ;
  assign n23597 = n23119 ^ n23083 ;
  assign n23598 = n23597 ^ n23312 ;
  assign n23596 = n23588 ^ n23312 ;
  assign n23599 = n23598 ^ n23596 ;
  assign n23600 = ~n23595 & ~n23599 ;
  assign n23601 = n23600 ^ n23596 ;
  assign n23602 = ~n23313 & n23601 ;
  assign n23603 = n23602 ^ n23312 ;
  assign n23604 = n23603 ^ n23307 ;
  assign n23605 = ~n23309 & n23604 ;
  assign n23606 = n23605 ^ n23308 ;
  assign n23609 = n23608 ^ n23606 ;
  assign n23610 = n23133 ^ n23129 ;
  assign n23611 = n23610 ^ n23128 ;
  assign n23614 = n23611 ^ n23606 ;
  assign n23615 = n23609 & n23614 ;
  assign n23612 = n23611 ^ n23303 ;
  assign n23616 = n23615 ^ n23612 ;
  assign n23617 = ~n23305 & n23616 ;
  assign n23618 = n23617 ^ n23304 ;
  assign n23619 = n23618 ^ n23300 ;
  assign n23620 = n23301 & n23619 ;
  assign n23621 = n23620 ^ n23300 ;
  assign n23622 = n23621 ^ n23291 ;
  assign n23623 = ~n23296 & ~n23622 ;
  assign n23292 = n23291 ^ n23289 ;
  assign n23624 = n23623 ^ n23292 ;
  assign n23625 = ~n23290 & ~n23624 ;
  assign n23626 = n23625 ^ n23289 ;
  assign n23627 = n23626 ^ n23283 ;
  assign n23628 = ~n23285 & ~n23627 ;
  assign n23629 = n23628 ^ n23284 ;
  assign n23630 = n23629 ^ n23277 ;
  assign n23631 = ~n23278 & ~n23630 ;
  assign n23279 = n23277 ^ n23271 ;
  assign n23632 = n23631 ^ n23279 ;
  assign n23633 = ~n23273 & ~n23632 ;
  assign n23635 = n23634 ^ n23633 ;
  assign n23636 = ~n23267 & n23635 ;
  assign n23637 = n23636 ^ n23266 ;
  assign n23638 = n23637 ^ n23261 ;
  assign n23639 = ~n23262 & n23638 ;
  assign n23641 = n23640 ^ n23639 ;
  assign n23642 = ~n23257 & ~n23641 ;
  assign n23644 = n23643 ^ n23642 ;
  assign n23645 = n23252 & ~n23644 ;
  assign n23646 = n23645 ^ n23251 ;
  assign n24017 = n23647 ^ n23646 ;
  assign n24018 = n23650 & ~n24017 ;
  assign n24019 = n24018 ^ n23647 ;
  assign n24024 = n24023 ^ n24019 ;
  assign n24025 = n24024 ^ n20941 ;
  assign n23653 = n23644 ^ n23248 ;
  assign n23654 = n23653 ^ n20952 ;
  assign n23780 = n23641 ^ n23255 ;
  assign n23655 = n23637 ^ n23262 ;
  assign n23656 = n23655 ^ n21485 ;
  assign n23657 = n23635 ^ n23265 ;
  assign n23658 = n23657 ^ n21372 ;
  assign n23659 = n23632 ^ n23272 ;
  assign n23660 = n23659 ^ n21365 ;
  assign n23661 = n23629 ^ n23278 ;
  assign n23662 = n23661 ^ n21357 ;
  assign n23663 = n23626 ^ n23285 ;
  assign n23664 = n23663 ^ n21347 ;
  assign n23665 = n23624 ^ n23288 ;
  assign n23666 = n23665 ^ n21282 ;
  assign n23667 = n23621 ^ n23296 ;
  assign n23668 = n23667 ^ n21278 ;
  assign n23753 = n23618 ^ n23301 ;
  assign n23669 = n23616 ^ n23304 ;
  assign n23670 = n23669 ^ n21289 ;
  assign n23744 = n23611 ^ n23608 ;
  assign n23745 = n23744 ^ n23606 ;
  assign n23671 = n23603 ^ n23309 ;
  assign n23672 = n23671 ^ n21256 ;
  assign n23673 = n23590 ^ n23586 ;
  assign n23674 = n23673 ^ n21308 ;
  assign n23675 = n23583 ^ n23578 ;
  assign n23676 = n23675 ^ n21314 ;
  assign n23678 = n23570 ^ n23321 ;
  assign n23679 = n23678 ^ n21133 ;
  assign n23681 = n23565 ^ n23328 ;
  assign n23682 = n23681 ^ n21015 ;
  assign n23683 = n23559 ^ n23531 ;
  assign n23684 = n23683 ^ n20438 ;
  assign n23686 = n23553 ^ n23537 ;
  assign n23687 = n23686 ^ n20450 ;
  assign n23688 = n23547 ^ n23545 ;
  assign n23689 = ~n20457 & ~n23688 ;
  assign n23690 = n23689 ^ n20452 ;
  assign n23691 = n23550 ^ n23549 ;
  assign n23692 = n23691 ^ n23689 ;
  assign n23693 = n23690 & ~n23692 ;
  assign n23694 = n23693 ^ n20452 ;
  assign n23695 = n23694 ^ n23686 ;
  assign n23696 = ~n23687 & ~n23695 ;
  assign n23697 = n23696 ^ n20450 ;
  assign n23685 = n23555 ^ n23536 ;
  assign n23698 = n23697 ^ n23685 ;
  assign n23699 = n23697 ^ n20443 ;
  assign n23700 = n23698 & ~n23699 ;
  assign n23701 = n23700 ^ n20443 ;
  assign n23702 = n23701 ^ n23683 ;
  assign n23703 = ~n23684 & ~n23702 ;
  assign n23704 = n23703 ^ n20438 ;
  assign n23705 = n23704 ^ n20433 ;
  assign n23706 = n23561 ^ n23333 ;
  assign n23707 = n23706 ^ n23704 ;
  assign n23708 = ~n23705 & n23707 ;
  assign n23709 = n23708 ^ n20433 ;
  assign n23710 = n23709 ^ n23681 ;
  assign n23711 = ~n23682 & n23710 ;
  assign n23712 = n23711 ^ n21015 ;
  assign n23680 = n23567 ^ n23325 ;
  assign n23713 = n23712 ^ n23680 ;
  assign n23714 = n23712 ^ n21125 ;
  assign n23715 = n23713 & n23714 ;
  assign n23716 = n23715 ^ n21125 ;
  assign n23717 = n23716 ^ n23678 ;
  assign n23718 = n23679 & n23717 ;
  assign n23719 = n23718 ^ n21133 ;
  assign n23677 = n23573 ^ n23317 ;
  assign n23720 = n23719 ^ n23677 ;
  assign n23721 = n23675 ^ n21248 ;
  assign n23722 = n23721 ^ n23675 ;
  assign n23723 = n23722 ^ n23677 ;
  assign n23724 = n23720 & n23723 ;
  assign n23725 = n23724 ^ n23721 ;
  assign n23726 = ~n23676 & ~n23725 ;
  assign n23727 = n23726 ^ n21314 ;
  assign n23728 = n23727 ^ n23673 ;
  assign n23729 = n23674 & n23728 ;
  assign n23730 = n23729 ^ n21308 ;
  assign n23731 = n23730 ^ n21306 ;
  assign n23732 = n23597 ^ n23595 ;
  assign n23733 = n23732 ^ n23730 ;
  assign n23734 = ~n23731 & ~n23733 ;
  assign n23735 = n23734 ^ n21306 ;
  assign n23736 = n23735 ^ n21300 ;
  assign n23737 = n23601 ^ n23311 ;
  assign n23738 = n23737 ^ n23735 ;
  assign n23739 = n23736 & ~n23738 ;
  assign n23740 = n23739 ^ n21300 ;
  assign n23741 = n23740 ^ n23671 ;
  assign n23742 = ~n23672 & ~n23741 ;
  assign n23743 = n23742 ^ n21256 ;
  assign n23746 = n23745 ^ n23743 ;
  assign n23747 = n23745 ^ n21295 ;
  assign n23748 = n23746 & ~n23747 ;
  assign n23749 = n23748 ^ n21295 ;
  assign n23750 = n23749 ^ n23669 ;
  assign n23751 = n23670 & n23750 ;
  assign n23752 = n23751 ^ n21289 ;
  assign n23754 = n23753 ^ n23752 ;
  assign n23755 = n23667 ^ n21285 ;
  assign n23756 = n23755 ^ n23667 ;
  assign n23757 = n23756 ^ n23752 ;
  assign n23758 = n23754 & n23757 ;
  assign n23759 = n23758 ^ n23755 ;
  assign n23760 = n23668 & ~n23759 ;
  assign n23761 = n23760 ^ n21278 ;
  assign n23762 = n23761 ^ n23665 ;
  assign n23763 = n23666 & n23762 ;
  assign n23764 = n23763 ^ n21282 ;
  assign n23765 = n23764 ^ n23663 ;
  assign n23766 = ~n23664 & n23765 ;
  assign n23767 = n23766 ^ n21347 ;
  assign n23768 = n23767 ^ n23661 ;
  assign n23769 = ~n23662 & ~n23768 ;
  assign n23770 = n23769 ^ n21357 ;
  assign n23771 = n23770 ^ n23659 ;
  assign n23772 = ~n23660 & ~n23771 ;
  assign n23773 = n23772 ^ n21365 ;
  assign n23774 = n23773 ^ n23657 ;
  assign n23775 = n23658 & ~n23774 ;
  assign n23776 = n23775 ^ n21372 ;
  assign n23777 = n23776 ^ n23655 ;
  assign n23778 = ~n23656 & ~n23777 ;
  assign n23779 = n23778 ^ n21485 ;
  assign n23781 = n23780 ^ n23779 ;
  assign n23782 = n23780 ^ n20947 ;
  assign n23783 = n23781 & n23782 ;
  assign n23784 = n23783 ^ n20947 ;
  assign n23785 = n23784 ^ n23653 ;
  assign n23786 = n23654 & ~n23785 ;
  assign n23787 = n23786 ^ n20952 ;
  assign n23651 = n23650 ^ n23646 ;
  assign n24013 = n23787 ^ n23651 ;
  assign n24014 = n23787 ^ n20950 ;
  assign n24015 = n24013 & n24014 ;
  assign n24016 = n24015 ^ n20950 ;
  assign n24026 = n24025 ^ n24016 ;
  assign n23652 = n23651 ^ n20950 ;
  assign n23788 = n23787 ^ n23652 ;
  assign n23789 = n23779 ^ n20947 ;
  assign n23790 = n23789 ^ n23780 ;
  assign n23791 = n23759 ^ n21278 ;
  assign n23792 = n23747 ^ n23743 ;
  assign n23793 = n23737 ^ n23736 ;
  assign n23794 = n23732 ^ n23731 ;
  assign n23795 = n23709 ^ n23682 ;
  assign n23796 = n23706 ^ n23705 ;
  assign n23797 = n23701 ^ n23684 ;
  assign n23798 = n23685 ^ n20443 ;
  assign n23799 = n23798 ^ n23697 ;
  assign n23800 = n23694 ^ n23687 ;
  assign n23801 = n23688 ^ n20457 ;
  assign n23802 = n23691 ^ n23690 ;
  assign n23803 = n23801 & n23802 ;
  assign n23804 = ~n23800 & n23803 ;
  assign n23805 = ~n23799 & n23804 ;
  assign n23806 = ~n23797 & n23805 ;
  assign n23807 = n23796 & ~n23806 ;
  assign n23808 = ~n23795 & ~n23807 ;
  assign n23809 = n23713 ^ n21125 ;
  assign n23810 = ~n23808 & n23809 ;
  assign n23811 = n23716 ^ n23679 ;
  assign n23812 = n23810 & ~n23811 ;
  assign n23813 = n23719 ^ n21248 ;
  assign n23814 = n23813 ^ n23677 ;
  assign n23815 = n23812 & n23814 ;
  assign n23816 = n23725 ^ n21314 ;
  assign n23817 = ~n23815 & ~n23816 ;
  assign n23818 = n23727 ^ n23674 ;
  assign n23819 = ~n23817 & n23818 ;
  assign n23820 = ~n23794 & ~n23819 ;
  assign n23821 = n23793 & ~n23820 ;
  assign n23822 = n23740 ^ n23672 ;
  assign n23823 = n23821 & ~n23822 ;
  assign n23824 = n23792 & n23823 ;
  assign n23825 = n23749 ^ n23670 ;
  assign n23826 = n23824 & ~n23825 ;
  assign n23827 = n23752 ^ n21285 ;
  assign n23828 = n23827 ^ n23753 ;
  assign n23829 = ~n23826 & n23828 ;
  assign n23830 = ~n23791 & n23829 ;
  assign n23831 = n23761 ^ n21282 ;
  assign n23832 = n23831 ^ n23665 ;
  assign n23833 = ~n23830 & n23832 ;
  assign n23834 = n23764 ^ n21347 ;
  assign n23835 = n23834 ^ n23663 ;
  assign n23836 = n23833 & n23835 ;
  assign n23837 = n23767 ^ n23662 ;
  assign n23838 = ~n23836 & ~n23837 ;
  assign n23839 = n23770 ^ n21365 ;
  assign n23840 = n23839 ^ n23659 ;
  assign n23841 = ~n23838 & ~n23840 ;
  assign n23842 = n23773 ^ n23658 ;
  assign n23843 = n23841 & ~n23842 ;
  assign n23844 = n23776 ^ n21485 ;
  assign n23845 = n23844 ^ n23655 ;
  assign n23846 = ~n23843 & ~n23845 ;
  assign n23847 = n23790 & ~n23846 ;
  assign n23848 = n23784 ^ n23654 ;
  assign n23849 = n23847 & ~n23848 ;
  assign n24027 = n23788 & n23849 ;
  assign n24054 = ~n24026 & ~n24027 ;
  assign n24055 = n24024 ^ n24016 ;
  assign n24063 = n23486 ^ n23473 ;
  assign n24056 = n22202 ^ n21576 ;
  assign n24057 = n24056 ^ n22862 ;
  assign n24058 = n24057 ^ n24022 ;
  assign n24059 = n24058 ^ n24057 ;
  assign n24060 = n24059 ^ n24019 ;
  assign n24061 = n24023 & n24060 ;
  assign n24062 = n24061 ^ n24058 ;
  assign n24064 = n24063 ^ n24062 ;
  assign n24065 = n24064 ^ n20941 ;
  assign n24066 = n24065 ^ n24064 ;
  assign n24067 = n24066 ^ n24016 ;
  assign n24068 = ~n24055 & ~n24067 ;
  assign n24069 = n24068 ^ n24065 ;
  assign n24070 = n24069 ^ n20988 ;
  assign n24120 = ~n24054 & ~n24070 ;
  assign n24116 = n24064 ^ n20988 ;
  assign n24117 = n24069 & ~n24116 ;
  assign n24118 = n24117 ^ n20988 ;
  assign n24112 = n21856 ^ n21271 ;
  assign n24113 = n24112 ^ n22854 ;
  assign n24106 = n23489 ^ n23468 ;
  assign n24108 = n24106 ^ n24057 ;
  assign n24107 = n24106 ^ n24063 ;
  assign n24109 = n24108 ^ n24107 ;
  assign n24110 = ~n24062 & n24109 ;
  assign n24111 = n24110 ^ n24108 ;
  assign n24114 = n24113 ^ n24111 ;
  assign n24115 = n24114 ^ n20467 ;
  assign n24119 = n24118 ^ n24115 ;
  assign n24121 = n24120 ^ n24119 ;
  assign n24028 = n24027 ^ n24026 ;
  assign n24029 = n24028 ^ n2633 ;
  assign n23850 = n23849 ^ n23788 ;
  assign n2587 = n2577 ^ n2490 ;
  assign n2591 = n2590 ^ n2587 ;
  assign n2592 = n2591 ^ n2586 ;
  assign n23851 = n23850 ^ n2592 ;
  assign n24000 = n2872 ^ n2569 ;
  assign n24001 = n24000 ^ n18780 ;
  assign n24002 = n24001 ^ n1829 ;
  assign n24003 = n24002 ^ n3110 ;
  assign n23852 = n23846 ^ n23790 ;
  assign n23853 = n23852 ^ n3110 ;
  assign n23854 = n23845 ^ n23843 ;
  assign n23855 = n23854 ^ n2849 ;
  assign n23983 = n23840 ^ n23838 ;
  assign n23856 = n23837 ^ n23836 ;
  assign n1736 = n1416 ^ n1305 ;
  assign n1737 = n1736 ^ n1055 ;
  assign n1738 = n1737 ^ n1244 ;
  assign n23857 = n23856 ^ n1738 ;
  assign n23858 = n23835 ^ n23833 ;
  assign n23859 = n23858 ^ n1064 ;
  assign n23860 = n23832 ^ n23830 ;
  assign n897 = n896 ^ n856 ;
  assign n904 = n903 ^ n897 ;
  assign n908 = n907 ^ n904 ;
  assign n23861 = n23860 ^ n908 ;
  assign n23862 = n23829 ^ n23791 ;
  assign n23973 = n23862 ^ n908 ;
  assign n23863 = n23862 ^ n919 ;
  assign n23970 = n23862 ^ n818 ;
  assign n23864 = n23825 ^ n23824 ;
  assign n23865 = n23864 ^ n806 ;
  assign n23868 = n23823 ^ n23792 ;
  assign n23869 = n23868 ^ n1559 ;
  assign n23870 = n23822 ^ n23821 ;
  assign n23871 = n23870 ^ n1570 ;
  assign n23872 = n23820 ^ n23793 ;
  assign n23873 = n23872 ^ n2951 ;
  assign n23874 = n23819 ^ n23794 ;
  assign n23878 = n23877 ^ n23874 ;
  assign n23879 = n23818 ^ n23817 ;
  assign n23880 = n23879 ^ n596 ;
  assign n23885 = n23814 ^ n23812 ;
  assign n23886 = n23885 ^ n23884 ;
  assign n23887 = n23811 ^ n23810 ;
  assign n23888 = n23887 ^ n2390 ;
  assign n23889 = n23809 ^ n23808 ;
  assign n23890 = n23889 ^ n2277 ;
  assign n23931 = n23889 ^ n2259 ;
  assign n23891 = n23807 ^ n23795 ;
  assign n23892 = n23891 ^ n2259 ;
  assign n23893 = n23806 ^ n23796 ;
  assign n2241 = n2177 ^ n2122 ;
  assign n2248 = n2247 ^ n2241 ;
  assign n2249 = n2248 ^ n2075 ;
  assign n23894 = n23893 ^ n2249 ;
  assign n23896 = n21801 ^ n2102 ;
  assign n23897 = n23896 ^ n1976 ;
  assign n23898 = n23897 ^ n2244 ;
  assign n23895 = n23805 ^ n23797 ;
  assign n23899 = n23898 ^ n23895 ;
  assign n23903 = n23804 ^ n23799 ;
  assign n23900 = n21805 ^ n2106 ;
  assign n23901 = n23900 ^ n18828 ;
  assign n23902 = n23901 ^ n1974 ;
  assign n23904 = n23903 ^ n23902 ;
  assign n1899 = n1898 ^ n1877 ;
  assign n1906 = n1905 ^ n1899 ;
  assign n1910 = n1909 ^ n1906 ;
  assign n23919 = n23902 ^ n1910 ;
  assign n23908 = n1863 & ~n23801 ;
  assign n23905 = n21810 ^ n14844 ;
  assign n23906 = n23905 ^ n1867 ;
  assign n23907 = n23906 ^ n1903 ;
  assign n23909 = n23908 ^ n23907 ;
  assign n23912 = n23802 ^ n23801 ;
  assign n23913 = n23912 ^ n23907 ;
  assign n23914 = n23909 & n23913 ;
  assign n23910 = n23907 ^ n1910 ;
  assign n23915 = n23914 ^ n23910 ;
  assign n23916 = n23803 ^ n23800 ;
  assign n23917 = n23916 ^ n1910 ;
  assign n23918 = n23915 & ~n23917 ;
  assign n23920 = n23919 ^ n23918 ;
  assign n23921 = ~n23904 & ~n23920 ;
  assign n23922 = n23921 ^ n23903 ;
  assign n23923 = n23922 ^ n23895 ;
  assign n23924 = ~n23899 & ~n23923 ;
  assign n23925 = n23924 ^ n23898 ;
  assign n23926 = n23925 ^ n23893 ;
  assign n23927 = n23894 & ~n23926 ;
  assign n23928 = n23927 ^ n2249 ;
  assign n23929 = n23928 ^ n2259 ;
  assign n23930 = n23892 & n23929 ;
  assign n23932 = n23931 ^ n23930 ;
  assign n23933 = n23890 & ~n23932 ;
  assign n23934 = n23933 ^ n2277 ;
  assign n23935 = n23934 ^ n2390 ;
  assign n23936 = n23888 & ~n23935 ;
  assign n23937 = n23936 ^ n23887 ;
  assign n23938 = n23937 ^ n23884 ;
  assign n23939 = ~n23886 & n23938 ;
  assign n23940 = n23939 ^ n23884 ;
  assign n23881 = n23816 ^ n23815 ;
  assign n23941 = n23940 ^ n23881 ;
  assign n24172 = n23944 ^ n23881 ;
  assign n23948 = ~n23941 & n24172 ;
  assign n23945 = n23944 ^ n596 ;
  assign n23949 = n23948 ^ n23945 ;
  assign n23950 = n23880 & n23949 ;
  assign n23951 = n23950 ^ n596 ;
  assign n23952 = n23951 ^ n23874 ;
  assign n23953 = n23878 & ~n23952 ;
  assign n23954 = n23953 ^ n23877 ;
  assign n23955 = n23954 ^ n23872 ;
  assign n23956 = ~n23873 & n23955 ;
  assign n23957 = n23956 ^ n23954 ;
  assign n23958 = n23957 ^ n1570 ;
  assign n23959 = n23871 & ~n23958 ;
  assign n23960 = n23959 ^ n23870 ;
  assign n23961 = n23960 ^ n1559 ;
  assign n23962 = ~n23869 & ~n23961 ;
  assign n23963 = n23962 ^ n23868 ;
  assign n23964 = n23963 ^ n806 ;
  assign n23965 = n23865 & ~n23964 ;
  assign n23866 = n818 ^ n806 ;
  assign n23966 = n23965 ^ n23866 ;
  assign n23967 = n23828 ^ n23826 ;
  assign n23968 = n23967 ^ n818 ;
  assign n23969 = n23966 & ~n23968 ;
  assign n23971 = n23970 ^ n23969 ;
  assign n23972 = ~n23863 & ~n23971 ;
  assign n23974 = n23973 ^ n23972 ;
  assign n23975 = n23861 & n23974 ;
  assign n23976 = n23975 ^ n23860 ;
  assign n23977 = n23976 ^ n23858 ;
  assign n23978 = ~n23859 & n23977 ;
  assign n23979 = n23978 ^ n1064 ;
  assign n23980 = n23979 ^ n1738 ;
  assign n23981 = n23857 & ~n23980 ;
  assign n23982 = n23981 ^ n23856 ;
  assign n23984 = n23983 ^ n23982 ;
  assign n1257 = n1256 ^ n1157 ;
  assign n1258 = n1257 ^ n1250 ;
  assign n1259 = n1258 ^ n1238 ;
  assign n23987 = n23982 ^ n1259 ;
  assign n23988 = n23984 & n23987 ;
  assign n23985 = n2837 ^ n1259 ;
  assign n23989 = n23988 ^ n23985 ;
  assign n23991 = n23842 ^ n23841 ;
  assign n23992 = n23991 ^ n23854 ;
  assign n23990 = n23854 ^ n2837 ;
  assign n23993 = n23992 ^ n23990 ;
  assign n23994 = n23989 & n23993 ;
  assign n23995 = n23994 ^ n23990 ;
  assign n23996 = n23855 & n23995 ;
  assign n23997 = n23996 ^ n23854 ;
  assign n23998 = n23997 ^ n3110 ;
  assign n23999 = n23853 & n23998 ;
  assign n24004 = n24003 ^ n23999 ;
  assign n24007 = n23848 ^ n23847 ;
  assign n24008 = n24007 ^ n24002 ;
  assign n24009 = n24004 & n24008 ;
  assign n24005 = n24002 ^ n2592 ;
  assign n24010 = n24009 ^ n24005 ;
  assign n24011 = ~n23851 & n24010 ;
  assign n24012 = n24011 ^ n2592 ;
  assign n24073 = n24028 ^ n24012 ;
  assign n24074 = n24029 & ~n24073 ;
  assign n24075 = n24074 ^ n2633 ;
  assign n24071 = n24070 ^ n24054 ;
  assign n24100 = n24075 ^ n24071 ;
  assign n24103 = n24075 ^ n2532 ;
  assign n24104 = n24100 & n24103 ;
  assign n24101 = n3197 ^ n2532 ;
  assign n24105 = n24104 ^ n24101 ;
  assign n24122 = n24121 ^ n24105 ;
  assign n24098 = n22413 ^ n22395 ;
  assign n24099 = n24098 ^ n23320 ;
  assign n24123 = n24122 ^ n24099 ;
  assign n24072 = n24071 ^ n2532 ;
  assign n24076 = n24075 ^ n24072 ;
  assign n24052 = n22397 ^ n22353 ;
  assign n24053 = n24052 ^ n23322 ;
  assign n24077 = n24076 ^ n24053 ;
  assign n24033 = n22410 ^ n22273 ;
  assign n24034 = n24033 ^ n23332 ;
  assign n24035 = n24010 ^ n23850 ;
  assign n24036 = ~n24034 & ~n24035 ;
  assign n24031 = n22402 ^ n22301 ;
  assign n24032 = n24031 ^ n23328 ;
  assign n24037 = n24036 ^ n24032 ;
  assign n24030 = n24029 ^ n24012 ;
  assign n24049 = n24032 ^ n24030 ;
  assign n24050 = n24037 & n24049 ;
  assign n24051 = n24050 ^ n24032 ;
  assign n24095 = n24053 ^ n24051 ;
  assign n24096 = n24077 & n24095 ;
  assign n24097 = n24096 ^ n24076 ;
  assign n24124 = n24123 ^ n24097 ;
  assign n24125 = n24124 ^ n21622 ;
  assign n24039 = n24035 ^ n24034 ;
  assign n24040 = ~n21265 & n24039 ;
  assign n24041 = n24040 ^ n21260 ;
  assign n24038 = n24037 ^ n24030 ;
  assign n24045 = n24040 ^ n24038 ;
  assign n24046 = ~n24041 & ~n24045 ;
  assign n24047 = n24046 ^ n21260 ;
  assign n24048 = n24047 ^ n21262 ;
  assign n24078 = n24077 ^ n24051 ;
  assign n24092 = n24078 ^ n24047 ;
  assign n24093 = ~n24048 & n24092 ;
  assign n24094 = n24093 ^ n21262 ;
  assign n24338 = n24124 ^ n24094 ;
  assign n24339 = ~n24125 & ~n24338 ;
  assign n24340 = n24339 ^ n21622 ;
  assign n24451 = n24340 ^ n21628 ;
  assign n24235 = n24121 ^ n3197 ;
  assign n24236 = n24105 & n24235 ;
  assign n24227 = n23492 ^ n23466 ;
  assign n24225 = n23518 ^ n2753 ;
  assign n24226 = n24225 ^ n21855 ;
  assign n24228 = n24227 ^ n24226 ;
  assign n24229 = n24228 ^ n22852 ;
  assign n24230 = n24229 ^ n24113 ;
  assign n24231 = n24230 ^ n3197 ;
  assign n24232 = n24231 ^ n20467 ;
  assign n24224 = ~n24119 & n24120 ;
  assign n24233 = n24232 ^ n24224 ;
  assign n24222 = n24113 ^ n24106 ;
  assign n24223 = ~n24111 & ~n24222 ;
  assign n24234 = n24233 ^ n24223 ;
  assign n24237 = n24236 ^ n24234 ;
  assign n24219 = n24118 ^ n24114 ;
  assign n24220 = n24118 ^ n20467 ;
  assign n24221 = n24219 & n24220 ;
  assign n24238 = n24237 ^ n24221 ;
  assign n24242 = n24238 ^ n24122 ;
  assign n24240 = n24122 ^ n24097 ;
  assign n24241 = ~n24123 & ~n24240 ;
  assign n24243 = n24242 ^ n24241 ;
  assign n24216 = n22482 ^ n22390 ;
  assign n24217 = n24216 ^ n23314 ;
  assign n24336 = n24243 ^ n24217 ;
  assign n24452 = n24451 ^ n24336 ;
  assign n24042 = n24041 ^ n24038 ;
  assign n24043 = n24039 ^ n21265 ;
  assign n24044 = ~n24042 & ~n24043 ;
  assign n24079 = n24078 ^ n24048 ;
  assign n24091 = n24044 & ~n24079 ;
  assign n24126 = n24125 ^ n24094 ;
  assign n24450 = n24091 & ~n24126 ;
  assign n24565 = n24452 ^ n24450 ;
  assign n2023 = n2019 ^ n1983 ;
  assign n2027 = n2026 ^ n2023 ;
  assign n2031 = n2030 ^ n2027 ;
  assign n24566 = n24565 ^ n2031 ;
  assign n24127 = n24126 ^ n24091 ;
  assign n1964 = n1942 ^ n1927 ;
  assign n1965 = n1964 ^ n1961 ;
  assign n1969 = n1968 ^ n1965 ;
  assign n24128 = n24127 ^ n1969 ;
  assign n24080 = n24079 ^ n24044 ;
  assign n1946 = n1936 ^ n1918 ;
  assign n1953 = n1952 ^ n1946 ;
  assign n1957 = n1956 ^ n1953 ;
  assign n24081 = n24080 ^ n1957 ;
  assign n3055 = n3030 ^ n1889 ;
  assign n3059 = n3058 ^ n3055 ;
  assign n3060 = n3059 ^ n1949 ;
  assign n24087 = n3060 ^ n1957 ;
  assign n24082 = n3022 & n24043 ;
  assign n24083 = n24082 ^ n3060 ;
  assign n24084 = n24043 ^ n24042 ;
  assign n24085 = n24084 ^ n3060 ;
  assign n24086 = n24083 & n24085 ;
  assign n24088 = n24087 ^ n24086 ;
  assign n24089 = ~n24081 & n24088 ;
  assign n24090 = n24089 ^ n1957 ;
  assign n24567 = n24090 ^ n1969 ;
  assign n24568 = ~n24128 & n24567 ;
  assign n24569 = n24568 ^ n1969 ;
  assign n24570 = n24569 ^ n2031 ;
  assign n24571 = n24566 & ~n24570 ;
  assign n24572 = n24571 ^ n24565 ;
  assign n24239 = n24238 ^ n24217 ;
  assign n24244 = ~n24239 & n24243 ;
  assign n24214 = n23801 ^ n1863 ;
  assign n24218 = n24217 ^ n24214 ;
  assign n24245 = n24244 ^ n24218 ;
  assign n24212 = n23576 ^ n22408 ;
  assign n24213 = n24212 ^ n22385 ;
  assign n24344 = n24245 ^ n24213 ;
  assign n24346 = n24344 ^ n21636 ;
  assign n24337 = n24336 ^ n21628 ;
  assign n24341 = n24340 ^ n24336 ;
  assign n24342 = ~n24337 & ~n24341 ;
  assign n24343 = n24342 ^ n21628 ;
  assign n24454 = n24346 ^ n24343 ;
  assign n24453 = n24450 & n24452 ;
  assign n24563 = n24454 ^ n24453 ;
  assign n24560 = n22319 ^ n2325 ;
  assign n24561 = n24560 ^ n2035 ;
  assign n24562 = n24561 ^ n2140 ;
  assign n24564 = n24563 ^ n24562 ;
  assign n24720 = n24572 ^ n24564 ;
  assign n24181 = n23932 ^ n2277 ;
  assign n25173 = n24720 ^ n24181 ;
  assign n25174 = n25173 ^ n23597 ;
  assign n24694 = n23528 ^ n3037 ;
  assign n24695 = n24694 ^ n20332 ;
  assign n24696 = n24695 ^ n1791 ;
  assign n24647 = n22741 ^ n3115 ;
  assign n24648 = n24647 ^ n2510 ;
  assign n24649 = n24648 ^ n3096 ;
  assign n24650 = n24649 ^ n24512 ;
  assign n24142 = n23967 ^ n23966 ;
  assign n24140 = n23647 ^ n23259 ;
  assign n24141 = n24140 ^ n22555 ;
  assign n24143 = n24142 ^ n24141 ;
  assign n24146 = n23963 ^ n23865 ;
  assign n24144 = n23264 ^ n22547 ;
  assign n24145 = n24144 ^ n23248 ;
  assign n24147 = n24146 ^ n24145 ;
  assign n24149 = n23270 ^ n22539 ;
  assign n24150 = n24149 ^ n23256 ;
  assign n24148 = n23960 ^ n23869 ;
  assign n24151 = n24150 ^ n24148 ;
  assign n24154 = n23957 ^ n23871 ;
  assign n24152 = n23275 ^ n22433 ;
  assign n24153 = n24152 ^ n23261 ;
  assign n24155 = n24154 ^ n24153 ;
  assign n24160 = n23954 ^ n23873 ;
  assign n24158 = n23266 ^ n22431 ;
  assign n24159 = n24158 ^ n23282 ;
  assign n24161 = n24160 ^ n24159 ;
  assign n24164 = n23951 ^ n23878 ;
  assign n24162 = n23272 ^ n22436 ;
  assign n24163 = n24162 ^ n23287 ;
  assign n24165 = n24164 ^ n24163 ;
  assign n24168 = n23949 ^ n23879 ;
  assign n24166 = n23294 ^ n23277 ;
  assign n24167 = n24166 ^ n22440 ;
  assign n24169 = n24168 ^ n24167 ;
  assign n24173 = n24172 ^ n23940 ;
  assign n24170 = n23284 ^ n22444 ;
  assign n24171 = n24170 ^ n23298 ;
  assign n24174 = n24173 ^ n24171 ;
  assign n24176 = n23232 ^ n22448 ;
  assign n24177 = n24176 ^ n23289 ;
  assign n24175 = n23937 ^ n23886 ;
  assign n24178 = n24177 ^ n24175 ;
  assign n24183 = n23934 ^ n23888 ;
  assign n24271 = n24183 ^ n24175 ;
  assign n24179 = n23300 ^ n21851 ;
  assign n24180 = n24179 ^ n23197 ;
  assign n24182 = n24181 ^ n24180 ;
  assign n24188 = n23928 ^ n23892 ;
  assign n24186 = n23304 ^ n23169 ;
  assign n24187 = n24186 ^ n22379 ;
  assign n24189 = n24188 ^ n24187 ;
  assign n24193 = n23925 ^ n23894 ;
  assign n24190 = n23611 ^ n22383 ;
  assign n24191 = n24190 ^ n23015 ;
  assign n24194 = n24193 ^ n24191 ;
  assign n24196 = n23308 ^ n23003 ;
  assign n24197 = n24196 ^ n22388 ;
  assign n24195 = n23922 ^ n23899 ;
  assign n24198 = n24197 ^ n24195 ;
  assign n24201 = n23312 ^ n22918 ;
  assign n24202 = n24201 ^ n22393 ;
  assign n24130 = n23920 ^ n23903 ;
  assign n24203 = n24202 ^ n24130 ;
  assign n24206 = n23916 ^ n23915 ;
  assign n24204 = n23597 ^ n22398 ;
  assign n24205 = n24204 ^ n22374 ;
  assign n24207 = n24206 ^ n24205 ;
  assign n24209 = n23579 ^ n22404 ;
  assign n24210 = n24209 ^ n22376 ;
  assign n24208 = n23912 ^ n23909 ;
  assign n24211 = n24210 ^ n24208 ;
  assign n24247 = n24214 ^ n24208 ;
  assign n24215 = n24214 ^ n24213 ;
  assign n24246 = n24215 & ~n24245 ;
  assign n24248 = n24247 ^ n24246 ;
  assign n24249 = ~n24211 & n24248 ;
  assign n24250 = n24249 ^ n24210 ;
  assign n24251 = n24250 ^ n24205 ;
  assign n24252 = ~n24207 & n24251 ;
  assign n24253 = n24252 ^ n24206 ;
  assign n24254 = n24253 ^ n24130 ;
  assign n24255 = n24203 & ~n24254 ;
  assign n24256 = n24255 ^ n24202 ;
  assign n24257 = n24256 ^ n24195 ;
  assign n24258 = ~n24198 & ~n24257 ;
  assign n24199 = n24195 ^ n24191 ;
  assign n24259 = n24258 ^ n24199 ;
  assign n24260 = ~n24194 & ~n24259 ;
  assign n24192 = n24191 ^ n24188 ;
  assign n24261 = n24260 ^ n24192 ;
  assign n24262 = ~n24189 & ~n24261 ;
  assign n24263 = n24262 ^ n24188 ;
  assign n24184 = n24183 ^ n24181 ;
  assign n24185 = n24184 ^ n24183 ;
  assign n24264 = n24263 ^ n24185 ;
  assign n24265 = ~n24182 & n24264 ;
  assign n24266 = n24265 ^ n24184 ;
  assign n24267 = n23291 ^ n22452 ;
  assign n24268 = n24267 ^ n23217 ;
  assign n24269 = n24268 ^ n24183 ;
  assign n24270 = n24266 & n24269 ;
  assign n24272 = n24271 ^ n24270 ;
  assign n24273 = n24178 & n24272 ;
  assign n24274 = n24273 ^ n24177 ;
  assign n24275 = n24274 ^ n24171 ;
  assign n24276 = ~n24174 & ~n24275 ;
  assign n24277 = n24276 ^ n24173 ;
  assign n24278 = n24277 ^ n24167 ;
  assign n24279 = n24169 & ~n24278 ;
  assign n24280 = n24279 ^ n24168 ;
  assign n24281 = n24280 ^ n24163 ;
  assign n24282 = n24165 & ~n24281 ;
  assign n24283 = n24282 ^ n24164 ;
  assign n24284 = n24283 ^ n24159 ;
  assign n24285 = n24161 & ~n24284 ;
  assign n24286 = n24285 ^ n24160 ;
  assign n24287 = n24286 ^ n24154 ;
  assign n24288 = ~n24155 & n24287 ;
  assign n24156 = n24154 ^ n24150 ;
  assign n24289 = n24288 ^ n24156 ;
  assign n24290 = n24151 & ~n24289 ;
  assign n24291 = n24290 ^ n24150 ;
  assign n24292 = n24291 ^ n24146 ;
  assign n24293 = ~n24147 & n24292 ;
  assign n24294 = n24293 ^ n24291 ;
  assign n24295 = n24294 ^ n24141 ;
  assign n24296 = n24143 & ~n24295 ;
  assign n24297 = n24296 ^ n24142 ;
  assign n24138 = n23971 ^ n919 ;
  assign n24136 = n23254 ^ n22563 ;
  assign n24137 = n24136 ^ n24022 ;
  assign n24139 = n24138 ^ n24137 ;
  assign n24311 = n24297 ^ n24139 ;
  assign n24312 = n24311 ^ n22053 ;
  assign n24313 = n24294 ^ n24143 ;
  assign n24314 = n24313 ^ n21965 ;
  assign n24315 = n24291 ^ n24147 ;
  assign n24316 = n24315 ^ n21957 ;
  assign n24318 = n24286 ^ n24155 ;
  assign n24319 = n24318 ^ n21940 ;
  assign n24321 = n24280 ^ n24165 ;
  assign n24322 = n24321 ^ n21922 ;
  assign n24324 = n24272 ^ n24177 ;
  assign n24325 = n24324 ^ n21255 ;
  assign n24376 = n24268 ^ n24266 ;
  assign n24327 = n24261 ^ n24187 ;
  assign n24328 = n24327 ^ n21882 ;
  assign n24363 = n24259 ^ n24193 ;
  assign n24329 = n24256 ^ n24198 ;
  assign n24330 = n24329 ^ n21891 ;
  assign n24332 = n24250 ^ n24207 ;
  assign n24333 = n24332 ^ n21753 ;
  assign n24334 = n24248 ^ n24210 ;
  assign n24335 = n24334 ^ n21736 ;
  assign n24345 = n24344 ^ n24343 ;
  assign n24347 = ~n24345 & n24346 ;
  assign n24348 = n24347 ^ n21636 ;
  assign n24349 = n24348 ^ n24334 ;
  assign n24350 = n24335 & ~n24349 ;
  assign n24351 = n24350 ^ n21736 ;
  assign n24352 = n24351 ^ n24332 ;
  assign n24353 = ~n24333 & ~n24352 ;
  assign n24354 = n24353 ^ n21753 ;
  assign n24331 = n24253 ^ n24203 ;
  assign n24355 = n24354 ^ n24331 ;
  assign n24356 = n24329 ^ n21893 ;
  assign n24357 = n24356 ^ n24329 ;
  assign n24358 = n24357 ^ n24331 ;
  assign n24359 = ~n24355 & n24358 ;
  assign n24360 = n24359 ^ n24356 ;
  assign n24361 = ~n24330 & n24360 ;
  assign n24362 = n24361 ^ n21891 ;
  assign n24364 = n24363 ^ n24362 ;
  assign n24365 = n24327 ^ n21884 ;
  assign n24366 = n24365 ^ n24327 ;
  assign n24367 = n24366 ^ n24362 ;
  assign n24368 = ~n24364 & n24367 ;
  assign n24369 = n24368 ^ n24365 ;
  assign n24370 = ~n24328 & n24369 ;
  assign n24371 = n24370 ^ n21882 ;
  assign n24326 = n24263 ^ n24182 ;
  assign n24372 = n24371 ^ n24326 ;
  assign n24373 = n24371 ^ n21875 ;
  assign n24374 = ~n24372 & n24373 ;
  assign n24375 = n24374 ^ n21875 ;
  assign n24377 = n24376 ^ n24375 ;
  assign n24378 = n24324 ^ n21873 ;
  assign n24379 = n24378 ^ n24324 ;
  assign n24380 = n24379 ^ n24375 ;
  assign n24381 = n24377 & ~n24380 ;
  assign n24382 = n24381 ^ n24378 ;
  assign n24383 = ~n24325 & ~n24382 ;
  assign n24384 = n24383 ^ n21255 ;
  assign n24323 = n24274 ^ n24174 ;
  assign n24385 = n24384 ^ n24323 ;
  assign n24386 = n24277 ^ n24169 ;
  assign n24387 = n24386 ^ n21863 ;
  assign n24388 = n24387 ^ n24323 ;
  assign n24389 = n24388 ^ n24386 ;
  assign n24390 = n24385 & n24389 ;
  assign n24391 = n24390 ^ n24387 ;
  assign n24393 = n24321 ^ n21865 ;
  assign n24392 = n24386 ^ n24321 ;
  assign n24394 = n24393 ^ n24392 ;
  assign n24395 = ~n24391 & ~n24394 ;
  assign n24396 = n24395 ^ n24393 ;
  assign n24397 = ~n24322 & n24396 ;
  assign n24398 = n24397 ^ n21922 ;
  assign n24320 = n24283 ^ n24161 ;
  assign n24399 = n24398 ^ n24320 ;
  assign n24400 = n24318 ^ n21932 ;
  assign n24401 = n24400 ^ n24318 ;
  assign n24402 = n24401 ^ n24320 ;
  assign n24403 = n24399 & n24402 ;
  assign n24404 = n24403 ^ n24400 ;
  assign n24405 = n24319 & n24404 ;
  assign n24406 = n24405 ^ n21940 ;
  assign n24317 = n24289 ^ n24148 ;
  assign n24407 = n24406 ^ n24317 ;
  assign n24408 = n24315 ^ n21949 ;
  assign n24409 = n24408 ^ n24317 ;
  assign n24410 = n24409 ^ n24315 ;
  assign n24411 = n24407 & ~n24410 ;
  assign n24412 = n24411 ^ n24408 ;
  assign n24413 = ~n24316 & ~n24412 ;
  assign n24414 = n24413 ^ n21957 ;
  assign n24415 = n24414 ^ n24313 ;
  assign n24416 = n24314 & n24415 ;
  assign n24417 = n24416 ^ n21965 ;
  assign n24418 = n24417 ^ n24311 ;
  assign n24419 = n24312 & ~n24418 ;
  assign n24420 = n24419 ^ n22053 ;
  assign n24422 = n24420 ^ n22196 ;
  assign n24298 = n24297 ^ n24137 ;
  assign n24299 = n24139 & ~n24298 ;
  assign n24300 = n24299 ^ n24138 ;
  assign n24134 = n23974 ^ n23860 ;
  assign n24132 = n24063 ^ n22421 ;
  assign n24133 = n24132 ^ n23250 ;
  assign n24135 = n24134 ^ n24133 ;
  assign n24310 = n24300 ^ n24135 ;
  assign n24488 = n24422 ^ n24310 ;
  assign n24439 = n24414 ^ n24314 ;
  assign n24440 = n24412 ^ n21957 ;
  assign n24441 = n24376 ^ n21873 ;
  assign n24442 = n24441 ^ n24375 ;
  assign n24443 = n24326 ^ n21875 ;
  assign n24444 = n24443 ^ n24371 ;
  assign n24445 = n24369 ^ n21882 ;
  assign n24446 = n24362 ^ n21884 ;
  assign n24447 = n24446 ^ n24363 ;
  assign n24448 = n24354 ^ n21893 ;
  assign n24449 = n24448 ^ n24331 ;
  assign n24455 = ~n24453 & ~n24454 ;
  assign n24456 = n24348 ^ n24335 ;
  assign n24457 = ~n24455 & n24456 ;
  assign n24458 = n24351 ^ n24333 ;
  assign n24459 = ~n24457 & n24458 ;
  assign n24460 = n24449 & n24459 ;
  assign n24461 = n24360 ^ n21891 ;
  assign n24462 = n24460 & ~n24461 ;
  assign n24463 = ~n24447 & ~n24462 ;
  assign n24464 = ~n24445 & ~n24463 ;
  assign n24465 = ~n24444 & ~n24464 ;
  assign n24466 = n24442 & ~n24465 ;
  assign n24467 = n24382 ^ n21255 ;
  assign n24468 = n24466 & n24467 ;
  assign n24469 = n24323 ^ n21863 ;
  assign n24470 = n24469 ^ n24384 ;
  assign n24471 = n24468 & n24470 ;
  assign n24472 = n24391 ^ n21865 ;
  assign n24473 = n24471 & n24472 ;
  assign n24474 = n24396 ^ n21922 ;
  assign n24475 = ~n24473 & n24474 ;
  assign n24476 = n24320 ^ n21932 ;
  assign n24477 = n24476 ^ n24398 ;
  assign n24478 = n24475 & ~n24477 ;
  assign n24479 = n24404 ^ n21940 ;
  assign n24480 = ~n24478 & ~n24479 ;
  assign n24481 = n24317 ^ n21949 ;
  assign n24482 = n24481 ^ n24406 ;
  assign n24483 = n24480 & ~n24482 ;
  assign n24484 = n24440 & ~n24483 ;
  assign n24485 = ~n24439 & ~n24484 ;
  assign n24486 = n24417 ^ n24312 ;
  assign n24487 = n24485 & n24486 ;
  assign n24508 = n24488 ^ n24487 ;
  assign n24509 = n24508 ^ n2642 ;
  assign n24515 = n24486 ^ n24485 ;
  assign n1377 = n1376 ^ n1241 ;
  assign n1378 = n1377 ^ n1340 ;
  assign n1379 = n1378 ^ n1373 ;
  assign n24516 = n24515 ^ n1379 ;
  assign n24517 = n24484 ^ n24439 ;
  assign n24518 = n24517 ^ n1346 ;
  assign n24519 = n24483 ^ n24440 ;
  assign n24520 = n24519 ^ n1175 ;
  assign n24521 = n24482 ^ n24480 ;
  assign n24522 = n24521 ^ n1047 ;
  assign n24523 = n24479 ^ n24478 ;
  assign n1024 = n990 ^ n948 ;
  assign n1025 = n1024 ^ n1021 ;
  assign n1029 = n1028 ^ n1025 ;
  assign n24524 = n24523 ^ n1029 ;
  assign n24525 = n24477 ^ n24475 ;
  assign n24526 = n24525 ^ n1017 ;
  assign n24622 = n1631 ^ n1017 ;
  assign n24527 = n24472 ^ n24471 ;
  assign n24528 = n24527 ^ n1625 ;
  assign n24531 = n24470 ^ n24468 ;
  assign n24532 = n24531 ^ n653 ;
  assign n24612 = n2965 ^ n653 ;
  assign n24533 = n24467 ^ n24466 ;
  assign n24534 = n24533 ^ n2965 ;
  assign n24539 = n24463 ^ n24445 ;
  assign n24540 = n24539 ^ n1487 ;
  assign n24541 = n24462 ^ n24447 ;
  assign n24545 = n24544 ^ n24541 ;
  assign n24547 = n2402 ^ n2353 ;
  assign n24548 = n24547 ^ n2282 ;
  assign n24549 = n24548 ^ n14260 ;
  assign n24546 = n24459 ^ n24449 ;
  assign n24550 = n24549 ^ n24546 ;
  assign n24554 = n24458 ^ n24457 ;
  assign n24558 = n24557 ^ n24554 ;
  assign n24573 = n24572 ^ n24562 ;
  assign n24574 = ~n24564 & n24573 ;
  assign n24575 = n24574 ^ n24562 ;
  assign n24579 = n24575 ^ n24557 ;
  assign n24559 = n24456 ^ n24455 ;
  assign n24576 = n24575 ^ n24559 ;
  assign n2136 = n2135 ^ n2081 ;
  assign n2143 = n2142 ^ n2136 ;
  assign n2147 = n2146 ^ n2143 ;
  assign n24577 = n24559 ^ n2147 ;
  assign n24578 = ~n24576 & n24577 ;
  assign n24580 = n24579 ^ n24578 ;
  assign n24581 = n24558 & n24580 ;
  assign n24582 = n24581 ^ n24557 ;
  assign n24551 = n24461 ^ n24460 ;
  assign n24552 = n24551 ^ n24549 ;
  assign n24553 = n24552 ^ n24551 ;
  assign n24583 = n24582 ^ n24553 ;
  assign n24584 = ~n24550 & n24583 ;
  assign n24585 = n24584 ^ n24552 ;
  assign n24587 = n2428 ^ n1454 ;
  assign n24588 = n24587 ^ n19513 ;
  assign n24589 = n24588 ^ n2906 ;
  assign n24590 = n24589 ^ n24544 ;
  assign n24586 = n24551 ^ n24544 ;
  assign n24591 = n24590 ^ n24586 ;
  assign n24592 = ~n24585 & n24591 ;
  assign n24593 = n24592 ^ n24590 ;
  assign n24594 = n24545 & n24593 ;
  assign n24595 = n24594 ^ n24544 ;
  assign n24596 = n24595 ^ n1487 ;
  assign n24597 = ~n24540 & n24596 ;
  assign n24538 = n24537 ^ n1487 ;
  assign n24598 = n24597 ^ n24538 ;
  assign n24602 = n24464 ^ n24444 ;
  assign n24599 = n24465 ^ n24442 ;
  assign n24600 = n24599 ^ n24537 ;
  assign n24601 = n24600 ^ n24599 ;
  assign n24603 = n24602 ^ n24601 ;
  assign n24604 = n24598 & n24603 ;
  assign n24605 = n24604 ^ n24600 ;
  assign n24607 = n24599 ^ n2965 ;
  assign n24606 = n2965 ^ n618 ;
  assign n24608 = n24607 ^ n24606 ;
  assign n24609 = ~n24605 & n24608 ;
  assign n24610 = n24609 ^ n24606 ;
  assign n24611 = ~n24534 & n24610 ;
  assign n24613 = n24612 ^ n24611 ;
  assign n24614 = ~n24532 & ~n24613 ;
  assign n24615 = n24614 ^ n24531 ;
  assign n24616 = n24615 ^ n1625 ;
  assign n24617 = ~n24528 & ~n24616 ;
  assign n24529 = n1631 ^ n1625 ;
  assign n24618 = n24617 ^ n24529 ;
  assign n24619 = n24474 ^ n24473 ;
  assign n24620 = n24619 ^ n1631 ;
  assign n24621 = n24618 & ~n24620 ;
  assign n24623 = n24622 ^ n24621 ;
  assign n24624 = ~n24526 & ~n24623 ;
  assign n24625 = n24624 ^ n24525 ;
  assign n24626 = n24625 ^ n1029 ;
  assign n24627 = ~n24524 & n24626 ;
  assign n24628 = n24627 ^ n24523 ;
  assign n24629 = n24628 ^ n1047 ;
  assign n24630 = n24522 & n24629 ;
  assign n24631 = n24630 ^ n24521 ;
  assign n24632 = n24631 ^ n1175 ;
  assign n24633 = ~n24520 & ~n24632 ;
  assign n24634 = n24633 ^ n24519 ;
  assign n24635 = n24634 ^ n24517 ;
  assign n24636 = ~n24518 & ~n24635 ;
  assign n24637 = n24636 ^ n1346 ;
  assign n24638 = n24637 ^ n24515 ;
  assign n24639 = ~n24516 & n24638 ;
  assign n24640 = n24639 ^ n1379 ;
  assign n24513 = n24512 ^ n2642 ;
  assign n24514 = n24513 ^ n24512 ;
  assign n24641 = n24640 ^ n24514 ;
  assign n24642 = ~n24509 & n24641 ;
  assign n24643 = n24642 ^ n24513 ;
  assign n24489 = ~n24487 & n24488 ;
  assign n24421 = n24420 ^ n24310 ;
  assign n24423 = ~n24421 & ~n24422 ;
  assign n24424 = n24423 ^ n22196 ;
  assign n24306 = n23976 ^ n23859 ;
  assign n24304 = n24106 ^ n22866 ;
  assign n24305 = n24304 ^ n22210 ;
  assign n24307 = n24306 ^ n24305 ;
  assign n24301 = n24300 ^ n24133 ;
  assign n24302 = n24135 & ~n24301 ;
  assign n24303 = n24302 ^ n24134 ;
  assign n24308 = n24307 ^ n24303 ;
  assign n24309 = n24308 ^ n21591 ;
  assign n24438 = n24424 ^ n24309 ;
  assign n24644 = n24489 ^ n24438 ;
  assign n24645 = n24644 ^ n24512 ;
  assign n24646 = n24643 & ~n24645 ;
  assign n24651 = n24650 ^ n24646 ;
  assign n24490 = ~n24438 & ~n24489 ;
  assign n24433 = n23979 ^ n23857 ;
  assign n24431 = n22872 ^ n22216 ;
  assign n24432 = n24431 ^ n24227 ;
  assign n24434 = n24433 ^ n24432 ;
  assign n24428 = n24305 ^ n24303 ;
  assign n24429 = n24307 & ~n24428 ;
  assign n24430 = n24429 ^ n24306 ;
  assign n24435 = n24434 ^ n24430 ;
  assign n24436 = n24435 ^ n21594 ;
  assign n24425 = n24424 ^ n24308 ;
  assign n24426 = n24309 & n24425 ;
  assign n24427 = n24426 ^ n21591 ;
  assign n24437 = n24436 ^ n24427 ;
  assign n24654 = n24490 ^ n24437 ;
  assign n24655 = n24654 ^ n24649 ;
  assign n24656 = n24651 & n24655 ;
  assign n24502 = n24435 ^ n24427 ;
  assign n24503 = ~n24436 & n24502 ;
  assign n24504 = n24503 ^ n21594 ;
  assign n24497 = n23983 ^ n1259 ;
  assign n24498 = n24497 ^ n23982 ;
  assign n24495 = n23547 ^ n22862 ;
  assign n24496 = n24495 ^ n22213 ;
  assign n24499 = n24498 ^ n24496 ;
  assign n24492 = n24432 ^ n24430 ;
  assign n24493 = ~n24434 & ~n24492 ;
  assign n24494 = n24493 ^ n24433 ;
  assign n24500 = n24499 ^ n24494 ;
  assign n24501 = n24500 ^ n21583 ;
  assign n24505 = n24504 ^ n24501 ;
  assign n24491 = ~n24437 & n24490 ;
  assign n24506 = n24505 ^ n24491 ;
  assign n24652 = n24649 ^ n24506 ;
  assign n24657 = n24656 ^ n24652 ;
  assign n24682 = n24657 ^ n3104 ;
  assign n24680 = n24214 ^ n22410 ;
  assign n24681 = n24680 ^ n23322 ;
  assign n24688 = n24682 ^ n24681 ;
  assign n24692 = n24688 ^ n22273 ;
  assign n25172 = n24696 ^ n24692 ;
  assign n25175 = n25174 ^ n25172 ;
  assign n24724 = n24569 ^ n24566 ;
  assign n25451 = n24724 ^ n23579 ;
  assign n25452 = n25451 ^ n24188 ;
  assign n3159 = n3157 ^ n2763 ;
  assign n3160 = n3159 ^ n2474 ;
  assign n3161 = n3160 ^ n1808 ;
  assign n25448 = n3161 ^ n1847 ;
  assign n25443 = n24654 ^ n24651 ;
  assign n25441 = n24238 ^ n23328 ;
  assign n25442 = n25441 ^ n22887 ;
  assign n25444 = n25443 ^ n25442 ;
  assign n25180 = n24644 ^ n24643 ;
  assign n25440 = n25180 ^ n21857 ;
  assign n25445 = n25444 ^ n25440 ;
  assign n25177 = n24076 ^ n23531 ;
  assign n25178 = n25177 ^ n22852 ;
  assign n25176 = n24640 ^ n24509 ;
  assign n25179 = n25178 ^ n25176 ;
  assign n25183 = n23533 ^ n22854 ;
  assign n25184 = n25183 ^ n24030 ;
  assign n25109 = n24637 ^ n24516 ;
  assign n25185 = n25184 ^ n25109 ;
  assign n25186 = n24035 ^ n23537 ;
  assign n25187 = n25186 ^ n22862 ;
  assign n25105 = n24634 ^ n24518 ;
  assign n25188 = n25187 ^ n25105 ;
  assign n25115 = n24631 ^ n24520 ;
  assign n25251 = n25115 ^ n25105 ;
  assign n24781 = n24007 ^ n24004 ;
  assign n25189 = n24781 ^ n23550 ;
  assign n25190 = n25189 ^ n22872 ;
  assign n25191 = n25190 ^ n25115 ;
  assign n24766 = n23997 ^ n23853 ;
  assign n25192 = n24766 ^ n22866 ;
  assign n25193 = n25192 ^ n23547 ;
  assign n25120 = n24628 ^ n24522 ;
  assign n25194 = n25193 ^ n25120 ;
  assign n24753 = n23995 ^ n2849 ;
  assign n25195 = n24753 ^ n23250 ;
  assign n25196 = n25195 ^ n24227 ;
  assign n25124 = n24625 ^ n24524 ;
  assign n25197 = n25196 ^ n25124 ;
  assign n25232 = n24623 ^ n24525 ;
  assign n25242 = n25232 ^ n25124 ;
  assign n25200 = n24615 ^ n24528 ;
  assign n25198 = n24022 ^ n23264 ;
  assign n25199 = n25198 ^ n24433 ;
  assign n25201 = n25200 ^ n25199 ;
  assign n25206 = n24306 ^ n23647 ;
  assign n25207 = n25206 ^ n23270 ;
  assign n25129 = n24613 ^ n24531 ;
  assign n25208 = n25207 ^ n25129 ;
  assign n25209 = n24134 ^ n23248 ;
  assign n25210 = n25209 ^ n23275 ;
  assign n25135 = n24610 ^ n24533 ;
  assign n25211 = n25210 ^ n25135 ;
  assign n25214 = n24138 ^ n23282 ;
  assign n25215 = n25214 ^ n23256 ;
  assign n25141 = n24605 ^ n618 ;
  assign n25216 = n25215 ^ n25141 ;
  assign n25091 = n24602 ^ n24598 ;
  assign n25089 = n24142 ^ n23261 ;
  assign n25090 = n25089 ^ n23287 ;
  assign n25092 = n25091 ^ n25090 ;
  assign n24861 = n24148 ^ n23298 ;
  assign n24862 = n24861 ^ n23272 ;
  assign n24860 = n24593 ^ n24541 ;
  assign n24863 = n24862 ^ n24860 ;
  assign n25067 = n24146 ^ n23266 ;
  assign n25068 = n25067 ^ n23294 ;
  assign n25069 = n25068 ^ n24860 ;
  assign n25070 = n25069 ^ n25068 ;
  assign n24706 = n24589 ^ n24585 ;
  assign n24704 = n24154 ^ n23277 ;
  assign n24705 = n24704 ^ n23232 ;
  assign n24707 = n24706 ^ n24705 ;
  assign n24710 = n24580 ^ n24554 ;
  assign n24708 = n24164 ^ n23197 ;
  assign n24709 = n24708 ^ n23289 ;
  assign n24711 = n24710 ^ n24709 ;
  assign n24717 = n23291 ^ n23169 ;
  assign n24718 = n24717 ^ n24168 ;
  assign n24716 = n24577 ^ n24575 ;
  assign n24719 = n24718 ^ n24716 ;
  assign n24721 = n24173 ^ n23015 ;
  assign n24722 = n24721 ^ n23300 ;
  assign n24723 = n24722 ^ n24720 ;
  assign n24725 = n24175 ^ n23003 ;
  assign n24726 = n24725 ^ n23304 ;
  assign n24727 = n24726 ^ n24724 ;
  assign n24730 = n24183 ^ n22918 ;
  assign n24731 = n24730 ^ n23611 ;
  assign n24129 = n24128 ^ n24090 ;
  assign n24732 = n24731 ^ n24129 ;
  assign n24734 = n24181 ^ n22374 ;
  assign n24735 = n24734 ^ n23308 ;
  assign n24733 = n24088 ^ n24080 ;
  assign n24736 = n24735 ^ n24733 ;
  assign n24739 = n24084 ^ n24083 ;
  assign n24737 = n24188 ^ n22376 ;
  assign n24738 = n24737 ^ n23312 ;
  assign n24740 = n24739 ^ n24738 ;
  assign n24743 = n24043 ^ n3022 ;
  assign n24831 = n24743 ^ n24738 ;
  assign n24741 = n23597 ^ n22385 ;
  assign n24742 = n24741 ^ n24193 ;
  assign n24744 = n24743 ^ n24742 ;
  assign n24668 = n23991 ^ n23989 ;
  assign n24666 = n23550 ^ n22854 ;
  assign n24667 = n24666 ^ n22222 ;
  assign n24669 = n24668 ^ n24667 ;
  assign n24663 = n24496 ^ n24494 ;
  assign n24664 = ~n24499 & ~n24663 ;
  assign n24665 = n24664 ^ n24498 ;
  assign n24670 = n24669 ^ n24665 ;
  assign n24671 = n24670 ^ n21578 ;
  assign n24660 = n24504 ^ n24500 ;
  assign n24661 = ~n24501 & ~n24660 ;
  assign n24662 = n24661 ^ n21583 ;
  assign n24755 = n24670 ^ n24662 ;
  assign n24756 = ~n24671 & ~n24755 ;
  assign n24757 = n24756 ^ n21578 ;
  assign n24750 = n22852 ^ n22202 ;
  assign n24751 = n24750 ^ n23537 ;
  assign n24747 = n24667 ^ n24665 ;
  assign n24748 = ~n24669 & ~n24747 ;
  assign n24749 = n24748 ^ n24668 ;
  assign n24752 = n24751 ^ n24749 ;
  assign n24754 = n24753 ^ n24752 ;
  assign n24758 = n24757 ^ n24754 ;
  assign n24759 = n24757 ^ n21576 ;
  assign n24760 = ~n24758 & n24759 ;
  assign n24761 = n24760 ^ n21576 ;
  assign n24793 = n24761 ^ n21271 ;
  assign n24772 = n22412 ^ n21856 ;
  assign n24773 = n24772 ^ n23533 ;
  assign n24767 = n24766 ^ n24753 ;
  assign n24768 = n24767 ^ n24766 ;
  assign n24769 = n24768 ^ n24749 ;
  assign n24770 = n24752 & n24769 ;
  assign n24771 = n24770 ^ n24767 ;
  assign n24774 = n24773 ^ n24771 ;
  assign n24794 = n24793 ^ n24774 ;
  assign n24672 = n24671 ^ n24662 ;
  assign n24673 = n24491 & ~n24505 ;
  assign n24762 = ~n24672 & ~n24673 ;
  assign n24763 = n24754 ^ n21576 ;
  assign n24764 = n24763 ^ n24757 ;
  assign n24765 = ~n24762 & n24764 ;
  assign n24795 = n24794 ^ n24765 ;
  assign n24796 = n24795 ^ n2723 ;
  assign n24797 = n24764 ^ n24762 ;
  assign n2715 = n2669 ^ n2615 ;
  assign n2716 = n2715 ^ n1838 ;
  assign n2717 = n2716 ^ n2711 ;
  assign n24798 = n24797 ^ n2717 ;
  assign n24675 = n22733 ^ n2601 ;
  assign n24676 = n24675 ^ n3127 ;
  assign n24677 = n24676 ^ n1814 ;
  assign n24674 = n24673 ^ n24672 ;
  assign n24678 = n24677 ^ n24674 ;
  assign n24507 = n24506 ^ n3104 ;
  assign n24658 = n24507 & ~n24657 ;
  assign n24659 = n24658 ^ n3104 ;
  assign n24799 = n24674 ^ n24659 ;
  assign n24800 = n24678 & ~n24799 ;
  assign n24801 = n24800 ^ n24677 ;
  assign n24802 = n24801 ^ n24797 ;
  assign n24803 = n24798 & ~n24802 ;
  assign n24804 = n24803 ^ n2717 ;
  assign n24805 = n24804 ^ n2723 ;
  assign n24806 = ~n24796 & n24805 ;
  assign n24791 = n3010 ^ n2723 ;
  assign n24787 = n24773 ^ n24766 ;
  assign n24788 = ~n24771 & ~n24787 ;
  assign n24782 = n23531 ^ n21855 ;
  assign n24783 = n24782 ^ n22887 ;
  assign n24784 = n24783 ^ n24773 ;
  assign n24785 = n24784 ^ n24781 ;
  assign n24786 = n24785 ^ n21610 ;
  assign n24789 = n24788 ^ n24786 ;
  assign n24775 = n24774 ^ n24765 ;
  assign n24778 = n24765 ^ n24761 ;
  assign n24779 = ~n24775 & ~n24778 ;
  assign n24776 = n24775 ^ n24761 ;
  assign n24777 = ~n21271 & n24776 ;
  assign n24780 = n24779 ^ n24777 ;
  assign n24790 = n24789 ^ n24780 ;
  assign n24792 = n24791 ^ n24790 ;
  assign n24807 = n24806 ^ n24792 ;
  assign n24745 = n23579 ^ n22390 ;
  assign n24746 = n24745 ^ n24195 ;
  assign n24808 = n24807 ^ n24746 ;
  assign n24811 = n24804 ^ n24796 ;
  assign n24809 = n24130 ^ n22395 ;
  assign n24810 = n24809 ^ n23576 ;
  assign n24812 = n24811 ^ n24810 ;
  assign n24815 = n24801 ^ n24798 ;
  assign n24822 = n24815 ^ n24811 ;
  assign n24813 = n24206 ^ n23314 ;
  assign n24814 = n24813 ^ n22397 ;
  assign n24816 = n24815 ^ n24814 ;
  assign n24684 = n24208 ^ n22402 ;
  assign n24685 = n24684 ^ n23320 ;
  assign n24819 = n24815 ^ n24685 ;
  assign n24683 = ~n24681 & n24682 ;
  assign n24686 = n24685 ^ n24683 ;
  assign n24679 = n24678 ^ n24659 ;
  assign n24817 = n24685 ^ n24679 ;
  assign n24818 = n24686 & n24817 ;
  assign n24820 = n24819 ^ n24818 ;
  assign n24821 = ~n24816 & n24820 ;
  assign n24823 = n24822 ^ n24821 ;
  assign n24824 = ~n24812 & ~n24823 ;
  assign n24825 = n24824 ^ n24811 ;
  assign n24826 = n24825 ^ n24746 ;
  assign n24827 = n24808 & n24826 ;
  assign n24828 = n24827 ^ n24807 ;
  assign n24829 = n24828 ^ n24743 ;
  assign n24830 = n24744 & n24829 ;
  assign n24832 = n24831 ^ n24830 ;
  assign n24833 = n24740 & ~n24832 ;
  assign n24834 = n24833 ^ n24739 ;
  assign n24835 = n24834 ^ n24733 ;
  assign n24836 = ~n24736 & n24835 ;
  assign n24837 = n24836 ^ n24735 ;
  assign n24838 = n24837 ^ n24129 ;
  assign n24839 = n24732 & n24838 ;
  assign n24840 = n24839 ^ n24731 ;
  assign n24728 = n24724 ^ n24722 ;
  assign n24729 = n24728 ^ n24722 ;
  assign n24841 = n24840 ^ n24729 ;
  assign n24842 = ~n24727 & ~n24841 ;
  assign n24843 = n24842 ^ n24728 ;
  assign n24844 = n24723 & ~n24843 ;
  assign n24845 = n24844 ^ n24722 ;
  assign n24846 = n24845 ^ n24716 ;
  assign n24847 = ~n24719 & ~n24846 ;
  assign n24848 = n24847 ^ n24718 ;
  assign n24712 = n24160 ^ n23217 ;
  assign n24713 = n24712 ^ n23284 ;
  assign n24714 = n24713 ^ n24710 ;
  assign n24715 = n24714 ^ n24713 ;
  assign n24849 = n24848 ^ n24715 ;
  assign n24850 = ~n24711 & n24849 ;
  assign n24851 = n24850 ^ n24714 ;
  assign n24854 = n24713 ^ n24706 ;
  assign n24852 = n24582 ^ n24550 ;
  assign n24853 = n24852 ^ n24706 ;
  assign n24855 = n24854 ^ n24853 ;
  assign n24856 = n24851 & ~n24855 ;
  assign n24857 = n24856 ^ n24854 ;
  assign n24858 = n24707 & n24857 ;
  assign n24859 = n24858 ^ n24706 ;
  assign n25071 = n25070 ^ n24859 ;
  assign n25072 = n24863 & n25071 ;
  assign n25073 = n25072 ^ n25069 ;
  assign n25074 = n24595 ^ n24540 ;
  assign n25093 = n25074 ^ n25068 ;
  assign n25094 = n25073 & ~n25093 ;
  assign n25095 = n25094 ^ n25068 ;
  assign n25217 = n25095 ^ n25091 ;
  assign n25218 = ~n25092 & n25217 ;
  assign n25219 = n25218 ^ n25095 ;
  assign n25220 = n25219 ^ n25215 ;
  assign n25221 = n25216 & ~n25220 ;
  assign n25222 = n25221 ^ n25141 ;
  assign n25223 = n25222 ^ n25135 ;
  assign n25224 = ~n25211 & ~n25223 ;
  assign n25212 = n25135 ^ n25129 ;
  assign n25225 = n25224 ^ n25212 ;
  assign n25226 = ~n25208 & ~n25225 ;
  assign n25227 = n25226 ^ n25207 ;
  assign n25202 = n24063 ^ n23259 ;
  assign n25203 = n25202 ^ n24498 ;
  assign n25204 = n25203 ^ n25200 ;
  assign n25205 = n25204 ^ n25203 ;
  assign n25228 = n25227 ^ n25205 ;
  assign n25229 = ~n25201 & n25228 ;
  assign n25230 = n25229 ^ n25204 ;
  assign n25234 = n25232 ^ n25203 ;
  assign n25231 = n24619 ^ n24618 ;
  assign n25233 = n25232 ^ n25231 ;
  assign n25235 = n25234 ^ n25233 ;
  assign n25236 = ~n25230 & n25235 ;
  assign n25237 = n25236 ^ n25234 ;
  assign n25238 = n24106 ^ n23254 ;
  assign n25239 = n25238 ^ n24668 ;
  assign n25240 = n25239 ^ n25232 ;
  assign n25241 = n25237 & ~n25240 ;
  assign n25243 = n25242 ^ n25241 ;
  assign n25244 = n25197 & ~n25243 ;
  assign n25245 = n25244 ^ n25124 ;
  assign n25246 = n25245 ^ n25193 ;
  assign n25247 = n25194 & n25246 ;
  assign n25248 = n25247 ^ n25120 ;
  assign n25249 = n25248 ^ n25115 ;
  assign n25250 = n25191 & n25249 ;
  assign n25252 = n25251 ^ n25250 ;
  assign n25253 = n25188 & ~n25252 ;
  assign n25254 = n25253 ^ n25105 ;
  assign n25255 = n25254 ^ n25184 ;
  assign n25256 = n25185 & n25255 ;
  assign n25257 = n25256 ^ n25109 ;
  assign n25181 = n25180 ^ n25176 ;
  assign n25182 = n25181 ^ n25180 ;
  assign n25258 = n25257 ^ n25182 ;
  assign n25259 = n25179 & n25258 ;
  assign n25260 = n25259 ^ n25181 ;
  assign n25261 = n24122 ^ n23332 ;
  assign n25262 = n25261 ^ n22412 ;
  assign n25438 = n25262 ^ n25180 ;
  assign n25439 = n25260 & ~n25438 ;
  assign n25446 = n25445 ^ n25439 ;
  assign n25323 = n25254 ^ n25185 ;
  assign n25266 = n25245 ^ n25194 ;
  assign n25267 = n25266 ^ n22210 ;
  assign n25305 = n25243 ^ n25196 ;
  assign n25268 = n25239 ^ n25237 ;
  assign n25269 = n25268 ^ n22563 ;
  assign n25270 = n25231 ^ n25230 ;
  assign n25271 = n25270 ^ n22555 ;
  assign n25281 = n25222 ^ n25211 ;
  assign n25272 = n25219 ^ n25216 ;
  assign n25273 = n25272 ^ n22431 ;
  assign n25075 = n25074 ^ n25073 ;
  assign n24866 = n24857 ^ n24705 ;
  assign n24867 = n24866 ^ n22448 ;
  assign n24869 = n24848 ^ n24711 ;
  assign n24870 = n24869 ^ n21851 ;
  assign n24872 = n24837 ^ n24732 ;
  assign n24873 = n24872 ^ n22393 ;
  assign n24874 = n24834 ^ n24736 ;
  assign n24875 = n24874 ^ n22398 ;
  assign n24891 = n24825 ^ n24808 ;
  assign n24878 = n24823 ^ n24810 ;
  assign n24879 = n24878 ^ n22413 ;
  assign n24689 = ~n22273 & ~n24688 ;
  assign n24690 = n24689 ^ n22301 ;
  assign n24687 = n24686 ^ n24679 ;
  assign n24881 = n24689 ^ n24687 ;
  assign n24882 = n24690 & ~n24881 ;
  assign n24883 = n24882 ^ n22301 ;
  assign n24880 = n24820 ^ n24814 ;
  assign n24884 = n24883 ^ n24880 ;
  assign n24885 = n24883 ^ n22353 ;
  assign n24886 = n24884 & ~n24885 ;
  assign n24887 = n24886 ^ n22353 ;
  assign n24888 = n24887 ^ n24878 ;
  assign n24889 = ~n24879 & ~n24888 ;
  assign n24890 = n24889 ^ n22413 ;
  assign n24892 = n24891 ^ n24890 ;
  assign n24893 = n24891 ^ n22482 ;
  assign n24894 = n24892 & n24893 ;
  assign n24895 = n24894 ^ n22482 ;
  assign n24877 = n24828 ^ n24744 ;
  assign n24896 = n24895 ^ n24877 ;
  assign n24897 = n24895 ^ n22408 ;
  assign n24898 = n24896 & n24897 ;
  assign n24899 = n24898 ^ n22408 ;
  assign n24876 = n24832 ^ n24739 ;
  assign n24900 = n24899 ^ n24876 ;
  assign n24901 = n24874 ^ n22404 ;
  assign n24902 = n24901 ^ n24874 ;
  assign n24903 = n24902 ^ n24876 ;
  assign n24904 = n24900 & ~n24903 ;
  assign n24905 = n24904 ^ n24901 ;
  assign n24906 = n24875 & ~n24905 ;
  assign n24907 = n24906 ^ n22398 ;
  assign n24908 = n24907 ^ n24872 ;
  assign n24909 = n24873 & n24908 ;
  assign n24910 = n24909 ^ n22393 ;
  assign n24911 = n24910 ^ n22388 ;
  assign n24912 = n24840 ^ n24727 ;
  assign n24913 = n24912 ^ n24910 ;
  assign n24914 = ~n24911 & ~n24913 ;
  assign n24915 = n24914 ^ n22388 ;
  assign n24916 = n24915 ^ n22383 ;
  assign n24917 = n24843 ^ n24720 ;
  assign n24918 = n24917 ^ n24915 ;
  assign n24919 = ~n24916 & n24918 ;
  assign n24920 = n24919 ^ n22383 ;
  assign n24871 = n24845 ^ n24719 ;
  assign n24921 = n24920 ^ n24871 ;
  assign n24922 = n24920 ^ n22379 ;
  assign n24923 = ~n24921 & n24922 ;
  assign n24924 = n24923 ^ n22379 ;
  assign n24925 = n24924 ^ n24869 ;
  assign n24926 = ~n24870 & n24925 ;
  assign n24927 = n24926 ^ n21851 ;
  assign n24868 = n24852 ^ n24851 ;
  assign n24928 = n24927 ^ n24868 ;
  assign n24929 = n24927 ^ n22452 ;
  assign n24930 = n24928 & n24929 ;
  assign n24931 = n24930 ^ n22452 ;
  assign n24932 = n24931 ^ n24866 ;
  assign n24933 = ~n24867 & ~n24932 ;
  assign n24934 = n24933 ^ n22448 ;
  assign n24864 = n24863 ^ n24859 ;
  assign n25063 = n24934 ^ n24864 ;
  assign n25064 = n24934 ^ n22444 ;
  assign n25065 = n25063 & ~n25064 ;
  assign n25066 = n25065 ^ n22444 ;
  assign n25088 = n25075 ^ n25066 ;
  assign n25096 = n25095 ^ n25092 ;
  assign n25097 = n25096 ^ n22440 ;
  assign n25098 = n25097 ^ n25096 ;
  assign n25099 = n25098 ^ n25066 ;
  assign n25100 = n25088 & n25099 ;
  assign n25101 = n25100 ^ n25097 ;
  assign n25275 = n25272 ^ n22436 ;
  assign n25274 = n25272 ^ n25096 ;
  assign n25276 = n25275 ^ n25274 ;
  assign n25277 = ~n25101 & ~n25276 ;
  assign n25278 = n25277 ^ n25275 ;
  assign n25279 = n25273 & n25278 ;
  assign n25280 = n25279 ^ n22431 ;
  assign n25282 = n25281 ^ n25280 ;
  assign n25283 = n25225 ^ n25207 ;
  assign n25284 = n25283 ^ n22433 ;
  assign n25285 = n25284 ^ n25280 ;
  assign n25286 = n25285 ^ n25283 ;
  assign n25287 = n25282 & n25286 ;
  assign n25288 = n25287 ^ n25284 ;
  assign n25289 = n25227 ^ n25201 ;
  assign n25291 = n25289 ^ n22539 ;
  assign n25290 = n25289 ^ n25283 ;
  assign n25292 = n25291 ^ n25290 ;
  assign n25293 = ~n25288 & n25292 ;
  assign n25294 = n25293 ^ n25291 ;
  assign n25296 = n25270 ^ n22547 ;
  assign n25295 = n25289 ^ n25270 ;
  assign n25297 = n25296 ^ n25295 ;
  assign n25298 = n25294 & n25297 ;
  assign n25299 = n25298 ^ n25296 ;
  assign n25300 = n25271 & n25299 ;
  assign n25301 = n25300 ^ n22555 ;
  assign n25302 = n25301 ^ n25268 ;
  assign n25303 = n25269 & ~n25302 ;
  assign n25304 = n25303 ^ n22563 ;
  assign n25306 = n25305 ^ n25304 ;
  assign n25307 = n25305 ^ n22421 ;
  assign n25308 = n25306 & n25307 ;
  assign n25309 = n25308 ^ n22421 ;
  assign n25310 = n25309 ^ n25266 ;
  assign n25311 = ~n25267 & n25310 ;
  assign n25312 = n25311 ^ n22210 ;
  assign n25313 = n25312 ^ n22216 ;
  assign n25314 = n25248 ^ n25191 ;
  assign n25315 = n25314 ^ n25312 ;
  assign n25316 = n25313 & ~n25315 ;
  assign n25317 = n25316 ^ n22216 ;
  assign n25318 = n25317 ^ n22213 ;
  assign n25319 = n25252 ^ n25187 ;
  assign n25320 = n25319 ^ n25317 ;
  assign n25321 = n25318 & ~n25320 ;
  assign n25322 = n25321 ^ n22213 ;
  assign n25324 = n25323 ^ n25322 ;
  assign n25325 = n25323 ^ n22222 ;
  assign n25326 = n25324 & n25325 ;
  assign n25327 = n25326 ^ n22222 ;
  assign n25329 = n25327 ^ n22202 ;
  assign n25265 = n25257 ^ n25179 ;
  assign n25333 = n25329 ^ n25265 ;
  assign n25334 = n25325 ^ n25322 ;
  assign n25335 = n25319 ^ n25318 ;
  assign n25336 = n25314 ^ n25313 ;
  assign n25337 = n25299 ^ n22555 ;
  assign n25338 = n25280 ^ n22433 ;
  assign n25339 = n25338 ^ n25281 ;
  assign n25076 = n25075 ^ n22440 ;
  assign n25077 = n25076 ^ n25066 ;
  assign n24865 = n24864 ^ n22444 ;
  assign n24935 = n24934 ^ n24865 ;
  assign n24936 = n24912 ^ n24911 ;
  assign n24937 = n24905 ^ n22398 ;
  assign n24938 = n24876 ^ n22404 ;
  assign n24939 = n24938 ^ n24899 ;
  assign n24691 = n24690 ^ n24687 ;
  assign n24940 = n24691 & n24692 ;
  assign n24941 = n24880 ^ n22353 ;
  assign n24942 = n24941 ^ n24883 ;
  assign n24943 = n24940 & n24942 ;
  assign n24944 = n24887 ^ n22413 ;
  assign n24945 = n24944 ^ n24878 ;
  assign n24946 = n24943 & n24945 ;
  assign n24947 = n24893 ^ n24890 ;
  assign n24948 = n24946 & n24947 ;
  assign n24949 = n24896 ^ n22408 ;
  assign n24950 = ~n24948 & ~n24949 ;
  assign n24951 = n24939 & ~n24950 ;
  assign n24952 = n24937 & ~n24951 ;
  assign n24953 = n24907 ^ n24873 ;
  assign n24954 = n24952 & n24953 ;
  assign n24955 = n24936 & n24954 ;
  assign n24956 = n24917 ^ n24916 ;
  assign n24957 = ~n24955 & ~n24956 ;
  assign n24958 = n24871 ^ n22379 ;
  assign n24959 = n24958 ^ n24920 ;
  assign n24960 = ~n24957 & ~n24959 ;
  assign n24961 = n24924 ^ n21851 ;
  assign n24962 = n24961 ^ n24869 ;
  assign n24963 = ~n24960 & ~n24962 ;
  assign n24964 = n24868 ^ n22452 ;
  assign n24965 = n24964 ^ n24927 ;
  assign n24966 = ~n24963 & n24965 ;
  assign n24967 = n24931 ^ n24867 ;
  assign n24968 = n24966 & n24967 ;
  assign n25078 = n24935 & n24968 ;
  assign n25087 = n25077 & n25078 ;
  assign n25102 = n25101 ^ n22436 ;
  assign n25340 = ~n25087 & ~n25102 ;
  assign n25341 = n25278 ^ n22431 ;
  assign n25342 = n25340 & ~n25341 ;
  assign n25343 = n25339 & ~n25342 ;
  assign n25344 = n25288 ^ n22539 ;
  assign n25345 = n25343 & ~n25344 ;
  assign n25346 = n25294 ^ n22547 ;
  assign n25347 = ~n25345 & n25346 ;
  assign n25348 = n25337 & ~n25347 ;
  assign n25349 = n25301 ^ n25269 ;
  assign n25350 = n25348 & ~n25349 ;
  assign n25351 = n25307 ^ n25304 ;
  assign n25352 = ~n25350 & n25351 ;
  assign n25353 = n25309 ^ n25267 ;
  assign n25354 = ~n25352 & ~n25353 ;
  assign n25355 = n25336 & n25354 ;
  assign n25356 = n25335 & n25355 ;
  assign n25357 = ~n25334 & ~n25356 ;
  assign n25358 = ~n25333 & ~n25357 ;
  assign n25328 = n25327 ^ n25265 ;
  assign n25330 = n25328 & ~n25329 ;
  assign n25331 = n25330 ^ n22202 ;
  assign n25432 = n25358 ^ n25331 ;
  assign n25263 = n25262 ^ n25260 ;
  assign n25435 = n25358 ^ n25263 ;
  assign n25436 = ~n25432 & n25435 ;
  assign n25433 = n25432 ^ n25263 ;
  assign n25434 = n21856 & n25433 ;
  assign n25437 = n25436 ^ n25434 ;
  assign n25447 = n25446 ^ n25437 ;
  assign n25449 = n25448 ^ n25447 ;
  assign n25264 = n25263 ^ n21856 ;
  assign n25332 = n25331 ^ n25264 ;
  assign n25359 = n25358 ^ n25332 ;
  assign n25360 = n25359 ^ n3161 ;
  assign n25412 = n25355 ^ n25335 ;
  assign n25361 = n25354 ^ n25336 ;
  assign n2559 = n2558 ^ n2480 ;
  assign n2566 = n2565 ^ n2559 ;
  assign n2570 = n2569 ^ n2566 ;
  assign n25362 = n25361 ^ n2570 ;
  assign n25363 = n25353 ^ n25352 ;
  assign n25367 = n25366 ^ n25363 ;
  assign n25368 = n25351 ^ n25350 ;
  assign n25369 = n25368 ^ n2822 ;
  assign n25370 = n25349 ^ n25348 ;
  assign n25371 = n25370 ^ n2797 ;
  assign n25399 = n25370 ^ n1321 ;
  assign n1301 = n1204 ^ n1133 ;
  assign n1302 = n1301 ^ n1067 ;
  assign n1306 = n1305 ^ n1302 ;
  assign n25394 = n1321 ^ n1306 ;
  assign n25372 = n25346 ^ n25345 ;
  assign n25373 = n25372 ^ n1306 ;
  assign n25374 = n25344 ^ n25343 ;
  assign n1292 = n1195 ^ n1102 ;
  assign n1296 = n1295 ^ n1292 ;
  assign n1297 = n1296 ^ n1061 ;
  assign n25375 = n25374 ^ n1297 ;
  assign n25376 = n25342 ^ n25339 ;
  assign n926 = n925 ^ n842 ;
  assign n927 = n926 ^ n915 ;
  assign n928 = n927 ^ n896 ;
  assign n25377 = n25376 ^ n928 ;
  assign n25079 = n25078 ^ n25077 ;
  assign n25080 = n25079 ^ n709 ;
  assign n24969 = n24968 ^ n24935 ;
  assign n24970 = n24969 ^ n709 ;
  assign n24974 = n24967 ^ n24966 ;
  assign n24975 = n24974 ^ n24973 ;
  assign n24976 = n24965 ^ n24963 ;
  assign n24977 = n24976 ^ n1530 ;
  assign n24983 = n24962 ^ n24960 ;
  assign n25054 = n24983 ^ n1530 ;
  assign n24978 = n24959 ^ n24957 ;
  assign n24982 = n24981 ^ n24978 ;
  assign n24986 = n24956 ^ n24955 ;
  assign n2916 = n2915 ^ n2909 ;
  assign n2917 = n2916 ^ n590 ;
  assign n2921 = n2920 ^ n2917 ;
  assign n24987 = n24986 ^ n2921 ;
  assign n24988 = n24954 ^ n24936 ;
  assign n24992 = n24991 ^ n24988 ;
  assign n24993 = n24953 ^ n24952 ;
  assign n25039 = n24993 ^ n24991 ;
  assign n2365 = n2292 ^ n584 ;
  assign n2369 = n2368 ^ n2365 ;
  assign n2373 = n2372 ^ n2369 ;
  assign n24994 = n24993 ^ n2373 ;
  assign n24995 = n24950 ^ n24939 ;
  assign n2219 = n2209 ^ n2155 ;
  assign n2220 = n2219 ^ n2130 ;
  assign n2224 = n2223 ^ n2220 ;
  assign n24996 = n24995 ^ n2224 ;
  assign n25000 = n24949 ^ n24948 ;
  assign n2118 = n2090 ^ n2063 ;
  assign n2119 = n2118 ^ n2115 ;
  assign n2123 = n2122 ^ n2119 ;
  assign n25001 = n25000 ^ n2123 ;
  assign n25002 = n24947 ^ n24946 ;
  assign n2109 = n2051 ^ n2013 ;
  assign n2110 = n2109 ^ n2108 ;
  assign n2111 = n2110 ^ n2102 ;
  assign n25003 = n25002 ^ n2111 ;
  assign n25007 = n23096 ^ n2001 ;
  assign n25008 = n25007 ^ n19844 ;
  assign n25009 = n25008 ^ n2106 ;
  assign n25006 = n24945 ^ n24943 ;
  assign n25010 = n25009 ^ n25006 ;
  assign n25014 = n24942 ^ n24940 ;
  assign n24698 = n3074 ^ n3051 ;
  assign n24699 = n24698 ^ n1793 ;
  assign n24700 = n24699 ^ n14844 ;
  assign n24697 = ~n24692 & n24696 ;
  assign n24701 = n24700 ^ n24697 ;
  assign n24693 = n24692 ^ n24691 ;
  assign n25011 = n24700 ^ n24693 ;
  assign n25012 = n24701 & n25011 ;
  assign n25013 = n25012 ^ n24700 ;
  assign n25015 = n25014 ^ n25013 ;
  assign n25016 = n3080 ^ n1994 ;
  assign n25017 = n25016 ^ n19851 ;
  assign n25018 = n25017 ^ n1898 ;
  assign n25019 = n25018 ^ n25013 ;
  assign n25020 = n25015 & n25019 ;
  assign n25021 = n25020 ^ n25013 ;
  assign n25022 = n25021 ^ n25006 ;
  assign n25023 = n25010 & ~n25022 ;
  assign n25024 = n25023 ^ n25009 ;
  assign n25004 = n2123 ^ n2111 ;
  assign n25005 = n25004 ^ n2123 ;
  assign n25025 = n25024 ^ n25005 ;
  assign n25026 = n25003 & n25025 ;
  assign n25027 = n25026 ^ n25004 ;
  assign n25028 = ~n25001 & ~n25027 ;
  assign n25029 = n25028 ^ n25000 ;
  assign n24997 = n24951 ^ n24937 ;
  assign n24998 = n24997 ^ n2224 ;
  assign n24999 = n24998 ^ n24997 ;
  assign n25030 = n25029 ^ n24999 ;
  assign n25031 = ~n24996 & ~n25030 ;
  assign n25032 = n25031 ^ n24998 ;
  assign n2231 = n2215 ^ n2164 ;
  assign n2232 = n2231 ^ n2228 ;
  assign n2233 = n2232 ^ n1460 ;
  assign n25034 = n24993 ^ n2233 ;
  assign n25033 = n24997 ^ n24993 ;
  assign n25035 = n25034 ^ n25033 ;
  assign n25036 = n25032 & n25035 ;
  assign n25037 = n25036 ^ n25033 ;
  assign n25038 = ~n24994 & ~n25037 ;
  assign n25040 = n25039 ^ n25038 ;
  assign n25041 = ~n24992 & ~n25040 ;
  assign n25042 = n25041 ^ n24991 ;
  assign n25043 = n25042 ^ n2921 ;
  assign n25044 = n24987 & ~n25043 ;
  assign n25045 = n25044 ^ n24986 ;
  assign n24984 = n24983 ^ n24981 ;
  assign n24985 = n24984 ^ n24983 ;
  assign n25046 = n25045 ^ n24985 ;
  assign n25047 = ~n24982 & n25046 ;
  assign n25048 = n25047 ^ n24984 ;
  assign n25052 = n25051 ^ n24983 ;
  assign n25053 = n25048 & n25052 ;
  assign n25055 = n25054 ^ n25053 ;
  assign n25056 = n24977 & ~n25055 ;
  assign n25057 = n25056 ^ n24976 ;
  assign n25058 = n25057 ^ n24973 ;
  assign n25059 = ~n24975 & ~n25058 ;
  assign n25060 = n25059 ^ n24974 ;
  assign n25061 = n25060 ^ n709 ;
  assign n25062 = ~n24970 & ~n25061 ;
  assign n25081 = n25080 ^ n25062 ;
  assign n25082 = n25079 ^ n786 ;
  assign n25083 = n25082 ^ n721 ;
  assign n25084 = n25083 ^ n786 ;
  assign n25085 = ~n25081 & ~n25084 ;
  assign n25086 = n25085 ^ n25082 ;
  assign n25103 = n25102 ^ n25087 ;
  assign n25379 = n25103 ^ n786 ;
  assign n25380 = ~n25086 & n25379 ;
  assign n25381 = n25380 ^ n786 ;
  assign n25385 = n25381 ^ n928 ;
  assign n25378 = n25341 ^ n25340 ;
  assign n25382 = n25381 ^ n25378 ;
  assign n1684 = n1664 ^ n1110 ;
  assign n1685 = n1684 ^ n790 ;
  assign n1686 = n1685 ^ n912 ;
  assign n25383 = n25378 ^ n1686 ;
  assign n25384 = ~n25382 & n25383 ;
  assign n25386 = n25385 ^ n25384 ;
  assign n25387 = n25377 & n25386 ;
  assign n25388 = n25387 ^ n928 ;
  assign n25389 = n25388 ^ n1297 ;
  assign n25390 = n25375 & ~n25389 ;
  assign n25391 = n25390 ^ n25374 ;
  assign n25392 = n25391 ^ n1306 ;
  assign n25393 = ~n25373 & n25392 ;
  assign n25395 = n25394 ^ n25393 ;
  assign n25396 = n25347 ^ n25337 ;
  assign n25397 = n25396 ^ n1321 ;
  assign n25398 = n25395 & n25397 ;
  assign n25400 = n25399 ^ n25398 ;
  assign n25401 = n25371 & n25400 ;
  assign n25402 = n25401 ^ n25370 ;
  assign n25403 = n25402 ^ n25368 ;
  assign n25404 = ~n25369 & n25403 ;
  assign n25405 = n25404 ^ n2822 ;
  assign n25406 = n25405 ^ n25363 ;
  assign n25407 = ~n25367 & n25406 ;
  assign n25408 = n25407 ^ n25366 ;
  assign n25409 = n25408 ^ n25361 ;
  assign n25410 = ~n25362 & n25409 ;
  assign n25411 = n25410 ^ n2570 ;
  assign n25413 = n25412 ^ n25411 ;
  assign n25416 = n25411 ^ n3215 ;
  assign n25417 = n25413 & n25416 ;
  assign n25414 = n3215 ^ n2519 ;
  assign n25418 = n25417 ^ n25414 ;
  assign n25421 = n3168 ^ n2519 ;
  assign n25419 = n25356 ^ n25334 ;
  assign n25420 = n25419 ^ n3168 ;
  assign n25422 = n25421 ^ n25420 ;
  assign n25423 = n25418 & n25422 ;
  assign n25424 = n25423 ^ n25421 ;
  assign n25427 = n3168 ^ n3161 ;
  assign n25425 = n25357 ^ n25333 ;
  assign n25426 = n25425 ^ n3161 ;
  assign n25428 = n25427 ^ n25426 ;
  assign n25429 = n25424 & ~n25428 ;
  assign n25430 = n25429 ^ n25427 ;
  assign n25431 = ~n25360 & n25430 ;
  assign n25450 = n25449 ^ n25431 ;
  assign n25453 = n25452 ^ n25450 ;
  assign n25456 = n25430 ^ n25359 ;
  assign n25454 = n24193 ^ n24129 ;
  assign n25455 = n25454 ^ n23576 ;
  assign n25457 = n25456 ^ n25455 ;
  assign n25460 = n25425 ^ n25424 ;
  assign n25476 = n25460 ^ n25455 ;
  assign n25458 = n24195 ^ n23314 ;
  assign n25459 = n25458 ^ n24733 ;
  assign n25461 = n25460 ^ n25459 ;
  assign n25464 = n24743 ^ n24206 ;
  assign n25465 = n25464 ^ n23322 ;
  assign n25466 = n25412 ^ n3215 ;
  assign n25467 = n25466 ^ n25411 ;
  assign n25468 = n25465 & ~n25467 ;
  assign n25462 = n24739 ^ n23320 ;
  assign n25463 = n25462 ^ n24130 ;
  assign n25469 = n25468 ^ n25463 ;
  assign n25470 = n25419 ^ n25418 ;
  assign n25471 = n25470 ^ n25463 ;
  assign n25472 = n25469 & n25471 ;
  assign n25473 = n25472 ^ n25463 ;
  assign n25474 = n25473 ^ n25460 ;
  assign n25475 = ~n25461 & ~n25474 ;
  assign n25477 = n25476 ^ n25475 ;
  assign n25478 = ~n25457 & n25477 ;
  assign n25479 = n25478 ^ n25456 ;
  assign n25480 = n25479 ^ n25450 ;
  assign n25481 = n25453 & n25480 ;
  assign n25482 = n25481 ^ n25452 ;
  assign n25483 = n25482 ^ n25172 ;
  assign n25484 = ~n25175 & n25483 ;
  assign n25485 = n25484 ^ n25174 ;
  assign n25169 = n24716 ^ n23312 ;
  assign n25170 = n25169 ^ n24183 ;
  assign n24702 = n24701 ^ n24693 ;
  assign n25171 = n25170 ^ n24702 ;
  assign n25578 = n25485 ^ n25171 ;
  assign n25579 = n25578 ^ n22376 ;
  assign n25581 = n25479 ^ n25453 ;
  assign n25582 = n25581 ^ n22390 ;
  assign n25583 = n25477 ^ n25456 ;
  assign n25584 = n25583 ^ n22395 ;
  assign n25587 = n25467 ^ n25465 ;
  assign n25588 = ~n22410 & ~n25587 ;
  assign n25586 = n25470 ^ n25469 ;
  assign n25589 = n25588 ^ n25586 ;
  assign n25590 = n25588 ^ n22402 ;
  assign n25591 = ~n25589 & ~n25590 ;
  assign n25592 = n25591 ^ n22402 ;
  assign n25585 = n25473 ^ n25461 ;
  assign n25593 = n25592 ^ n25585 ;
  assign n25594 = n25583 ^ n22397 ;
  assign n25595 = n25594 ^ n25583 ;
  assign n25596 = n25595 ^ n25585 ;
  assign n25597 = ~n25593 & n25596 ;
  assign n25598 = n25597 ^ n25594 ;
  assign n25599 = n25584 & n25598 ;
  assign n25600 = n25599 ^ n22395 ;
  assign n25601 = n25600 ^ n25581 ;
  assign n25602 = ~n25582 & n25601 ;
  assign n25603 = n25602 ^ n22390 ;
  assign n25580 = n25482 ^ n25175 ;
  assign n25604 = n25603 ^ n25580 ;
  assign n25605 = n25578 ^ n22385 ;
  assign n25606 = n25605 ^ n25578 ;
  assign n25607 = n25606 ^ n25580 ;
  assign n25608 = n25604 & n25607 ;
  assign n25609 = n25608 ^ n25605 ;
  assign n25610 = ~n25579 & ~n25609 ;
  assign n25611 = n25610 ^ n22376 ;
  assign n25721 = n25611 ^ n22374 ;
  assign n25165 = n25018 ^ n25015 ;
  assign n25488 = n25165 ^ n24702 ;
  assign n25486 = n25485 ^ n24702 ;
  assign n25487 = ~n25171 & n25486 ;
  assign n25489 = n25488 ^ n25487 ;
  assign n25166 = n24710 ^ n23308 ;
  assign n25167 = n25166 ^ n24175 ;
  assign n25577 = n25489 ^ n25167 ;
  assign n25722 = n25721 ^ n25577 ;
  assign n25705 = n25598 ^ n22395 ;
  assign n25706 = n25585 ^ n22397 ;
  assign n25707 = n25706 ^ n25592 ;
  assign n25708 = n25590 ^ n25586 ;
  assign n25709 = n25587 ^ n22410 ;
  assign n25710 = ~n25708 & n25709 ;
  assign n25711 = ~n25707 & n25710 ;
  assign n25712 = ~n25705 & n25711 ;
  assign n25713 = n25600 ^ n22390 ;
  assign n25714 = n25713 ^ n25581 ;
  assign n25715 = n25712 & ~n25714 ;
  assign n25716 = n25603 ^ n22385 ;
  assign n25717 = n25716 ^ n25580 ;
  assign n25718 = ~n25715 & ~n25717 ;
  assign n25719 = n25609 ^ n22376 ;
  assign n25720 = ~n25718 & n25719 ;
  assign n25837 = n25722 ^ n25720 ;
  assign n25838 = n25837 ^ n2340 ;
  assign n25875 = n25719 ^ n25718 ;
  assign n25840 = n23898 ^ n2171 ;
  assign n25841 = n25840 ^ n2021 ;
  assign n25842 = n25841 ^ n2325 ;
  assign n25839 = n25717 ^ n25715 ;
  assign n25843 = n25842 ^ n25839 ;
  assign n25864 = n25714 ^ n25712 ;
  assign n25844 = n25711 ^ n25705 ;
  assign n1932 = n1931 ^ n1910 ;
  assign n1939 = n1938 ^ n1932 ;
  assign n1943 = n1942 ^ n1939 ;
  assign n25845 = n25844 ^ n1943 ;
  assign n25848 = n23907 ^ n16729 ;
  assign n25849 = n25848 ^ n1894 ;
  assign n25850 = n25849 ^ n1936 ;
  assign n25860 = n25850 ^ n1943 ;
  assign n25846 = n25709 ^ n25708 ;
  assign n1879 = n1875 ^ n1863 ;
  assign n1886 = n1885 ^ n1879 ;
  assign n1890 = n1889 ^ n1886 ;
  assign n25847 = n25846 ^ n1890 ;
  assign n25851 = n3002 & ~n25709 ;
  assign n25852 = n25851 ^ n25850 ;
  assign n25853 = n25852 ^ n1890 ;
  assign n25854 = n25853 ^ n25850 ;
  assign n25855 = n25847 & n25854 ;
  assign n25856 = n25855 ^ n25852 ;
  assign n25857 = n25710 ^ n25707 ;
  assign n25858 = n25857 ^ n25850 ;
  assign n25859 = n25856 & ~n25858 ;
  assign n25861 = n25860 ^ n25859 ;
  assign n25862 = ~n25845 & ~n25861 ;
  assign n25863 = n25862 ^ n25844 ;
  assign n25865 = n25864 ^ n25863 ;
  assign n25866 = n23902 ^ n2175 ;
  assign n25867 = n25866 ^ n20390 ;
  assign n25868 = n25867 ^ n2019 ;
  assign n25869 = n25868 ^ n25863 ;
  assign n25870 = ~n25865 & ~n25869 ;
  assign n25871 = n25870 ^ n25868 ;
  assign n25872 = n25871 ^ n25839 ;
  assign n25873 = ~n25843 & n25872 ;
  assign n25874 = n25873 ^ n25842 ;
  assign n25876 = n25875 ^ n25874 ;
  assign n2322 = n2249 ^ n2191 ;
  assign n2329 = n2328 ^ n2322 ;
  assign n2330 = n2329 ^ n2135 ;
  assign n25877 = n25874 ^ n2330 ;
  assign n25878 = n25876 & n25877 ;
  assign n25879 = n25878 ^ n2330 ;
  assign n25880 = n25879 ^ n2340 ;
  assign n25881 = n25838 & n25880 ;
  assign n25883 = n25882 ^ n25881 ;
  assign n25612 = n25611 ^ n25577 ;
  assign n25168 = n25167 ^ n25165 ;
  assign n25490 = ~n25168 & ~n25489 ;
  assign n25491 = n25490 ^ n25167 ;
  assign n25163 = n25021 ^ n25010 ;
  assign n25161 = n24173 ^ n23611 ;
  assign n25162 = n25161 ^ n24852 ;
  assign n25164 = n25163 ^ n25162 ;
  assign n25613 = n25491 ^ n25164 ;
  assign n25614 = n25613 ^ n22374 ;
  assign n25615 = n25614 ^ n25577 ;
  assign n25616 = n25615 ^ n25613 ;
  assign n25617 = n25612 & ~n25616 ;
  assign n25618 = n25617 ^ n25614 ;
  assign n25724 = n25618 ^ n22918 ;
  assign n25723 = ~n25720 & n25722 ;
  assign n25835 = n25724 ^ n25723 ;
  assign n26169 = n25883 ^ n25835 ;
  assign n25535 = n25055 ^ n24976 ;
  assign n26167 = n25535 ^ n25129 ;
  assign n26168 = n26167 ^ n24148 ;
  assign n26170 = n26169 ^ n26168 ;
  assign n26171 = n25135 ^ n24154 ;
  assign n25520 = n25051 ^ n25048 ;
  assign n26172 = n26171 ^ n25520 ;
  assign n26133 = n25879 ^ n25838 ;
  assign n26173 = n26172 ^ n26133 ;
  assign n26176 = n25876 ^ n2330 ;
  assign n26174 = n25141 ^ n24160 ;
  assign n25134 = n25045 ^ n24982 ;
  assign n26175 = n26174 ^ n25134 ;
  assign n26177 = n26176 ^ n26175 ;
  assign n26180 = n25871 ^ n25843 ;
  assign n25132 = n25042 ^ n24987 ;
  assign n26178 = n25132 ^ n24164 ;
  assign n26179 = n26178 ^ n25091 ;
  assign n26181 = n26180 ^ n26179 ;
  assign n26184 = n25868 ^ n25865 ;
  assign n26213 = n26184 ^ n26180 ;
  assign n26182 = n25074 ^ n24168 ;
  assign n25138 = n25040 ^ n24988 ;
  assign n26183 = n26182 ^ n25138 ;
  assign n26185 = n26184 ^ n26183 ;
  assign n26188 = n25861 ^ n25844 ;
  assign n26186 = n24860 ^ n24173 ;
  assign n25140 = n25037 ^ n2373 ;
  assign n26187 = n26186 ^ n25140 ;
  assign n26189 = n26188 ^ n26187 ;
  assign n26192 = n25857 ^ n25856 ;
  assign n25147 = n25032 ^ n2233 ;
  assign n26190 = n25147 ^ n24706 ;
  assign n26191 = n26190 ^ n24175 ;
  assign n26193 = n26192 ^ n26191 ;
  assign n26196 = n25851 ^ n1890 ;
  assign n26197 = n26196 ^ n25846 ;
  assign n26194 = n24852 ^ n24183 ;
  assign n25151 = n25029 ^ n24996 ;
  assign n26195 = n26194 ^ n25151 ;
  assign n26198 = n26197 ^ n26195 ;
  assign n26102 = n25709 ^ n3002 ;
  assign n26201 = n26197 ^ n26102 ;
  assign n25153 = n25027 ^ n25000 ;
  assign n26100 = n25153 ^ n24181 ;
  assign n26101 = n26100 ^ n24710 ;
  assign n26103 = n26102 ^ n26101 ;
  assign n26035 = n25405 ^ n25367 ;
  assign n26033 = n24214 ^ n23332 ;
  assign n26034 = n26033 ^ n24811 ;
  assign n26036 = n26035 ^ n26034 ;
  assign n25989 = n25402 ^ n25369 ;
  assign n25987 = n24238 ^ n23531 ;
  assign n25988 = n25987 ^ n24815 ;
  assign n25990 = n25989 ^ n25988 ;
  assign n25780 = n24076 ^ n23537 ;
  assign n25781 = n25780 ^ n24682 ;
  assign n25779 = n25396 ^ n25395 ;
  assign n25782 = n25781 ^ n25779 ;
  assign n25961 = n25400 ^ n2797 ;
  assign n25962 = n25961 ^ n25779 ;
  assign n25963 = n25962 ^ n25961 ;
  assign n25106 = n25105 ^ n24063 ;
  assign n25107 = n25106 ^ n24753 ;
  assign n25104 = n25103 ^ n25086 ;
  assign n25108 = n25107 ^ n25104 ;
  assign n25116 = n25115 ^ n24022 ;
  assign n25117 = n25116 ^ n24668 ;
  assign n25114 = n25081 ^ n721 ;
  assign n25118 = n25117 ^ n25114 ;
  assign n25121 = n25120 ^ n24498 ;
  assign n25122 = n25121 ^ n23647 ;
  assign n25119 = n25060 ^ n24970 ;
  assign n25123 = n25122 ^ n25119 ;
  assign n25127 = n25057 ^ n24975 ;
  assign n25541 = n25127 ^ n25119 ;
  assign n25125 = n25124 ^ n24433 ;
  assign n25126 = n25125 ^ n23248 ;
  assign n25128 = n25127 ^ n25126 ;
  assign n25528 = n25232 ^ n24306 ;
  assign n25529 = n25528 ^ n23256 ;
  assign n25538 = n25529 ^ n25126 ;
  assign n25130 = n25129 ^ n24142 ;
  assign n25131 = n25130 ^ n23272 ;
  assign n25133 = n25132 ^ n25131 ;
  assign n25136 = n25135 ^ n23277 ;
  assign n25137 = n25136 ^ n24146 ;
  assign n25139 = n25138 ^ n25137 ;
  assign n25142 = n24148 ^ n23284 ;
  assign n25143 = n25142 ^ n25141 ;
  assign n25144 = n25143 ^ n25140 ;
  assign n25145 = n25091 ^ n23289 ;
  assign n25146 = n25145 ^ n24154 ;
  assign n25148 = n25147 ^ n25146 ;
  assign n25503 = n25151 ^ n25146 ;
  assign n25149 = n24160 ^ n23291 ;
  assign n25150 = n25149 ^ n25074 ;
  assign n25152 = n25151 ^ n25150 ;
  assign n25154 = n24860 ^ n23300 ;
  assign n25155 = n25154 ^ n24164 ;
  assign n25156 = n25155 ^ n25153 ;
  assign n25157 = n25024 ^ n25003 ;
  assign n25497 = n25157 ^ n25153 ;
  assign n25158 = n24168 ^ n23304 ;
  assign n25159 = n25158 ^ n24706 ;
  assign n25160 = n25159 ^ n25157 ;
  assign n25492 = n25491 ^ n25162 ;
  assign n25493 = ~n25164 & ~n25492 ;
  assign n25494 = n25493 ^ n25163 ;
  assign n25495 = n25494 ^ n25157 ;
  assign n25496 = n25160 & n25495 ;
  assign n25498 = n25497 ^ n25496 ;
  assign n25499 = ~n25156 & n25498 ;
  assign n25500 = n25499 ^ n25155 ;
  assign n25501 = n25500 ^ n25151 ;
  assign n25502 = n25152 & n25501 ;
  assign n25504 = n25503 ^ n25502 ;
  assign n25505 = n25148 & ~n25504 ;
  assign n25506 = n25505 ^ n25147 ;
  assign n25507 = n25506 ^ n25140 ;
  assign n25508 = ~n25144 & ~n25507 ;
  assign n25509 = n25508 ^ n25140 ;
  assign n25510 = n25509 ^ n25138 ;
  assign n25511 = n25139 & ~n25510 ;
  assign n25512 = n25511 ^ n25138 ;
  assign n25515 = n25512 ^ n25131 ;
  assign n25516 = n25133 & ~n25515 ;
  assign n25513 = n25512 ^ n25134 ;
  assign n25517 = n25516 ^ n25513 ;
  assign n25522 = n25520 ^ n25134 ;
  assign n25518 = n25200 ^ n23266 ;
  assign n25519 = n25518 ^ n24138 ;
  assign n25521 = n25520 ^ n25519 ;
  assign n25523 = n25522 ^ n25521 ;
  assign n25524 = ~n25517 & ~n25523 ;
  assign n25525 = n25524 ^ n25522 ;
  assign n25531 = n25529 ^ n25520 ;
  assign n25526 = n25231 ^ n23261 ;
  assign n25527 = n25526 ^ n24134 ;
  assign n25530 = n25529 ^ n25527 ;
  assign n25532 = n25531 ^ n25530 ;
  assign n25533 = ~n25525 & ~n25532 ;
  assign n25534 = n25533 ^ n25531 ;
  assign n25536 = n25535 ^ n25529 ;
  assign n25537 = n25534 & n25536 ;
  assign n25539 = n25538 ^ n25537 ;
  assign n25540 = n25128 & n25539 ;
  assign n25542 = n25541 ^ n25540 ;
  assign n25543 = n25123 & n25542 ;
  assign n25544 = n25543 ^ n25122 ;
  assign n25545 = n25544 ^ n25114 ;
  assign n25546 = n25118 & n25545 ;
  assign n25547 = n25546 ^ n25117 ;
  assign n25110 = n25109 ^ n24766 ;
  assign n25111 = n25110 ^ n24106 ;
  assign n25112 = n25111 ^ n25104 ;
  assign n25113 = n25112 ^ n25111 ;
  assign n25548 = n25547 ^ n25113 ;
  assign n25549 = n25108 & n25548 ;
  assign n25550 = n25549 ^ n25112 ;
  assign n25554 = n25383 ^ n25381 ;
  assign n25551 = n25176 ^ n24227 ;
  assign n25552 = n25551 ^ n24781 ;
  assign n25555 = n25554 ^ n25552 ;
  assign n25553 = n25552 ^ n25111 ;
  assign n25556 = n25555 ^ n25553 ;
  assign n25557 = ~n25550 & ~n25556 ;
  assign n25558 = n25557 ^ n25553 ;
  assign n25687 = n24035 ^ n23547 ;
  assign n25688 = n25687 ^ n25180 ;
  assign n25559 = n25386 ^ n25376 ;
  assign n25690 = n25688 ^ n25559 ;
  assign n25689 = n25688 ^ n25552 ;
  assign n25691 = n25690 ^ n25689 ;
  assign n25692 = n25558 & n25691 ;
  assign n25693 = n25692 ^ n25689 ;
  assign n25760 = n25443 ^ n24030 ;
  assign n25761 = n25760 ^ n23550 ;
  assign n25694 = n25388 ^ n25375 ;
  assign n25763 = n25761 ^ n25694 ;
  assign n25762 = n25761 ^ n25688 ;
  assign n25764 = n25763 ^ n25762 ;
  assign n25765 = n25693 & n25764 ;
  assign n25766 = n25765 ^ n25762 ;
  assign n25767 = n25391 ^ n25373 ;
  assign n25776 = n25767 ^ n25761 ;
  assign n25777 = n25766 & ~n25776 ;
  assign n25778 = n25777 ^ n25761 ;
  assign n25964 = n25963 ^ n25778 ;
  assign n25965 = ~n25782 & n25964 ;
  assign n25966 = n25965 ^ n25962 ;
  assign n25967 = n24122 ^ n23533 ;
  assign n25968 = n25967 ^ n24679 ;
  assign n25984 = n25968 ^ n25961 ;
  assign n25985 = n25966 & n25984 ;
  assign n25986 = n25985 ^ n25961 ;
  assign n26030 = n25988 ^ n25986 ;
  assign n26031 = n25990 & n26030 ;
  assign n26032 = n26031 ^ n25989 ;
  assign n26037 = n26036 ^ n26032 ;
  assign n25969 = n25968 ^ n25966 ;
  assign n25970 = n25969 ^ n22854 ;
  assign n25561 = n25554 ^ n25550 ;
  assign n25562 = n25561 ^ n23254 ;
  assign n25564 = n25542 ^ n25122 ;
  assign n25565 = n25564 ^ n23270 ;
  assign n25566 = n25539 ^ n25127 ;
  assign n25567 = n25566 ^ n23275 ;
  assign n25570 = n25519 ^ n25517 ;
  assign n25571 = n25570 ^ n23294 ;
  assign n25649 = n25512 ^ n25133 ;
  assign n25572 = n25500 ^ n25152 ;
  assign n25573 = n25572 ^ n23169 ;
  assign n25575 = n25494 ^ n25160 ;
  assign n25576 = n25575 ^ n23003 ;
  assign n25620 = n25575 ^ n22918 ;
  assign n25619 = n25613 ^ n25575 ;
  assign n25621 = n25620 ^ n25619 ;
  assign n25622 = ~n25618 & ~n25621 ;
  assign n25623 = n25622 ^ n25620 ;
  assign n25624 = n25576 & n25623 ;
  assign n25625 = n25624 ^ n23003 ;
  assign n25574 = n25498 ^ n25155 ;
  assign n25626 = n25625 ^ n25574 ;
  assign n25627 = n25572 ^ n23015 ;
  assign n25628 = n25627 ^ n25572 ;
  assign n25629 = n25628 ^ n25574 ;
  assign n25630 = n25626 & n25629 ;
  assign n25631 = n25630 ^ n25627 ;
  assign n25632 = ~n25573 & n25631 ;
  assign n25633 = n25632 ^ n23169 ;
  assign n25634 = n25633 ^ n23197 ;
  assign n25635 = n25504 ^ n25147 ;
  assign n25636 = n25635 ^ n25633 ;
  assign n25637 = n25634 & n25636 ;
  assign n25638 = n25637 ^ n23197 ;
  assign n25639 = n25638 ^ n23217 ;
  assign n25640 = n25506 ^ n25144 ;
  assign n25641 = n25640 ^ n25638 ;
  assign n25642 = n25639 & ~n25641 ;
  assign n25643 = n25642 ^ n23217 ;
  assign n25644 = n25643 ^ n23232 ;
  assign n25645 = n25509 ^ n25139 ;
  assign n25646 = n25645 ^ n25643 ;
  assign n25647 = ~n25644 & ~n25646 ;
  assign n25648 = n25647 ^ n23232 ;
  assign n25650 = n25649 ^ n25648 ;
  assign n25651 = n25570 ^ n23298 ;
  assign n25652 = n25651 ^ n25570 ;
  assign n25653 = n25652 ^ n25648 ;
  assign n25654 = n25650 & n25653 ;
  assign n25655 = n25654 ^ n25651 ;
  assign n25656 = ~n25571 & n25655 ;
  assign n25657 = n25656 ^ n23294 ;
  assign n25569 = n25527 ^ n25525 ;
  assign n25658 = n25657 ^ n25569 ;
  assign n25659 = n25657 ^ n23287 ;
  assign n25660 = ~n25658 & n25659 ;
  assign n25661 = n25660 ^ n23287 ;
  assign n25568 = n25535 ^ n25534 ;
  assign n25662 = n25661 ^ n25568 ;
  assign n25663 = n25661 ^ n23282 ;
  assign n25664 = ~n25662 & ~n25663 ;
  assign n25665 = n25664 ^ n23282 ;
  assign n25666 = n25665 ^ n25566 ;
  assign n25667 = n25567 & n25666 ;
  assign n25668 = n25667 ^ n23275 ;
  assign n25669 = n25668 ^ n25564 ;
  assign n25670 = n25565 & n25669 ;
  assign n25671 = n25670 ^ n23270 ;
  assign n25563 = n25544 ^ n25118 ;
  assign n25672 = n25671 ^ n25563 ;
  assign n25673 = n25547 ^ n25108 ;
  assign n25674 = n25673 ^ n23264 ;
  assign n25675 = n25674 ^ n25563 ;
  assign n25676 = n25675 ^ n25673 ;
  assign n25677 = n25672 & ~n25676 ;
  assign n25678 = n25677 ^ n25674 ;
  assign n25680 = n25561 ^ n23259 ;
  assign n25679 = n25673 ^ n25561 ;
  assign n25681 = n25680 ^ n25679 ;
  assign n25682 = ~n25678 & n25681 ;
  assign n25683 = n25682 ^ n25680 ;
  assign n25684 = ~n25562 & n25683 ;
  assign n25685 = n25684 ^ n23254 ;
  assign n25560 = n25559 ^ n25558 ;
  assign n25686 = n25685 ^ n25560 ;
  assign n25695 = n25694 ^ n25693 ;
  assign n25696 = n25695 ^ n23250 ;
  assign n25697 = n25696 ^ n25560 ;
  assign n25698 = n25697 ^ n25695 ;
  assign n25699 = n25686 & ~n25698 ;
  assign n25700 = n25699 ^ n25696 ;
  assign n25768 = n25767 ^ n25766 ;
  assign n25770 = n25768 ^ n22866 ;
  assign n25769 = n25768 ^ n25695 ;
  assign n25771 = n25770 ^ n25769 ;
  assign n25772 = n25700 & ~n25771 ;
  assign n25773 = n25772 ^ n25770 ;
  assign n25785 = n25768 ^ n22872 ;
  assign n25786 = ~n25773 & n25785 ;
  assign n25787 = n25786 ^ n22872 ;
  assign n25783 = n25782 ^ n25778 ;
  assign n25957 = n25787 ^ n25783 ;
  assign n25958 = n25787 ^ n22862 ;
  assign n25959 = ~n25957 & n25958 ;
  assign n25960 = n25959 ^ n22862 ;
  assign n25993 = n25969 ^ n25960 ;
  assign n25994 = ~n25970 & n25993 ;
  assign n25995 = n25994 ^ n22854 ;
  assign n25991 = n25990 ^ n25986 ;
  assign n26025 = n25995 ^ n25991 ;
  assign n26026 = n25995 ^ n22852 ;
  assign n26027 = n26025 & ~n26026 ;
  assign n26028 = n26027 ^ n22852 ;
  assign n26029 = n26028 ^ n22412 ;
  assign n26038 = n26037 ^ n26029 ;
  assign n25992 = n25991 ^ n22852 ;
  assign n25996 = n25995 ^ n25992 ;
  assign n25971 = n25970 ^ n25960 ;
  assign n25701 = n25700 ^ n22866 ;
  assign n25702 = n25574 ^ n23015 ;
  assign n25703 = n25702 ^ n25625 ;
  assign n25704 = n25623 ^ n23003 ;
  assign n25725 = n25723 & n25724 ;
  assign n25726 = n25704 & n25725 ;
  assign n25727 = n25703 & ~n25726 ;
  assign n25728 = n25631 ^ n23169 ;
  assign n25729 = ~n25727 & ~n25728 ;
  assign n25730 = n25635 ^ n25634 ;
  assign n25731 = ~n25729 & n25730 ;
  assign n25732 = n25640 ^ n25639 ;
  assign n25733 = ~n25731 & n25732 ;
  assign n25734 = n25645 ^ n25644 ;
  assign n25735 = n25733 & ~n25734 ;
  assign n25736 = n25648 ^ n23298 ;
  assign n25737 = n25736 ^ n25649 ;
  assign n25738 = n25735 & n25737 ;
  assign n25739 = n25655 ^ n23294 ;
  assign n25740 = n25738 & n25739 ;
  assign n25741 = n25659 ^ n25569 ;
  assign n25742 = ~n25740 & n25741 ;
  assign n25743 = n25663 ^ n25568 ;
  assign n25744 = n25742 & ~n25743 ;
  assign n25745 = n25665 ^ n25567 ;
  assign n25746 = ~n25744 & n25745 ;
  assign n25747 = n25668 ^ n25565 ;
  assign n25748 = n25746 & ~n25747 ;
  assign n25749 = n25563 ^ n23264 ;
  assign n25750 = n25749 ^ n25671 ;
  assign n25751 = ~n25748 & n25750 ;
  assign n25752 = n25678 ^ n23259 ;
  assign n25753 = ~n25751 & n25752 ;
  assign n25754 = n25683 ^ n23254 ;
  assign n25755 = n25753 & ~n25754 ;
  assign n25756 = n25560 ^ n23250 ;
  assign n25757 = n25756 ^ n25685 ;
  assign n25758 = ~n25755 & n25757 ;
  assign n25759 = ~n25701 & ~n25758 ;
  assign n25774 = n25773 ^ n22872 ;
  assign n25775 = n25759 & n25774 ;
  assign n25784 = n25783 ^ n22862 ;
  assign n25788 = n25787 ^ n25784 ;
  assign n25972 = n25775 & n25788 ;
  assign n25997 = n25971 & ~n25972 ;
  assign n26039 = n25996 & ~n25997 ;
  assign n26079 = ~n26038 & n26039 ;
  assign n26073 = n22887 ^ n22412 ;
  assign n26069 = n24807 ^ n24208 ;
  assign n26070 = n26069 ^ n23328 ;
  assign n26071 = n26070 ^ n26034 ;
  assign n26068 = n25408 ^ n25362 ;
  assign n26072 = n26071 ^ n26068 ;
  assign n26074 = n26073 ^ n26072 ;
  assign n26075 = n26074 ^ n2703 ;
  assign n26076 = n26075 ^ n3200 ;
  assign n26065 = n26037 ^ n26028 ;
  assign n26066 = n26037 ^ n22412 ;
  assign n26067 = n26065 & n26066 ;
  assign n26077 = n26076 ^ n26067 ;
  assign n26063 = n26034 ^ n26032 ;
  assign n26064 = n26036 & n26063 ;
  assign n26078 = n26077 ^ n26064 ;
  assign n26080 = n26079 ^ n26078 ;
  assign n25998 = n25997 ^ n25996 ;
  assign n25999 = n25998 ^ n2636 ;
  assign n26040 = n26039 ^ n26038 ;
  assign n26041 = n26040 ^ n2636 ;
  assign n25973 = n25972 ^ n25971 ;
  assign n2602 = n2592 ^ n2496 ;
  assign n2606 = n2605 ^ n2602 ;
  assign n2607 = n2606 ^ n2601 ;
  assign n25974 = n25973 ^ n2607 ;
  assign n25947 = n24002 ^ n2581 ;
  assign n25948 = n25947 ^ n20871 ;
  assign n25949 = n25948 ^ n1832 ;
  assign n3111 = n3110 ^ n2575 ;
  assign n3112 = n3111 ^ n2901 ;
  assign n3116 = n3115 ^ n3112 ;
  assign n25950 = n25949 ^ n3116 ;
  assign n25790 = n25774 ^ n25759 ;
  assign n25791 = n25790 ^ n3116 ;
  assign n25792 = n25758 ^ n25701 ;
  assign n2889 = n2866 ^ n2849 ;
  assign n2890 = n2889 ^ n2886 ;
  assign n2894 = n2893 ^ n2890 ;
  assign n25793 = n25792 ^ n2894 ;
  assign n25794 = n25757 ^ n25755 ;
  assign n25795 = n25794 ^ n2882 ;
  assign n25921 = n25750 ^ n25748 ;
  assign n25796 = n25747 ^ n25746 ;
  assign n998 = n968 ^ n908 ;
  assign n999 = n998 ^ n995 ;
  assign n1003 = n1002 ^ n999 ;
  assign n25797 = n25796 ^ n1003 ;
  assign n25798 = n25745 ^ n25744 ;
  assign n25799 = n25798 ^ n991 ;
  assign n25802 = n25743 ^ n25742 ;
  assign n25914 = n25802 ^ n25798 ;
  assign n25800 = n25741 ^ n25740 ;
  assign n25801 = n25800 ^ n872 ;
  assign n25805 = n25739 ^ n25738 ;
  assign n25806 = n25805 ^ n1594 ;
  assign n25807 = n25737 ^ n25735 ;
  assign n25808 = n25807 ^ n1585 ;
  assign n25809 = n25734 ^ n25733 ;
  assign n25810 = n25809 ^ n2960 ;
  assign n25811 = n25732 ^ n25731 ;
  assign n25815 = n25814 ^ n25811 ;
  assign n25816 = n25730 ^ n25729 ;
  assign n25817 = n25816 ^ n599 ;
  assign n25820 = n25728 ^ n25727 ;
  assign n25824 = n25823 ^ n25820 ;
  assign n25828 = n25726 ^ n25703 ;
  assign n25891 = n25828 ^ n25820 ;
  assign n25829 = n25828 ^ n25827 ;
  assign n25888 = n25832 ^ n25828 ;
  assign n25833 = n25725 ^ n25704 ;
  assign n25834 = n25833 ^ n25832 ;
  assign n25836 = n25835 ^ n2356 ;
  assign n25884 = ~n25836 & n25883 ;
  assign n25885 = n25884 ^ n2356 ;
  assign n25886 = n25885 ^ n25832 ;
  assign n25887 = ~n25834 & n25886 ;
  assign n25889 = n25888 ^ n25887 ;
  assign n25890 = ~n25829 & ~n25889 ;
  assign n25892 = n25891 ^ n25890 ;
  assign n25893 = ~n25824 & ~n25892 ;
  assign n25894 = n25893 ^ n25823 ;
  assign n25895 = n25894 ^ n599 ;
  assign n25896 = ~n25817 & n25895 ;
  assign n25818 = n25814 ^ n599 ;
  assign n25897 = n25896 ^ n25818 ;
  assign n25898 = n25815 & n25897 ;
  assign n25899 = n25898 ^ n25814 ;
  assign n25900 = n25899 ^ n2960 ;
  assign n25901 = n25810 & ~n25900 ;
  assign n25902 = n25901 ^ n25809 ;
  assign n25903 = n25902 ^ n1585 ;
  assign n25904 = ~n25808 & ~n25903 ;
  assign n25905 = n25904 ^ n25807 ;
  assign n25906 = n25905 ^ n1594 ;
  assign n25907 = ~n25806 & n25906 ;
  assign n25908 = n25907 ^ n25805 ;
  assign n25803 = n25802 ^ n872 ;
  assign n25804 = n25803 ^ n25802 ;
  assign n25909 = n25908 ^ n25804 ;
  assign n25910 = ~n25801 & ~n25909 ;
  assign n25911 = n25910 ^ n25803 ;
  assign n25912 = n25802 ^ n884 ;
  assign n25913 = ~n25911 & ~n25912 ;
  assign n25915 = n25914 ^ n25913 ;
  assign n25916 = n25799 & ~n25915 ;
  assign n25917 = n25916 ^ n25798 ;
  assign n25918 = n25917 ^ n1003 ;
  assign n25919 = n25797 & ~n25918 ;
  assign n25920 = n25919 ^ n25796 ;
  assign n25922 = n25921 ^ n25920 ;
  assign n25923 = n25752 ^ n25751 ;
  assign n25924 = n25923 ^ n1151 ;
  assign n25925 = n25924 ^ n25923 ;
  assign n25926 = n25925 ^ n25920 ;
  assign n25927 = n25922 & n25926 ;
  assign n25928 = n25927 ^ n25924 ;
  assign n25929 = n25754 ^ n25753 ;
  assign n1763 = n1738 ^ n1409 ;
  assign n1764 = n1763 ^ n1142 ;
  assign n1765 = n1764 ^ n1343 ;
  assign n25931 = n25929 ^ n1765 ;
  assign n25930 = n25929 ^ n25923 ;
  assign n25932 = n25931 ^ n25930 ;
  assign n25933 = n25928 & n25932 ;
  assign n25934 = n25933 ^ n25930 ;
  assign n25936 = n25929 ^ n25794 ;
  assign n1383 = n1382 ^ n1259 ;
  assign n1384 = n1383 ^ n1349 ;
  assign n1385 = n1384 ^ n1376 ;
  assign n25935 = n25794 ^ n1385 ;
  assign n25937 = n25936 ^ n25935 ;
  assign n25938 = ~n25934 & n25937 ;
  assign n25939 = n25938 ^ n25935 ;
  assign n25940 = ~n25795 & n25939 ;
  assign n25941 = n25940 ^ n2882 ;
  assign n25942 = n25941 ^ n2894 ;
  assign n25943 = ~n25793 & ~n25942 ;
  assign n25944 = n25943 ^ n25792 ;
  assign n25945 = n25944 ^ n3116 ;
  assign n25946 = ~n25791 & ~n25945 ;
  assign n25951 = n25950 ^ n25946 ;
  assign n25789 = n25788 ^ n25775 ;
  assign n25975 = n25949 ^ n25789 ;
  assign n25976 = n25951 & ~n25975 ;
  assign n25977 = n25976 ^ n25949 ;
  assign n26000 = n25977 ^ n2607 ;
  assign n26001 = ~n25974 & n26000 ;
  assign n26002 = n26001 ^ n2607 ;
  assign n26042 = n26041 ^ n26002 ;
  assign n26043 = n26042 ^ n26040 ;
  assign n26044 = n25999 & n26043 ;
  assign n26045 = n26044 ^ n26041 ;
  assign n26061 = n26040 ^ n2703 ;
  assign n26062 = ~n26045 & n26061 ;
  assign n26081 = n26080 ^ n26062 ;
  assign n26059 = n25157 ^ n24716 ;
  assign n26060 = n26059 ^ n24188 ;
  assign n26082 = n26081 ^ n26060 ;
  assign n26003 = n26002 ^ n25999 ;
  assign n25982 = n25165 ^ n24724 ;
  assign n25983 = n25982 ^ n24195 ;
  assign n26004 = n26003 ^ n25983 ;
  assign n26018 = n25163 ^ n24193 ;
  assign n26019 = n26018 ^ n24720 ;
  assign n26020 = n26019 ^ n26003 ;
  assign n26021 = n26020 ^ n26019 ;
  assign n25952 = n25951 ^ n25789 ;
  assign n25953 = n25172 ^ n24733 ;
  assign n25954 = n25953 ^ n24206 ;
  assign n25955 = ~n25952 & ~n25954 ;
  assign n24131 = n24130 ^ n24129 ;
  assign n24703 = n24702 ^ n24131 ;
  assign n25956 = n25955 ^ n24703 ;
  assign n25978 = n25977 ^ n25974 ;
  assign n25979 = n25978 ^ n25955 ;
  assign n25980 = ~n25956 & ~n25979 ;
  assign n25981 = n25980 ^ n25978 ;
  assign n26022 = n26021 ^ n25981 ;
  assign n26023 = n26004 & ~n26022 ;
  assign n26024 = n26023 ^ n26020 ;
  assign n26046 = n26045 ^ n2703 ;
  assign n26056 = n26046 ^ n26019 ;
  assign n26057 = ~n26024 & ~n26056 ;
  assign n26058 = n26057 ^ n26019 ;
  assign n26097 = n26060 ^ n26058 ;
  assign n26098 = ~n26082 & ~n26097 ;
  assign n26099 = n26098 ^ n26081 ;
  assign n26199 = n26102 ^ n26099 ;
  assign n26200 = n26103 & ~n26199 ;
  assign n26202 = n26201 ^ n26200 ;
  assign n26203 = n26198 & n26202 ;
  assign n26204 = n26203 ^ n26197 ;
  assign n26205 = n26204 ^ n26191 ;
  assign n26206 = n26193 & ~n26205 ;
  assign n26207 = n26206 ^ n26192 ;
  assign n26208 = n26207 ^ n26187 ;
  assign n26209 = n26189 & ~n26208 ;
  assign n26210 = n26209 ^ n26188 ;
  assign n26211 = n26210 ^ n26183 ;
  assign n26212 = ~n26185 & ~n26211 ;
  assign n26214 = n26213 ^ n26212 ;
  assign n26215 = ~n26181 & ~n26214 ;
  assign n26216 = n26215 ^ n26180 ;
  assign n26217 = n26216 ^ n26175 ;
  assign n26218 = n26177 & ~n26217 ;
  assign n26219 = n26218 ^ n26176 ;
  assign n26220 = n26219 ^ n26172 ;
  assign n26221 = ~n26173 & ~n26220 ;
  assign n26222 = n26221 ^ n26133 ;
  assign n26223 = n26222 ^ n26168 ;
  assign n26224 = ~n26170 & ~n26223 ;
  assign n26225 = n26224 ^ n26169 ;
  assign n26165 = n25885 ^ n25834 ;
  assign n26163 = n25200 ^ n24146 ;
  assign n26164 = n26163 ^ n25127 ;
  assign n26166 = n26165 ^ n26164 ;
  assign n26269 = n26225 ^ n26166 ;
  assign n26270 = n26269 ^ n23277 ;
  assign n26271 = n26222 ^ n26170 ;
  assign n26272 = n26271 ^ n23284 ;
  assign n26273 = n26219 ^ n26173 ;
  assign n26274 = n26273 ^ n23289 ;
  assign n26275 = n26214 ^ n26179 ;
  assign n26276 = n26275 ^ n23300 ;
  assign n26279 = n26204 ^ n26193 ;
  assign n26280 = n26279 ^ n23308 ;
  assign n26285 = n26202 ^ n26195 ;
  assign n26104 = n26103 ^ n26099 ;
  assign n26005 = n26004 ^ n25981 ;
  assign n26006 = n26005 ^ n23314 ;
  assign n26009 = n25978 ^ n25956 ;
  assign n26007 = n25954 ^ n25952 ;
  assign n26008 = ~n23322 & n26007 ;
  assign n26010 = n26009 ^ n26008 ;
  assign n26011 = n26009 ^ n23320 ;
  assign n26012 = n26010 & n26011 ;
  assign n26013 = n26012 ^ n23320 ;
  assign n26014 = n26013 ^ n26005 ;
  assign n26015 = n26006 & ~n26014 ;
  assign n26016 = n26015 ^ n23314 ;
  assign n26017 = n26016 ^ n23576 ;
  assign n26047 = n26046 ^ n26024 ;
  assign n26085 = n26047 ^ n26016 ;
  assign n26086 = n26017 & ~n26085 ;
  assign n26087 = n26086 ^ n23576 ;
  assign n26083 = n26082 ^ n26058 ;
  assign n26092 = n26087 ^ n26083 ;
  assign n26093 = n26087 ^ n23579 ;
  assign n26094 = n26092 & ~n26093 ;
  assign n26095 = n26094 ^ n23579 ;
  assign n26281 = n26104 ^ n26095 ;
  assign n26282 = n26104 ^ n23597 ;
  assign n26283 = ~n26281 & ~n26282 ;
  assign n26284 = n26283 ^ n23597 ;
  assign n26286 = n26285 ^ n26284 ;
  assign n26287 = n26285 ^ n23312 ;
  assign n26288 = ~n26286 & ~n26287 ;
  assign n26289 = n26288 ^ n23312 ;
  assign n26290 = n26289 ^ n26279 ;
  assign n26291 = ~n26280 & n26290 ;
  assign n26292 = n26291 ^ n23308 ;
  assign n26278 = n26207 ^ n26189 ;
  assign n26293 = n26292 ^ n26278 ;
  assign n26294 = n26292 ^ n23611 ;
  assign n26295 = n26293 & n26294 ;
  assign n26296 = n26295 ^ n23611 ;
  assign n26277 = n26210 ^ n26185 ;
  assign n26297 = n26296 ^ n26277 ;
  assign n26366 = n26277 ^ n23304 ;
  assign n26301 = ~n26297 & n26366 ;
  assign n26298 = n26275 ^ n23304 ;
  assign n26302 = n26301 ^ n26298 ;
  assign n26303 = ~n26276 & n26302 ;
  assign n26304 = n26303 ^ n23300 ;
  assign n26305 = n26304 ^ n23291 ;
  assign n26306 = n26216 ^ n26177 ;
  assign n26307 = n26306 ^ n26304 ;
  assign n26308 = ~n26305 & n26307 ;
  assign n26309 = n26308 ^ n23291 ;
  assign n26310 = n26309 ^ n26273 ;
  assign n26311 = n26274 & n26310 ;
  assign n26312 = n26311 ^ n23289 ;
  assign n26313 = n26312 ^ n26271 ;
  assign n26314 = n26272 & n26313 ;
  assign n26315 = n26314 ^ n23284 ;
  assign n26316 = n26315 ^ n26269 ;
  assign n26317 = n26270 & n26316 ;
  assign n26318 = n26317 ^ n23277 ;
  assign n26159 = n25231 ^ n25119 ;
  assign n26160 = n26159 ^ n24142 ;
  assign n26228 = n26165 ^ n26160 ;
  assign n26226 = n26225 ^ n26165 ;
  assign n26227 = ~n26166 & n26226 ;
  assign n26229 = n26228 ^ n26227 ;
  assign n26161 = n25889 ^ n25827 ;
  assign n26267 = n26229 ^ n26161 ;
  assign n26268 = n26267 ^ n23272 ;
  assign n26378 = n26318 ^ n26268 ;
  assign n26356 = n26306 ^ n26305 ;
  assign n26357 = n26302 ^ n23300 ;
  assign n26358 = n26284 ^ n23312 ;
  assign n26359 = n26358 ^ n26285 ;
  assign n26048 = n26047 ^ n26017 ;
  assign n26049 = n26013 ^ n26006 ;
  assign n26050 = n26007 ^ n23322 ;
  assign n26051 = n26008 ^ n23320 ;
  assign n26052 = n26051 ^ n26009 ;
  assign n26053 = ~n26050 & n26052 ;
  assign n26054 = ~n26049 & n26053 ;
  assign n26055 = ~n26048 & n26054 ;
  assign n26084 = n26083 ^ n23579 ;
  assign n26088 = n26087 ^ n26084 ;
  assign n26091 = n26055 & ~n26088 ;
  assign n26096 = n26095 ^ n23597 ;
  assign n26105 = n26104 ^ n26096 ;
  assign n26360 = ~n26091 & n26105 ;
  assign n26361 = n26359 & ~n26360 ;
  assign n26362 = n26289 ^ n26280 ;
  assign n26363 = ~n26361 & n26362 ;
  assign n26364 = n26294 ^ n26278 ;
  assign n26365 = n26363 & n26364 ;
  assign n26367 = n26366 ^ n26296 ;
  assign n26368 = n26365 & ~n26367 ;
  assign n26369 = ~n26357 & ~n26368 ;
  assign n26370 = ~n26356 & ~n26369 ;
  assign n26371 = n26309 ^ n26274 ;
  assign n26372 = ~n26370 & ~n26371 ;
  assign n26373 = n26312 ^ n26272 ;
  assign n26374 = ~n26372 & ~n26373 ;
  assign n26375 = n26315 ^ n23277 ;
  assign n26376 = n26375 ^ n26269 ;
  assign n26377 = n26374 & n26376 ;
  assign n26539 = n26378 ^ n26377 ;
  assign n26468 = n26376 ^ n26374 ;
  assign n26469 = n26468 ^ n633 ;
  assign n26535 = n26525 ^ n26468 ;
  assign n26473 = n26368 ^ n26357 ;
  assign n26470 = n24589 ^ n1473 ;
  assign n26471 = n26470 ^ n21165 ;
  assign n26472 = n26471 ^ n2909 ;
  assign n26474 = n26473 ^ n26472 ;
  assign n26479 = n24549 ^ n2436 ;
  assign n26480 = n26479 ^ n2363 ;
  assign n26481 = n26480 ^ n16155 ;
  assign n26478 = n26367 ^ n26365 ;
  assign n26482 = n26481 ^ n26478 ;
  assign n26483 = n26364 ^ n26363 ;
  assign n26487 = n26486 ^ n26483 ;
  assign n2205 = n2204 ^ n2147 ;
  assign n2212 = n2211 ^ n2205 ;
  assign n2216 = n2215 ^ n2212 ;
  assign n26505 = n26486 ^ n2216 ;
  assign n26089 = n26088 ^ n26055 ;
  assign n2009 = n1987 ^ n1969 ;
  assign n2010 = n2009 ^ n2006 ;
  assign n2014 = n2013 ^ n2010 ;
  assign n26090 = n26089 ^ n2014 ;
  assign n26107 = n26054 ^ n26048 ;
  assign n1991 = n1981 ^ n1957 ;
  assign n1998 = n1997 ^ n1991 ;
  assign n2002 = n2001 ^ n1998 ;
  assign n26108 = n26107 ^ n2002 ;
  assign n26110 = n3060 ^ n1922 ;
  assign n26111 = n26110 ^ n21195 ;
  assign n26112 = n26111 ^ n1994 ;
  assign n26109 = n26053 ^ n26049 ;
  assign n26113 = n26112 ^ n26109 ;
  assign n3038 = n3028 ^ n3010 ;
  assign n3039 = n3038 ^ n2781 ;
  assign n3040 = n3039 ^ n3037 ;
  assign n26114 = n3040 & n26050 ;
  assign n3047 = n3022 ^ n1916 ;
  assign n3048 = n3047 ^ n3044 ;
  assign n3052 = n3051 ^ n3048 ;
  assign n26115 = n26114 ^ n3052 ;
  assign n26116 = n26052 ^ n26050 ;
  assign n26117 = n26116 ^ n3052 ;
  assign n26118 = n26115 & n26117 ;
  assign n26119 = n26118 ^ n26114 ;
  assign n26120 = n26119 ^ n26109 ;
  assign n26121 = ~n26113 & n26120 ;
  assign n26122 = n26121 ^ n26112 ;
  assign n26123 = n26122 ^ n2002 ;
  assign n26124 = ~n26108 & n26123 ;
  assign n26125 = n26124 ^ n2002 ;
  assign n26607 = n26125 ^ n2014 ;
  assign n26129 = n26090 & n26607 ;
  assign n26106 = n26105 ^ n26091 ;
  assign n26126 = n26125 ^ n26106 ;
  assign n26130 = n26129 ^ n26126 ;
  assign n26488 = n26360 ^ n26359 ;
  assign n2083 = n2079 ^ n2031 ;
  assign n2087 = n2086 ^ n2083 ;
  assign n2091 = n2090 ^ n2087 ;
  assign n26490 = n26488 ^ n2091 ;
  assign n26489 = n26488 ^ n26106 ;
  assign n26491 = n26490 ^ n26489 ;
  assign n26492 = n26130 & n26491 ;
  assign n26493 = n26492 ^ n26489 ;
  assign n26495 = n24562 ^ n2406 ;
  assign n26496 = n26495 ^ n2095 ;
  assign n26497 = n26496 ^ n2209 ;
  assign n26498 = n26497 ^ n2216 ;
  assign n26494 = n26488 ^ n2216 ;
  assign n26499 = n26498 ^ n26494 ;
  assign n26500 = ~n26493 & ~n26499 ;
  assign n26501 = n26500 ^ n26494 ;
  assign n26502 = n26362 ^ n26361 ;
  assign n26503 = n26502 ^ n2216 ;
  assign n26504 = ~n26501 & n26503 ;
  assign n26506 = n26505 ^ n26504 ;
  assign n26507 = ~n26487 & n26506 ;
  assign n26508 = n26507 ^ n26486 ;
  assign n26509 = n26508 ^ n26478 ;
  assign n26510 = n26482 & ~n26509 ;
  assign n26511 = n26510 ^ n26481 ;
  assign n26475 = n26369 ^ n26356 ;
  assign n26476 = n26475 ^ n26472 ;
  assign n26477 = n26476 ^ n26475 ;
  assign n26512 = n26511 ^ n26477 ;
  assign n26513 = n26474 & n26512 ;
  assign n26514 = n26513 ^ n26476 ;
  assign n26519 = n26475 ^ n1499 ;
  assign n26518 = n26517 ^ n1499 ;
  assign n26520 = n26519 ^ n26518 ;
  assign n26521 = ~n26514 & ~n26520 ;
  assign n26522 = n26521 ^ n26519 ;
  assign n26528 = n26525 ^ n1499 ;
  assign n26526 = n26371 ^ n26370 ;
  assign n26527 = n26526 ^ n26525 ;
  assign n26529 = n26528 ^ n26527 ;
  assign n26530 = ~n26522 & n26529 ;
  assign n26531 = n26530 ^ n26528 ;
  assign n26532 = n26373 ^ n26372 ;
  assign n26533 = n26532 ^ n26525 ;
  assign n26534 = n26531 & ~n26533 ;
  assign n26536 = n26535 ^ n26534 ;
  assign n26537 = ~n26469 & ~n26536 ;
  assign n26538 = n26537 ^ n26468 ;
  assign n26540 = n26539 ^ n26538 ;
  assign n26541 = n26538 ^ n2974 ;
  assign n26542 = ~n26540 & ~n26541 ;
  assign n26543 = n26542 ^ n2974 ;
  assign n26653 = n26543 ^ n695 ;
  assign n26319 = n26318 ^ n26267 ;
  assign n26320 = ~n26268 & ~n26319 ;
  assign n26321 = n26320 ^ n23272 ;
  assign n26162 = n26161 ^ n26160 ;
  assign n26230 = ~n26162 & n26229 ;
  assign n26231 = n26230 ^ n26161 ;
  assign n26156 = n25114 ^ n24138 ;
  assign n26157 = n26156 ^ n25232 ;
  assign n26155 = n25892 ^ n25823 ;
  assign n26158 = n26157 ^ n26155 ;
  assign n26265 = n26231 ^ n26158 ;
  assign n26266 = n26265 ^ n23266 ;
  assign n26380 = n26321 ^ n26266 ;
  assign n26379 = n26377 & n26378 ;
  assign n26467 = n26380 ^ n26379 ;
  assign n26654 = n26653 ^ n26467 ;
  assign n26651 = n25961 ^ n25109 ;
  assign n26428 = n25920 ^ n1151 ;
  assign n26429 = n26428 ^ n25921 ;
  assign n26652 = n26651 ^ n26429 ;
  assign n26655 = n26654 ^ n26652 ;
  assign n26658 = n26540 ^ n2974 ;
  assign n26413 = n25917 ^ n25797 ;
  assign n26656 = n26413 ^ n25779 ;
  assign n26657 = n26656 ^ n25105 ;
  assign n26659 = n26658 ^ n26657 ;
  assign n26662 = n26506 ^ n26483 ;
  assign n26147 = n25897 ^ n25811 ;
  assign n26660 = n26147 ^ n25119 ;
  assign n26661 = n26660 ^ n25129 ;
  assign n26663 = n26662 ^ n26661 ;
  assign n26669 = n26502 ^ n26501 ;
  assign n26667 = n25135 ^ n25127 ;
  assign n26151 = n25894 ^ n25817 ;
  assign n26668 = n26667 ^ n26151 ;
  assign n26670 = n26669 ^ n26668 ;
  assign n26672 = n26155 ^ n25141 ;
  assign n26673 = n26672 ^ n25535 ;
  assign n26671 = n26497 ^ n26493 ;
  assign n26674 = n26673 ^ n26671 ;
  assign n26675 = n26161 ^ n25091 ;
  assign n26676 = n26675 ^ n25520 ;
  assign n26131 = n26130 ^ n2091 ;
  assign n26677 = n26676 ^ n26131 ;
  assign n26678 = n26165 ^ n25134 ;
  assign n26679 = n26678 ^ n25074 ;
  assign n26608 = n26607 ^ n26089 ;
  assign n26680 = n26679 ^ n26608 ;
  assign n26683 = n26122 ^ n26108 ;
  assign n26817 = n26683 ^ n26608 ;
  assign n26681 = n25132 ^ n24860 ;
  assign n26682 = n26681 ^ n26169 ;
  assign n26684 = n26683 ^ n26682 ;
  assign n26687 = n26119 ^ n26113 ;
  assign n26685 = n26133 ^ n24706 ;
  assign n26686 = n26685 ^ n25138 ;
  assign n26688 = n26687 ^ n26686 ;
  assign n26691 = n26116 ^ n26115 ;
  assign n26689 = n26176 ^ n25140 ;
  assign n26690 = n26689 ^ n24852 ;
  assign n26692 = n26691 ^ n26690 ;
  assign n26694 = n26180 ^ n24710 ;
  assign n26695 = n26694 ^ n25147 ;
  assign n26808 = n26695 ^ n26690 ;
  assign n26693 = n26050 ^ n3040 ;
  assign n26696 = n26695 ^ n26693 ;
  assign n26717 = n25460 ^ n24238 ;
  assign n26718 = n26717 ^ n24807 ;
  assign n26637 = n25939 ^ n2882 ;
  assign n26719 = n26718 ^ n26637 ;
  assign n26702 = n25470 ^ n24122 ;
  assign n26703 = n26702 ^ n24811 ;
  assign n26646 = n25934 ^ n1385 ;
  assign n26704 = n26703 ^ n26646 ;
  assign n26430 = n26068 ^ n24030 ;
  assign n26431 = n26430 ^ n24679 ;
  assign n26432 = n26431 ^ n26429 ;
  assign n26583 = n25928 ^ n1765 ;
  assign n26584 = n26583 ^ n26429 ;
  assign n26585 = n26584 ^ n26583 ;
  assign n26414 = n26035 ^ n24035 ;
  assign n26415 = n26414 ^ n24682 ;
  assign n26416 = n26415 ^ n26413 ;
  assign n26399 = n25989 ^ n25443 ;
  assign n26400 = n26399 ^ n24781 ;
  assign n26398 = n25915 ^ n991 ;
  assign n26401 = n26400 ^ n26398 ;
  assign n26350 = n25911 ^ n884 ;
  assign n26348 = n25961 ^ n25180 ;
  assign n26349 = n26348 ^ n24766 ;
  assign n26351 = n26350 ^ n26349 ;
  assign n26249 = n25908 ^ n25801 ;
  assign n26137 = n25905 ^ n25806 ;
  assign n26250 = n26249 ^ n26137 ;
  assign n26135 = n25767 ^ n24668 ;
  assign n26136 = n26135 ^ n25109 ;
  assign n26138 = n26137 ^ n26136 ;
  assign n26140 = n25105 ^ n24498 ;
  assign n26141 = n26140 ^ n25694 ;
  assign n26139 = n25902 ^ n25808 ;
  assign n26142 = n26141 ^ n26139 ;
  assign n26145 = n25899 ^ n25810 ;
  assign n26143 = n25559 ^ n24433 ;
  assign n26144 = n26143 ^ n25115 ;
  assign n26146 = n26145 ^ n26144 ;
  assign n26148 = n25120 ^ n24306 ;
  assign n26149 = n26148 ^ n25554 ;
  assign n26150 = n26149 ^ n26147 ;
  assign n26152 = n25124 ^ n24134 ;
  assign n26153 = n26152 ^ n25104 ;
  assign n26154 = n26153 ^ n26151 ;
  assign n26232 = n26231 ^ n26155 ;
  assign n26233 = ~n26158 & n26232 ;
  assign n26234 = n26233 ^ n26157 ;
  assign n26235 = n26234 ^ n26151 ;
  assign n26236 = ~n26154 & ~n26235 ;
  assign n26237 = n26236 ^ n26153 ;
  assign n26238 = n26237 ^ n26147 ;
  assign n26239 = ~n26150 & ~n26238 ;
  assign n26240 = n26239 ^ n26149 ;
  assign n26241 = n26240 ^ n26144 ;
  assign n26242 = ~n26146 & ~n26241 ;
  assign n26243 = n26242 ^ n26145 ;
  assign n26244 = n26243 ^ n26139 ;
  assign n26245 = n26142 & n26244 ;
  assign n26246 = n26245 ^ n26141 ;
  assign n26247 = n26246 ^ n26137 ;
  assign n26248 = n26138 & ~n26247 ;
  assign n26251 = n26250 ^ n26248 ;
  assign n26252 = n25779 ^ n24753 ;
  assign n26253 = n26252 ^ n25176 ;
  assign n26345 = n26253 ^ n26249 ;
  assign n26346 = ~n26251 & ~n26345 ;
  assign n26347 = n26346 ^ n26253 ;
  assign n26395 = n26349 ^ n26347 ;
  assign n26396 = n26351 & ~n26395 ;
  assign n26397 = n26396 ^ n26350 ;
  assign n26410 = n26398 ^ n26397 ;
  assign n26411 = n26401 & ~n26410 ;
  assign n26412 = n26411 ^ n26400 ;
  assign n26425 = n26413 ^ n26412 ;
  assign n26426 = n26416 & n26425 ;
  assign n26427 = n26426 ^ n26415 ;
  assign n26586 = n26585 ^ n26427 ;
  assign n26587 = n26432 & ~n26586 ;
  assign n26588 = n26587 ^ n26584 ;
  assign n26589 = n25467 ^ n24815 ;
  assign n26590 = n26589 ^ n24076 ;
  assign n26699 = n26590 ^ n26583 ;
  assign n26700 = ~n26588 & n26699 ;
  assign n26701 = n26700 ^ n26583 ;
  assign n26714 = n26701 ^ n26646 ;
  assign n26715 = ~n26704 & n26714 ;
  assign n26716 = n26715 ^ n26646 ;
  assign n26720 = n26719 ^ n26716 ;
  assign n26721 = n26720 ^ n23531 ;
  assign n26705 = n26704 ^ n26701 ;
  assign n26706 = n26705 ^ n23533 ;
  assign n26352 = n26351 ^ n26347 ;
  assign n26353 = n26352 ^ n24106 ;
  assign n26254 = n26253 ^ n26251 ;
  assign n26255 = n26254 ^ n24063 ;
  assign n26257 = n26243 ^ n26142 ;
  assign n26258 = n26257 ^ n23647 ;
  assign n26259 = n26240 ^ n26146 ;
  assign n26260 = n26259 ^ n23248 ;
  assign n26261 = n26237 ^ n26150 ;
  assign n26262 = n26261 ^ n23256 ;
  assign n26263 = n26234 ^ n26154 ;
  assign n26264 = n26263 ^ n23261 ;
  assign n26322 = n26321 ^ n26265 ;
  assign n26323 = ~n26266 & n26322 ;
  assign n26324 = n26323 ^ n23266 ;
  assign n26325 = n26324 ^ n26263 ;
  assign n26326 = ~n26264 & n26325 ;
  assign n26327 = n26326 ^ n23261 ;
  assign n26328 = n26327 ^ n26261 ;
  assign n26329 = ~n26262 & ~n26328 ;
  assign n26330 = n26329 ^ n23256 ;
  assign n26331 = n26330 ^ n26259 ;
  assign n26332 = ~n26260 & ~n26331 ;
  assign n26333 = n26332 ^ n23248 ;
  assign n26334 = n26333 ^ n26257 ;
  assign n26335 = n26258 & n26334 ;
  assign n26336 = n26335 ^ n23647 ;
  assign n26256 = n26246 ^ n26138 ;
  assign n26337 = n26336 ^ n26256 ;
  assign n26338 = n26254 ^ n24022 ;
  assign n26339 = n26338 ^ n26254 ;
  assign n26340 = n26339 ^ n26256 ;
  assign n26341 = n26337 & ~n26340 ;
  assign n26342 = n26341 ^ n26338 ;
  assign n26343 = n26255 & n26342 ;
  assign n26344 = n26343 ^ n24063 ;
  assign n26404 = n26352 ^ n26344 ;
  assign n26405 = n26353 & ~n26404 ;
  assign n26406 = n26405 ^ n24106 ;
  assign n26402 = n26401 ^ n26397 ;
  assign n26409 = n26406 ^ n26402 ;
  assign n26417 = n26416 ^ n26412 ;
  assign n26418 = n26417 ^ n24227 ;
  assign n26419 = n26418 ^ n26402 ;
  assign n26420 = n26419 ^ n26417 ;
  assign n26421 = ~n26409 & n26420 ;
  assign n26422 = n26421 ^ n26418 ;
  assign n26433 = n26432 ^ n26427 ;
  assign n26435 = n26433 ^ n23547 ;
  assign n26434 = n26433 ^ n26417 ;
  assign n26436 = n26435 ^ n26434 ;
  assign n26437 = ~n26422 & ~n26436 ;
  assign n26438 = n26437 ^ n26435 ;
  assign n26591 = n26590 ^ n26588 ;
  assign n26593 = n26591 ^ n23550 ;
  assign n26592 = n26591 ^ n26433 ;
  assign n26594 = n26593 ^ n26592 ;
  assign n26595 = ~n26438 & n26594 ;
  assign n26596 = n26595 ^ n26593 ;
  assign n26708 = n26705 ^ n23537 ;
  assign n26707 = n26705 ^ n26591 ;
  assign n26709 = n26708 ^ n26707 ;
  assign n26710 = n26596 & ~n26709 ;
  assign n26711 = n26710 ^ n26708 ;
  assign n26712 = ~n26706 & n26711 ;
  assign n26713 = n26712 ^ n23533 ;
  assign n26722 = n26721 ^ n26713 ;
  assign n26597 = n26596 ^ n23537 ;
  assign n26354 = n26353 ^ n26344 ;
  assign n26355 = n26342 ^ n24063 ;
  assign n26381 = n26379 & ~n26380 ;
  assign n26382 = n26324 ^ n26264 ;
  assign n26383 = ~n26381 & n26382 ;
  assign n26384 = n26327 ^ n26262 ;
  assign n26385 = n26383 & n26384 ;
  assign n26386 = n26330 ^ n26260 ;
  assign n26387 = ~n26385 & n26386 ;
  assign n26388 = n26333 ^ n26258 ;
  assign n26389 = n26387 & n26388 ;
  assign n26390 = n26256 ^ n24022 ;
  assign n26391 = n26390 ^ n26336 ;
  assign n26392 = ~n26389 & ~n26391 ;
  assign n26393 = ~n26355 & ~n26392 ;
  assign n26394 = n26354 & n26393 ;
  assign n26403 = n26402 ^ n24227 ;
  assign n26407 = n26406 ^ n26403 ;
  assign n26408 = ~n26394 & ~n26407 ;
  assign n26423 = n26422 ^ n23547 ;
  assign n26424 = ~n26408 & ~n26423 ;
  assign n26439 = n26438 ^ n23550 ;
  assign n26598 = n26424 & ~n26439 ;
  assign n26723 = n26597 & n26598 ;
  assign n26724 = n26711 ^ n23533 ;
  assign n26725 = ~n26723 & ~n26724 ;
  assign n26726 = n26722 & ~n26725 ;
  assign n26733 = n26716 ^ n26637 ;
  assign n26734 = ~n26719 & ~n26733 ;
  assign n26735 = n26734 ^ n26637 ;
  assign n26730 = n25456 ^ n24214 ;
  assign n26731 = n26730 ^ n24743 ;
  assign n26633 = n25941 ^ n25793 ;
  assign n26732 = n26731 ^ n26633 ;
  assign n26736 = n26735 ^ n26732 ;
  assign n26737 = n26736 ^ n23332 ;
  assign n26727 = n26720 ^ n26713 ;
  assign n26728 = ~n26721 & n26727 ;
  assign n26729 = n26728 ^ n23531 ;
  assign n26738 = n26737 ^ n26729 ;
  assign n26775 = n26726 & n26738 ;
  assign n26769 = n23332 ^ n23328 ;
  assign n26765 = n25450 ^ n24739 ;
  assign n26766 = n26765 ^ n24208 ;
  assign n26626 = n25944 ^ n25791 ;
  assign n26767 = n26766 ^ n26626 ;
  assign n26768 = n26767 ^ n26731 ;
  assign n26770 = n26769 ^ n26768 ;
  assign n26771 = n26770 ^ n2767 ;
  assign n2770 = n2717 ^ n2680 ;
  assign n2771 = n2770 ^ n1841 ;
  assign n2772 = n2771 ^ n2763 ;
  assign n26772 = n26771 ^ n2772 ;
  assign n26763 = n26736 ^ n26729 ;
  assign n26764 = ~n26737 & ~n26763 ;
  assign n26773 = n26772 ^ n26764 ;
  assign n26761 = n26735 ^ n26731 ;
  assign n26762 = ~n26732 & ~n26761 ;
  assign n26774 = n26773 ^ n26762 ;
  assign n26776 = n26775 ^ n26774 ;
  assign n26739 = n26738 ^ n26726 ;
  assign n26740 = n26739 ^ n2772 ;
  assign n26751 = n26725 ^ n26722 ;
  assign n26741 = n26724 ^ n26723 ;
  assign n26742 = n26741 ^ n3138 ;
  assign n26579 = n24649 ^ n3121 ;
  assign n26580 = n26579 ^ n2513 ;
  assign n26581 = n26580 ^ n3133 ;
  assign n26440 = n26439 ^ n26424 ;
  assign n26444 = n26443 ^ n26440 ;
  assign n26445 = n26423 ^ n26408 ;
  assign n26446 = n26445 ^ n2645 ;
  assign n26448 = n3203 ^ n1379 ;
  assign n26449 = n26448 ^ n21516 ;
  assign n26450 = n26449 ^ n2544 ;
  assign n26447 = n26407 ^ n26394 ;
  assign n26451 = n26450 ^ n26447 ;
  assign n26452 = n26392 ^ n26355 ;
  assign n26453 = n26452 ^ n1277 ;
  assign n26457 = n26391 ^ n26389 ;
  assign n26458 = n26457 ^ n1134 ;
  assign n26459 = n26388 ^ n26387 ;
  assign n1095 = n1077 ^ n1029 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1103 = n1102 ^ n1099 ;
  assign n26460 = n26459 ^ n1103 ;
  assign n26461 = n26386 ^ n26385 ;
  assign n26462 = n26461 ^ n1114 ;
  assign n26463 = n26384 ^ n26383 ;
  assign n26464 = n26463 ^ n1652 ;
  assign n26465 = n26382 ^ n26381 ;
  assign n26466 = n26465 ^ n1646 ;
  assign n26547 = n26543 ^ n26465 ;
  assign n26544 = n26543 ^ n26467 ;
  assign n26545 = n26467 ^ n695 ;
  assign n26546 = n26544 & ~n26545 ;
  assign n26548 = n26547 ^ n26546 ;
  assign n26549 = ~n26466 & ~n26548 ;
  assign n26550 = n26549 ^ n26465 ;
  assign n26551 = n26550 ^ n1652 ;
  assign n26552 = n26464 & n26551 ;
  assign n26553 = n26552 ^ n26463 ;
  assign n26554 = n26553 ^ n1114 ;
  assign n26555 = n26462 & ~n26554 ;
  assign n26556 = n26555 ^ n26461 ;
  assign n26557 = n26556 ^ n1103 ;
  assign n26558 = ~n26460 & ~n26557 ;
  assign n26559 = n26558 ^ n26459 ;
  assign n26560 = n26559 ^ n1134 ;
  assign n26561 = n26458 & n26560 ;
  assign n26562 = n26561 ^ n26457 ;
  assign n26454 = n26393 ^ n26354 ;
  assign n26455 = n26454 ^ n1277 ;
  assign n26456 = n26455 ^ n26454 ;
  assign n26563 = n26562 ^ n26456 ;
  assign n26564 = ~n26453 & n26563 ;
  assign n26565 = n26564 ^ n26455 ;
  assign n26567 = n26447 ^ n2789 ;
  assign n26566 = n26454 ^ n26447 ;
  assign n26568 = n26567 ^ n26566 ;
  assign n26569 = n26565 & ~n26568 ;
  assign n26570 = n26569 ^ n26567 ;
  assign n26571 = n26451 & ~n26570 ;
  assign n26572 = n26571 ^ n26450 ;
  assign n26573 = n26572 ^ n26445 ;
  assign n26574 = ~n26446 & n26573 ;
  assign n26575 = n26574 ^ n2645 ;
  assign n26576 = n26575 ^ n26440 ;
  assign n26577 = n26444 & ~n26576 ;
  assign n26578 = n26577 ^ n26443 ;
  assign n26582 = n26581 ^ n26578 ;
  assign n26599 = n26598 ^ n26597 ;
  assign n26743 = n26599 ^ n26578 ;
  assign n26747 = n26582 & n26743 ;
  assign n26744 = n26581 ^ n3138 ;
  assign n26748 = n26747 ^ n26744 ;
  assign n26749 = n26742 & n26748 ;
  assign n26750 = n26749 ^ n3138 ;
  assign n26752 = n26751 ^ n26750 ;
  assign n26753 = n24677 ^ n2665 ;
  assign n26754 = n26753 ^ n3142 ;
  assign n26755 = n26754 ^ n1817 ;
  assign n26756 = n26755 ^ n26751 ;
  assign n26757 = ~n26752 & n26756 ;
  assign n26758 = n26757 ^ n26755 ;
  assign n26759 = n26758 ^ n2772 ;
  assign n26760 = ~n26740 & n26759 ;
  assign n26777 = n26776 ^ n26760 ;
  assign n26697 = n26184 ^ n24716 ;
  assign n26698 = n26697 ^ n25151 ;
  assign n26778 = n26777 ^ n26698 ;
  assign n26792 = n26188 ^ n24720 ;
  assign n26793 = n26792 ^ n25153 ;
  assign n26802 = n26793 ^ n26698 ;
  assign n26600 = n26599 ^ n26582 ;
  assign n26601 = n26102 ^ n24733 ;
  assign n26602 = n26601 ^ n25165 ;
  assign n26781 = ~n26600 & n26602 ;
  assign n26779 = n26197 ^ n25163 ;
  assign n26780 = n26779 ^ n24129 ;
  assign n26782 = n26781 ^ n26780 ;
  assign n26787 = n26748 ^ n26741 ;
  assign n26783 = n25157 ^ n24724 ;
  assign n26784 = n26783 ^ n26192 ;
  assign n26785 = n26784 ^ n26780 ;
  assign n26786 = n26785 ^ n26784 ;
  assign n26788 = n26787 ^ n26786 ;
  assign n26789 = n26782 & n26788 ;
  assign n26790 = n26789 ^ n26785 ;
  assign n26795 = n26793 ^ n26784 ;
  assign n26791 = n26756 ^ n26750 ;
  assign n26794 = n26793 ^ n26791 ;
  assign n26796 = n26795 ^ n26794 ;
  assign n26797 = ~n26790 & ~n26796 ;
  assign n26798 = n26797 ^ n26795 ;
  assign n26799 = n26758 ^ n26740 ;
  assign n26800 = n26799 ^ n26793 ;
  assign n26801 = n26798 & n26800 ;
  assign n26803 = n26802 ^ n26801 ;
  assign n26804 = n26778 & ~n26803 ;
  assign n26805 = n26804 ^ n26777 ;
  assign n26806 = n26805 ^ n26693 ;
  assign n26807 = ~n26696 & n26806 ;
  assign n26809 = n26808 ^ n26807 ;
  assign n26810 = n26692 & ~n26809 ;
  assign n26811 = n26810 ^ n26691 ;
  assign n26812 = n26811 ^ n26686 ;
  assign n26813 = ~n26688 & n26812 ;
  assign n26814 = n26813 ^ n26687 ;
  assign n26815 = n26814 ^ n26683 ;
  assign n26816 = n26684 & n26815 ;
  assign n26818 = n26817 ^ n26816 ;
  assign n26819 = n26680 & n26818 ;
  assign n26820 = n26819 ^ n26608 ;
  assign n26821 = n26820 ^ n26676 ;
  assign n26822 = ~n26677 & ~n26821 ;
  assign n26823 = n26822 ^ n26131 ;
  assign n26824 = n26823 ^ n26671 ;
  assign n26825 = ~n26674 & n26824 ;
  assign n26826 = n26825 ^ n26673 ;
  assign n26827 = n26826 ^ n26668 ;
  assign n26828 = n26670 & n26827 ;
  assign n26829 = n26828 ^ n26669 ;
  assign n26664 = n26508 ^ n26482 ;
  assign n26665 = n26664 ^ n26662 ;
  assign n26666 = n26665 ^ n26664 ;
  assign n26830 = n26829 ^ n26666 ;
  assign n26831 = n26663 & n26830 ;
  assign n26832 = n26831 ^ n26665 ;
  assign n26833 = n26511 ^ n26474 ;
  assign n26837 = n26833 ^ n26664 ;
  assign n26834 = n26145 ^ n25200 ;
  assign n26835 = n26834 ^ n25114 ;
  assign n26836 = n26835 ^ n26833 ;
  assign n26838 = n26837 ^ n26836 ;
  assign n26839 = ~n26832 & ~n26838 ;
  assign n26840 = n26839 ^ n26837 ;
  assign n26841 = n26517 ^ n26514 ;
  assign n26845 = n26841 ^ n26833 ;
  assign n26842 = n26139 ^ n25104 ;
  assign n26843 = n26842 ^ n25231 ;
  assign n26844 = n26843 ^ n26841 ;
  assign n26846 = n26845 ^ n26844 ;
  assign n26847 = n26840 & ~n26846 ;
  assign n26848 = n26847 ^ n26845 ;
  assign n26849 = n26249 ^ n25559 ;
  assign n26850 = n26849 ^ n25124 ;
  assign n26854 = n26850 ^ n26841 ;
  assign n26851 = n25554 ^ n25232 ;
  assign n26852 = n26851 ^ n26137 ;
  assign n26853 = n26852 ^ n26850 ;
  assign n26855 = n26854 ^ n26853 ;
  assign n26856 = ~n26848 & ~n26855 ;
  assign n26857 = n26856 ^ n26854 ;
  assign n26858 = n26350 ^ n25120 ;
  assign n26859 = n26858 ^ n25694 ;
  assign n26862 = n26859 ^ n26850 ;
  assign n26860 = n26526 ^ n26522 ;
  assign n26861 = n26860 ^ n26859 ;
  assign n26863 = n26862 ^ n26861 ;
  assign n26864 = ~n26857 & ~n26863 ;
  assign n26865 = n26864 ^ n26862 ;
  assign n26866 = n26398 ^ n25115 ;
  assign n26867 = n26866 ^ n25767 ;
  assign n26870 = n26867 ^ n26859 ;
  assign n26868 = n26532 ^ n26531 ;
  assign n26869 = n26868 ^ n26867 ;
  assign n26871 = n26870 ^ n26869 ;
  assign n26872 = n26865 & ~n26871 ;
  assign n26873 = n26872 ^ n26870 ;
  assign n26876 = n26867 ^ n26658 ;
  assign n26874 = n26536 ^ n633 ;
  assign n26875 = n26874 ^ n26658 ;
  assign n26877 = n26876 ^ n26875 ;
  assign n26878 = ~n26873 & n26877 ;
  assign n26879 = n26878 ^ n26876 ;
  assign n26880 = n26659 & ~n26879 ;
  assign n26881 = n26880 ^ n26658 ;
  assign n26882 = n26881 ^ n26652 ;
  assign n26883 = n26655 & ~n26882 ;
  assign n26884 = n26883 ^ n26654 ;
  assign n26644 = n26548 ^ n1646 ;
  assign n26642 = n25989 ^ n25176 ;
  assign n26643 = n26642 ^ n26583 ;
  assign n26645 = n26644 ^ n26643 ;
  assign n26925 = n26884 ^ n26645 ;
  assign n27117 = n26925 ^ n24753 ;
  assign n26926 = n26881 ^ n26655 ;
  assign n26927 = n26926 ^ n24668 ;
  assign n27029 = n26879 ^ n26657 ;
  assign n26929 = n26868 ^ n26865 ;
  assign n26930 = n26929 ^ n24306 ;
  assign n27016 = n26860 ^ n26857 ;
  assign n26931 = n26843 ^ n26840 ;
  assign n26932 = n26931 ^ n24142 ;
  assign n26934 = n26823 ^ n26674 ;
  assign n26935 = n26934 ^ n24160 ;
  assign n26936 = n26820 ^ n26677 ;
  assign n26937 = n26936 ^ n24164 ;
  assign n26939 = n26814 ^ n26684 ;
  assign n26940 = n26939 ^ n24173 ;
  assign n26941 = n26811 ^ n26688 ;
  assign n26942 = n26941 ^ n24175 ;
  assign n26944 = n26805 ^ n26696 ;
  assign n26945 = n26944 ^ n24181 ;
  assign n26946 = n26803 ^ n26777 ;
  assign n26947 = n26946 ^ n24188 ;
  assign n26959 = n26799 ^ n26798 ;
  assign n26603 = n26602 ^ n26600 ;
  assign n26948 = ~n24206 & ~n26603 ;
  assign n26949 = n26948 ^ n24130 ;
  assign n26950 = n26787 ^ n26782 ;
  assign n26951 = n26950 ^ n26948 ;
  assign n26952 = ~n26949 & ~n26951 ;
  assign n26953 = n26952 ^ n24130 ;
  assign n26954 = n26953 ^ n24195 ;
  assign n26955 = n26791 ^ n26790 ;
  assign n26956 = n26955 ^ n26953 ;
  assign n26957 = ~n26954 & ~n26956 ;
  assign n26958 = n26957 ^ n24195 ;
  assign n26960 = n26959 ^ n26958 ;
  assign n26961 = n26959 ^ n24193 ;
  assign n26962 = n26960 & ~n26961 ;
  assign n26963 = n26962 ^ n24193 ;
  assign n26964 = n26963 ^ n26946 ;
  assign n26965 = ~n26947 & n26964 ;
  assign n26966 = n26965 ^ n24188 ;
  assign n26967 = n26966 ^ n26944 ;
  assign n26968 = n26945 & ~n26967 ;
  assign n26969 = n26968 ^ n24181 ;
  assign n26943 = n26809 ^ n26691 ;
  assign n26970 = n26969 ^ n26943 ;
  assign n26971 = n26941 ^ n24183 ;
  assign n26972 = n26971 ^ n26941 ;
  assign n26973 = n26972 ^ n26943 ;
  assign n26974 = n26970 & ~n26973 ;
  assign n26975 = n26974 ^ n26971 ;
  assign n26976 = ~n26942 & ~n26975 ;
  assign n26977 = n26976 ^ n24175 ;
  assign n26978 = n26977 ^ n26939 ;
  assign n26979 = ~n26940 & ~n26978 ;
  assign n26980 = n26979 ^ n24173 ;
  assign n26938 = n26818 ^ n26679 ;
  assign n26981 = n26980 ^ n26938 ;
  assign n26982 = n26936 ^ n24168 ;
  assign n26983 = n26982 ^ n26936 ;
  assign n26984 = n26983 ^ n26938 ;
  assign n26985 = n26981 & ~n26984 ;
  assign n26986 = n26985 ^ n26982 ;
  assign n26987 = n26937 & ~n26986 ;
  assign n26988 = n26987 ^ n24164 ;
  assign n26989 = n26988 ^ n26934 ;
  assign n26990 = ~n26935 & n26989 ;
  assign n26991 = n26990 ^ n24160 ;
  assign n26992 = n26991 ^ n24154 ;
  assign n26993 = n26826 ^ n26670 ;
  assign n26994 = n26993 ^ n26991 ;
  assign n26995 = n26992 & ~n26994 ;
  assign n26996 = n26995 ^ n24154 ;
  assign n26933 = n26829 ^ n26663 ;
  assign n26997 = n26996 ^ n26933 ;
  assign n26998 = n26835 ^ n26832 ;
  assign n26999 = n26998 ^ n24148 ;
  assign n27000 = n26999 ^ n26933 ;
  assign n27001 = n27000 ^ n26998 ;
  assign n27002 = n26997 & n27001 ;
  assign n27003 = n27002 ^ n26999 ;
  assign n27005 = n26931 ^ n24146 ;
  assign n27004 = n26998 ^ n26931 ;
  assign n27006 = n27005 ^ n27004 ;
  assign n27007 = n27003 & ~n27006 ;
  assign n27008 = n27007 ^ n27005 ;
  assign n27009 = n26932 & ~n27008 ;
  assign n27010 = n27009 ^ n24142 ;
  assign n27011 = n27010 ^ n24138 ;
  assign n27012 = n26852 ^ n26848 ;
  assign n27013 = n27012 ^ n27010 ;
  assign n27014 = n27011 & ~n27013 ;
  assign n27015 = n27014 ^ n24138 ;
  assign n27017 = n27016 ^ n27015 ;
  assign n27018 = n26929 ^ n24134 ;
  assign n27019 = n27018 ^ n27015 ;
  assign n27020 = n27019 ^ n26929 ;
  assign n27021 = n27017 & n27020 ;
  assign n27022 = n27021 ^ n27018 ;
  assign n27023 = n26930 & ~n27022 ;
  assign n27024 = n27023 ^ n24306 ;
  assign n26928 = n26874 ^ n26873 ;
  assign n27025 = n27024 ^ n26928 ;
  assign n27026 = n27024 ^ n24433 ;
  assign n27027 = n27025 & ~n27026 ;
  assign n27028 = n27027 ^ n24433 ;
  assign n27030 = n27029 ^ n27028 ;
  assign n27031 = n27029 ^ n24498 ;
  assign n27032 = n27030 & n27031 ;
  assign n27033 = n27032 ^ n24498 ;
  assign n27034 = n27033 ^ n26926 ;
  assign n27035 = n26927 & n27034 ;
  assign n27036 = n27035 ^ n24668 ;
  assign n27118 = n27117 ^ n27036 ;
  assign n27067 = n26928 ^ n24433 ;
  assign n27068 = n27067 ^ n27024 ;
  assign n27069 = n27022 ^ n24306 ;
  assign n27070 = n27003 ^ n24146 ;
  assign n27071 = n26996 ^ n24148 ;
  assign n27072 = n27071 ^ n26933 ;
  assign n27073 = n26993 ^ n26992 ;
  assign n27074 = n26963 ^ n24188 ;
  assign n27075 = n27074 ^ n26946 ;
  assign n27076 = n26961 ^ n26958 ;
  assign n26604 = n26603 ^ n24206 ;
  assign n27077 = n26950 ^ n26949 ;
  assign n27078 = n26604 & ~n27077 ;
  assign n27079 = n26955 ^ n26954 ;
  assign n27080 = n27078 & n27079 ;
  assign n27081 = ~n27076 & n27080 ;
  assign n27082 = ~n27075 & n27081 ;
  assign n27083 = n26966 ^ n24181 ;
  assign n27084 = n27083 ^ n26944 ;
  assign n27085 = ~n27082 & ~n27084 ;
  assign n27086 = n26969 ^ n24183 ;
  assign n27087 = n27086 ^ n26943 ;
  assign n27088 = ~n27085 & ~n27087 ;
  assign n27089 = n26975 ^ n24175 ;
  assign n27090 = ~n27088 & n27089 ;
  assign n27091 = n26977 ^ n26940 ;
  assign n27092 = n27090 & ~n27091 ;
  assign n27093 = n26938 ^ n24168 ;
  assign n27094 = n27093 ^ n26980 ;
  assign n27095 = n27092 & n27094 ;
  assign n27096 = n26986 ^ n24164 ;
  assign n27097 = ~n27095 & n27096 ;
  assign n27098 = n26988 ^ n26935 ;
  assign n27099 = ~n27097 & n27098 ;
  assign n27100 = n27073 & ~n27099 ;
  assign n27101 = ~n27072 & ~n27100 ;
  assign n27102 = ~n27070 & n27101 ;
  assign n27103 = n27008 ^ n24142 ;
  assign n27104 = n27102 & n27103 ;
  assign n27105 = n27012 ^ n27011 ;
  assign n27106 = n27104 & n27105 ;
  assign n27107 = n27016 ^ n24134 ;
  assign n27108 = n27107 ^ n27015 ;
  assign n27109 = ~n27106 & n27108 ;
  assign n27110 = ~n27069 & n27109 ;
  assign n27111 = n27068 & ~n27110 ;
  assign n27112 = n27028 ^ n24498 ;
  assign n27113 = n27112 ^ n27029 ;
  assign n27114 = n27111 & ~n27113 ;
  assign n27115 = n27033 ^ n26927 ;
  assign n27116 = ~n27114 & ~n27115 ;
  assign n27312 = n27118 ^ n27116 ;
  assign n27176 = n27115 ^ n27114 ;
  assign n1413 = n1297 ^ n1211 ;
  assign n1417 = n1416 ^ n1413 ;
  assign n1418 = n1417 ^ n1148 ;
  assign n27177 = n27176 ^ n1418 ;
  assign n1705 = n1686 ^ n1193 ;
  assign n1706 = n1705 ^ n856 ;
  assign n1707 = n1706 ^ n971 ;
  assign n981 = n980 ^ n928 ;
  assign n982 = n981 ^ n977 ;
  assign n983 = n982 ^ n968 ;
  assign n27302 = n1707 ^ n983 ;
  assign n27178 = n27110 ^ n27068 ;
  assign n27179 = n27178 ^ n1707 ;
  assign n27180 = n27109 ^ n27069 ;
  assign n27181 = n27180 ^ n852 ;
  assign n27296 = n27180 ^ n769 ;
  assign n27182 = n27105 ^ n27104 ;
  assign n27183 = n27182 ^ n757 ;
  assign n27189 = n27103 ^ n27102 ;
  assign n27190 = n27189 ^ n27188 ;
  assign n27286 = n27189 ^ n1548 ;
  assign n27191 = n27101 ^ n27070 ;
  assign n27192 = n27191 ^ n1548 ;
  assign n27196 = n27100 ^ n27072 ;
  assign n27197 = n27196 ^ n27195 ;
  assign n27198 = n27099 ^ n27073 ;
  assign n27202 = n27201 ^ n27198 ;
  assign n2925 = n2924 ^ n2921 ;
  assign n2926 = n2925 ^ n593 ;
  assign n2930 = n2929 ^ n2926 ;
  assign n27277 = n27198 ^ n2930 ;
  assign n27203 = n27098 ^ n27097 ;
  assign n27204 = n27203 ^ n2930 ;
  assign n27205 = n27096 ^ n27095 ;
  assign n27209 = n27208 ^ n27205 ;
  assign n27213 = n27094 ^ n27092 ;
  assign n27210 = n2373 ^ n587 ;
  assign n27211 = n27210 ^ n21785 ;
  assign n27212 = n27211 ^ n16711 ;
  assign n27214 = n27213 ^ n27212 ;
  assign n2312 = n2296 ^ n2233 ;
  assign n2313 = n2312 ^ n2309 ;
  assign n2314 = n2313 ^ n1463 ;
  assign n27268 = n27212 ^ n2314 ;
  assign n27215 = n27087 ^ n27085 ;
  assign n2187 = n2159 ^ n2123 ;
  assign n2188 = n2187 ^ n2184 ;
  assign n2192 = n2191 ^ n2188 ;
  assign n27216 = n27215 ^ n2192 ;
  assign n27217 = n27084 ^ n27082 ;
  assign n2178 = n2111 ^ n2070 ;
  assign n2179 = n2178 ^ n2177 ;
  assign n2180 = n2179 ^ n2171 ;
  assign n27218 = n27217 ^ n2180 ;
  assign n27220 = n25009 ^ n2055 ;
  assign n27221 = n27220 ^ n21801 ;
  assign n27222 = n27221 ^ n2175 ;
  assign n27251 = n27222 ^ n2180 ;
  assign n27219 = n27081 ^ n27075 ;
  assign n27223 = n27222 ^ n27219 ;
  assign n27236 = n27079 ^ n27078 ;
  assign n27228 = n24696 ^ n3070 ;
  assign n27229 = n27228 ^ n21810 ;
  assign n27230 = n27229 ^ n1875 ;
  assign n27227 = n1850 & ~n26604 ;
  assign n27231 = n27230 ^ n27227 ;
  assign n27232 = n27077 ^ n26604 ;
  assign n27233 = n27232 ^ n27227 ;
  assign n27234 = n27231 & n27233 ;
  assign n27235 = n27234 ^ n27230 ;
  assign n27237 = n27236 ^ n27235 ;
  assign n27238 = n24700 ^ n3087 ;
  assign n27239 = n27238 ^ n1877 ;
  assign n27240 = n27239 ^ n16729 ;
  assign n27241 = n27240 ^ n27235 ;
  assign n27242 = ~n27237 & n27241 ;
  assign n27243 = n27242 ^ n27240 ;
  assign n27224 = n25018 ^ n2048 ;
  assign n27225 = n27224 ^ n21805 ;
  assign n27226 = n27225 ^ n1931 ;
  assign n27244 = n27243 ^ n27226 ;
  assign n27245 = n27080 ^ n27076 ;
  assign n27246 = n27245 ^ n27226 ;
  assign n27247 = n27244 & n27246 ;
  assign n27248 = n27247 ^ n27243 ;
  assign n27249 = n27248 ^ n27222 ;
  assign n27250 = ~n27223 & n27249 ;
  assign n27252 = n27251 ^ n27250 ;
  assign n27253 = ~n27218 & n27252 ;
  assign n27254 = n27253 ^ n2180 ;
  assign n27255 = n27254 ^ n2192 ;
  assign n27256 = n27216 & ~n27255 ;
  assign n27257 = n27256 ^ n27215 ;
  assign n2300 = n2286 ^ n2224 ;
  assign n2301 = n2300 ^ n2199 ;
  assign n2305 = n2304 ^ n2301 ;
  assign n27258 = n27257 ^ n2305 ;
  assign n27259 = n27089 ^ n27088 ;
  assign n27262 = n27259 ^ n27257 ;
  assign n27263 = ~n27258 & n27262 ;
  assign n27260 = n27259 ^ n2314 ;
  assign n27264 = n27263 ^ n27260 ;
  assign n27265 = n27091 ^ n27090 ;
  assign n27266 = n27265 ^ n2314 ;
  assign n27267 = n27264 & n27266 ;
  assign n27269 = n27268 ^ n27267 ;
  assign n27270 = ~n27214 & ~n27269 ;
  assign n27271 = n27270 ^ n27213 ;
  assign n27272 = n27271 ^ n27205 ;
  assign n27273 = ~n27209 & ~n27272 ;
  assign n27274 = n27273 ^ n27208 ;
  assign n27275 = n27274 ^ n2930 ;
  assign n27276 = n27204 & n27275 ;
  assign n27278 = n27277 ^ n27276 ;
  assign n27279 = ~n27202 & n27278 ;
  assign n27280 = n27279 ^ n27201 ;
  assign n27281 = n27280 ^ n27195 ;
  assign n27282 = ~n27197 & ~n27281 ;
  assign n27283 = n27282 ^ n27196 ;
  assign n27284 = n27283 ^ n1548 ;
  assign n27285 = n27192 & ~n27284 ;
  assign n27287 = n27286 ^ n27285 ;
  assign n27288 = ~n27190 & ~n27287 ;
  assign n27289 = n27288 ^ n27189 ;
  assign n27290 = n27289 ^ n757 ;
  assign n27291 = ~n27183 & ~n27290 ;
  assign n27184 = n769 ^ n757 ;
  assign n27292 = n27291 ^ n27184 ;
  assign n27293 = n27108 ^ n27106 ;
  assign n27294 = n27293 ^ n769 ;
  assign n27295 = n27292 & ~n27294 ;
  assign n27297 = n27296 ^ n27295 ;
  assign n27298 = ~n27181 & ~n27297 ;
  assign n27299 = n27298 ^ n27180 ;
  assign n27300 = n27299 ^ n1707 ;
  assign n27301 = n27179 & ~n27300 ;
  assign n27303 = n27302 ^ n27301 ;
  assign n27305 = n27113 ^ n27111 ;
  assign n27304 = n1418 ^ n983 ;
  assign n27306 = n27305 ^ n27304 ;
  assign n27307 = n27306 ^ n1418 ;
  assign n27308 = n27303 & n27307 ;
  assign n27309 = n27308 ^ n27304 ;
  assign n27310 = n27177 & ~n27309 ;
  assign n27311 = n27310 ^ n27176 ;
  assign n27313 = n27312 ^ n27311 ;
  assign n1405 = n1306 ^ n1229 ;
  assign n1406 = n1405 ^ n1157 ;
  assign n1410 = n1409 ^ n1406 ;
  assign n27892 = n27313 ^ n1410 ;
  assign n26907 = n26570 ^ n26450 ;
  assign n28128 = n27892 ^ n26907 ;
  assign n27831 = n1615 ^ n1606 ;
  assign n27412 = n27240 ^ n27237 ;
  assign n27410 = n26165 ^ n25138 ;
  assign n27411 = n27410 ^ n26669 ;
  assign n27413 = n27412 ^ n27411 ;
  assign n27373 = n27232 ^ n27231 ;
  assign n27371 = n26671 ^ n26169 ;
  assign n27372 = n27371 ^ n25140 ;
  assign n27374 = n27373 ^ n27372 ;
  assign n26605 = n26604 ^ n1850 ;
  assign n26132 = n26131 ^ n25147 ;
  assign n26134 = n26133 ^ n26132 ;
  assign n26606 = n26605 ^ n26134 ;
  assign n26619 = n26565 ^ n2789 ;
  assign n26617 = n25978 ^ n25456 ;
  assign n26618 = n26617 ^ n24811 ;
  assign n26620 = n26619 ^ n26618 ;
  assign n26623 = n26562 ^ n26453 ;
  assign n26621 = n25460 ^ n24815 ;
  assign n26622 = n26621 ^ n25952 ;
  assign n26624 = n26623 ^ n26622 ;
  assign n26628 = n26559 ^ n26458 ;
  assign n26625 = n25470 ^ n24679 ;
  assign n26627 = n26626 ^ n26625 ;
  assign n26629 = n26628 ^ n26627 ;
  assign n26635 = n26556 ^ n26460 ;
  assign n26632 = n25467 ^ n24682 ;
  assign n26634 = n26633 ^ n26632 ;
  assign n26636 = n26635 ^ n26634 ;
  assign n26640 = n26553 ^ n26462 ;
  assign n26638 = n26637 ^ n25443 ;
  assign n26639 = n26638 ^ n26068 ;
  assign n26641 = n26640 ^ n26639 ;
  assign n26888 = n26550 ^ n26464 ;
  assign n26891 = n26888 ^ n26640 ;
  assign n26647 = n26646 ^ n25180 ;
  assign n26648 = n26647 ^ n26035 ;
  assign n26649 = n26648 ^ n26644 ;
  assign n26650 = n26649 ^ n26648 ;
  assign n26885 = n26884 ^ n26650 ;
  assign n26886 = ~n26645 & ~n26885 ;
  assign n26887 = n26886 ^ n26649 ;
  assign n26889 = n26888 ^ n26648 ;
  assign n26890 = n26887 & ~n26889 ;
  assign n26892 = n26891 ^ n26890 ;
  assign n26893 = n26641 & ~n26892 ;
  assign n26894 = n26893 ^ n26640 ;
  assign n26895 = n26894 ^ n26634 ;
  assign n26896 = ~n26636 & ~n26895 ;
  assign n26897 = n26896 ^ n26635 ;
  assign n26630 = n26628 ^ n26622 ;
  assign n26631 = n26630 ^ n26622 ;
  assign n26898 = n26897 ^ n26631 ;
  assign n26899 = ~n26629 & n26898 ;
  assign n26900 = n26899 ^ n26630 ;
  assign n26901 = ~n26624 & n26900 ;
  assign n26902 = n26901 ^ n26623 ;
  assign n26903 = n26902 ^ n26619 ;
  assign n26904 = n26620 & n26903 ;
  assign n26905 = n26904 ^ n26619 ;
  assign n26615 = n25450 ^ n24807 ;
  assign n26616 = n26615 ^ n26003 ;
  assign n26906 = n26905 ^ n26616 ;
  assign n26908 = n26907 ^ n26905 ;
  assign n26909 = n26906 & ~n26908 ;
  assign n26910 = n26909 ^ n26907 ;
  assign n26613 = n26572 ^ n26446 ;
  assign n26611 = n25172 ^ n24743 ;
  assign n26612 = n26611 ^ n26046 ;
  assign n26614 = n26613 ^ n26612 ;
  assign n27134 = n26910 ^ n26614 ;
  assign n27151 = n27134 ^ n24214 ;
  assign n26913 = n26907 ^ n26616 ;
  assign n26914 = n26913 ^ n26905 ;
  assign n26915 = n26914 ^ n24238 ;
  assign n26917 = n26900 ^ n26623 ;
  assign n26918 = n26917 ^ n24076 ;
  assign n26919 = n26897 ^ n26629 ;
  assign n26920 = n26919 ^ n24030 ;
  assign n26921 = n26894 ^ n26636 ;
  assign n26922 = n26921 ^ n24035 ;
  assign n26923 = n26892 ^ n26639 ;
  assign n26924 = n26923 ^ n24781 ;
  assign n27037 = n27036 ^ n26925 ;
  assign n27038 = n26888 ^ n26887 ;
  assign n27039 = n27038 ^ n24753 ;
  assign n27040 = n27039 ^ n26925 ;
  assign n27041 = n27040 ^ n27038 ;
  assign n27042 = n27037 & ~n27041 ;
  assign n27043 = n27042 ^ n27039 ;
  assign n27045 = n26923 ^ n24766 ;
  assign n27044 = n27038 ^ n26923 ;
  assign n27046 = n27045 ^ n27044 ;
  assign n27047 = ~n27043 & n27046 ;
  assign n27048 = n27047 ^ n27045 ;
  assign n27049 = ~n26924 & n27048 ;
  assign n27050 = n27049 ^ n24781 ;
  assign n27051 = n27050 ^ n26921 ;
  assign n27052 = n26922 & n27051 ;
  assign n27053 = n27052 ^ n24035 ;
  assign n27054 = n27053 ^ n26919 ;
  assign n27055 = n26920 & n27054 ;
  assign n27056 = n27055 ^ n24030 ;
  assign n27057 = n27056 ^ n26917 ;
  assign n27058 = ~n26918 & ~n27057 ;
  assign n27059 = n27058 ^ n24076 ;
  assign n26916 = n26902 ^ n26620 ;
  assign n27060 = n27059 ^ n26916 ;
  assign n27061 = n27059 ^ n24122 ;
  assign n27062 = ~n27060 & ~n27061 ;
  assign n27063 = n27062 ^ n24242 ;
  assign n27064 = n26915 & n27063 ;
  assign n27065 = n27064 ^ n26914 ;
  assign n27152 = n27151 ^ n27065 ;
  assign n27066 = n27061 ^ n26916 ;
  assign n27119 = ~n27116 & n27118 ;
  assign n27120 = n27043 ^ n24766 ;
  assign n27121 = n27119 & ~n27120 ;
  assign n27122 = n27048 ^ n24781 ;
  assign n27123 = ~n27121 & ~n27122 ;
  assign n27124 = n27050 ^ n26922 ;
  assign n27125 = ~n27123 & ~n27124 ;
  assign n27126 = n27053 ^ n24030 ;
  assign n27127 = n27126 ^ n26919 ;
  assign n27128 = n27125 & n27127 ;
  assign n27129 = n27056 ^ n26918 ;
  assign n27130 = n27128 & n27129 ;
  assign n27131 = n27066 & ~n27130 ;
  assign n27132 = n27063 ^ n26914 ;
  assign n27133 = ~n27131 & ~n27132 ;
  assign n27153 = n27152 ^ n27133 ;
  assign n27154 = n27153 ^ n3190 ;
  assign n27155 = n27132 ^ n27131 ;
  assign n27156 = n27155 ^ n2522 ;
  assign n27159 = n27130 ^ n27066 ;
  assign n27160 = n27159 ^ n3218 ;
  assign n27161 = n27129 ^ n27128 ;
  assign n2571 = n2570 ^ n2486 ;
  assign n2578 = n2577 ^ n2571 ;
  assign n2582 = n2581 ^ n2578 ;
  assign n27162 = n27161 ^ n2582 ;
  assign n27166 = n25366 ^ n2624 ;
  assign n27167 = n27166 ^ n2872 ;
  assign n27168 = n27167 ^ n2575 ;
  assign n27165 = n27127 ^ n27125 ;
  assign n27169 = n27168 ^ n27165 ;
  assign n27170 = n27124 ^ n27123 ;
  assign n2862 = n2822 ^ n2553 ;
  assign n2863 = n2862 ^ n2861 ;
  assign n2867 = n2866 ^ n2863 ;
  assign n27171 = n27170 ^ n2867 ;
  assign n27172 = n27122 ^ n27121 ;
  assign n27173 = n27172 ^ n2811 ;
  assign n27174 = n27120 ^ n27119 ;
  assign n27175 = n27174 ^ n1435 ;
  assign n27314 = n27311 ^ n1410 ;
  assign n27315 = ~n27313 & n27314 ;
  assign n27316 = n27315 ^ n1410 ;
  assign n27317 = n27316 ^ n1435 ;
  assign n27318 = n27175 & ~n27317 ;
  assign n27319 = n27318 ^ n27174 ;
  assign n27320 = n27319 ^ n2811 ;
  assign n27321 = n27173 & ~n27320 ;
  assign n27322 = n27321 ^ n27172 ;
  assign n27323 = n27322 ^ n27170 ;
  assign n27324 = ~n27171 & n27323 ;
  assign n27325 = n27324 ^ n2867 ;
  assign n27326 = n27325 ^ n27165 ;
  assign n27327 = ~n27169 & n27326 ;
  assign n27328 = n27327 ^ n27168 ;
  assign n27163 = n27159 ^ n2582 ;
  assign n27164 = n27163 ^ n27159 ;
  assign n27329 = n27328 ^ n27164 ;
  assign n27330 = ~n27162 & n27329 ;
  assign n27331 = n27330 ^ n27163 ;
  assign n27332 = ~n27160 & n27331 ;
  assign n27333 = n27332 ^ n3218 ;
  assign n27157 = n27153 ^ n2522 ;
  assign n27158 = n27157 ^ n27153 ;
  assign n27334 = n27333 ^ n27158 ;
  assign n27335 = ~n27156 & n27334 ;
  assign n27336 = n27335 ^ n27157 ;
  assign n27337 = n27154 & ~n27336 ;
  assign n27145 = n26575 ^ n26444 ;
  assign n27143 = n24739 ^ n24702 ;
  assign n27144 = n27143 ^ n26081 ;
  assign n27146 = n27145 ^ n27144 ;
  assign n27142 = n26612 ^ n24247 ;
  assign n27147 = n27146 ^ n27142 ;
  assign n27135 = n27134 ^ n27133 ;
  assign n27138 = n27133 ^ n27065 ;
  assign n27139 = n27135 & ~n27138 ;
  assign n27136 = n27135 ^ n27065 ;
  assign n27137 = ~n24214 & n27136 ;
  assign n27140 = n27139 ^ n27137 ;
  assign n3181 = n3176 ^ n3161 ;
  assign n3182 = n3181 ^ n2696 ;
  assign n3183 = n3182 ^ n1811 ;
  assign n27141 = n27140 ^ n3183 ;
  assign n27148 = n27147 ^ n27141 ;
  assign n27149 = n27148 ^ n3190 ;
  assign n26911 = n26910 ^ n26612 ;
  assign n26912 = n26614 & ~n26911 ;
  assign n27150 = n27149 ^ n26912 ;
  assign n27338 = n27337 ^ n27150 ;
  assign n26609 = n26608 ^ n25151 ;
  assign n26610 = n26609 ^ n26176 ;
  assign n27339 = n27338 ^ n26610 ;
  assign n27342 = n27336 ^ n3190 ;
  assign n27340 = n26683 ^ n25153 ;
  assign n27341 = n27340 ^ n26180 ;
  assign n27343 = n27342 ^ n27341 ;
  assign n27345 = n26687 ^ n25157 ;
  assign n27346 = n27345 ^ n26184 ;
  assign n27361 = n27346 ^ n27341 ;
  assign n27344 = n27333 ^ n27156 ;
  assign n27347 = n27346 ^ n27344 ;
  assign n27352 = n27331 ^ n3218 ;
  assign n27358 = n27352 ^ n27344 ;
  assign n27348 = n26693 ^ n26192 ;
  assign n27349 = n27348 ^ n25165 ;
  assign n27350 = n27328 ^ n27162 ;
  assign n27351 = ~n27349 & ~n27350 ;
  assign n27353 = n27352 ^ n27351 ;
  assign n27354 = n26691 ^ n25163 ;
  assign n27355 = n27354 ^ n26188 ;
  assign n27356 = n27355 ^ n27351 ;
  assign n27357 = ~n27353 & ~n27356 ;
  assign n27359 = n27358 ^ n27357 ;
  assign n27360 = n27347 & ~n27359 ;
  assign n27362 = n27361 ^ n27360 ;
  assign n27363 = ~n27343 & ~n27362 ;
  assign n27364 = n27363 ^ n27342 ;
  assign n27365 = n27364 ^ n26610 ;
  assign n27366 = ~n27339 & ~n27365 ;
  assign n27367 = n27366 ^ n27338 ;
  assign n27368 = n27367 ^ n26134 ;
  assign n27369 = ~n26606 & n27368 ;
  assign n27370 = n27369 ^ n26605 ;
  assign n27407 = n27372 ^ n27370 ;
  assign n27408 = n27374 & ~n27407 ;
  assign n27409 = n27408 ^ n27373 ;
  assign n27414 = n27413 ^ n27409 ;
  assign n27415 = n27414 ^ n24706 ;
  assign n27375 = n27374 ^ n27370 ;
  assign n27376 = n27375 ^ n24852 ;
  assign n27399 = n27367 ^ n26606 ;
  assign n27377 = n27364 ^ n27339 ;
  assign n27378 = n27377 ^ n24716 ;
  assign n27379 = n27362 ^ n27342 ;
  assign n27380 = n27379 ^ n24720 ;
  assign n27388 = n27359 ^ n27346 ;
  assign n27381 = n27350 ^ n27349 ;
  assign n27382 = ~n24733 & n27381 ;
  assign n27383 = n27382 ^ n24129 ;
  assign n27384 = n27356 ^ n27352 ;
  assign n27385 = n27384 ^ n27382 ;
  assign n27386 = ~n27383 & n27385 ;
  assign n27387 = n27386 ^ n24129 ;
  assign n27389 = n27388 ^ n27387 ;
  assign n27390 = n27388 ^ n24724 ;
  assign n27391 = ~n27389 & ~n27390 ;
  assign n27392 = n27391 ^ n24724 ;
  assign n27393 = n27392 ^ n27379 ;
  assign n27394 = ~n27380 & ~n27393 ;
  assign n27395 = n27394 ^ n24720 ;
  assign n27396 = n27395 ^ n27377 ;
  assign n27397 = n27378 & ~n27396 ;
  assign n27398 = n27397 ^ n24716 ;
  assign n27400 = n27399 ^ n27398 ;
  assign n27401 = n27399 ^ n24710 ;
  assign n27402 = n27400 & n27401 ;
  assign n27403 = n27402 ^ n24710 ;
  assign n27404 = n27403 ^ n27375 ;
  assign n27405 = n27376 & n27404 ;
  assign n27406 = n27405 ^ n24852 ;
  assign n27488 = n27414 ^ n27406 ;
  assign n27489 = ~n27415 & ~n27488 ;
  assign n27490 = n27489 ^ n24706 ;
  assign n27485 = n27246 ^ n27243 ;
  assign n27481 = n26662 ^ n26161 ;
  assign n27482 = n27481 ^ n25132 ;
  assign n27483 = n27482 ^ n27412 ;
  assign n27479 = n27412 ^ n27409 ;
  assign n27480 = n27413 & ~n27479 ;
  assign n27484 = n27483 ^ n27480 ;
  assign n27486 = n27485 ^ n27484 ;
  assign n27487 = n27486 ^ n24860 ;
  assign n27491 = n27490 ^ n27487 ;
  assign n27416 = n27415 ^ n27406 ;
  assign n27417 = n27398 ^ n24710 ;
  assign n27418 = n27417 ^ n27399 ;
  assign n27419 = n27381 ^ n24733 ;
  assign n27420 = n27384 ^ n27383 ;
  assign n27421 = ~n27419 & n27420 ;
  assign n27422 = n27390 ^ n27387 ;
  assign n27423 = n27421 & n27422 ;
  assign n27424 = n27392 ^ n27380 ;
  assign n27425 = n27423 & ~n27424 ;
  assign n27426 = n27395 ^ n27378 ;
  assign n27427 = n27425 & ~n27426 ;
  assign n27428 = n27418 & ~n27427 ;
  assign n27429 = n27403 ^ n27376 ;
  assign n27430 = ~n27428 & n27429 ;
  assign n27492 = ~n27416 & ~n27430 ;
  assign n27497 = n27491 & n27492 ;
  assign n27498 = n27490 ^ n27486 ;
  assign n27503 = n26664 ^ n26155 ;
  assign n27504 = n27503 ^ n25134 ;
  assign n27502 = n27248 ^ n27223 ;
  assign n27505 = n27504 ^ n27502 ;
  assign n27499 = n27485 ^ n27482 ;
  assign n27500 = n27484 & ~n27499 ;
  assign n27501 = n27500 ^ n27482 ;
  assign n27506 = n27505 ^ n27501 ;
  assign n27507 = n27506 ^ n24860 ;
  assign n27508 = n27507 ^ n27486 ;
  assign n27509 = n27508 ^ n27506 ;
  assign n27510 = n27498 & ~n27509 ;
  assign n27511 = n27510 ^ n27507 ;
  assign n27512 = n27511 ^ n25074 ;
  assign n27715 = n27497 & n27512 ;
  assign n27576 = n27252 ^ n27217 ;
  assign n27569 = n26833 ^ n25520 ;
  assign n27570 = n27569 ^ n26151 ;
  assign n27571 = n27570 ^ n27502 ;
  assign n27572 = n27571 ^ n27570 ;
  assign n27573 = n27572 ^ n27501 ;
  assign n27574 = n27505 & ~n27573 ;
  assign n27575 = n27574 ^ n27571 ;
  assign n27644 = n27576 ^ n27575 ;
  assign n27647 = n27644 ^ n25074 ;
  assign n27646 = n27644 ^ n27506 ;
  assign n27648 = n27647 ^ n27646 ;
  assign n27649 = ~n27511 & ~n27648 ;
  assign n27650 = n27649 ^ n27647 ;
  assign n27716 = n27650 ^ n25091 ;
  assign n27717 = ~n27715 & n27716 ;
  assign n27645 = n27644 ^ n25091 ;
  assign n27651 = ~n27645 & ~n27650 ;
  assign n27652 = n27651 ^ n25091 ;
  assign n27718 = n27652 ^ n25141 ;
  assign n27583 = n26841 ^ n26147 ;
  assign n27584 = n27583 ^ n25535 ;
  assign n27577 = n27254 ^ n27216 ;
  assign n27579 = n27577 ^ n27570 ;
  assign n27578 = n27577 ^ n27576 ;
  assign n27580 = n27579 ^ n27578 ;
  assign n27581 = n27575 & n27580 ;
  assign n27582 = n27581 ^ n27579 ;
  assign n27642 = n27584 ^ n27582 ;
  assign n27719 = n27718 ^ n27642 ;
  assign n27720 = ~n27717 & ~n27719 ;
  assign n27643 = n27642 ^ n25141 ;
  assign n27653 = n27652 ^ n27642 ;
  assign n27654 = n27643 & ~n27653 ;
  assign n27655 = n27654 ^ n25141 ;
  assign n27564 = n26860 ^ n25127 ;
  assign n27565 = n27564 ^ n26145 ;
  assign n27587 = n27577 ^ n27565 ;
  assign n27585 = n27584 ^ n27577 ;
  assign n27586 = ~n27582 & ~n27585 ;
  assign n27588 = n27587 ^ n27586 ;
  assign n27566 = n27259 ^ n2305 ;
  assign n27567 = n27566 ^ n27257 ;
  assign n27640 = n27588 ^ n27567 ;
  assign n27641 = n27640 ^ n25135 ;
  assign n27721 = n27655 ^ n27641 ;
  assign n27722 = ~n27720 & ~n27721 ;
  assign n27562 = n27265 ^ n27264 ;
  assign n27590 = n27567 ^ n27562 ;
  assign n27568 = n27567 ^ n27565 ;
  assign n27589 = n27568 & ~n27588 ;
  assign n27591 = n27590 ^ n27589 ;
  assign n27560 = n26868 ^ n26139 ;
  assign n27561 = n27560 ^ n25119 ;
  assign n27639 = n27591 ^ n27561 ;
  assign n27723 = n27639 ^ n25129 ;
  assign n27656 = n27655 ^ n27640 ;
  assign n27657 = ~n27641 & ~n27656 ;
  assign n27658 = n27657 ^ n25135 ;
  assign n27724 = n27723 ^ n27658 ;
  assign n27725 = ~n27722 & ~n27724 ;
  assign n27659 = n27658 ^ n27639 ;
  assign n27558 = n27269 ^ n27213 ;
  assign n27593 = n27562 ^ n27558 ;
  assign n27563 = n27562 ^ n27561 ;
  assign n27592 = n27563 & n27591 ;
  assign n27594 = n27593 ^ n27592 ;
  assign n27556 = n26874 ^ n26137 ;
  assign n27557 = n27556 ^ n25114 ;
  assign n27637 = n27594 ^ n27557 ;
  assign n27660 = n27637 ^ n25129 ;
  assign n27661 = n27660 ^ n27637 ;
  assign n27662 = n27661 ^ n27639 ;
  assign n27663 = n27659 & ~n27662 ;
  assign n27664 = n27663 ^ n27660 ;
  assign n27726 = n27664 ^ n25200 ;
  assign n27727 = n27725 & ~n27726 ;
  assign n27638 = n27637 ^ n25200 ;
  assign n27665 = ~n27638 & ~n27664 ;
  assign n27666 = n27665 ^ n25200 ;
  assign n27559 = n27558 ^ n27557 ;
  assign n27595 = ~n27559 & ~n27594 ;
  assign n27596 = n27595 ^ n27558 ;
  assign n27554 = n27271 ^ n27209 ;
  assign n27552 = n26658 ^ n26249 ;
  assign n27553 = n27552 ^ n25104 ;
  assign n27555 = n27554 ^ n27553 ;
  assign n27635 = n27596 ^ n27555 ;
  assign n27636 = n27635 ^ n25231 ;
  assign n27728 = n27666 ^ n27636 ;
  assign n27729 = n27727 & n27728 ;
  assign n27597 = n27596 ^ n27553 ;
  assign n27598 = ~n27555 & ~n27597 ;
  assign n27599 = n27598 ^ n27554 ;
  assign n27549 = n26350 ^ n25554 ;
  assign n27550 = n27549 ^ n26654 ;
  assign n27517 = n27274 ^ n27204 ;
  assign n27551 = n27550 ^ n27517 ;
  assign n27670 = n27599 ^ n27551 ;
  assign n27672 = n27670 ^ n25232 ;
  assign n27667 = n27666 ^ n27635 ;
  assign n27668 = ~n27636 & ~n27667 ;
  assign n27669 = n27668 ^ n25231 ;
  assign n27714 = n27672 ^ n27669 ;
  assign n27782 = n27729 ^ n27714 ;
  assign n27783 = n27782 ^ n1606 ;
  assign n27828 = n2969 ^ n1606 ;
  assign n27824 = n27728 ^ n27727 ;
  assign n27787 = n27726 ^ n27725 ;
  assign n27788 = n27787 ^ n27786 ;
  assign n27789 = n27724 ^ n27722 ;
  assign n27790 = n27789 ^ n608 ;
  assign n27791 = n27721 ^ n27720 ;
  assign n27795 = n27794 ^ n27791 ;
  assign n27796 = n27719 ^ n27717 ;
  assign n27800 = n27799 ^ n27796 ;
  assign n27804 = n27716 ^ n27715 ;
  assign n27805 = n27804 ^ n27803 ;
  assign n27513 = n27512 ^ n27497 ;
  assign n2416 = n2385 ^ n2340 ;
  assign n2417 = n2416 ^ n2402 ;
  assign n2421 = n2420 ^ n2417 ;
  assign n27514 = n27513 ^ n2421 ;
  assign n27493 = n27492 ^ n27491 ;
  assign n27431 = n27430 ^ n27416 ;
  assign n2403 = n2330 ^ n2266 ;
  assign n2410 = n2409 ^ n2403 ;
  assign n2411 = n2410 ^ n2204 ;
  assign n27432 = n27431 ^ n2411 ;
  assign n27434 = n25842 ^ n2240 ;
  assign n27435 = n27434 ^ n2081 ;
  assign n27436 = n27435 ^ n2406 ;
  assign n27433 = n27429 ^ n27428 ;
  assign n27437 = n27436 ^ n27433 ;
  assign n27460 = n27427 ^ n27418 ;
  assign n27472 = n27460 ^ n27433 ;
  assign n1912 = n1905 ^ n1890 ;
  assign n1919 = n1918 ^ n1912 ;
  assign n1923 = n1922 ^ n1919 ;
  assign n27443 = n3032 ^ n1923 ;
  assign n27438 = n27420 ^ n27419 ;
  assign n27439 = n27438 ^ n3032 ;
  assign n27440 = n3240 & n27419 ;
  assign n27441 = n27440 ^ n27438 ;
  assign n27442 = ~n27439 & n27441 ;
  assign n27444 = n27443 ^ n27442 ;
  assign n27446 = n25850 ^ n18828 ;
  assign n27447 = n27446 ^ n1927 ;
  assign n27448 = n27447 ^ n1981 ;
  assign n27450 = n27448 ^ n1923 ;
  assign n27445 = n27422 ^ n27421 ;
  assign n27449 = n27448 ^ n27445 ;
  assign n27451 = n27450 ^ n27449 ;
  assign n27452 = n27444 & n27451 ;
  assign n27453 = n27452 ^ n27450 ;
  assign n1977 = n1976 ^ n1943 ;
  assign n1984 = n1983 ^ n1977 ;
  assign n1988 = n1987 ^ n1984 ;
  assign n27456 = n27448 ^ n1988 ;
  assign n27454 = n27424 ^ n27423 ;
  assign n27455 = n27454 ^ n1988 ;
  assign n27457 = n27456 ^ n27455 ;
  assign n27458 = n27453 & ~n27457 ;
  assign n27459 = n27458 ^ n27456 ;
  assign n27463 = n27460 ^ n1988 ;
  assign n27461 = n27426 ^ n27425 ;
  assign n27462 = n27461 ^ n27460 ;
  assign n27464 = n27463 ^ n27462 ;
  assign n27465 = n27459 & ~n27464 ;
  assign n27466 = n27465 ^ n27463 ;
  assign n27467 = n25868 ^ n2247 ;
  assign n27468 = n27467 ^ n22319 ;
  assign n27469 = n27468 ^ n2079 ;
  assign n27470 = n27469 ^ n27460 ;
  assign n27471 = n27466 & n27470 ;
  assign n27473 = n27472 ^ n27471 ;
  assign n27474 = ~n27437 & n27473 ;
  assign n27475 = n27474 ^ n27436 ;
  assign n27476 = n27475 ^ n27431 ;
  assign n27477 = ~n27432 & n27476 ;
  assign n27478 = n27477 ^ n2411 ;
  assign n27494 = n27493 ^ n27478 ;
  assign n27495 = n27478 ^ n2421 ;
  assign n27496 = n27494 & n27495 ;
  assign n27515 = n27514 ^ n27496 ;
  assign n2437 = n2356 ^ n1466 ;
  assign n2438 = n2437 ^ n2428 ;
  assign n2439 = n2438 ^ n2436 ;
  assign n27806 = n27513 ^ n2439 ;
  assign n27807 = n27515 & ~n27806 ;
  assign n27808 = n27807 ^ n2439 ;
  assign n27809 = n27808 ^ n27803 ;
  assign n27810 = ~n27805 & ~n27809 ;
  assign n27811 = n27810 ^ n27804 ;
  assign n27812 = n27811 ^ n27796 ;
  assign n27813 = ~n27800 & ~n27812 ;
  assign n27814 = n27813 ^ n27799 ;
  assign n27815 = n27814 ^ n27791 ;
  assign n27816 = n27795 & ~n27815 ;
  assign n27817 = n27816 ^ n27794 ;
  assign n27818 = n27817 ^ n27789 ;
  assign n27819 = ~n27790 & n27818 ;
  assign n27820 = n27819 ^ n608 ;
  assign n27821 = n27820 ^ n27786 ;
  assign n27822 = n27788 & ~n27821 ;
  assign n27823 = n27822 ^ n27787 ;
  assign n27825 = n27824 ^ n27823 ;
  assign n27826 = n27823 ^ n2969 ;
  assign n27827 = n27825 & n27826 ;
  assign n27829 = n27828 ^ n27827 ;
  assign n27830 = n27783 & n27829 ;
  assign n27832 = n27831 ^ n27830 ;
  assign n27730 = ~n27714 & n27729 ;
  assign n27671 = n27670 ^ n27669 ;
  assign n27673 = n27671 & ~n27672 ;
  assign n27674 = n27673 ^ n25232 ;
  assign n27547 = n27278 ^ n27201 ;
  assign n27602 = n27547 ^ n27517 ;
  assign n27600 = n27599 ^ n27550 ;
  assign n27601 = n27551 & ~n27600 ;
  assign n27603 = n27602 ^ n27601 ;
  assign n27545 = n26644 ^ n26398 ;
  assign n27546 = n27545 ^ n25559 ;
  assign n27633 = n27603 ^ n27546 ;
  assign n27634 = n27633 ^ n25124 ;
  assign n27713 = n27674 ^ n27634 ;
  assign n27780 = n27730 ^ n27713 ;
  assign n28129 = n27832 ^ n27780 ;
  assign n28130 = n28129 ^ n26637 ;
  assign n28131 = n28130 ^ n27892 ;
  assign n28132 = n28131 ^ n28129 ;
  assign n28133 = ~n28128 & ~n28132 ;
  assign n28134 = n28133 ^ n28130 ;
  assign n27917 = n27316 ^ n27175 ;
  assign n28297 = n27917 ^ n26613 ;
  assign n28298 = n26633 ^ n26613 ;
  assign n28299 = n28297 & n28298 ;
  assign n28300 = n28299 ^ n26633 ;
  assign n28302 = n28300 ^ n28129 ;
  assign n28136 = n26646 ^ n26619 ;
  assign n27766 = n27309 ^ n27176 ;
  assign n28137 = n27766 ^ n26619 ;
  assign n28138 = ~n28136 & n28137 ;
  assign n28139 = n28138 ^ n26646 ;
  assign n28135 = n27829 ^ n27782 ;
  assign n28140 = n28139 ^ n28135 ;
  assign n27750 = n27305 ^ n27303 ;
  assign n28141 = n27750 ^ n26623 ;
  assign n28142 = n27825 ^ n2969 ;
  assign n28143 = n28142 ^ n26583 ;
  assign n28144 = n28143 ^ n26623 ;
  assign n28145 = n28144 ^ n28142 ;
  assign n28146 = n28141 & ~n28145 ;
  assign n28147 = n28146 ^ n28143 ;
  assign n28282 = n27820 ^ n27788 ;
  assign n27621 = n27297 ^ n852 ;
  assign n28150 = n27621 ^ n26635 ;
  assign n28155 = n27814 ^ n27795 ;
  assign n27525 = n27293 ^ n27292 ;
  assign n28151 = n27525 ^ n26640 ;
  assign n28152 = n27525 ^ n26398 ;
  assign n28153 = n28151 & n28152 ;
  assign n28154 = n28153 ^ n26398 ;
  assign n28156 = n28155 ^ n28154 ;
  assign n27527 = n27289 ^ n27183 ;
  assign n28159 = n27527 ^ n26888 ;
  assign n28160 = n27527 ^ n26350 ;
  assign n28161 = n28159 & ~n28160 ;
  assign n28162 = n28161 ^ n26350 ;
  assign n28157 = n27811 ^ n27800 ;
  assign n28163 = n28162 ^ n28157 ;
  assign n27536 = n27283 ^ n27192 ;
  assign n28164 = n27536 ^ n26654 ;
  assign n27516 = n27515 ^ n2439 ;
  assign n28165 = n27516 ^ n26137 ;
  assign n28166 = n28165 ^ n26654 ;
  assign n28167 = n28166 ^ n27516 ;
  assign n28168 = n28164 & n28167 ;
  assign n28169 = n28168 ^ n28165 ;
  assign n28177 = n27494 ^ n2421 ;
  assign n27543 = n27280 ^ n27197 ;
  assign n28173 = n27543 ^ n26658 ;
  assign n28174 = n26658 ^ n26139 ;
  assign n28175 = n28173 & ~n28174 ;
  assign n28176 = n28175 ^ n26139 ;
  assign n28178 = n28177 ^ n28176 ;
  assign n28179 = n27547 ^ n26874 ;
  assign n28180 = n26874 ^ n26145 ;
  assign n28181 = ~n28179 & ~n28180 ;
  assign n28182 = n28181 ^ n26145 ;
  assign n28075 = n27475 ^ n27432 ;
  assign n28183 = n28182 ^ n28075 ;
  assign n28184 = n26868 ^ n26147 ;
  assign n28185 = n27517 ^ n26868 ;
  assign n28186 = ~n28184 & n28185 ;
  assign n28187 = n28186 ^ n26147 ;
  assign n28082 = n27473 ^ n27436 ;
  assign n28188 = n28187 ^ n28082 ;
  assign n28189 = n27554 ^ n26860 ;
  assign n28090 = n27469 ^ n27466 ;
  assign n28190 = n28090 ^ n26151 ;
  assign n28191 = n28190 ^ n27554 ;
  assign n28192 = n28191 ^ n28090 ;
  assign n28193 = n28189 & ~n28192 ;
  assign n28194 = n28193 ^ n28190 ;
  assign n28195 = n26841 ^ n26155 ;
  assign n28196 = n27558 ^ n26841 ;
  assign n28197 = ~n28195 & ~n28196 ;
  assign n28198 = n28197 ^ n26155 ;
  assign n28100 = n27461 ^ n27459 ;
  assign n28199 = n28198 ^ n28100 ;
  assign n28201 = n27454 ^ n27453 ;
  assign n28241 = n28201 ^ n28100 ;
  assign n28200 = n27562 ^ n26833 ;
  assign n28202 = n28201 ^ n26161 ;
  assign n28203 = n28202 ^ n27562 ;
  assign n28204 = n28203 ^ n28201 ;
  assign n28205 = ~n28200 & ~n28204 ;
  assign n28206 = n28205 ^ n28202 ;
  assign n28211 = n27445 ^ n27444 ;
  assign n28207 = n26664 ^ n26165 ;
  assign n28208 = n27567 ^ n26664 ;
  assign n28209 = ~n28207 & ~n28208 ;
  assign n28210 = n28209 ^ n26165 ;
  assign n28212 = n28211 ^ n28210 ;
  assign n28225 = n27440 ^ n3032 ;
  assign n28226 = n28225 ^ n27438 ;
  assign n28217 = n27419 ^ n3240 ;
  assign n28213 = n26669 ^ n26133 ;
  assign n28214 = n27576 ^ n26669 ;
  assign n28215 = ~n28213 & ~n28214 ;
  assign n28216 = n28215 ^ n26133 ;
  assign n28218 = n28217 ^ n28216 ;
  assign n27975 = n27485 ^ n26131 ;
  assign n27519 = n27373 ^ n26683 ;
  assign n27748 = n25952 ^ n25467 ;
  assign n27749 = n27748 ^ n26613 ;
  assign n27751 = n27750 ^ n27749 ;
  assign n27759 = n27145 ^ n25978 ;
  assign n27760 = n27759 ^ n25470 ;
  assign n27761 = n27760 ^ n27750 ;
  assign n27762 = n27761 ^ n27760 ;
  assign n27700 = n27299 ^ n27179 ;
  assign n27701 = n27700 ^ n27621 ;
  assign n27619 = n26633 ^ n26035 ;
  assign n27620 = n27619 ^ n26619 ;
  assign n27622 = n27621 ^ n27620 ;
  assign n27523 = n26623 ^ n25989 ;
  assign n27524 = n27523 ^ n26637 ;
  assign n27526 = n27525 ^ n27524 ;
  assign n27529 = n26646 ^ n26628 ;
  assign n27530 = n27529 ^ n25961 ;
  assign n27531 = n27530 ^ n27527 ;
  assign n27534 = n27287 ^ n27188 ;
  assign n27532 = n26635 ^ n26583 ;
  assign n27533 = n27532 ^ n25779 ;
  assign n27535 = n27534 ^ n27533 ;
  assign n27538 = n26429 ^ n25767 ;
  assign n27539 = n27538 ^ n26640 ;
  assign n27540 = n27539 ^ n27536 ;
  assign n27541 = n26888 ^ n26413 ;
  assign n27542 = n27541 ^ n25694 ;
  assign n27544 = n27543 ^ n27542 ;
  assign n27548 = n27547 ^ n27546 ;
  assign n27604 = ~n27548 & ~n27603 ;
  assign n27605 = n27604 ^ n27547 ;
  assign n27606 = n27605 ^ n27542 ;
  assign n27607 = n27544 & ~n27606 ;
  assign n27608 = n27607 ^ n27543 ;
  assign n27609 = n27608 ^ n27536 ;
  assign n27610 = ~n27540 & n27609 ;
  assign n27537 = n27536 ^ n27534 ;
  assign n27611 = n27610 ^ n27537 ;
  assign n27612 = n27535 & n27611 ;
  assign n27613 = n27612 ^ n27534 ;
  assign n27614 = n27613 ^ n27527 ;
  assign n27615 = ~n27531 & ~n27614 ;
  assign n27528 = n27527 ^ n27525 ;
  assign n27616 = n27615 ^ n27528 ;
  assign n27617 = n27526 & ~n27616 ;
  assign n27618 = n27617 ^ n27525 ;
  assign n27698 = n27621 ^ n27618 ;
  assign n27699 = n27622 & n27698 ;
  assign n27702 = n27701 ^ n27699 ;
  assign n27703 = n26626 ^ n26068 ;
  assign n27704 = n27703 ^ n26907 ;
  assign n27745 = n27704 ^ n27700 ;
  assign n27746 = ~n27702 & n27745 ;
  assign n27747 = n27746 ^ n27704 ;
  assign n27763 = n27762 ^ n27747 ;
  assign n27764 = ~n27751 & ~n27763 ;
  assign n27765 = n27764 ^ n27761 ;
  assign n27885 = n26003 ^ n25460 ;
  assign n27886 = n27885 ^ n26600 ;
  assign n27888 = n27886 ^ n27760 ;
  assign n27887 = n27886 ^ n27766 ;
  assign n27889 = n27888 ^ n27887 ;
  assign n27890 = ~n27765 & ~n27889 ;
  assign n27891 = n27890 ^ n27888 ;
  assign n27893 = n27892 ^ n27891 ;
  assign n27894 = n27893 ^ n24815 ;
  assign n27767 = n27766 ^ n27765 ;
  assign n27768 = n27767 ^ n24679 ;
  assign n27752 = n27751 ^ n27747 ;
  assign n27753 = n27752 ^ n24682 ;
  assign n27705 = n27704 ^ n27702 ;
  assign n27706 = n27705 ^ n25443 ;
  assign n27624 = n27616 ^ n27524 ;
  assign n27625 = n27624 ^ n25176 ;
  assign n27627 = n27611 ^ n27533 ;
  assign n27628 = n27627 ^ n25105 ;
  assign n27629 = n27608 ^ n27540 ;
  assign n27630 = n27629 ^ n25115 ;
  assign n27631 = n27605 ^ n27544 ;
  assign n27632 = n27631 ^ n25120 ;
  assign n27675 = n27674 ^ n27633 ;
  assign n27676 = ~n27634 & ~n27675 ;
  assign n27677 = n27676 ^ n25124 ;
  assign n27678 = n27677 ^ n27631 ;
  assign n27679 = n27632 & n27678 ;
  assign n27680 = n27679 ^ n25120 ;
  assign n27681 = n27680 ^ n27629 ;
  assign n27682 = ~n27630 & n27681 ;
  assign n27683 = n27682 ^ n25115 ;
  assign n27684 = n27683 ^ n27627 ;
  assign n27685 = ~n27628 & ~n27684 ;
  assign n27686 = n27685 ^ n25105 ;
  assign n27626 = n27613 ^ n27531 ;
  assign n27687 = n27686 ^ n27626 ;
  assign n27688 = n27686 ^ n25109 ;
  assign n27689 = ~n27687 & ~n27688 ;
  assign n27690 = n27689 ^ n25109 ;
  assign n27691 = n27690 ^ n27624 ;
  assign n27692 = ~n27625 & n27691 ;
  assign n27693 = n27692 ^ n25176 ;
  assign n27623 = n27622 ^ n27618 ;
  assign n27694 = n27693 ^ n27623 ;
  assign n27695 = n27693 ^ n25180 ;
  assign n27696 = ~n27694 & n27695 ;
  assign n27697 = n27696 ^ n25180 ;
  assign n27742 = n27705 ^ n27697 ;
  assign n27743 = ~n27706 & ~n27742 ;
  assign n27744 = n27743 ^ n25443 ;
  assign n27756 = n27752 ^ n27744 ;
  assign n27757 = n27753 & ~n27756 ;
  assign n27758 = n27757 ^ n24682 ;
  assign n27882 = n27767 ^ n27758 ;
  assign n27883 = ~n27768 & n27882 ;
  assign n27884 = n27883 ^ n24679 ;
  assign n27895 = n27894 ^ n27884 ;
  assign n27707 = n27706 ^ n27697 ;
  assign n27708 = n27623 ^ n25180 ;
  assign n27709 = n27708 ^ n27693 ;
  assign n27710 = n27690 ^ n27625 ;
  assign n27711 = n27626 ^ n25109 ;
  assign n27712 = n27711 ^ n27686 ;
  assign n27731 = n27713 & ~n27730 ;
  assign n27732 = n27677 ^ n27632 ;
  assign n27733 = n27731 & n27732 ;
  assign n27734 = n27680 ^ n27630 ;
  assign n27735 = ~n27733 & ~n27734 ;
  assign n27736 = n27683 ^ n27628 ;
  assign n27737 = n27735 & ~n27736 ;
  assign n27738 = ~n27712 & ~n27737 ;
  assign n27739 = ~n27710 & ~n27738 ;
  assign n27740 = n27709 & n27739 ;
  assign n27741 = n27707 & ~n27740 ;
  assign n27754 = n27753 ^ n27744 ;
  assign n27755 = ~n27741 & ~n27754 ;
  assign n27769 = n27768 ^ n27758 ;
  assign n27881 = n27755 & n27769 ;
  assign n27896 = n27895 ^ n27881 ;
  assign n27770 = n27769 ^ n27755 ;
  assign n27520 = n18780 ^ n2894 ;
  assign n27521 = n27520 ^ n22741 ;
  assign n27522 = n27521 ^ n3092 ;
  assign n27771 = n27770 ^ n27522 ;
  assign n27859 = n2841 ^ n1385 ;
  assign n27860 = n27859 ^ n2639 ;
  assign n27861 = n27860 ^ n3203 ;
  assign n27847 = n27738 ^ n27710 ;
  assign n27772 = n27737 ^ n27712 ;
  assign n1085 = n1055 ^ n1003 ;
  assign n1086 = n1085 ^ n1082 ;
  assign n1090 = n1089 ^ n1086 ;
  assign n27773 = n27772 ^ n1090 ;
  assign n27843 = n27772 ^ n1078 ;
  assign n27774 = n27736 ^ n27735 ;
  assign n27775 = n27774 ^ n1078 ;
  assign n27776 = n27734 ^ n27733 ;
  assign n27777 = n27776 ^ n956 ;
  assign n27837 = n956 ^ n944 ;
  assign n27778 = n27732 ^ n27731 ;
  assign n27779 = n27778 ^ n944 ;
  assign n27781 = n27780 ^ n1615 ;
  assign n27833 = ~n27781 & ~n27832 ;
  assign n27834 = n27833 ^ n27780 ;
  assign n27835 = n27834 ^ n944 ;
  assign n27836 = n27779 & ~n27835 ;
  assign n27838 = n27837 ^ n27836 ;
  assign n27839 = ~n27777 & ~n27838 ;
  assign n27840 = n27839 ^ n27776 ;
  assign n27841 = n27840 ^ n1078 ;
  assign n27842 = n27775 & ~n27841 ;
  assign n27844 = n27843 ^ n27842 ;
  assign n27845 = n27773 & n27844 ;
  assign n27846 = n27845 ^ n27772 ;
  assign n27848 = n27847 ^ n27846 ;
  assign n27849 = n27846 ^ n1253 ;
  assign n27850 = n27848 & n27849 ;
  assign n27851 = n27850 ^ n1253 ;
  assign n27862 = n27861 ^ n27851 ;
  assign n27852 = n27739 ^ n27709 ;
  assign n27853 = n27852 ^ n27851 ;
  assign n27854 = n2834 ^ n1765 ;
  assign n27855 = n27854 ^ n1241 ;
  assign n27856 = n27855 ^ n2537 ;
  assign n27857 = n27856 ^ n27851 ;
  assign n27858 = ~n27853 & n27857 ;
  assign n27863 = n27862 ^ n27858 ;
  assign n27869 = n27867 ^ n27861 ;
  assign n27864 = n27740 ^ n27707 ;
  assign n27868 = n27867 ^ n27864 ;
  assign n27870 = n27869 ^ n27868 ;
  assign n27871 = n27863 & ~n27870 ;
  assign n27872 = n27871 ^ n27869 ;
  assign n27875 = n27867 ^ n27522 ;
  assign n27873 = n27754 ^ n27741 ;
  assign n27874 = n27873 ^ n27522 ;
  assign n27876 = n27875 ^ n27874 ;
  assign n27877 = n27872 & ~n27876 ;
  assign n27878 = n27877 ^ n27875 ;
  assign n27879 = ~n27771 & ~n27878 ;
  assign n27880 = n27879 ^ n27770 ;
  assign n27897 = n27896 ^ n27880 ;
  assign n3117 = n3116 ^ n2590 ;
  assign n3118 = n3117 ^ n3101 ;
  assign n3122 = n3121 ^ n3118 ;
  assign n27898 = n27897 ^ n3122 ;
  assign n27899 = n26687 ^ n26192 ;
  assign n27900 = n26605 ^ n26192 ;
  assign n27901 = n27899 & ~n27900 ;
  assign n27902 = n27901 ^ n26687 ;
  assign n27903 = n27898 & ~n27902 ;
  assign n27904 = n27903 ^ n26188 ;
  assign n27905 = n27904 ^ n27373 ;
  assign n27906 = n27905 ^ n27903 ;
  assign n27907 = ~n27519 & n27906 ;
  assign n27908 = n27907 ^ n27904 ;
  assign n27919 = n27893 ^ n27884 ;
  assign n27920 = ~n27894 & n27919 ;
  assign n27921 = n27920 ^ n24815 ;
  assign n27922 = n27921 ^ n24811 ;
  assign n27910 = n26787 ^ n25456 ;
  assign n27911 = n27910 ^ n26046 ;
  assign n27913 = n27911 ^ n27886 ;
  assign n27912 = n27911 ^ n27892 ;
  assign n27914 = n27913 ^ n27912 ;
  assign n27915 = ~n27891 & n27914 ;
  assign n27916 = n27915 ^ n27913 ;
  assign n27918 = n27917 ^ n27916 ;
  assign n27945 = n27921 ^ n27918 ;
  assign n27946 = ~n27922 & n27945 ;
  assign n27947 = n27946 ^ n24811 ;
  assign n27940 = n27917 ^ n27911 ;
  assign n27941 = ~n27916 & ~n27940 ;
  assign n27942 = n27941 ^ n27911 ;
  assign n27938 = n27319 ^ n27173 ;
  assign n27936 = n26081 ^ n25450 ;
  assign n27937 = n27936 ^ n26791 ;
  assign n27939 = n27938 ^ n27937 ;
  assign n27943 = n27942 ^ n27939 ;
  assign n27944 = n27943 ^ n24807 ;
  assign n27948 = n27947 ^ n27944 ;
  assign n27909 = n27881 & n27895 ;
  assign n27923 = n27922 ^ n27918 ;
  assign n27935 = ~n27909 & n27923 ;
  assign n27949 = n27948 ^ n27935 ;
  assign n27925 = n25949 ^ n2596 ;
  assign n27926 = n27925 ^ n22733 ;
  assign n27927 = n27926 ^ n1835 ;
  assign n27924 = n27923 ^ n27909 ;
  assign n27928 = n27927 ^ n27924 ;
  assign n27929 = n27880 ^ n3122 ;
  assign n27930 = ~n27897 & ~n27929 ;
  assign n27931 = n27930 ^ n3122 ;
  assign n27932 = n27931 ^ n27924 ;
  assign n27933 = ~n27928 & n27932 ;
  assign n27934 = n27933 ^ n27927 ;
  assign n27950 = n27949 ^ n27934 ;
  assign n2666 = n2607 ^ n2530 ;
  assign n2670 = n2669 ^ n2666 ;
  assign n2671 = n2670 ^ n2665 ;
  assign n27951 = n27950 ^ n2671 ;
  assign n27954 = n27951 ^ n27903 ;
  assign n27952 = n27931 ^ n27928 ;
  assign n27953 = n27952 ^ n27951 ;
  assign n27955 = n27954 ^ n27953 ;
  assign n27956 = ~n27908 & ~n27955 ;
  assign n27957 = n27956 ^ n27954 ;
  assign n27958 = n26608 ^ n26184 ;
  assign n27959 = n27412 ^ n26608 ;
  assign n27960 = ~n27958 & n27959 ;
  assign n27961 = n27960 ^ n26184 ;
  assign n27976 = n27961 ^ n27951 ;
  assign n27977 = n27957 & ~n27976 ;
  assign n27978 = n27977 ^ n27961 ;
  assign n27979 = n27978 ^ n26180 ;
  assign n27980 = n27979 ^ n27485 ;
  assign n27981 = n27980 ^ n27978 ;
  assign n27982 = n27975 & n27981 ;
  assign n27983 = n27982 ^ n27979 ;
  assign n27997 = ~n27935 & ~n27948 ;
  assign n27992 = n27947 ^ n24807 ;
  assign n27993 = ~n27944 & ~n27992 ;
  assign n27994 = n27993 ^ n24807 ;
  assign n27995 = n27994 ^ n24743 ;
  assign n27989 = n27322 ^ n27171 ;
  assign n27987 = n26799 ^ n25172 ;
  assign n27988 = n27987 ^ n26102 ;
  assign n27990 = n27989 ^ n27988 ;
  assign n27984 = n27942 ^ n27938 ;
  assign n27985 = ~n27939 & ~n27984 ;
  assign n27986 = n27985 ^ n27942 ;
  assign n27991 = n27990 ^ n27986 ;
  assign n27996 = n27995 ^ n27991 ;
  assign n27998 = n27997 ^ n27996 ;
  assign n27999 = n27998 ^ n2671 ;
  assign n28000 = n27999 ^ n27934 ;
  assign n28001 = n28000 ^ n27998 ;
  assign n28002 = n27950 & n28001 ;
  assign n28003 = n28002 ^ n27999 ;
  assign n28004 = n28003 ^ n2683 ;
  assign n28061 = n28004 ^ n27978 ;
  assign n28062 = n27983 & ~n28061 ;
  assign n28063 = n28062 ^ n28004 ;
  assign n28221 = n28217 ^ n28063 ;
  assign n28036 = n27502 ^ n26671 ;
  assign n28052 = n27998 ^ n2683 ;
  assign n28053 = n28003 & ~n28052 ;
  assign n28049 = n27994 ^ n27991 ;
  assign n28050 = n27995 & n28049 ;
  assign n28043 = n27325 ^ n27169 ;
  assign n28040 = n27143 ^ n2750 ;
  assign n28041 = n28040 ^ n26777 ;
  assign n28042 = n28041 ^ n26197 ;
  assign n28044 = n28043 ^ n28042 ;
  assign n28045 = n28044 ^ n24743 ;
  assign n28046 = n28045 ^ n2683 ;
  assign n28047 = n28046 ^ n27988 ;
  assign n28039 = n27996 & n27997 ;
  assign n28048 = n28047 ^ n28039 ;
  assign n28051 = n28050 ^ n28048 ;
  assign n28054 = n28053 ^ n28051 ;
  assign n28037 = n27988 ^ n27986 ;
  assign n28038 = n27990 & n28037 ;
  assign n28055 = n28054 ^ n28038 ;
  assign n28056 = n28055 ^ n26176 ;
  assign n28057 = n28056 ^ n27502 ;
  assign n28058 = n28057 ^ n28055 ;
  assign n28059 = ~n28036 & n28058 ;
  assign n28060 = n28059 ^ n28056 ;
  assign n28219 = n28063 ^ n28055 ;
  assign n28220 = ~n28060 & n28219 ;
  assign n28222 = n28221 ^ n28220 ;
  assign n28223 = n28218 & ~n28222 ;
  assign n28224 = n28223 ^ n28217 ;
  assign n28227 = n28226 ^ n28224 ;
  assign n28228 = n27577 ^ n26662 ;
  assign n28229 = n28226 ^ n26169 ;
  assign n28230 = n28229 ^ n27577 ;
  assign n28231 = n28230 ^ n28226 ;
  assign n28232 = n28228 & ~n28231 ;
  assign n28233 = n28232 ^ n28229 ;
  assign n28234 = ~n28227 & n28233 ;
  assign n28235 = n28234 ^ n28226 ;
  assign n28236 = n28235 ^ n28210 ;
  assign n28237 = ~n28212 & ~n28236 ;
  assign n28238 = n28237 ^ n28211 ;
  assign n28239 = n28238 ^ n28201 ;
  assign n28240 = n28206 & ~n28239 ;
  assign n28242 = n28241 ^ n28240 ;
  assign n28243 = ~n28199 & ~n28242 ;
  assign n28244 = n28243 ^ n28198 ;
  assign n28245 = n28244 ^ n28090 ;
  assign n28246 = ~n28194 & n28245 ;
  assign n28247 = n28246 ^ n28090 ;
  assign n28248 = n28247 ^ n28187 ;
  assign n28249 = ~n28188 & ~n28248 ;
  assign n28250 = n28249 ^ n28082 ;
  assign n28251 = n28250 ^ n28182 ;
  assign n28252 = ~n28183 & n28251 ;
  assign n28253 = n28252 ^ n28075 ;
  assign n28254 = n28253 ^ n28176 ;
  assign n28255 = n28178 & ~n28254 ;
  assign n28256 = n28255 ^ n28177 ;
  assign n28170 = n27808 ^ n27805 ;
  assign n28171 = n28170 ^ n27516 ;
  assign n28172 = n28171 ^ n28170 ;
  assign n28257 = n28256 ^ n28172 ;
  assign n28258 = ~n28169 & n28257 ;
  assign n28259 = n28258 ^ n28171 ;
  assign n28265 = n28170 ^ n28157 ;
  assign n28260 = n27534 ^ n26644 ;
  assign n28261 = n27534 ^ n26249 ;
  assign n28262 = ~n28260 & ~n28261 ;
  assign n28263 = n28262 ^ n26249 ;
  assign n28264 = n28263 ^ n28157 ;
  assign n28266 = n28265 ^ n28264 ;
  assign n28267 = n28259 & ~n28266 ;
  assign n28268 = n28267 ^ n28265 ;
  assign n28269 = ~n28163 & ~n28268 ;
  assign n28158 = n28157 ^ n28155 ;
  assign n28270 = n28269 ^ n28158 ;
  assign n28271 = ~n28156 & n28270 ;
  assign n28272 = n28271 ^ n28155 ;
  assign n28273 = n28272 ^ n26413 ;
  assign n28274 = n28273 ^ n26635 ;
  assign n28275 = n28274 ^ n28272 ;
  assign n28276 = ~n28150 & ~n28275 ;
  assign n28277 = n28276 ^ n28273 ;
  assign n28278 = n27817 ^ n27790 ;
  assign n28279 = n28278 ^ n28272 ;
  assign n28280 = ~n28277 & ~n28279 ;
  assign n28281 = n28280 ^ n28278 ;
  assign n28283 = n28282 ^ n28281 ;
  assign n28284 = n27700 ^ n26628 ;
  assign n28285 = n28282 ^ n26429 ;
  assign n28286 = n28285 ^ n26628 ;
  assign n28287 = n28286 ^ n28282 ;
  assign n28288 = ~n28284 & n28287 ;
  assign n28289 = n28288 ^ n28285 ;
  assign n28290 = ~n28283 & ~n28289 ;
  assign n28291 = n28290 ^ n28282 ;
  assign n28292 = n28291 ^ n28142 ;
  assign n28293 = ~n28147 & ~n28292 ;
  assign n28148 = n28142 ^ n28139 ;
  assign n28294 = n28293 ^ n28148 ;
  assign n28295 = n28140 & ~n28294 ;
  assign n28296 = n28295 ^ n28139 ;
  assign n28301 = n28300 ^ n28296 ;
  assign n28303 = n28302 ^ n28301 ;
  assign n28304 = n28134 & ~n28303 ;
  assign n28305 = n28304 ^ n28302 ;
  assign n28306 = n27938 ^ n27145 ;
  assign n28307 = n27145 ^ n26626 ;
  assign n28308 = ~n28306 & n28307 ;
  assign n28309 = n28308 ^ n26626 ;
  assign n28312 = n28309 ^ n28300 ;
  assign n28310 = n27834 ^ n27779 ;
  assign n28311 = n28310 ^ n28309 ;
  assign n28313 = n28312 ^ n28311 ;
  assign n28314 = n28305 & n28313 ;
  assign n28315 = n28314 ^ n28312 ;
  assign n28126 = n27840 ^ n27775 ;
  assign n28318 = n28309 ^ n28126 ;
  assign n28316 = n27838 ^ n27776 ;
  assign n28317 = n28316 ^ n28126 ;
  assign n28319 = n28318 ^ n28317 ;
  assign n28320 = ~n28315 & ~n28319 ;
  assign n28321 = n28320 ^ n28318 ;
  assign n28122 = n26600 ^ n25952 ;
  assign n28123 = n27989 ^ n26600 ;
  assign n28124 = n28122 & ~n28123 ;
  assign n28125 = n28124 ^ n25952 ;
  assign n28348 = n28321 ^ n28125 ;
  assign n28349 = n28348 ^ n25467 ;
  assign n28350 = n28316 ^ n28315 ;
  assign n28351 = n28350 ^ n26068 ;
  assign n28451 = n28310 ^ n28305 ;
  assign n28442 = n28294 ^ n28135 ;
  assign n28353 = n28291 ^ n28147 ;
  assign n28354 = n28353 ^ n25779 ;
  assign n28355 = n28289 ^ n28281 ;
  assign n28356 = n28355 ^ n25767 ;
  assign n28358 = n28263 ^ n28259 ;
  assign n28359 = n28358 ^ n25104 ;
  assign n28361 = n28253 ^ n28178 ;
  assign n28362 = n28361 ^ n25119 ;
  assign n28363 = n28250 ^ n28183 ;
  assign n28364 = n28363 ^ n25127 ;
  assign n28400 = n28247 ^ n28188 ;
  assign n28365 = n28244 ^ n28194 ;
  assign n28366 = n28365 ^ n25520 ;
  assign n28367 = n28242 ^ n28198 ;
  assign n28368 = n28367 ^ n25134 ;
  assign n28369 = n28235 ^ n28212 ;
  assign n28370 = n28369 ^ n25138 ;
  assign n28376 = n28222 ^ n28216 ;
  assign n28064 = n28063 ^ n28060 ;
  assign n28372 = n28064 ^ n25151 ;
  assign n28005 = n28004 ^ n27983 ;
  assign n28006 = n28005 ^ n25153 ;
  assign n27962 = n27961 ^ n27957 ;
  assign n27963 = n27962 ^ n25157 ;
  assign n27965 = n27902 ^ n27898 ;
  assign n27966 = n25165 & ~n27965 ;
  assign n27964 = n27952 ^ n27908 ;
  assign n27967 = n27966 ^ n27964 ;
  assign n27968 = n27962 ^ n25163 ;
  assign n27969 = n27968 ^ n27964 ;
  assign n27970 = n27969 ^ n27962 ;
  assign n27971 = ~n27967 & n27970 ;
  assign n27972 = n27971 ^ n27968 ;
  assign n27973 = ~n27963 & n27972 ;
  assign n27974 = n27973 ^ n25157 ;
  assign n28032 = n28005 ^ n27974 ;
  assign n28033 = ~n28006 & ~n28032 ;
  assign n28034 = n28033 ^ n25153 ;
  assign n28373 = n28064 ^ n28034 ;
  assign n28374 = ~n28372 & ~n28373 ;
  assign n28375 = n28374 ^ n25151 ;
  assign n28377 = n28376 ^ n28375 ;
  assign n28378 = n28376 ^ n25147 ;
  assign n28379 = n28377 & ~n28378 ;
  assign n28380 = n28379 ^ n25147 ;
  assign n28371 = n28233 ^ n28224 ;
  assign n28381 = n28380 ^ n28371 ;
  assign n28382 = n28369 ^ n25140 ;
  assign n28383 = n28382 ^ n28369 ;
  assign n28384 = n28383 ^ n28371 ;
  assign n28385 = ~n28381 & ~n28384 ;
  assign n28386 = n28385 ^ n28382 ;
  assign n28387 = n28370 & n28386 ;
  assign n28388 = n28387 ^ n25138 ;
  assign n28389 = n28388 ^ n25132 ;
  assign n28390 = n28238 ^ n28206 ;
  assign n28391 = n28390 ^ n28388 ;
  assign n28392 = n28389 & ~n28391 ;
  assign n28393 = n28392 ^ n25132 ;
  assign n28394 = n28393 ^ n28367 ;
  assign n28395 = ~n28368 & ~n28394 ;
  assign n28396 = n28395 ^ n25134 ;
  assign n28397 = n28396 ^ n28365 ;
  assign n28398 = ~n28366 & ~n28397 ;
  assign n28399 = n28398 ^ n25520 ;
  assign n28401 = n28400 ^ n28399 ;
  assign n28402 = n28400 ^ n25535 ;
  assign n28403 = n28401 & ~n28402 ;
  assign n28404 = n28403 ^ n25535 ;
  assign n28405 = n28404 ^ n28363 ;
  assign n28406 = ~n28364 & ~n28405 ;
  assign n28407 = n28406 ^ n25127 ;
  assign n28408 = n28407 ^ n28361 ;
  assign n28409 = ~n28362 & ~n28408 ;
  assign n28410 = n28409 ^ n25119 ;
  assign n28360 = n28256 ^ n28169 ;
  assign n28411 = n28410 ^ n28360 ;
  assign n28412 = n28358 ^ n25114 ;
  assign n28413 = n28412 ^ n28358 ;
  assign n28414 = n28413 ^ n28360 ;
  assign n28415 = ~n28411 & ~n28414 ;
  assign n28416 = n28415 ^ n28412 ;
  assign n28417 = ~n28359 & n28416 ;
  assign n28418 = n28417 ^ n25104 ;
  assign n28357 = n28268 ^ n28162 ;
  assign n28419 = n28418 ^ n28357 ;
  assign n28420 = n28270 ^ n28154 ;
  assign n28421 = n28420 ^ n25554 ;
  assign n28422 = n28421 ^ n28357 ;
  assign n28423 = n28422 ^ n28420 ;
  assign n28424 = n28419 & ~n28423 ;
  assign n28425 = n28424 ^ n28421 ;
  assign n28426 = n28278 ^ n28277 ;
  assign n28428 = n28426 ^ n25559 ;
  assign n28427 = n28426 ^ n28420 ;
  assign n28429 = n28428 ^ n28427 ;
  assign n28430 = ~n28425 & ~n28429 ;
  assign n28431 = n28430 ^ n28428 ;
  assign n28433 = n28355 ^ n25694 ;
  assign n28432 = n28426 ^ n28355 ;
  assign n28434 = n28433 ^ n28432 ;
  assign n28435 = n28431 & ~n28434 ;
  assign n28436 = n28435 ^ n28433 ;
  assign n28437 = ~n28356 & ~n28436 ;
  assign n28438 = n28437 ^ n25767 ;
  assign n28439 = n28438 ^ n28353 ;
  assign n28440 = ~n28354 & ~n28439 ;
  assign n28441 = n28440 ^ n25779 ;
  assign n28443 = n28442 ^ n28441 ;
  assign n28444 = n28442 ^ n25961 ;
  assign n28445 = n28443 & ~n28444 ;
  assign n28446 = n28445 ^ n25961 ;
  assign n28352 = n28296 ^ n28134 ;
  assign n28447 = n28446 ^ n28352 ;
  assign n28448 = n28446 ^ n25989 ;
  assign n28449 = ~n28447 & ~n28448 ;
  assign n28450 = n28449 ^ n25989 ;
  assign n28452 = n28451 ^ n28450 ;
  assign n28453 = n28350 ^ n26035 ;
  assign n28454 = n28453 ^ n28350 ;
  assign n28455 = n28454 ^ n28450 ;
  assign n28456 = ~n28452 & n28455 ;
  assign n28457 = n28456 ^ n28453 ;
  assign n28458 = ~n28351 & n28457 ;
  assign n28459 = n28458 ^ n26068 ;
  assign n28460 = n28459 ^ n28348 ;
  assign n28461 = ~n28349 & n28460 ;
  assign n28462 = n28461 ^ n25467 ;
  assign n28127 = n28126 ^ n28125 ;
  assign n28322 = n28127 & ~n28321 ;
  assign n28323 = n28322 ^ n28126 ;
  assign n28111 = n28043 ^ n26787 ;
  assign n28112 = n27844 ^ n1090 ;
  assign n28113 = n28112 ^ n25978 ;
  assign n28114 = n28113 ^ n28043 ;
  assign n28115 = n28114 ^ n28112 ;
  assign n28116 = n28111 & n28115 ;
  assign n28117 = n28116 ^ n28113 ;
  assign n28346 = n28323 ^ n28117 ;
  assign n28347 = n28346 ^ n25470 ;
  assign n28543 = n28462 ^ n28347 ;
  assign n28494 = n28352 ^ n25989 ;
  assign n28495 = n28494 ^ n28446 ;
  assign n28496 = n28444 ^ n28441 ;
  assign n28497 = n28431 ^ n25694 ;
  assign n28498 = n28416 ^ n25104 ;
  assign n28499 = n28360 ^ n25114 ;
  assign n28500 = n28499 ^ n28410 ;
  assign n28501 = n28404 ^ n28364 ;
  assign n28502 = n28402 ^ n28399 ;
  assign n28503 = n28390 ^ n28389 ;
  assign n28504 = n28386 ^ n25138 ;
  assign n28505 = n28378 ^ n28375 ;
  assign n28035 = n28034 ^ n25151 ;
  assign n28065 = n28064 ^ n28035 ;
  assign n28007 = n28006 ^ n27974 ;
  assign n28008 = n27972 ^ n25157 ;
  assign n28066 = n28007 & n28008 ;
  assign n28506 = ~n28065 & n28066 ;
  assign n28507 = ~n28505 & ~n28506 ;
  assign n28508 = n28371 ^ n25140 ;
  assign n28509 = n28508 ^ n28380 ;
  assign n28510 = ~n28507 & n28509 ;
  assign n28511 = n28504 & n28510 ;
  assign n28512 = n28503 & ~n28511 ;
  assign n28513 = n28393 ^ n28368 ;
  assign n28514 = n28512 & ~n28513 ;
  assign n28515 = n28396 ^ n28366 ;
  assign n28516 = ~n28514 & ~n28515 ;
  assign n28517 = n28502 & n28516 ;
  assign n28518 = n28501 & n28517 ;
  assign n28519 = n28407 ^ n28362 ;
  assign n28520 = n28518 & ~n28519 ;
  assign n28521 = ~n28500 & ~n28520 ;
  assign n28522 = ~n28498 & ~n28521 ;
  assign n28523 = n28418 ^ n25554 ;
  assign n28524 = n28523 ^ n28357 ;
  assign n28525 = n28522 & ~n28524 ;
  assign n28526 = n28425 ^ n25559 ;
  assign n28527 = n28525 & ~n28526 ;
  assign n28528 = ~n28497 & ~n28527 ;
  assign n28529 = n28436 ^ n25767 ;
  assign n28530 = ~n28528 & n28529 ;
  assign n28531 = n28438 ^ n25779 ;
  assign n28532 = n28531 ^ n28353 ;
  assign n28533 = n28530 & ~n28532 ;
  assign n28534 = ~n28496 & ~n28533 ;
  assign n28535 = ~n28495 & n28534 ;
  assign n28536 = n28450 ^ n26035 ;
  assign n28537 = n28536 ^ n28451 ;
  assign n28538 = n28535 & ~n28537 ;
  assign n28539 = n28457 ^ n26068 ;
  assign n28540 = ~n28538 & ~n28539 ;
  assign n28541 = n28459 ^ n28349 ;
  assign n28542 = n28540 & ~n28541 ;
  assign n28591 = n28543 ^ n28542 ;
  assign n2646 = n2645 ^ n2510 ;
  assign n2647 = n2646 ^ n2558 ;
  assign n2648 = n2647 ^ n2624 ;
  assign n28592 = n28591 ^ n2648 ;
  assign n28596 = n26450 ^ n3206 ;
  assign n28597 = n28596 ^ n23472 ;
  assign n28598 = n28597 ^ n2553 ;
  assign n28595 = n28541 ^ n28540 ;
  assign n28599 = n28598 ^ n28595 ;
  assign n28600 = n28539 ^ n28538 ;
  assign n28601 = n28600 ^ n2804 ;
  assign n28602 = n28537 ^ n28535 ;
  assign n28603 = n28602 ^ n1369 ;
  assign n28604 = n28534 ^ n28495 ;
  assign n28605 = n28604 ^ n1230 ;
  assign n28606 = n28533 ^ n28496 ;
  assign n1207 = n1167 ^ n1103 ;
  assign n1208 = n1207 ^ n1204 ;
  assign n1212 = n1211 ^ n1208 ;
  assign n28607 = n28606 ^ n1212 ;
  assign n1189 = n1114 ^ n1036 ;
  assign n1196 = n1195 ^ n1189 ;
  assign n1197 = n1196 ^ n980 ;
  assign n28710 = n1212 ^ n1197 ;
  assign n28608 = n28532 ^ n28530 ;
  assign n28609 = n28608 ^ n1197 ;
  assign n28610 = n28529 ^ n28528 ;
  assign n1671 = n1652 ^ n1021 ;
  assign n1672 = n1671 ^ n842 ;
  assign n1673 = n1672 ^ n1193 ;
  assign n28611 = n28610 ^ n1673 ;
  assign n28612 = n28527 ^ n28497 ;
  assign n1661 = n1646 ^ n1015 ;
  assign n1665 = n1664 ^ n1661 ;
  assign n1666 = n1665 ^ n836 ;
  assign n28613 = n28612 ^ n1666 ;
  assign n729 = n728 ^ n695 ;
  assign n739 = n738 ^ n729 ;
  assign n743 = n742 ^ n739 ;
  assign n28701 = n1666 ^ n743 ;
  assign n28614 = n28524 ^ n28522 ;
  assign n2981 = n2974 ^ n1623 ;
  assign n2982 = n2981 ^ n679 ;
  assign n2983 = n2982 ^ n733 ;
  assign n28615 = n28614 ^ n2983 ;
  assign n28618 = n28521 ^ n28498 ;
  assign n28619 = n28618 ^ n672 ;
  assign n28623 = n28520 ^ n28500 ;
  assign n28624 = n28623 ^ n28622 ;
  assign n28688 = n28623 ^ n1517 ;
  assign n28625 = n28519 ^ n28518 ;
  assign n28626 = n28625 ^ n1517 ;
  assign n28630 = n28517 ^ n28501 ;
  assign n28631 = n28630 ^ n28629 ;
  assign n28634 = n26481 ^ n19526 ;
  assign n28635 = n28634 ^ n2915 ;
  assign n28636 = n28635 ^ n18027 ;
  assign n28633 = n28515 ^ n28514 ;
  assign n28637 = n28636 ^ n28633 ;
  assign n28642 = n28510 ^ n28504 ;
  assign n28639 = n26497 ^ n19489 ;
  assign n28640 = n28639 ^ n2164 ;
  assign n28641 = n28640 ^ n2286 ;
  assign n28643 = n28642 ^ n28641 ;
  assign n28644 = n28509 ^ n28507 ;
  assign n2149 = n2142 ^ n2091 ;
  assign n2156 = n2155 ^ n2149 ;
  assign n2160 = n2159 ^ n2156 ;
  assign n28645 = n28644 ^ n2160 ;
  assign n28067 = n28066 ^ n28065 ;
  assign n2039 = n2026 ^ n2002 ;
  assign n2052 = n2051 ^ n2039 ;
  assign n2056 = n2055 ^ n2052 ;
  assign n28068 = n28067 ^ n2056 ;
  assign n28010 = n26112 ^ n1961 ;
  assign n28011 = n28010 ^ n23096 ;
  assign n28012 = n28011 ^ n2048 ;
  assign n28009 = n28008 ^ n28007 ;
  assign n28013 = n28012 ^ n28009 ;
  assign n3083 = n3052 ^ n1952 ;
  assign n3084 = n3083 ^ n3080 ;
  assign n3088 = n3087 ^ n3084 ;
  assign n28014 = n28008 ^ n3088 ;
  assign n28015 = n3014 ^ n2767 ;
  assign n28016 = n28015 ^ n23528 ;
  assign n28017 = n28016 ^ n1787 ;
  assign n28018 = n27965 ^ n25165 ;
  assign n28019 = n28017 & ~n28018 ;
  assign n3071 = n3058 ^ n3040 ;
  assign n3075 = n3074 ^ n3071 ;
  assign n3076 = n3075 ^ n3070 ;
  assign n28020 = n28019 ^ n3076 ;
  assign n28021 = n27966 ^ n25163 ;
  assign n28022 = n28021 ^ n27964 ;
  assign n28023 = n28022 ^ n28019 ;
  assign n28024 = n28020 & ~n28023 ;
  assign n28025 = n28024 ^ n3076 ;
  assign n28026 = n28025 ^ n28008 ;
  assign n28027 = n28014 & ~n28026 ;
  assign n28028 = n28027 ^ n3088 ;
  assign n28029 = n28028 ^ n28009 ;
  assign n28030 = ~n28013 & n28029 ;
  assign n28031 = n28030 ^ n28012 ;
  assign n28647 = n28031 ^ n2056 ;
  assign n28648 = n28068 & n28647 ;
  assign n28649 = n28648 ^ n2056 ;
  assign n28653 = n28649 ^ n2160 ;
  assign n28646 = n28506 ^ n28505 ;
  assign n28650 = n28649 ^ n28646 ;
  assign n2066 = n2035 ^ n2014 ;
  assign n2067 = n2066 ^ n2063 ;
  assign n2071 = n2070 ^ n2067 ;
  assign n28651 = n28646 ^ n2071 ;
  assign n28652 = n28650 & ~n28651 ;
  assign n28654 = n28653 ^ n28652 ;
  assign n28655 = n28645 & ~n28654 ;
  assign n28656 = n28655 ^ n28644 ;
  assign n28657 = n28656 ^ n28641 ;
  assign n28658 = ~n28643 & n28657 ;
  assign n28659 = n28658 ^ n28641 ;
  assign n28666 = n28665 ^ n28659 ;
  assign n28638 = n28511 ^ n28503 ;
  assign n28660 = n28659 ^ n28638 ;
  assign n2283 = n2282 ^ n2216 ;
  assign n2293 = n2292 ^ n2283 ;
  assign n2297 = n2296 ^ n2293 ;
  assign n28661 = n28638 ^ n2297 ;
  assign n28662 = ~n28660 & n28661 ;
  assign n28667 = n28666 ^ n28662 ;
  assign n28670 = n28665 ^ n28636 ;
  assign n28668 = n28513 ^ n28512 ;
  assign n28669 = n28668 ^ n28636 ;
  assign n28671 = n28670 ^ n28669 ;
  assign n28672 = n28667 & ~n28671 ;
  assign n28673 = n28672 ^ n28670 ;
  assign n28674 = ~n28637 & n28673 ;
  assign n28675 = n28674 ^ n28636 ;
  assign n28682 = n28675 ^ n28629 ;
  assign n28632 = n28516 ^ n28502 ;
  assign n28676 = n28675 ^ n28632 ;
  assign n28677 = n26472 ^ n1482 ;
  assign n28678 = n28677 ^ n23133 ;
  assign n28679 = n28678 ^ n2924 ;
  assign n28680 = n28679 ^ n28675 ;
  assign n28681 = ~n28676 & n28680 ;
  assign n28683 = n28682 ^ n28681 ;
  assign n28684 = ~n28631 & ~n28683 ;
  assign n28685 = n28684 ^ n28630 ;
  assign n28686 = n28685 ^ n1517 ;
  assign n28687 = n28626 & ~n28686 ;
  assign n28689 = n28688 ^ n28687 ;
  assign n28690 = n28624 & n28689 ;
  assign n28691 = n28690 ^ n28623 ;
  assign n28692 = n28691 ^ n672 ;
  assign n28693 = ~n28619 & ~n28692 ;
  assign n28694 = n28693 ^ n28618 ;
  assign n28616 = n2983 ^ n743 ;
  assign n28617 = n28616 ^ n743 ;
  assign n28695 = n28694 ^ n28617 ;
  assign n28696 = n28615 & ~n28695 ;
  assign n28697 = n28696 ^ n28616 ;
  assign n28698 = n28526 ^ n28525 ;
  assign n28699 = n28698 ^ n743 ;
  assign n28700 = n28697 & n28699 ;
  assign n28702 = n28701 ^ n28700 ;
  assign n28703 = n28613 & ~n28702 ;
  assign n28704 = n28703 ^ n28612 ;
  assign n28705 = n28704 ^ n1673 ;
  assign n28706 = n28611 & ~n28705 ;
  assign n28707 = n28706 ^ n28610 ;
  assign n28708 = n28707 ^ n1197 ;
  assign n28709 = n28609 & n28708 ;
  assign n28711 = n28710 ^ n28709 ;
  assign n28712 = n28607 & ~n28711 ;
  assign n28713 = n28712 ^ n28606 ;
  assign n28714 = n28713 ^ n1230 ;
  assign n28715 = ~n28605 & ~n28714 ;
  assign n28716 = n28715 ^ n28604 ;
  assign n28717 = n28716 ^ n1369 ;
  assign n28718 = ~n28603 & n28717 ;
  assign n28719 = n28718 ^ n28602 ;
  assign n28720 = n28719 ^ n28600 ;
  assign n28721 = ~n28601 & ~n28720 ;
  assign n28722 = n28721 ^ n2804 ;
  assign n28723 = n28722 ^ n28595 ;
  assign n28724 = n28599 & ~n28723 ;
  assign n28725 = n28724 ^ n28598 ;
  assign n28329 = n27848 ^ n1253 ;
  assign n28118 = n26791 ^ n26003 ;
  assign n28119 = n27350 ^ n26791 ;
  assign n28120 = n28118 & n28119 ;
  assign n28121 = n28120 ^ n26003 ;
  assign n28325 = n28121 ^ n28112 ;
  assign n28324 = n28323 ^ n28121 ;
  assign n28326 = n28325 ^ n28324 ;
  assign n28327 = ~n28117 & ~n28326 ;
  assign n28328 = n28327 ^ n28325 ;
  assign n28345 = n28329 ^ n28328 ;
  assign n28545 = n28345 ^ n25460 ;
  assign n28463 = n28462 ^ n28346 ;
  assign n28464 = n28347 & n28463 ;
  assign n28465 = n28464 ^ n25470 ;
  assign n28546 = n28545 ^ n28465 ;
  assign n28544 = n28542 & n28543 ;
  assign n28586 = n28546 ^ n28544 ;
  assign n28593 = n28586 ^ n2648 ;
  assign n28594 = n28593 ^ n28586 ;
  assign n28726 = n28725 ^ n28594 ;
  assign n28727 = ~n28592 & n28726 ;
  assign n28728 = n28727 ^ n28593 ;
  assign n28754 = n28728 ^ n28589 ;
  assign n28750 = n27412 ^ n26687 ;
  assign n28751 = n28217 ^ n27412 ;
  assign n28752 = ~n28750 & ~n28751 ;
  assign n28753 = n28752 ^ n26687 ;
  assign n28803 = n28754 ^ n28753 ;
  assign n28905 = n28803 ^ n26192 ;
  assign n28902 = n20332 ^ n3183 ;
  assign n28903 = n28902 ^ n2753 ;
  assign n28904 = n28903 ^ n1858 ;
  assign n29021 = n28905 ^ n28904 ;
  assign n30279 = n29021 ^ n28211 ;
  assign n28080 = n28025 ^ n28014 ;
  assign n30280 = n28211 ^ n28080 ;
  assign n30281 = ~n30279 & n30280 ;
  assign n30282 = n30281 ^ n28080 ;
  assign n29092 = n28656 ^ n28643 ;
  assign n28946 = n27543 ^ n26868 ;
  assign n28947 = n28157 ^ n27543 ;
  assign n28948 = n28946 & n28947 ;
  assign n28949 = n28948 ^ n26868 ;
  assign n28945 = n28654 ^ n28644 ;
  assign n28950 = n28949 ^ n28945 ;
  assign n28845 = n27547 ^ n26860 ;
  assign n28846 = n28170 ^ n27547 ;
  assign n28847 = n28845 & ~n28846 ;
  assign n28848 = n28847 ^ n26860 ;
  assign n28844 = n28651 ^ n28649 ;
  assign n28849 = n28848 ^ n28844 ;
  assign n27518 = n27517 ^ n27516 ;
  assign n28069 = n28068 ^ n28031 ;
  assign n28070 = n28069 ^ n26841 ;
  assign n28071 = n28070 ^ n27516 ;
  assign n28072 = n28071 ^ n28069 ;
  assign n28073 = n27518 & n28072 ;
  assign n28074 = n28073 ^ n28070 ;
  assign n28783 = n28028 ^ n28013 ;
  assign n28076 = n28075 ^ n27558 ;
  assign n28077 = n27558 ^ n26664 ;
  assign n28078 = ~n28076 & ~n28077 ;
  assign n28079 = n28078 ^ n26664 ;
  assign n28081 = n28080 ^ n28079 ;
  assign n28088 = n28022 ^ n28020 ;
  assign n28083 = n28082 ^ n27562 ;
  assign n28084 = n27562 ^ n26662 ;
  assign n28085 = n28083 & ~n28084 ;
  assign n28086 = n28085 ^ n26662 ;
  assign n28089 = n28088 ^ n28086 ;
  assign n28091 = n28090 ^ n27567 ;
  assign n28092 = n28018 ^ n28017 ;
  assign n28093 = n28092 ^ n26669 ;
  assign n28094 = n28093 ^ n28090 ;
  assign n28095 = n28094 ^ n28092 ;
  assign n28096 = ~n28091 & ~n28095 ;
  assign n28097 = n28096 ^ n28093 ;
  assign n28341 = n27864 ^ n27863 ;
  assign n28337 = n26777 ^ n26081 ;
  assign n28338 = n27344 ^ n26777 ;
  assign n28339 = ~n28337 & ~n28338 ;
  assign n28340 = n28339 ^ n26081 ;
  assign n28342 = n28341 ^ n28340 ;
  assign n28106 = n26799 ^ n26046 ;
  assign n28107 = n27352 ^ n26799 ;
  assign n28108 = ~n28106 & ~n28107 ;
  assign n28109 = n28108 ^ n26046 ;
  assign n28105 = n27856 ^ n27853 ;
  assign n28110 = n28109 ^ n28105 ;
  assign n28331 = n28121 ^ n28109 ;
  assign n28330 = n28329 ^ n28109 ;
  assign n28332 = n28331 ^ n28330 ;
  assign n28333 = n28328 & ~n28332 ;
  assign n28334 = n28333 ^ n28331 ;
  assign n28335 = ~n28110 & n28334 ;
  assign n28336 = n28335 ^ n28109 ;
  assign n28486 = n28340 ^ n28336 ;
  assign n28487 = ~n28342 & ~n28486 ;
  assign n28488 = n28487 ^ n28341 ;
  assign n28479 = n27342 ^ n26693 ;
  assign n28480 = n27873 ^ n27872 ;
  assign n28481 = n28480 ^ n26102 ;
  assign n28482 = n28481 ^ n27342 ;
  assign n28483 = n28482 ^ n28480 ;
  assign n28484 = ~n28479 & ~n28483 ;
  assign n28485 = n28484 ^ n28481 ;
  assign n28489 = n28488 ^ n28485 ;
  assign n28573 = n28489 ^ n25172 ;
  assign n28343 = n28342 ^ n28336 ;
  assign n28344 = n28343 ^ n25450 ;
  assign n28470 = n28334 ^ n28105 ;
  assign n28466 = n28465 ^ n28345 ;
  assign n28467 = n28465 ^ n25460 ;
  assign n28468 = n28466 & ~n28467 ;
  assign n28469 = n28468 ^ n25460 ;
  assign n28471 = n28470 ^ n28469 ;
  assign n28472 = n28343 ^ n25456 ;
  assign n28473 = n28472 ^ n28343 ;
  assign n28474 = n28473 ^ n28469 ;
  assign n28475 = ~n28471 & n28474 ;
  assign n28476 = n28475 ^ n28472 ;
  assign n28477 = ~n28344 & ~n28476 ;
  assign n28478 = n28477 ^ n25450 ;
  assign n28574 = n28573 ^ n28478 ;
  assign n28492 = n28469 ^ n25456 ;
  assign n28493 = n28492 ^ n28470 ;
  assign n28547 = n28544 & ~n28546 ;
  assign n28548 = ~n28493 & ~n28547 ;
  assign n28549 = n28476 ^ n25450 ;
  assign n28550 = n28548 & n28549 ;
  assign n28575 = n28574 ^ n28550 ;
  assign n28569 = n26755 ^ n2713 ;
  assign n28570 = n28569 ^ n3157 ;
  assign n28571 = n28570 ^ n1820 ;
  assign n28576 = n28575 ^ n28571 ;
  assign n28577 = n28549 ^ n28548 ;
  assign n28578 = n28577 ^ n3153 ;
  assign n28580 = n26581 ^ n3127 ;
  assign n28581 = n28580 ^ n2516 ;
  assign n28582 = n28581 ^ n3148 ;
  assign n28579 = n28547 ^ n28493 ;
  assign n28583 = n28582 ^ n28579 ;
  assign n28590 = n28589 ^ n28586 ;
  assign n28729 = n28590 & ~n28728 ;
  assign n28730 = n28729 ^ n28589 ;
  assign n28584 = n28582 ^ n3153 ;
  assign n28585 = n28584 ^ n3153 ;
  assign n28731 = n28730 ^ n28585 ;
  assign n28732 = n28583 & n28731 ;
  assign n28733 = n28732 ^ n28584 ;
  assign n28734 = n28578 & n28733 ;
  assign n28735 = n28734 ^ n3153 ;
  assign n28736 = n28735 ^ n28571 ;
  assign n28737 = n28576 & n28736 ;
  assign n28563 = n26691 ^ n26197 ;
  assign n28564 = n27338 ^ n26691 ;
  assign n28565 = n28563 & ~n28564 ;
  assign n28559 = n28488 ^ n26197 ;
  assign n28558 = n27878 ^ n27770 ;
  assign n28560 = n28559 ^ n28558 ;
  assign n28561 = n28560 ^ n24702 ;
  assign n28556 = n28488 ^ n28480 ;
  assign n28557 = ~n28485 & n28556 ;
  assign n28562 = n28561 ^ n28557 ;
  assign n28566 = n28565 ^ n28562 ;
  assign n28490 = n28489 ^ n28478 ;
  assign n28551 = n28550 ^ n28478 ;
  assign n28554 = n28490 & ~n28551 ;
  assign n28552 = n28551 ^ n28489 ;
  assign n28553 = n25172 & ~n28552 ;
  assign n28555 = n28554 ^ n28553 ;
  assign n28567 = n28566 ^ n28555 ;
  assign n3177 = n2772 ^ n2730 ;
  assign n3178 = n3177 ^ n1844 ;
  assign n3179 = n3178 ^ n3176 ;
  assign n28568 = n28567 ^ n3179 ;
  assign n28572 = n28571 ^ n28568 ;
  assign n28738 = n28737 ^ n28572 ;
  assign n28101 = n28100 ^ n27577 ;
  assign n28102 = n27577 ^ n26671 ;
  assign n28103 = n28101 & ~n28102 ;
  assign n28104 = n28103 ^ n26671 ;
  assign n28739 = n28738 ^ n28104 ;
  assign n28744 = n28735 ^ n28576 ;
  assign n28740 = n28201 ^ n27576 ;
  assign n28741 = n27576 ^ n26131 ;
  assign n28742 = ~n28740 & ~n28741 ;
  assign n28743 = n28742 ^ n26131 ;
  assign n28745 = n28744 ^ n28743 ;
  assign n28761 = n27502 ^ n26608 ;
  assign n28762 = n28211 ^ n27502 ;
  assign n28763 = n28761 & n28762 ;
  assign n28764 = n28763 ^ n26608 ;
  assign n28755 = ~n28753 & n28754 ;
  assign n28746 = n27485 ^ n26683 ;
  assign n28747 = n28226 ^ n27485 ;
  assign n28748 = n28746 & ~n28747 ;
  assign n28749 = n28748 ^ n26683 ;
  assign n28756 = n28755 ^ n28749 ;
  assign n28757 = n28730 ^ n28583 ;
  assign n28758 = n28757 ^ n28749 ;
  assign n28759 = ~n28756 & n28758 ;
  assign n28760 = n28759 ^ n28755 ;
  assign n28765 = n28764 ^ n28760 ;
  assign n28766 = n28733 ^ n28577 ;
  assign n28767 = n28766 ^ n28764 ;
  assign n28768 = n28765 & ~n28767 ;
  assign n28769 = n28768 ^ n28766 ;
  assign n28770 = n28769 ^ n28743 ;
  assign n28771 = n28745 & ~n28770 ;
  assign n28772 = n28771 ^ n28744 ;
  assign n28773 = n28772 ^ n28104 ;
  assign n28774 = n28739 & n28773 ;
  assign n28775 = n28774 ^ n28738 ;
  assign n28776 = n28775 ^ n28092 ;
  assign n28777 = n28097 & n28776 ;
  assign n28098 = n28092 ^ n28086 ;
  assign n28778 = n28777 ^ n28098 ;
  assign n28779 = ~n28089 & n28778 ;
  assign n28087 = n28086 ^ n28079 ;
  assign n28780 = n28779 ^ n28087 ;
  assign n28781 = n28081 & n28780 ;
  assign n28782 = n28781 ^ n28080 ;
  assign n28784 = n28783 ^ n28782 ;
  assign n28785 = n28177 ^ n27554 ;
  assign n28786 = n28783 ^ n26833 ;
  assign n28787 = n28786 ^ n28177 ;
  assign n28788 = n28787 ^ n28783 ;
  assign n28789 = n28785 & ~n28788 ;
  assign n28790 = n28789 ^ n28786 ;
  assign n28791 = ~n28784 & ~n28790 ;
  assign n28792 = n28791 ^ n28783 ;
  assign n28841 = n28792 ^ n28069 ;
  assign n28842 = n28074 & ~n28841 ;
  assign n28843 = n28842 ^ n28792 ;
  assign n28942 = n28844 ^ n28843 ;
  assign n28943 = ~n28849 & n28942 ;
  assign n28944 = n28943 ^ n28848 ;
  assign n29089 = n28945 ^ n28944 ;
  assign n29090 = ~n28950 & n29089 ;
  assign n29091 = n29090 ^ n28949 ;
  assign n29093 = n29092 ^ n29091 ;
  assign n29094 = n28155 ^ n27536 ;
  assign n29095 = n29092 ^ n26874 ;
  assign n29096 = n29095 ^ n28155 ;
  assign n29097 = n29096 ^ n29092 ;
  assign n29098 = n29094 & ~n29097 ;
  assign n29099 = n29098 ^ n29095 ;
  assign n29100 = n29093 & n29099 ;
  assign n29101 = n29100 ^ n29092 ;
  assign n29084 = n27534 ^ n26658 ;
  assign n29085 = n28278 ^ n27534 ;
  assign n29086 = ~n29084 & ~n29085 ;
  assign n29087 = n29086 ^ n26658 ;
  assign n29004 = n28661 ^ n28659 ;
  assign n29088 = n29087 ^ n29004 ;
  assign n29223 = n29101 ^ n29088 ;
  assign n29309 = n29223 ^ n26139 ;
  assign n29224 = n29099 ^ n29091 ;
  assign n29225 = n29224 ^ n26145 ;
  assign n28850 = n28849 ^ n28843 ;
  assign n28851 = n28850 ^ n26151 ;
  assign n28794 = n28790 ^ n28782 ;
  assign n28795 = n28794 ^ n26161 ;
  assign n28797 = n28778 ^ n28088 ;
  assign n28798 = n28797 ^ n26169 ;
  assign n28799 = n28775 ^ n28097 ;
  assign n28800 = n28799 ^ n26133 ;
  assign n28818 = n28772 ^ n28739 ;
  assign n28801 = n28769 ^ n28745 ;
  assign n28802 = n28801 ^ n26180 ;
  assign n28810 = n28767 ^ n28760 ;
  assign n28804 = ~n26192 & ~n28803 ;
  assign n28805 = n28804 ^ n26188 ;
  assign n28806 = n28757 ^ n28756 ;
  assign n28807 = n28806 ^ n28804 ;
  assign n28808 = ~n28805 & n28807 ;
  assign n28809 = n28808 ^ n26188 ;
  assign n28811 = n28810 ^ n28809 ;
  assign n28812 = n28810 ^ n26184 ;
  assign n28813 = ~n28811 & ~n28812 ;
  assign n28814 = n28813 ^ n26184 ;
  assign n28815 = n28814 ^ n28801 ;
  assign n28816 = ~n28802 & ~n28815 ;
  assign n28817 = n28816 ^ n26180 ;
  assign n28819 = n28818 ^ n28817 ;
  assign n28820 = n28799 ^ n26176 ;
  assign n28821 = n28820 ^ n28799 ;
  assign n28822 = n28821 ^ n28817 ;
  assign n28823 = n28819 & n28822 ;
  assign n28824 = n28823 ^ n28820 ;
  assign n28825 = ~n28800 & ~n28824 ;
  assign n28826 = n28825 ^ n26133 ;
  assign n28827 = n28826 ^ n28797 ;
  assign n28828 = ~n28798 & ~n28827 ;
  assign n28829 = n28828 ^ n26169 ;
  assign n28796 = n28780 ^ n28080 ;
  assign n28830 = n28829 ^ n28796 ;
  assign n28831 = n28829 ^ n26165 ;
  assign n28832 = ~n28830 & n28831 ;
  assign n28833 = n28832 ^ n26165 ;
  assign n28834 = n28833 ^ n28794 ;
  assign n28835 = n28795 & ~n28834 ;
  assign n28836 = n28835 ^ n26161 ;
  assign n28793 = n28792 ^ n28074 ;
  assign n28837 = n28836 ^ n28793 ;
  assign n28838 = n28836 ^ n26155 ;
  assign n28839 = n28837 & ~n28838 ;
  assign n28840 = n28839 ^ n26155 ;
  assign n28953 = n28850 ^ n28840 ;
  assign n28954 = ~n28851 & ~n28953 ;
  assign n28955 = n28954 ^ n26151 ;
  assign n28951 = n28950 ^ n28944 ;
  assign n29226 = n28955 ^ n28951 ;
  assign n29227 = n28955 ^ n26147 ;
  assign n29228 = n29226 & ~n29227 ;
  assign n29229 = n29228 ^ n26147 ;
  assign n29230 = n29229 ^ n29224 ;
  assign n29231 = ~n29225 & n29230 ;
  assign n29232 = n29231 ^ n26145 ;
  assign n29310 = n29309 ^ n29232 ;
  assign n28952 = n28951 ^ n26147 ;
  assign n28956 = n28955 ^ n28952 ;
  assign n28852 = n28851 ^ n28840 ;
  assign n28853 = n28809 ^ n26184 ;
  assign n28854 = n28853 ^ n28810 ;
  assign n28855 = n28814 ^ n28802 ;
  assign n28856 = ~n28854 & n28855 ;
  assign n28857 = n28818 ^ n26176 ;
  assign n28858 = n28857 ^ n28817 ;
  assign n28859 = n28856 & ~n28858 ;
  assign n28860 = n28824 ^ n26133 ;
  assign n28861 = ~n28859 & n28860 ;
  assign n28862 = n28826 ^ n28798 ;
  assign n28863 = ~n28861 & n28862 ;
  assign n28864 = n28796 ^ n26165 ;
  assign n28865 = n28864 ^ n28829 ;
  assign n28866 = n28863 & n28865 ;
  assign n28867 = n28833 ^ n28795 ;
  assign n28868 = ~n28866 & ~n28867 ;
  assign n28869 = n28793 ^ n26155 ;
  assign n28870 = n28869 ^ n28836 ;
  assign n28871 = n28868 & ~n28870 ;
  assign n28957 = n28852 & ~n28871 ;
  assign n29311 = n28956 & n28957 ;
  assign n29312 = n29229 ^ n29225 ;
  assign n29313 = n29311 & n29312 ;
  assign n29314 = n29310 & n29313 ;
  assign n29233 = n29232 ^ n29223 ;
  assign n29234 = n29232 ^ n26139 ;
  assign n29235 = ~n29233 & ~n29234 ;
  assign n29236 = n29235 ^ n26139 ;
  assign n29315 = n29236 ^ n26137 ;
  assign n29102 = n29101 ^ n29087 ;
  assign n29103 = ~n29088 & n29102 ;
  assign n29104 = n29103 ^ n29004 ;
  assign n29072 = n28282 ^ n26654 ;
  assign n28998 = n28668 ^ n28667 ;
  assign n29073 = n28998 ^ n27527 ;
  assign n29074 = n29073 ^ n28282 ;
  assign n29075 = n29074 ^ n28998 ;
  assign n29076 = ~n29072 & n29075 ;
  assign n29077 = n29076 ^ n29073 ;
  assign n29237 = n29104 ^ n29077 ;
  assign n29316 = n29315 ^ n29237 ;
  assign n29317 = ~n29314 & ~n29316 ;
  assign n29238 = n29237 ^ n29236 ;
  assign n29108 = n28673 ^ n28633 ;
  assign n29078 = n27525 ^ n26644 ;
  assign n29079 = n28142 ^ n26644 ;
  assign n29080 = n29078 & ~n29079 ;
  assign n29081 = n29080 ^ n27525 ;
  assign n29082 = n29081 ^ n28998 ;
  assign n29083 = n29082 ^ n29081 ;
  assign n29105 = n29104 ^ n29083 ;
  assign n29106 = ~n29077 & n29105 ;
  assign n29107 = n29106 ^ n29082 ;
  assign n29221 = n29108 ^ n29107 ;
  assign n29239 = n29221 ^ n26137 ;
  assign n29240 = n29239 ^ n29221 ;
  assign n29241 = n29240 ^ n29236 ;
  assign n29242 = n29238 & ~n29241 ;
  assign n29243 = n29242 ^ n29239 ;
  assign n29318 = n29243 ^ n26249 ;
  assign n29319 = ~n29317 & n29318 ;
  assign n29222 = n29221 ^ n26249 ;
  assign n29244 = ~n29222 & n29243 ;
  assign n29245 = n29244 ^ n26249 ;
  assign n29307 = n29245 ^ n26350 ;
  assign n29070 = n28679 ^ n28676 ;
  assign n29111 = n29108 ^ n29070 ;
  assign n29109 = n29108 ^ n29081 ;
  assign n29110 = ~n29107 & n29109 ;
  assign n29112 = n29111 ^ n29110 ;
  assign n29066 = n27621 ^ n26888 ;
  assign n29067 = n28135 ^ n26888 ;
  assign n29068 = n29066 & n29067 ;
  assign n29069 = n29068 ^ n27621 ;
  assign n29246 = n29112 ^ n29069 ;
  assign n29308 = n29307 ^ n29246 ;
  assign n29404 = n29319 ^ n29308 ;
  assign n29405 = n29404 ^ n29403 ;
  assign n29436 = n29403 ^ n1572 ;
  assign n29406 = n29318 ^ n29317 ;
  assign n29407 = n29406 ^ n1572 ;
  assign n29408 = n29316 ^ n29314 ;
  assign n29412 = n29411 ^ n29408 ;
  assign n29413 = n29313 ^ n29310 ;
  assign n29417 = n29416 ^ n29413 ;
  assign n29420 = n29312 ^ n29311 ;
  assign n2934 = n2933 ^ n2930 ;
  assign n2935 = n2934 ^ n596 ;
  assign n2939 = n2938 ^ n2935 ;
  assign n29421 = n29420 ^ n2939 ;
  assign n28958 = n28957 ^ n28956 ;
  assign n28873 = n27212 ^ n590 ;
  assign n28874 = n28873 ^ n23884 ;
  assign n28875 = n28874 ^ n18811 ;
  assign n28959 = n28958 ^ n28875 ;
  assign n28872 = n28871 ^ n28852 ;
  assign n28876 = n28875 ^ n28872 ;
  assign n2393 = n2377 ^ n2314 ;
  assign n2394 = n2393 ^ n2390 ;
  assign n2395 = n2394 ^ n1466 ;
  assign n28939 = n28872 ^ n2395 ;
  assign n28877 = n28870 ^ n28868 ;
  assign n28878 = n28877 ^ n2395 ;
  assign n28879 = n28867 ^ n28866 ;
  assign n2381 = n2368 ^ n2305 ;
  assign n2382 = n2381 ^ n2277 ;
  assign n2386 = n2385 ^ n2382 ;
  assign n28880 = n28879 ^ n2386 ;
  assign n28881 = n28865 ^ n28863 ;
  assign n2262 = n2228 ^ n2192 ;
  assign n2263 = n2262 ^ n2259 ;
  assign n2267 = n2266 ^ n2263 ;
  assign n28882 = n28881 ^ n2267 ;
  assign n28883 = n28862 ^ n28861 ;
  assign n2250 = n2180 ^ n2130 ;
  assign n2251 = n2250 ^ n2249 ;
  assign n2252 = n2251 ^ n2240 ;
  assign n28884 = n28883 ^ n2252 ;
  assign n28888 = n27222 ^ n2115 ;
  assign n28889 = n28888 ^ n23898 ;
  assign n28890 = n28889 ^ n2247 ;
  assign n28887 = n28860 ^ n28859 ;
  assign n28891 = n28890 ^ n28887 ;
  assign n28895 = n28858 ^ n28856 ;
  assign n28892 = n27226 ^ n2108 ;
  assign n28893 = n28892 ^ n23902 ;
  assign n28894 = n28893 ^ n1976 ;
  assign n28896 = n28895 ^ n28894 ;
  assign n28900 = n28855 ^ n28854 ;
  assign n28922 = n28900 ^ n28894 ;
  assign n28897 = n27240 ^ n19844 ;
  assign n28898 = n28897 ^ n1910 ;
  assign n28899 = n28898 ^ n18828 ;
  assign n28901 = n28900 ^ n28899 ;
  assign n28907 = n28806 ^ n28805 ;
  assign n28911 = n28907 ^ n28854 ;
  assign n28906 = n28904 & n28905 ;
  assign n28908 = n28907 ^ n28906 ;
  assign n28909 = n28906 ^ n1868 ;
  assign n28910 = n28908 & ~n28909 ;
  assign n28912 = n28911 ^ n28910 ;
  assign n28917 = n28899 ^ n28854 ;
  assign n28913 = n27230 ^ n19851 ;
  assign n28914 = n28913 ^ n23907 ;
  assign n28915 = n28914 ^ n1905 ;
  assign n28916 = n28915 ^ n28899 ;
  assign n28918 = n28917 ^ n28916 ;
  assign n28919 = ~n28912 & ~n28918 ;
  assign n28920 = n28919 ^ n28917 ;
  assign n28921 = n28901 & n28920 ;
  assign n28923 = n28922 ^ n28921 ;
  assign n28924 = n28896 & ~n28923 ;
  assign n28925 = n28924 ^ n28895 ;
  assign n28926 = n28925 ^ n28887 ;
  assign n28927 = ~n28891 & n28926 ;
  assign n28928 = n28927 ^ n28890 ;
  assign n28885 = n2267 ^ n2252 ;
  assign n28886 = n28885 ^ n2267 ;
  assign n28929 = n28928 ^ n28886 ;
  assign n28930 = n28884 & n28929 ;
  assign n28931 = n28930 ^ n28885 ;
  assign n28932 = ~n28882 & ~n28931 ;
  assign n28933 = n28932 ^ n28881 ;
  assign n28934 = n28933 ^ n2386 ;
  assign n28935 = n28880 & n28934 ;
  assign n28936 = n28935 ^ n28879 ;
  assign n28937 = n28936 ^ n2395 ;
  assign n28938 = ~n28878 & n28937 ;
  assign n28940 = n28939 ^ n28938 ;
  assign n28941 = n28876 & ~n28940 ;
  assign n28960 = n28959 ^ n28941 ;
  assign n29423 = n28958 ^ n2939 ;
  assign n29422 = n28963 ^ n2939 ;
  assign n29424 = n29423 ^ n29422 ;
  assign n29425 = n28960 & ~n29424 ;
  assign n29426 = n29425 ^ n29422 ;
  assign n29427 = ~n29421 & ~n29426 ;
  assign n29428 = n29427 ^ n29420 ;
  assign n29429 = n29428 ^ n29416 ;
  assign n29430 = ~n29417 & ~n29429 ;
  assign n29418 = n29416 ^ n29411 ;
  assign n29431 = n29430 ^ n29418 ;
  assign n29432 = n29412 & n29431 ;
  assign n29433 = n29432 ^ n29411 ;
  assign n29434 = n29433 ^ n29406 ;
  assign n29435 = n29407 & ~n29434 ;
  assign n29437 = n29436 ^ n29435 ;
  assign n29438 = n29405 & ~n29437 ;
  assign n29439 = n29438 ^ n29404 ;
  assign n29247 = n29246 ^ n29245 ;
  assign n29248 = n29246 ^ n26350 ;
  assign n29249 = n29247 & n29248 ;
  assign n29250 = n29249 ^ n26350 ;
  assign n29071 = n29070 ^ n29069 ;
  assign n29113 = n29071 & n29112 ;
  assign n29114 = n29113 ^ n29070 ;
  assign n29060 = n28129 ^ n26640 ;
  assign n28992 = n28683 ^ n28630 ;
  assign n29061 = n28992 ^ n27700 ;
  assign n29062 = n29061 ^ n28129 ;
  assign n29063 = n29062 ^ n28992 ;
  assign n29064 = n29060 & n29063 ;
  assign n29065 = n29064 ^ n29061 ;
  assign n29219 = n29114 ^ n29065 ;
  assign n29220 = n29219 ^ n26398 ;
  assign n29321 = n29250 ^ n29220 ;
  assign n29320 = ~n29308 & n29319 ;
  assign n29399 = n29321 ^ n29320 ;
  assign n29400 = n29399 ^ n811 ;
  assign n30028 = n29439 ^ n29400 ;
  assign n29178 = n28713 ^ n28605 ;
  assign n30010 = n29178 ^ n28341 ;
  assign n30015 = n29437 ^ n29404 ;
  assign n29039 = n28711 ^ n28606 ;
  assign n30011 = n29039 ^ n28105 ;
  assign n30012 = n28105 ^ n27917 ;
  assign n30013 = n30011 & ~n30012 ;
  assign n30014 = n30013 ^ n27917 ;
  assign n30016 = n30015 ^ n30014 ;
  assign n29890 = n29433 ^ n29407 ;
  assign n29709 = n29431 ^ n29408 ;
  assign n29891 = n29890 ^ n29709 ;
  assign n29163 = n28704 ^ n28611 ;
  assign n29708 = n29163 ^ n28112 ;
  assign n29710 = n29709 ^ n27766 ;
  assign n29711 = n29710 ^ n29163 ;
  assign n29712 = n29711 ^ n29709 ;
  assign n29713 = ~n29708 & n29712 ;
  assign n29714 = n29713 ^ n29710 ;
  assign n29159 = n28702 ^ n28612 ;
  assign n29604 = n29159 ^ n28126 ;
  assign n29605 = n28126 ^ n27750 ;
  assign n29606 = n29604 & ~n29605 ;
  assign n29607 = n29606 ^ n27750 ;
  assign n29603 = n29428 ^ n29417 ;
  assign n29608 = n29607 ^ n29603 ;
  assign n29593 = n29426 ^ n29420 ;
  assign n28965 = n28694 ^ n28615 ;
  assign n28966 = n28965 ^ n28310 ;
  assign n28967 = n28310 ^ n27621 ;
  assign n28968 = ~n28966 & n28967 ;
  assign n28969 = n28968 ^ n27621 ;
  assign n28964 = n28963 ^ n28960 ;
  assign n28970 = n28969 ^ n28964 ;
  assign n28972 = n28691 ^ n28619 ;
  assign n28973 = n28972 ^ n28129 ;
  assign n28974 = n28129 ^ n27525 ;
  assign n28975 = ~n28973 & n28974 ;
  assign n28976 = n28975 ^ n27525 ;
  assign n28971 = n28940 ^ n28875 ;
  assign n28977 = n28976 ^ n28971 ;
  assign n28979 = n28135 ^ n27527 ;
  assign n28980 = n28689 ^ n28622 ;
  assign n28981 = n28980 ^ n28135 ;
  assign n28982 = n28979 & ~n28981 ;
  assign n28983 = n28982 ^ n27527 ;
  assign n28978 = n28936 ^ n28878 ;
  assign n28984 = n28983 ^ n28978 ;
  assign n28986 = n28685 ^ n28626 ;
  assign n28987 = n28986 ^ n28142 ;
  assign n28988 = n28142 ^ n27534 ;
  assign n28989 = ~n28987 & n28988 ;
  assign n28990 = n28989 ^ n27534 ;
  assign n29583 = n28990 ^ n28983 ;
  assign n28985 = n28933 ^ n28880 ;
  assign n28991 = n28990 ^ n28985 ;
  assign n28993 = n28992 ^ n28282 ;
  assign n28994 = n28282 ^ n27536 ;
  assign n28995 = n28993 & ~n28994 ;
  assign n28996 = n28995 ^ n27536 ;
  assign n29580 = n28996 ^ n28990 ;
  assign n29567 = n28928 ^ n28884 ;
  assign n29555 = n28925 ^ n28891 ;
  assign n28999 = n28998 ^ n28157 ;
  assign n29000 = n28157 ^ n27517 ;
  assign n29001 = n28999 & n29000 ;
  assign n29002 = n29001 ^ n27517 ;
  assign n28997 = n28923 ^ n28895 ;
  assign n29003 = n29002 ^ n28997 ;
  assign n29009 = n28920 ^ n28900 ;
  assign n29005 = n29004 ^ n28170 ;
  assign n29006 = n28170 ^ n27554 ;
  assign n29007 = ~n29005 & ~n29006 ;
  assign n29008 = n29007 ^ n27554 ;
  assign n29010 = n29009 ^ n29008 ;
  assign n29018 = n28915 ^ n28912 ;
  assign n29548 = n29018 ^ n29008 ;
  assign n29011 = n28945 ^ n28177 ;
  assign n29012 = n28909 ^ n28907 ;
  assign n29013 = n29012 ^ n27562 ;
  assign n29014 = n29013 ^ n28945 ;
  assign n29015 = n29014 ^ n29012 ;
  assign n29016 = n29011 & n29015 ;
  assign n29017 = n29016 ^ n29013 ;
  assign n29020 = n28844 ^ n28075 ;
  assign n29022 = n29021 ^ n27567 ;
  assign n29023 = n29022 ^ n29021 ;
  assign n29024 = n29023 ^ n28844 ;
  assign n29025 = n29020 & n29024 ;
  assign n29026 = n29025 ^ n29022 ;
  assign n29490 = n28082 ^ n27577 ;
  assign n29491 = n28082 ^ n28069 ;
  assign n29492 = ~n29490 & n29491 ;
  assign n29493 = n29492 ^ n27577 ;
  assign n29206 = n28722 ^ n28599 ;
  assign n29027 = n28004 ^ n26693 ;
  assign n29028 = n27951 ^ n27338 ;
  assign n29029 = n28719 ^ n28601 ;
  assign n29030 = n29029 ^ n26777 ;
  assign n29031 = n29030 ^ n27951 ;
  assign n29032 = n29031 ^ n29029 ;
  assign n29033 = ~n29028 & n29032 ;
  assign n29034 = n29033 ^ n29030 ;
  assign n29188 = n28716 ^ n28603 ;
  assign n29035 = n27352 ^ n26787 ;
  assign n29036 = n28558 ^ n27352 ;
  assign n29037 = ~n29035 & ~n29036 ;
  assign n29038 = n29037 ^ n26787 ;
  assign n29040 = n29039 ^ n29038 ;
  assign n29041 = n28480 ^ n27350 ;
  assign n29042 = n28707 ^ n28609 ;
  assign n29043 = n29042 ^ n26600 ;
  assign n29044 = n29043 ^ n28480 ;
  assign n29045 = n29044 ^ n29042 ;
  assign n29046 = ~n29041 & n29045 ;
  assign n29047 = n29046 ^ n29043 ;
  assign n29125 = n28980 ^ n28972 ;
  assign n29050 = n28310 ^ n26635 ;
  assign n29051 = n28986 ^ n27750 ;
  assign n29052 = n29051 ^ n28310 ;
  assign n29053 = n29052 ^ n28986 ;
  assign n29054 = ~n29050 & ~n29053 ;
  assign n29055 = n29054 ^ n29051 ;
  assign n29056 = n27766 ^ n26628 ;
  assign n29057 = n28316 ^ n27766 ;
  assign n29058 = ~n29056 & n29057 ;
  assign n29059 = n29058 ^ n26628 ;
  assign n29119 = n29059 ^ n28986 ;
  assign n29115 = n29114 ^ n28992 ;
  assign n29116 = n29065 & n29115 ;
  assign n29117 = n29116 ^ n28992 ;
  assign n29118 = n29117 ^ n29059 ;
  assign n29120 = n29119 ^ n29118 ;
  assign n29121 = ~n29055 & n29120 ;
  assign n29122 = n29121 ^ n29119 ;
  assign n29123 = n29059 ^ n28980 ;
  assign n29124 = ~n29122 & ~n29123 ;
  assign n29126 = n29125 ^ n29124 ;
  assign n29132 = n27892 ^ n26623 ;
  assign n29133 = n28126 ^ n27892 ;
  assign n29134 = ~n29132 & n29133 ;
  assign n29135 = n29134 ^ n26623 ;
  assign n29127 = n27917 ^ n26619 ;
  assign n29128 = n28112 ^ n27917 ;
  assign n29129 = ~n29127 & ~n29128 ;
  assign n29130 = n29129 ^ n26619 ;
  assign n29131 = n29130 ^ n28972 ;
  assign n29136 = n29135 ^ n29131 ;
  assign n29137 = n29136 ^ n29130 ;
  assign n29138 = ~n29126 & n29137 ;
  assign n29139 = n29138 ^ n29131 ;
  assign n29140 = n27938 ^ n26907 ;
  assign n29141 = n28329 ^ n27938 ;
  assign n29142 = n29140 & n29141 ;
  assign n29143 = n29142 ^ n26907 ;
  assign n29144 = n29143 ^ n28965 ;
  assign n29145 = n29144 ^ n29130 ;
  assign n29146 = n29145 ^ n29143 ;
  assign n29147 = ~n29139 & n29146 ;
  assign n29148 = n29147 ^ n29144 ;
  assign n29154 = n28698 ^ n28697 ;
  assign n29149 = n27989 ^ n26613 ;
  assign n29150 = n28105 ^ n27989 ;
  assign n29151 = n29149 & ~n29150 ;
  assign n29152 = n29151 ^ n26613 ;
  assign n29155 = n29154 ^ n29152 ;
  assign n29153 = n29152 ^ n29143 ;
  assign n29156 = n29155 ^ n29153 ;
  assign n29157 = n29148 & n29156 ;
  assign n29158 = n29157 ^ n29155 ;
  assign n29160 = n29159 ^ n29152 ;
  assign n29161 = n29158 & ~n29160 ;
  assign n29162 = n29161 ^ n29159 ;
  assign n29164 = n29163 ^ n29162 ;
  assign n29165 = n28341 ^ n28043 ;
  assign n29166 = n29163 ^ n27145 ;
  assign n29167 = n29166 ^ n28341 ;
  assign n29168 = n29167 ^ n29163 ;
  assign n29169 = ~n29165 & ~n29168 ;
  assign n29170 = n29169 ^ n29166 ;
  assign n29171 = n29164 & n29170 ;
  assign n29172 = n29171 ^ n29163 ;
  assign n29173 = n29172 ^ n29042 ;
  assign n29174 = ~n29047 & n29173 ;
  assign n29048 = n29042 ^ n29038 ;
  assign n29175 = n29174 ^ n29048 ;
  assign n29176 = n29040 & ~n29175 ;
  assign n29177 = n29176 ^ n29039 ;
  assign n29179 = n29178 ^ n29177 ;
  assign n29180 = n27898 ^ n27344 ;
  assign n29181 = n29178 ^ n26791 ;
  assign n29182 = n29181 ^ n27898 ;
  assign n29183 = n29182 ^ n29178 ;
  assign n29184 = n29180 & n29183 ;
  assign n29185 = n29184 ^ n29181 ;
  assign n29186 = ~n29179 & ~n29185 ;
  assign n29187 = n29186 ^ n29178 ;
  assign n29189 = n29188 ^ n29187 ;
  assign n29190 = n27952 ^ n27342 ;
  assign n29191 = n29188 ^ n26799 ;
  assign n29192 = n29191 ^ n27952 ;
  assign n29193 = n29192 ^ n29188 ;
  assign n29194 = n29190 & n29193 ;
  assign n29195 = n29194 ^ n29191 ;
  assign n29196 = ~n29189 & ~n29195 ;
  assign n29197 = n29196 ^ n29188 ;
  assign n29198 = n29197 ^ n29029 ;
  assign n29199 = ~n29034 & n29198 ;
  assign n29200 = n29199 ^ n29029 ;
  assign n29201 = n29200 ^ n26605 ;
  assign n29202 = n29201 ^ n28004 ;
  assign n29203 = n29202 ^ n29200 ;
  assign n29204 = n29027 & n29203 ;
  assign n29205 = n29204 ^ n29201 ;
  assign n29207 = n29206 ^ n29205 ;
  assign n29368 = n29207 ^ n26102 ;
  assign n29208 = n29195 ^ n29187 ;
  assign n29209 = n29208 ^ n26046 ;
  assign n29210 = n29185 ^ n29177 ;
  assign n29211 = n29210 ^ n26003 ;
  assign n29284 = n29172 ^ n29047 ;
  assign n29213 = n29170 ^ n29162 ;
  assign n29214 = n29213 ^ n26626 ;
  assign n29216 = n29154 ^ n29148 ;
  assign n29217 = n29216 ^ n26637 ;
  assign n29264 = n29135 ^ n29126 ;
  assign n29259 = n29122 ^ n28980 ;
  assign n29251 = n29250 ^ n29219 ;
  assign n29252 = n29220 & ~n29251 ;
  assign n29253 = n29252 ^ n26398 ;
  assign n29254 = n29253 ^ n26413 ;
  assign n29255 = n29117 ^ n29055 ;
  assign n29256 = n29255 ^ n29253 ;
  assign n29257 = ~n29254 & n29256 ;
  assign n29258 = n29257 ^ n26413 ;
  assign n29260 = n29259 ^ n29258 ;
  assign n29261 = n29259 ^ n26429 ;
  assign n29262 = ~n29260 & ~n29261 ;
  assign n29263 = n29262 ^ n26429 ;
  assign n29265 = n29264 ^ n29263 ;
  assign n29266 = n29264 ^ n26583 ;
  assign n29267 = n29265 & n29266 ;
  assign n29268 = n29267 ^ n26583 ;
  assign n29218 = n29139 ^ n28965 ;
  assign n29269 = n29268 ^ n29218 ;
  assign n29270 = n29268 ^ n26646 ;
  assign n29271 = n29269 & n29270 ;
  assign n29272 = n29271 ^ n26646 ;
  assign n29273 = n29272 ^ n29216 ;
  assign n29274 = n29217 & n29273 ;
  assign n29275 = n29274 ^ n26637 ;
  assign n29215 = n29159 ^ n29158 ;
  assign n29276 = n29275 ^ n29215 ;
  assign n29277 = n29213 ^ n26633 ;
  assign n29278 = n29277 ^ n29213 ;
  assign n29279 = n29278 ^ n29215 ;
  assign n29280 = ~n29276 & n29279 ;
  assign n29281 = n29280 ^ n29277 ;
  assign n29282 = n29214 & n29281 ;
  assign n29283 = n29282 ^ n26626 ;
  assign n29285 = n29284 ^ n29283 ;
  assign n29286 = n29284 ^ n25952 ;
  assign n29287 = n29285 & n29286 ;
  assign n29288 = n29287 ^ n25952 ;
  assign n29212 = n29175 ^ n29039 ;
  assign n29289 = n29288 ^ n29212 ;
  assign n29290 = n29288 ^ n25978 ;
  assign n29291 = n29289 & n29290 ;
  assign n29292 = n29291 ^ n25978 ;
  assign n29293 = n29292 ^ n29210 ;
  assign n29294 = ~n29211 & ~n29293 ;
  assign n29295 = n29294 ^ n26003 ;
  assign n29296 = n29295 ^ n29208 ;
  assign n29297 = n29209 & ~n29296 ;
  assign n29298 = n29297 ^ n26046 ;
  assign n29299 = n29298 ^ n26081 ;
  assign n29300 = n29197 ^ n29034 ;
  assign n29301 = n29300 ^ n29298 ;
  assign n29302 = n29299 & n29301 ;
  assign n29303 = n29302 ^ n26081 ;
  assign n29369 = n29368 ^ n29303 ;
  assign n29306 = n29295 ^ n29209 ;
  assign n29322 = n29320 & n29321 ;
  assign n29323 = n29255 ^ n29254 ;
  assign n29324 = ~n29322 & ~n29323 ;
  assign n29325 = n29258 ^ n26429 ;
  assign n29326 = n29325 ^ n29259 ;
  assign n29327 = ~n29324 & n29326 ;
  assign n29328 = n29263 ^ n26583 ;
  assign n29329 = n29328 ^ n29264 ;
  assign n29330 = n29327 & n29329 ;
  assign n29331 = n29270 ^ n29218 ;
  assign n29332 = ~n29330 & ~n29331 ;
  assign n29333 = n29272 ^ n29217 ;
  assign n29334 = n29332 & n29333 ;
  assign n29335 = n29215 ^ n26633 ;
  assign n29336 = n29335 ^ n29275 ;
  assign n29337 = n29334 & ~n29336 ;
  assign n29338 = n29281 ^ n26626 ;
  assign n29339 = ~n29337 & n29338 ;
  assign n29340 = n29286 ^ n29283 ;
  assign n29341 = n29339 & ~n29340 ;
  assign n29342 = n29290 ^ n29212 ;
  assign n29343 = n29341 & ~n29342 ;
  assign n29344 = n29292 ^ n29211 ;
  assign n29345 = n29343 & ~n29344 ;
  assign n29346 = n29306 & ~n29345 ;
  assign n29347 = n29300 ^ n29299 ;
  assign n29348 = n29346 & ~n29347 ;
  assign n29370 = n29369 ^ n29348 ;
  assign n29371 = n29370 ^ n2534 ;
  assign n29373 = n29345 ^ n29306 ;
  assign n2583 = n2582 ^ n2492 ;
  assign n2593 = n2592 ^ n2583 ;
  assign n2597 = n2596 ^ n2593 ;
  assign n29374 = n29373 ^ n2597 ;
  assign n29376 = n27168 ^ n2627 ;
  assign n29377 = n29376 ^ n24002 ;
  assign n29378 = n29377 ^ n2590 ;
  assign n29375 = n29344 ^ n29343 ;
  assign n29379 = n29378 ^ n29375 ;
  assign n29467 = n2867 ^ n2565 ;
  assign n29468 = n29467 ^ n3110 ;
  assign n29469 = n29468 ^ n18780 ;
  assign n29470 = n29469 ^ n2857 ;
  assign n29380 = n29338 ^ n29337 ;
  assign n29381 = n29380 ^ n2842 ;
  assign n29385 = n1410 ^ n1331 ;
  assign n29386 = n29385 ^ n1259 ;
  assign n29387 = n29386 ^ n2834 ;
  assign n29384 = n29336 ^ n29334 ;
  assign n29388 = n29387 ^ n29384 ;
  assign n29389 = n29333 ^ n29332 ;
  assign n1744 = n1418 ^ n1313 ;
  assign n1745 = n1744 ^ n1738 ;
  assign n1746 = n1745 ^ n1250 ;
  assign n29390 = n29389 ^ n1746 ;
  assign n29391 = n29331 ^ n29330 ;
  assign n1068 = n1067 ^ n983 ;
  assign n1069 = n1068 ^ n1064 ;
  assign n1070 = n1069 ^ n1055 ;
  assign n29392 = n29391 ^ n1070 ;
  assign n29393 = n29329 ^ n29327 ;
  assign n1726 = n1707 ^ n1295 ;
  assign n1727 = n1726 ^ n908 ;
  assign n1728 = n1727 ^ n1058 ;
  assign n29394 = n29393 ^ n1728 ;
  assign n29395 = n29326 ^ n29324 ;
  assign n29396 = n29395 ^ n921 ;
  assign n29397 = n29323 ^ n29322 ;
  assign n29398 = n29397 ^ n826 ;
  assign n29440 = n29439 ^ n811 ;
  assign n29441 = ~n29400 & ~n29440 ;
  assign n29442 = n29441 ^ n29399 ;
  assign n29443 = n29442 ^ n826 ;
  assign n29444 = n29398 & n29443 ;
  assign n29445 = n29444 ^ n29397 ;
  assign n29446 = n29445 ^ n921 ;
  assign n29447 = n29396 & ~n29446 ;
  assign n29448 = n29447 ^ n29395 ;
  assign n29449 = n29448 ^ n1728 ;
  assign n29450 = ~n29394 & ~n29449 ;
  assign n29451 = n29450 ^ n29393 ;
  assign n29452 = n29451 ^ n29391 ;
  assign n29453 = n29392 & n29452 ;
  assign n29454 = n29453 ^ n1070 ;
  assign n29455 = n29454 ^ n1746 ;
  assign n29456 = n29390 & ~n29455 ;
  assign n29457 = n29456 ^ n29389 ;
  assign n29458 = n29457 ^ n29384 ;
  assign n29459 = ~n29388 & n29458 ;
  assign n29460 = n29459 ^ n29387 ;
  assign n29461 = n29460 ^ n2842 ;
  assign n29462 = n29381 & n29461 ;
  assign n29382 = n2857 ^ n2842 ;
  assign n29463 = n29462 ^ n29382 ;
  assign n29464 = n29340 ^ n29339 ;
  assign n29465 = n29464 ^ n2857 ;
  assign n29466 = n29463 & n29465 ;
  assign n29471 = n29470 ^ n29466 ;
  assign n29474 = n29342 ^ n29341 ;
  assign n29475 = n29474 ^ n29469 ;
  assign n29476 = n29471 & n29475 ;
  assign n29472 = n29469 ^ n29375 ;
  assign n29477 = n29476 ^ n29472 ;
  assign n29478 = n29379 & ~n29477 ;
  assign n29479 = n29478 ^ n29378 ;
  assign n29480 = n29479 ^ n29373 ;
  assign n29481 = ~n29374 & n29480 ;
  assign n29482 = n29481 ^ n2597 ;
  assign n29372 = n29347 ^ n29346 ;
  assign n29483 = n29482 ^ n29372 ;
  assign n29484 = n29482 ^ n3221 ;
  assign n29485 = n29483 & n29484 ;
  assign n29486 = n29485 ^ n3221 ;
  assign n29487 = n29486 ^ n2534 ;
  assign n29488 = n29371 & n29487 ;
  assign n29366 = n3233 ^ n2534 ;
  assign n29360 = n29200 ^ n26691 ;
  assign n29359 = n28725 ^ n28592 ;
  assign n29361 = n29360 ^ n29359 ;
  assign n29362 = n29361 ^ n26201 ;
  assign n29357 = n29206 ^ n29200 ;
  assign n29358 = ~n29205 & n29357 ;
  assign n29363 = n29362 ^ n29358 ;
  assign n29354 = n28055 ^ n27373 ;
  assign n29355 = n27373 ^ n26691 ;
  assign n29356 = ~n29354 & n29355 ;
  assign n29364 = n29363 ^ n29356 ;
  assign n29304 = n29303 ^ n29207 ;
  assign n29349 = n29348 ^ n29207 ;
  assign n29352 = n29304 & n29349 ;
  assign n29350 = n29349 ^ n29303 ;
  assign n29351 = n26102 & n29350 ;
  assign n29353 = n29352 ^ n29351 ;
  assign n29365 = n29364 ^ n29353 ;
  assign n29367 = n29366 ^ n29365 ;
  assign n29489 = n29488 ^ n29367 ;
  assign n29494 = n29493 ^ n29489 ;
  assign n29495 = n28100 ^ n28080 ;
  assign n29496 = n29372 ^ n3221 ;
  assign n29497 = n29496 ^ n29482 ;
  assign n29498 = n29497 ^ n27502 ;
  assign n29499 = n29498 ^ n28100 ;
  assign n29500 = n29499 ^ n29497 ;
  assign n29501 = n29495 & n29500 ;
  assign n29502 = n29501 ^ n29498 ;
  assign n29518 = n28090 ^ n27576 ;
  assign n29519 = n28783 ^ n28090 ;
  assign n29520 = ~n29518 & n29519 ;
  assign n29521 = n29520 ^ n27576 ;
  assign n29523 = n29521 ^ n29497 ;
  assign n29507 = n29477 ^ n29378 ;
  assign n29508 = n28211 ^ n27412 ;
  assign n29509 = n28211 ^ n28092 ;
  assign n29510 = n29508 & n29509 ;
  assign n29511 = n29510 ^ n27412 ;
  assign n29512 = n29507 & n29511 ;
  assign n29503 = n28201 ^ n27485 ;
  assign n29504 = n28201 ^ n28088 ;
  assign n29505 = n29503 & n29504 ;
  assign n29506 = n29505 ^ n27485 ;
  assign n29513 = n29512 ^ n29506 ;
  assign n29514 = n29479 ^ n29374 ;
  assign n29515 = n29514 ^ n29506 ;
  assign n29516 = ~n29513 & n29515 ;
  assign n29517 = n29516 ^ n29506 ;
  assign n29522 = n29521 ^ n29517 ;
  assign n29524 = n29523 ^ n29522 ;
  assign n29525 = n29502 & n29524 ;
  assign n29526 = n29525 ^ n29523 ;
  assign n29528 = n29486 ^ n29371 ;
  assign n29529 = n29528 ^ n29493 ;
  assign n29527 = n29521 ^ n29493 ;
  assign n29530 = n29529 ^ n29527 ;
  assign n29531 = n29526 & ~n29530 ;
  assign n29532 = n29531 ^ n29527 ;
  assign n29533 = ~n29494 & ~n29532 ;
  assign n29534 = n29533 ^ n29493 ;
  assign n29535 = n29534 ^ n29021 ;
  assign n29536 = n29026 & n29535 ;
  assign n29537 = n29536 ^ n29021 ;
  assign n29538 = n29537 ^ n29018 ;
  assign n29019 = n29018 ^ n29012 ;
  assign n29539 = n29538 ^ n29019 ;
  assign n29540 = n29017 & n29539 ;
  assign n29541 = n29540 ^ n29019 ;
  assign n29542 = n27558 ^ n27516 ;
  assign n29543 = n29092 ^ n27516 ;
  assign n29544 = n29542 & ~n29543 ;
  assign n29545 = n29544 ^ n27558 ;
  assign n29546 = n29545 ^ n29018 ;
  assign n29547 = ~n29541 & n29546 ;
  assign n29549 = n29548 ^ n29547 ;
  assign n29550 = ~n29010 & n29549 ;
  assign n29551 = n29550 ^ n29009 ;
  assign n29552 = n29551 ^ n28997 ;
  assign n29553 = n29003 & n29552 ;
  assign n29554 = n29553 ^ n29002 ;
  assign n29556 = n29555 ^ n29554 ;
  assign n29557 = n29108 ^ n28155 ;
  assign n29558 = n29555 ^ n27547 ;
  assign n29559 = n29558 ^ n29108 ;
  assign n29560 = n29559 ^ n29555 ;
  assign n29561 = n29557 & n29560 ;
  assign n29562 = n29561 ^ n29558 ;
  assign n29563 = ~n29556 & n29562 ;
  assign n29564 = n29563 ^ n29555 ;
  assign n29568 = n29567 ^ n29564 ;
  assign n29569 = n29070 ^ n28278 ;
  assign n29570 = n29567 ^ n27543 ;
  assign n29571 = n29570 ^ n29070 ;
  assign n29572 = n29571 ^ n29567 ;
  assign n29573 = ~n29569 & n29572 ;
  assign n29574 = n29573 ^ n29570 ;
  assign n29575 = ~n29568 & n29574 ;
  assign n29565 = n29564 ^ n28996 ;
  assign n29576 = n29575 ^ n29565 ;
  assign n29577 = n28931 ^ n28881 ;
  assign n29578 = n29577 ^ n28996 ;
  assign n29579 = n29576 & n29578 ;
  assign n29581 = n29580 ^ n29579 ;
  assign n29582 = n28991 & n29581 ;
  assign n29584 = n29583 ^ n29582 ;
  assign n29585 = ~n28984 & ~n29584 ;
  assign n29586 = n29585 ^ n28983 ;
  assign n29587 = n29586 ^ n28971 ;
  assign n29588 = ~n28977 & ~n29587 ;
  assign n29589 = n29588 ^ n28976 ;
  assign n29590 = n29589 ^ n28964 ;
  assign n29591 = n28970 & ~n29590 ;
  assign n29592 = n29591 ^ n28969 ;
  assign n29594 = n29593 ^ n29592 ;
  assign n29595 = n29154 ^ n28316 ;
  assign n29596 = n29593 ^ n27700 ;
  assign n29597 = n29596 ^ n29154 ;
  assign n29598 = n29597 ^ n29593 ;
  assign n29599 = n29595 & ~n29598 ;
  assign n29600 = n29599 ^ n29596 ;
  assign n29601 = n29594 & n29600 ;
  assign n29602 = n29601 ^ n29593 ;
  assign n29705 = n29603 ^ n29602 ;
  assign n29706 = n29608 & n29705 ;
  assign n29707 = n29706 ^ n29607 ;
  assign n29888 = n29709 ^ n29707 ;
  assign n29889 = n29714 & n29888 ;
  assign n29892 = n29891 ^ n29889 ;
  assign n29893 = n29042 ^ n28329 ;
  assign n29894 = n28329 ^ n27892 ;
  assign n29895 = n29893 & ~n29894 ;
  assign n29896 = n29895 ^ n27892 ;
  assign n30017 = n29896 ^ n29890 ;
  assign n30018 = n29892 & n30017 ;
  assign n30019 = n30018 ^ n29890 ;
  assign n30020 = n30019 ^ n30014 ;
  assign n30021 = n30016 & ~n30020 ;
  assign n30022 = n30021 ^ n30015 ;
  assign n30023 = n30022 ^ n27938 ;
  assign n30024 = n30023 ^ n29178 ;
  assign n30025 = n30024 ^ n30022 ;
  assign n30026 = ~n30010 & ~n30025 ;
  assign n30027 = n30026 ^ n30023 ;
  assign n30058 = n30028 ^ n30027 ;
  assign n30059 = n30058 ^ n26907 ;
  assign n29897 = n29896 ^ n29892 ;
  assign n29898 = n29897 ^ n26623 ;
  assign n29715 = n29714 ^ n29707 ;
  assign n29716 = n29715 ^ n26628 ;
  assign n29609 = n29608 ^ n29602 ;
  assign n29610 = n29609 ^ n26635 ;
  assign n29611 = n29600 ^ n29592 ;
  assign n29612 = n29611 ^ n26640 ;
  assign n29613 = n29589 ^ n28970 ;
  assign n29614 = n29613 ^ n26888 ;
  assign n29615 = n29586 ^ n28977 ;
  assign n29616 = n29615 ^ n26644 ;
  assign n29617 = n29584 ^ n28978 ;
  assign n29618 = n29617 ^ n26654 ;
  assign n29620 = n29577 ^ n29576 ;
  assign n29621 = n29620 ^ n26874 ;
  assign n29622 = n29574 ^ n29564 ;
  assign n29623 = n29622 ^ n26868 ;
  assign n29624 = n29562 ^ n29554 ;
  assign n29625 = n29624 ^ n26860 ;
  assign n29626 = n29551 ^ n29003 ;
  assign n29627 = n29626 ^ n26841 ;
  assign n29628 = n29549 ^ n29009 ;
  assign n29629 = n29628 ^ n26833 ;
  assign n29630 = n29545 ^ n29541 ;
  assign n29631 = n29630 ^ n26664 ;
  assign n29651 = n29532 ^ n29489 ;
  assign n29633 = n29528 ^ n29526 ;
  assign n29634 = n29633 ^ n26131 ;
  assign n29635 = n29517 ^ n29502 ;
  assign n29636 = n29635 ^ n26608 ;
  assign n29638 = n29511 ^ n29507 ;
  assign n29639 = ~n26687 & n29638 ;
  assign n29637 = n29514 ^ n29513 ;
  assign n29640 = n29639 ^ n29637 ;
  assign n29641 = n29635 ^ n26683 ;
  assign n29642 = n29641 ^ n29635 ;
  assign n29643 = n29642 ^ n29637 ;
  assign n29644 = ~n29640 & ~n29643 ;
  assign n29645 = n29644 ^ n29641 ;
  assign n29646 = n29636 & ~n29645 ;
  assign n29647 = n29646 ^ n26608 ;
  assign n29648 = n29647 ^ n29633 ;
  assign n29649 = n29634 & n29648 ;
  assign n29650 = n29649 ^ n26131 ;
  assign n29652 = n29651 ^ n29650 ;
  assign n29653 = n29651 ^ n26671 ;
  assign n29654 = ~n29652 & ~n29653 ;
  assign n29655 = n29654 ^ n26671 ;
  assign n29632 = n29534 ^ n29026 ;
  assign n29656 = n29655 ^ n29632 ;
  assign n29657 = n29537 ^ n29017 ;
  assign n29658 = n29657 ^ n26669 ;
  assign n29659 = n29658 ^ n29632 ;
  assign n29660 = n29659 ^ n29657 ;
  assign n29661 = n29656 & ~n29660 ;
  assign n29662 = n29661 ^ n29658 ;
  assign n29664 = n29630 ^ n26662 ;
  assign n29663 = n29657 ^ n29630 ;
  assign n29665 = n29664 ^ n29663 ;
  assign n29666 = n29662 & ~n29665 ;
  assign n29667 = n29666 ^ n29664 ;
  assign n29668 = n29631 & n29667 ;
  assign n29669 = n29668 ^ n26664 ;
  assign n29670 = n29669 ^ n29628 ;
  assign n29671 = n29629 & ~n29670 ;
  assign n29672 = n29671 ^ n26833 ;
  assign n29673 = n29672 ^ n29626 ;
  assign n29674 = n29627 & n29673 ;
  assign n29675 = n29674 ^ n26841 ;
  assign n29676 = n29675 ^ n29624 ;
  assign n29677 = ~n29625 & n29676 ;
  assign n29678 = n29677 ^ n26860 ;
  assign n29679 = n29678 ^ n29622 ;
  assign n29680 = ~n29623 & n29679 ;
  assign n29681 = n29680 ^ n26868 ;
  assign n29682 = n29681 ^ n29620 ;
  assign n29683 = n29621 & ~n29682 ;
  assign n29684 = n29683 ^ n26874 ;
  assign n29619 = n29581 ^ n28985 ;
  assign n29685 = n29684 ^ n29619 ;
  assign n29686 = n29617 ^ n26658 ;
  assign n29687 = n29686 ^ n29617 ;
  assign n29688 = n29687 ^ n29619 ;
  assign n29689 = ~n29685 & ~n29688 ;
  assign n29690 = n29689 ^ n29686 ;
  assign n29691 = n29618 & ~n29690 ;
  assign n29692 = n29691 ^ n26654 ;
  assign n29693 = n29692 ^ n29615 ;
  assign n29694 = n29616 & n29693 ;
  assign n29695 = n29694 ^ n26644 ;
  assign n29696 = n29695 ^ n29613 ;
  assign n29697 = n29614 & ~n29696 ;
  assign n29698 = n29697 ^ n26888 ;
  assign n29699 = n29698 ^ n29611 ;
  assign n29700 = ~n29612 & ~n29699 ;
  assign n29701 = n29700 ^ n26640 ;
  assign n29702 = n29701 ^ n29609 ;
  assign n29703 = n29610 & n29702 ;
  assign n29704 = n29703 ^ n26635 ;
  assign n29885 = n29715 ^ n29704 ;
  assign n29886 = ~n29716 & n29885 ;
  assign n29887 = n29886 ^ n26628 ;
  assign n30061 = n29897 ^ n29887 ;
  assign n30062 = ~n29898 & n30061 ;
  assign n30063 = n30062 ^ n26623 ;
  assign n30060 = n30019 ^ n30016 ;
  assign n30064 = n30063 ^ n30060 ;
  assign n30065 = n30058 ^ n26619 ;
  assign n30066 = n30065 ^ n30058 ;
  assign n30067 = n30066 ^ n30060 ;
  assign n30068 = n30064 & ~n30067 ;
  assign n30069 = n30068 ^ n30065 ;
  assign n30070 = ~n30059 & ~n30069 ;
  assign n30071 = n30070 ^ n26907 ;
  assign n30008 = n29442 ^ n29398 ;
  assign n30031 = n30028 ^ n30008 ;
  assign n30029 = n30028 ^ n30022 ;
  assign n30030 = ~n30027 & ~n30029 ;
  assign n30032 = n30031 ^ n30030 ;
  assign n30004 = n28480 ^ n27989 ;
  assign n30005 = n29188 ^ n28480 ;
  assign n30006 = n30004 & n30005 ;
  assign n30007 = n30006 ^ n27989 ;
  assign n30056 = n30032 ^ n30007 ;
  assign n30057 = n30056 ^ n26613 ;
  assign n30133 = n30071 ^ n30057 ;
  assign n30134 = n30069 ^ n26907 ;
  assign n29717 = n29716 ^ n29704 ;
  assign n29718 = n29667 ^ n26664 ;
  assign n29719 = n29662 ^ n26662 ;
  assign n29720 = n29645 ^ n26608 ;
  assign n29721 = n29647 ^ n29634 ;
  assign n29722 = n29720 & n29721 ;
  assign n29723 = n29653 ^ n29650 ;
  assign n29724 = n29722 & n29723 ;
  assign n29725 = n29632 ^ n26669 ;
  assign n29726 = n29725 ^ n29655 ;
  assign n29727 = ~n29724 & n29726 ;
  assign n29728 = ~n29719 & ~n29727 ;
  assign n29729 = n29718 & n29728 ;
  assign n29730 = n29669 ^ n29629 ;
  assign n29731 = ~n29729 & n29730 ;
  assign n29732 = n29672 ^ n29627 ;
  assign n29733 = n29731 & n29732 ;
  assign n29734 = n29675 ^ n29625 ;
  assign n29735 = ~n29733 & ~n29734 ;
  assign n29736 = n29678 ^ n29623 ;
  assign n29737 = n29735 & ~n29736 ;
  assign n29738 = n29681 ^ n29621 ;
  assign n29739 = n29737 & n29738 ;
  assign n29740 = n29619 ^ n26658 ;
  assign n29741 = n29740 ^ n29684 ;
  assign n29742 = n29739 & ~n29741 ;
  assign n29743 = n29690 ^ n26654 ;
  assign n29744 = ~n29742 & n29743 ;
  assign n29745 = n29692 ^ n29616 ;
  assign n29746 = ~n29744 & ~n29745 ;
  assign n29747 = n29695 ^ n29614 ;
  assign n29748 = n29746 & n29747 ;
  assign n29749 = n29698 ^ n29612 ;
  assign n29750 = n29748 & ~n29749 ;
  assign n29751 = n29701 ^ n29610 ;
  assign n29752 = ~n29750 & n29751 ;
  assign n29884 = ~n29717 & ~n29752 ;
  assign n29899 = n29898 ^ n29887 ;
  assign n30135 = n29884 & ~n29899 ;
  assign n30136 = n30060 ^ n26619 ;
  assign n30137 = n30136 ^ n30063 ;
  assign n30138 = ~n30135 & n30137 ;
  assign n30139 = n30134 & n30138 ;
  assign n30140 = n30133 & n30139 ;
  assign n30009 = n30008 ^ n30007 ;
  assign n30033 = n30009 & n30032 ;
  assign n30034 = n30033 ^ n30008 ;
  assign n29998 = n29029 ^ n28558 ;
  assign n29929 = n29445 ^ n29396 ;
  assign n29999 = n29929 ^ n28043 ;
  assign n30000 = n29999 ^ n29029 ;
  assign n30001 = n30000 ^ n29929 ;
  assign n30002 = n29998 & ~n30001 ;
  assign n30003 = n30002 ^ n29999 ;
  assign n30075 = n30034 ^ n30003 ;
  assign n30141 = n30075 ^ n27145 ;
  assign n30072 = n30071 ^ n30056 ;
  assign n30073 = n30057 & n30072 ;
  assign n30074 = n30073 ^ n26613 ;
  assign n30142 = n30141 ^ n30074 ;
  assign n30143 = ~n30140 & n30142 ;
  assign n30076 = n30075 ^ n30074 ;
  assign n30035 = n27898 ^ n27350 ;
  assign n30036 = n29206 ^ n27898 ;
  assign n30037 = ~n30035 & ~n30036 ;
  assign n30038 = n30037 ^ n27350 ;
  assign n30040 = n30038 ^ n29929 ;
  assign n30039 = n30038 ^ n30034 ;
  assign n30041 = n30040 ^ n30039 ;
  assign n30042 = ~n30003 & ~n30041 ;
  assign n30043 = n30042 ^ n30040 ;
  assign n29923 = n29448 ^ n29394 ;
  assign n30077 = n30043 ^ n29923 ;
  assign n30078 = n30077 ^ n27145 ;
  assign n30079 = n30078 ^ n30074 ;
  assign n30080 = n30079 ^ n30077 ;
  assign n30081 = n30076 & ~n30080 ;
  assign n30082 = n30081 ^ n30078 ;
  assign n30144 = n30082 ^ n26600 ;
  assign n30145 = n30143 & n30144 ;
  assign n30053 = n29451 ^ n29392 ;
  assign n30044 = n27952 ^ n27352 ;
  assign n30045 = n29359 ^ n27952 ;
  assign n30046 = n30044 & ~n30045 ;
  assign n30047 = n30046 ^ n27352 ;
  assign n30049 = n30047 ^ n30038 ;
  assign n30048 = n30047 ^ n29923 ;
  assign n30050 = n30049 ^ n30048 ;
  assign n30051 = ~n30043 & n30050 ;
  assign n30052 = n30051 ^ n30049 ;
  assign n30054 = n30053 ^ n30052 ;
  assign n30084 = n30054 ^ n26600 ;
  assign n30083 = n30077 ^ n30054 ;
  assign n30085 = n30084 ^ n30083 ;
  assign n30086 = ~n30082 & ~n30085 ;
  assign n30087 = n30086 ^ n30084 ;
  assign n30132 = n30087 ^ n26787 ;
  assign n30203 = n30145 ^ n30132 ;
  assign n30207 = n30206 ^ n30203 ;
  assign n30209 = n27861 ^ n2886 ;
  assign n30210 = n30209 ^ n2642 ;
  assign n30211 = n30210 ^ n3206 ;
  assign n30208 = n30144 ^ n30143 ;
  assign n30212 = n30211 ^ n30208 ;
  assign n30216 = n30142 ^ n30140 ;
  assign n30213 = n27856 ^ n2879 ;
  assign n30214 = n30213 ^ n1379 ;
  assign n30215 = n30214 ^ n2540 ;
  assign n30217 = n30216 ^ n30215 ;
  assign n30220 = n30138 ^ n30134 ;
  assign n30231 = n30220 ^ n1352 ;
  assign n30218 = n30137 ^ n30135 ;
  assign n30219 = n30218 ^ n1168 ;
  assign n29900 = n29899 ^ n29884 ;
  assign n1032 = n995 ^ n956 ;
  assign n1033 = n1032 ^ n1029 ;
  assign n1037 = n1036 ^ n1033 ;
  assign n29901 = n29900 ^ n1037 ;
  assign n29753 = n29752 ^ n29717 ;
  assign n1008 = n944 ^ n891 ;
  assign n1018 = n1017 ^ n1008 ;
  assign n1022 = n1021 ^ n1018 ;
  assign n29754 = n29753 ^ n1022 ;
  assign n29755 = n29751 ^ n29750 ;
  assign n29756 = n29755 ^ n1636 ;
  assign n29757 = n29749 ^ n29748 ;
  assign n29877 = n29757 ^ n1636 ;
  assign n29758 = n29757 ^ n1627 ;
  assign n29759 = n29747 ^ n29746 ;
  assign n29760 = n29759 ^ n2978 ;
  assign n29764 = n29745 ^ n29744 ;
  assign n29765 = n29764 ^ n29763 ;
  assign n29766 = n29743 ^ n29742 ;
  assign n29767 = n29766 ^ n620 ;
  assign n29768 = n29741 ^ n29739 ;
  assign n29772 = n29771 ^ n29768 ;
  assign n29776 = n29738 ^ n29737 ;
  assign n29777 = n29776 ^ n29775 ;
  assign n29781 = n29736 ^ n29735 ;
  assign n29782 = n29781 ^ n29780 ;
  assign n29784 = n2439 ^ n1469 ;
  assign n29785 = n29784 ^ n24589 ;
  assign n29786 = n29785 ^ n19526 ;
  assign n29783 = n29734 ^ n29733 ;
  assign n29787 = n29786 ^ n29783 ;
  assign n29848 = n20768 ^ n2421 ;
  assign n29849 = n29848 ^ n24549 ;
  assign n29850 = n29849 ^ n19513 ;
  assign n29853 = n29850 ^ n29783 ;
  assign n29846 = n29732 ^ n29731 ;
  assign n29789 = n2411 ^ n2347 ;
  assign n29790 = n29789 ^ n24557 ;
  assign n29791 = n29790 ^ n2282 ;
  assign n29788 = n29730 ^ n29729 ;
  assign n29792 = n29791 ^ n29788 ;
  assign n29796 = n29728 ^ n29718 ;
  assign n29793 = n27436 ^ n2321 ;
  assign n29794 = n29793 ^ n2147 ;
  assign n29795 = n29794 ^ n19489 ;
  assign n29797 = n29796 ^ n29795 ;
  assign n29798 = n27469 ^ n2328 ;
  assign n29799 = n29798 ^ n24562 ;
  assign n29800 = n29799 ^ n2142 ;
  assign n29839 = n29800 ^ n29795 ;
  assign n29801 = n29727 ^ n29719 ;
  assign n29802 = n29801 ^ n29800 ;
  assign n29803 = n29726 ^ n29724 ;
  assign n2022 = n2021 ^ n1988 ;
  assign n2032 = n2031 ^ n2022 ;
  assign n2036 = n2035 ^ n2032 ;
  assign n29804 = n29803 ^ n2036 ;
  assign n29808 = n29723 ^ n29722 ;
  assign n29805 = n27448 ^ n20390 ;
  assign n29806 = n29805 ^ n1969 ;
  assign n29807 = n29806 ^ n2026 ;
  assign n29809 = n29808 ^ n29807 ;
  assign n1945 = n1938 ^ n1923 ;
  assign n1958 = n1957 ^ n1945 ;
  assign n1962 = n1961 ^ n1958 ;
  assign n29830 = n29807 ^ n1962 ;
  assign n29810 = n29721 ^ n29720 ;
  assign n29811 = n29810 ^ n1962 ;
  assign n29814 = n3240 ^ n1885 ;
  assign n29815 = n29814 ^ n3022 ;
  assign n29816 = n29815 ^ n3058 ;
  assign n29812 = n29638 ^ n26687 ;
  assign n29813 = n3015 & ~n29812 ;
  assign n29817 = n29816 ^ n29813 ;
  assign n29818 = n29639 ^ n26683 ;
  assign n29819 = n29818 ^ n29637 ;
  assign n29820 = n29819 ^ n29813 ;
  assign n29821 = n29817 & n29820 ;
  assign n29822 = n29821 ^ n29816 ;
  assign n3054 = n3032 ^ n1894 ;
  assign n3061 = n3060 ^ n3054 ;
  assign n3062 = n3061 ^ n1952 ;
  assign n29823 = n29822 ^ n3062 ;
  assign n29826 = n29822 ^ n29720 ;
  assign n29827 = ~n29823 & n29826 ;
  assign n29824 = n29720 ^ n1962 ;
  assign n29828 = n29827 ^ n29824 ;
  assign n29829 = ~n29811 & n29828 ;
  assign n29831 = n29830 ^ n29829 ;
  assign n29832 = ~n29809 & ~n29831 ;
  assign n29833 = n29832 ^ n29808 ;
  assign n29834 = n29833 ^ n2036 ;
  assign n29835 = ~n29804 & n29834 ;
  assign n29836 = n29835 ^ n29803 ;
  assign n29837 = n29836 ^ n29800 ;
  assign n29838 = ~n29802 & ~n29837 ;
  assign n29840 = n29839 ^ n29838 ;
  assign n29841 = ~n29797 & ~n29840 ;
  assign n29842 = n29841 ^ n29796 ;
  assign n29843 = n29842 ^ n29788 ;
  assign n29844 = ~n29792 & ~n29843 ;
  assign n29845 = n29844 ^ n29791 ;
  assign n29847 = n29846 ^ n29845 ;
  assign n29851 = n29850 ^ n29845 ;
  assign n29852 = ~n29847 & n29851 ;
  assign n29854 = n29853 ^ n29852 ;
  assign n29855 = ~n29787 & n29854 ;
  assign n29856 = n29855 ^ n29786 ;
  assign n29857 = n29856 ^ n29780 ;
  assign n29858 = n29782 & ~n29857 ;
  assign n29859 = n29858 ^ n29781 ;
  assign n29860 = n29859 ^ n29775 ;
  assign n29861 = ~n29777 & ~n29860 ;
  assign n29862 = n29861 ^ n29776 ;
  assign n29863 = n29862 ^ n29768 ;
  assign n29864 = n29772 & n29863 ;
  assign n29865 = n29864 ^ n29771 ;
  assign n29866 = n29865 ^ n620 ;
  assign n29867 = ~n29767 & n29866 ;
  assign n29868 = n29867 ^ n620 ;
  assign n29869 = n29868 ^ n29763 ;
  assign n29870 = ~n29765 & ~n29869 ;
  assign n29871 = n29870 ^ n29764 ;
  assign n29872 = n29871 ^ n2978 ;
  assign n29873 = ~n29760 & n29872 ;
  assign n29874 = n29873 ^ n29759 ;
  assign n29875 = n29874 ^ n1627 ;
  assign n29876 = n29758 & n29875 ;
  assign n29878 = n29877 ^ n29876 ;
  assign n29879 = ~n29756 & ~n29878 ;
  assign n29880 = n29879 ^ n29755 ;
  assign n29881 = n29880 ^ n1022 ;
  assign n29882 = ~n29754 & n29881 ;
  assign n29883 = n29882 ^ n29753 ;
  assign n30223 = n29883 ^ n1037 ;
  assign n30224 = n29901 & n30223 ;
  assign n30225 = n30224 ^ n29900 ;
  assign n30221 = n30220 ^ n1168 ;
  assign n30222 = n30221 ^ n30220 ;
  assign n30226 = n30225 ^ n30222 ;
  assign n30227 = ~n30219 & n30226 ;
  assign n30228 = n30227 ^ n30221 ;
  assign n1178 = n1142 ^ n1090 ;
  assign n1179 = n1178 ^ n1175 ;
  assign n1183 = n1182 ^ n1179 ;
  assign n30229 = n30220 ^ n1183 ;
  assign n30230 = n30228 & n30229 ;
  assign n30232 = n30231 ^ n30230 ;
  assign n30235 = n30215 ^ n1352 ;
  assign n30233 = n30139 ^ n30133 ;
  assign n30234 = n30233 ^ n30215 ;
  assign n30236 = n30235 ^ n30234 ;
  assign n30237 = n30232 & n30236 ;
  assign n30238 = n30237 ^ n30235 ;
  assign n30239 = n30217 & ~n30238 ;
  assign n30240 = n30239 ^ n30216 ;
  assign n30241 = n30240 ^ n30208 ;
  assign n30242 = ~n30212 & n30241 ;
  assign n30243 = n30242 ^ n30211 ;
  assign n30244 = n30243 ^ n30203 ;
  assign n30245 = n30207 & ~n30244 ;
  assign n30246 = n30245 ^ n30206 ;
  assign n30055 = n30054 ^ n26787 ;
  assign n30088 = ~n30055 & ~n30087 ;
  assign n30089 = n30088 ^ n26787 ;
  assign n30147 = n30089 ^ n26791 ;
  assign n30090 = n28754 ^ n27951 ;
  assign n30091 = n30053 ^ n30047 ;
  assign n30092 = n30052 & n30091 ;
  assign n30093 = n30092 ^ n30047 ;
  assign n30094 = n30093 ^ n27344 ;
  assign n30095 = n30094 ^ n28754 ;
  assign n30096 = n30095 ^ n30093 ;
  assign n30097 = n30090 & ~n30096 ;
  assign n30098 = n30097 ^ n30094 ;
  assign n29909 = n29454 ^ n29390 ;
  assign n30099 = n30098 ^ n29909 ;
  assign n30148 = n30147 ^ n30099 ;
  assign n30146 = ~n30132 & n30145 ;
  assign n30201 = n30148 ^ n30146 ;
  assign n30198 = n27522 ^ n20871 ;
  assign n30199 = n30198 ^ n24649 ;
  assign n30200 = n30199 ^ n3098 ;
  assign n30202 = n30201 ^ n30200 ;
  assign n30278 = n30246 ^ n30202 ;
  assign n30451 = n30282 ^ n30278 ;
  assign n30722 = n30451 ^ n27412 ;
  assign n30719 = n3179 ^ n2781 ;
  assign n30720 = n30719 ^ n1847 ;
  assign n30721 = n30720 ^ n20332 ;
  assign n31013 = n30722 ^ n30721 ;
  assign n29980 = n29720 ^ n3062 ;
  assign n29981 = n29980 ^ n29822 ;
  assign n31581 = n31013 ^ n29981 ;
  assign n31582 = n29981 ^ n29018 ;
  assign n31583 = ~n31581 & ~n31582 ;
  assign n31584 = n31583 ^ n29018 ;
  assign n31575 = n29469 ^ n2577 ;
  assign n31576 = n31575 ^ n3116 ;
  assign n31577 = n31576 ^ n20871 ;
  assign n31024 = n30240 ^ n30212 ;
  assign n31285 = n31024 ^ n29507 ;
  assign n30358 = n29859 ^ n29777 ;
  assign n30348 = n29856 ^ n29782 ;
  assign n29938 = n29890 ^ n29154 ;
  assign n29939 = n29854 ^ n29786 ;
  assign n29940 = n29939 ^ n28129 ;
  assign n29941 = n29940 ^ n29154 ;
  assign n29942 = n29941 ^ n29939 ;
  assign n29943 = ~n29938 & ~n29942 ;
  assign n29944 = n29943 ^ n29940 ;
  assign n30335 = n29850 ^ n29847 ;
  assign n30325 = n29842 ^ n29792 ;
  assign n29946 = n29593 ^ n28980 ;
  assign n29947 = n29593 ^ n28282 ;
  assign n29948 = n29946 & ~n29947 ;
  assign n29949 = n29948 ^ n28282 ;
  assign n29945 = n29840 ^ n29796 ;
  assign n29950 = n29949 ^ n29945 ;
  assign n29952 = n28986 ^ n28964 ;
  assign n29953 = n28986 ^ n28278 ;
  assign n29954 = ~n29952 & n29953 ;
  assign n29955 = n29954 ^ n28278 ;
  assign n29951 = n29836 ^ n29802 ;
  assign n29956 = n29955 ^ n29951 ;
  assign n29957 = n28992 ^ n28971 ;
  assign n29958 = n29833 ^ n29804 ;
  assign n29959 = n29958 ^ n28155 ;
  assign n29960 = n29959 ^ n28971 ;
  assign n29961 = n29960 ^ n29958 ;
  assign n29962 = n29957 & n29961 ;
  assign n29963 = n29962 ^ n29959 ;
  assign n29968 = n29831 ^ n29808 ;
  assign n29964 = n29070 ^ n28978 ;
  assign n29965 = n29070 ^ n28157 ;
  assign n29966 = ~n29964 & ~n29965 ;
  assign n29967 = n29966 ^ n28157 ;
  assign n29969 = n29968 ^ n29967 ;
  assign n29974 = n29828 ^ n29810 ;
  assign n29970 = n29108 ^ n28985 ;
  assign n29971 = n29108 ^ n28170 ;
  assign n29972 = ~n29970 & n29971 ;
  assign n29973 = n29972 ^ n28170 ;
  assign n29975 = n29974 ^ n29973 ;
  assign n29976 = n28998 ^ n27516 ;
  assign n29977 = n29577 ^ n28998 ;
  assign n29978 = n29976 & ~n29977 ;
  assign n29979 = n29978 ^ n27516 ;
  assign n29982 = n29981 ^ n29979 ;
  assign n29987 = n29819 ^ n29817 ;
  assign n30306 = n29987 ^ n29981 ;
  assign n29983 = n29004 ^ n28177 ;
  assign n29984 = n29567 ^ n29004 ;
  assign n29985 = n29983 & n29984 ;
  assign n29986 = n29985 ^ n28177 ;
  assign n29988 = n29987 ^ n29986 ;
  assign n29989 = n29555 ^ n29092 ;
  assign n29990 = n29812 ^ n3015 ;
  assign n29991 = n29990 ^ n28075 ;
  assign n29992 = n29991 ^ n29555 ;
  assign n29993 = n29992 ^ n29990 ;
  assign n29994 = ~n29989 & n29993 ;
  assign n29995 = n29994 ^ n29991 ;
  assign n30259 = n28945 ^ n28082 ;
  assign n30260 = n28997 ^ n28945 ;
  assign n30261 = ~n30259 & ~n30260 ;
  assign n30262 = n30261 ^ n28082 ;
  assign n29918 = n29457 ^ n29388 ;
  assign n30105 = n29918 ^ n29909 ;
  assign n30104 = n30093 ^ n29918 ;
  assign n30106 = n30105 ^ n30104 ;
  assign n30107 = ~n30098 & ~n30106 ;
  assign n30108 = n30107 ^ n30105 ;
  assign n30115 = n29460 ^ n29381 ;
  assign n30117 = n30115 ^ n29918 ;
  assign n30109 = n28004 ^ n27342 ;
  assign n30110 = n28757 ^ n28004 ;
  assign n30111 = ~n30109 & n30110 ;
  assign n30112 = n30111 ^ n27342 ;
  assign n30116 = n30115 ^ n30112 ;
  assign n30118 = n30117 ^ n30116 ;
  assign n30119 = n30108 & ~n30118 ;
  assign n30120 = n30119 ^ n30116 ;
  assign n30157 = n28217 ^ n26605 ;
  assign n30158 = n28744 ^ n28217 ;
  assign n30159 = ~n30157 & ~n30158 ;
  assign n30160 = n30159 ^ n26605 ;
  assign n30162 = n30160 ^ n30115 ;
  assign n30121 = n28766 ^ n28055 ;
  assign n30122 = n28766 ^ n27338 ;
  assign n30123 = n30121 & ~n30122 ;
  assign n30124 = n30123 ^ n27338 ;
  assign n30161 = n30160 ^ n30124 ;
  assign n30163 = n30162 ^ n30161 ;
  assign n30164 = n30120 & ~n30163 ;
  assign n30165 = n30164 ^ n30162 ;
  assign n29904 = n29464 ^ n29463 ;
  assign n30166 = n30165 ^ n29904 ;
  assign n30167 = n30166 ^ n26693 ;
  assign n30113 = n30112 ^ n30108 ;
  assign n30100 = n30099 ^ n30089 ;
  assign n30101 = n30099 ^ n26791 ;
  assign n30102 = ~n30100 & n30101 ;
  assign n30103 = n30102 ^ n26791 ;
  assign n30114 = n30113 ^ n30103 ;
  assign n30125 = n30124 ^ n30120 ;
  assign n30126 = n30125 ^ n26799 ;
  assign n30127 = n30126 ^ n30125 ;
  assign n30128 = n30127 ^ n30103 ;
  assign n30129 = n30114 & ~n30128 ;
  assign n30130 = n30129 ^ n30126 ;
  assign n30154 = n30125 ^ n26777 ;
  assign n30155 = ~n30130 & n30154 ;
  assign n30156 = n30155 ^ n26777 ;
  assign n30168 = n30167 ^ n30156 ;
  assign n30131 = n30130 ^ n26777 ;
  assign n30149 = n30146 & ~n30148 ;
  assign n30150 = n30113 ^ n26799 ;
  assign n30151 = n30150 ^ n30103 ;
  assign n30152 = ~n30149 & n30151 ;
  assign n30153 = ~n30131 & n30152 ;
  assign n30188 = n30168 ^ n30153 ;
  assign n2714 = n2701 ^ n2671 ;
  assign n2718 = n2717 ^ n2714 ;
  assign n2719 = n2718 ^ n2713 ;
  assign n30189 = n30188 ^ n2719 ;
  assign n30191 = n27927 ^ n2611 ;
  assign n30192 = n30191 ^ n24677 ;
  assign n30193 = n30192 ^ n1838 ;
  assign n30190 = n30152 ^ n30131 ;
  assign n30194 = n30193 ^ n30190 ;
  assign n30196 = n30151 ^ n30149 ;
  assign n3123 = n3122 ^ n2605 ;
  assign n3124 = n3123 ^ n3104 ;
  assign n3128 = n3127 ^ n3124 ;
  assign n30197 = n30196 ^ n3128 ;
  assign n30247 = n30246 ^ n30200 ;
  assign n30248 = n30202 & ~n30247 ;
  assign n30249 = n30248 ^ n30201 ;
  assign n30250 = n30249 ^ n30196 ;
  assign n30251 = ~n30197 & n30250 ;
  assign n30252 = n30251 ^ n3128 ;
  assign n30195 = n30193 ^ n30188 ;
  assign n30253 = n30252 ^ n30195 ;
  assign n30254 = n30253 ^ n30188 ;
  assign n30255 = ~n30194 & n30254 ;
  assign n30256 = n30255 ^ n30195 ;
  assign n30257 = n30189 & ~n30256 ;
  assign n30180 = n30160 ^ n29904 ;
  assign n30181 = ~n30165 & ~n30180 ;
  assign n30178 = n30160 ^ n27373 ;
  assign n30177 = n29474 ^ n29471 ;
  assign n30179 = n30178 ^ n30177 ;
  assign n30182 = n30181 ^ n30179 ;
  assign n30176 = n26693 ^ n26691 ;
  assign n30183 = n30182 ^ n30176 ;
  assign n30175 = n2731 ^ n2719 ;
  assign n30184 = n30183 ^ n30175 ;
  assign n30173 = n30166 ^ n30156 ;
  assign n30174 = ~n30167 & ~n30173 ;
  assign n30185 = n30184 ^ n30174 ;
  assign n30170 = n28738 ^ n28226 ;
  assign n30171 = n28226 ^ n27373 ;
  assign n30172 = ~n30170 & n30171 ;
  assign n30186 = n30185 ^ n30172 ;
  assign n30169 = n30153 & n30168 ;
  assign n30187 = n30186 ^ n30169 ;
  assign n30258 = n30257 ^ n30187 ;
  assign n30263 = n30262 ^ n30258 ;
  assign n30265 = n30256 ^ n2719 ;
  assign n30298 = n30265 ^ n30258 ;
  assign n30264 = n29009 ^ n28844 ;
  assign n30266 = n30265 ^ n28090 ;
  assign n30267 = n30266 ^ n29009 ;
  assign n30268 = n30267 ^ n30265 ;
  assign n30269 = n30264 & ~n30268 ;
  assign n30270 = n30269 ^ n30266 ;
  assign n30272 = n28100 ^ n28069 ;
  assign n30273 = n29018 ^ n28069 ;
  assign n30274 = ~n30272 & n30273 ;
  assign n30275 = n30274 ^ n28100 ;
  assign n30271 = n30252 ^ n30194 ;
  assign n30276 = n30275 ^ n30271 ;
  assign n30283 = n30278 & n30282 ;
  assign n30277 = n30249 ^ n30197 ;
  assign n30284 = n30283 ^ n30277 ;
  assign n30285 = n29012 ^ n28783 ;
  assign n30286 = n30283 ^ n28201 ;
  assign n30287 = n30286 ^ n29012 ;
  assign n30288 = n30287 ^ n30283 ;
  assign n30289 = n30285 & ~n30288 ;
  assign n30290 = n30289 ^ n30286 ;
  assign n30291 = ~n30284 & ~n30290 ;
  assign n30292 = n30291 ^ n30283 ;
  assign n30293 = n30292 ^ n30271 ;
  assign n30294 = n30276 & n30293 ;
  assign n30295 = n30294 ^ n30275 ;
  assign n30296 = n30295 ^ n30265 ;
  assign n30297 = n30270 & ~n30296 ;
  assign n30299 = n30298 ^ n30297 ;
  assign n30300 = ~n30263 & ~n30299 ;
  assign n30301 = n30300 ^ n30262 ;
  assign n30302 = n30301 ^ n29990 ;
  assign n30303 = n29995 & n30302 ;
  assign n29996 = n29990 ^ n29987 ;
  assign n30304 = n30303 ^ n29996 ;
  assign n30305 = n29988 & n30304 ;
  assign n30307 = n30306 ^ n30305 ;
  assign n30308 = ~n29982 & ~n30307 ;
  assign n30309 = n30308 ^ n29981 ;
  assign n30310 = n30309 ^ n29973 ;
  assign n30311 = n29975 & n30310 ;
  assign n30312 = n30311 ^ n29974 ;
  assign n30313 = n30312 ^ n29967 ;
  assign n30314 = ~n29969 & n30313 ;
  assign n30315 = n30314 ^ n29968 ;
  assign n30316 = n30315 ^ n29958 ;
  assign n30317 = n29963 & ~n30316 ;
  assign n30318 = n30317 ^ n29958 ;
  assign n30319 = n30318 ^ n29951 ;
  assign n30320 = ~n29956 & ~n30319 ;
  assign n30321 = n30320 ^ n29955 ;
  assign n30322 = n30321 ^ n29945 ;
  assign n30323 = ~n29950 & ~n30322 ;
  assign n30324 = n30323 ^ n29949 ;
  assign n30326 = n30325 ^ n30324 ;
  assign n30327 = n29603 ^ n28972 ;
  assign n30328 = n30325 ^ n28142 ;
  assign n30329 = n30328 ^ n28972 ;
  assign n30330 = n30329 ^ n30325 ;
  assign n30331 = n30327 & n30330 ;
  assign n30332 = n30331 ^ n30328 ;
  assign n30333 = n30326 & ~n30332 ;
  assign n30334 = n30333 ^ n30325 ;
  assign n30336 = n30335 ^ n30334 ;
  assign n30337 = n29709 ^ n28965 ;
  assign n30338 = n30334 ^ n28135 ;
  assign n30339 = n30338 ^ n28965 ;
  assign n30340 = n30339 ^ n30334 ;
  assign n30341 = n30337 & ~n30340 ;
  assign n30342 = n30341 ^ n30338 ;
  assign n30343 = n30336 & ~n30342 ;
  assign n30344 = n30343 ^ n30335 ;
  assign n30345 = n30344 ^ n29939 ;
  assign n30346 = n29944 & ~n30345 ;
  assign n30347 = n30346 ^ n29939 ;
  assign n30349 = n30348 ^ n30347 ;
  assign n30350 = n30015 ^ n29159 ;
  assign n30351 = n30347 ^ n28310 ;
  assign n30352 = n30351 ^ n29159 ;
  assign n30353 = n30352 ^ n30347 ;
  assign n30354 = ~n30350 & ~n30353 ;
  assign n30355 = n30354 ^ n30351 ;
  assign n30356 = ~n30349 & ~n30355 ;
  assign n30357 = n30356 ^ n30348 ;
  assign n30359 = n30358 ^ n30357 ;
  assign n30360 = n30028 ^ n29163 ;
  assign n30361 = n30358 ^ n28316 ;
  assign n30362 = n30361 ^ n30028 ;
  assign n30363 = n30362 ^ n30358 ;
  assign n30364 = n30360 & n30363 ;
  assign n30365 = n30364 ^ n30361 ;
  assign n30366 = ~n30359 & n30365 ;
  assign n30367 = n30366 ^ n30358 ;
  assign n29937 = n29862 ^ n29772 ;
  assign n30368 = n30367 ^ n29937 ;
  assign n30369 = n30008 ^ n29042 ;
  assign n30370 = n29937 ^ n28126 ;
  assign n30371 = n30370 ^ n29042 ;
  assign n30372 = n30371 ^ n29937 ;
  assign n30373 = n30369 & ~n30372 ;
  assign n30374 = n30373 ^ n30370 ;
  assign n30375 = n30368 & ~n30374 ;
  assign n30376 = n30375 ^ n30367 ;
  assign n29930 = n29929 ^ n29039 ;
  assign n29931 = n29865 ^ n29767 ;
  assign n29932 = n29931 ^ n28112 ;
  assign n29933 = n29932 ^ n29929 ;
  assign n29934 = n29933 ^ n29931 ;
  assign n29935 = ~n29930 & n29934 ;
  assign n29936 = n29935 ^ n29932 ;
  assign n30527 = n30376 ^ n29936 ;
  assign n30431 = n30374 ^ n30367 ;
  assign n30432 = n30431 ^ n27750 ;
  assign n30514 = n30355 ^ n30348 ;
  assign n30434 = n30344 ^ n29944 ;
  assign n30435 = n30434 ^ n27525 ;
  assign n30505 = n30342 ^ n30335 ;
  assign n30437 = n30321 ^ n29950 ;
  assign n30438 = n30437 ^ n27536 ;
  assign n30440 = n30315 ^ n29963 ;
  assign n30441 = n30440 ^ n27547 ;
  assign n30443 = n30309 ^ n29975 ;
  assign n30444 = n30443 ^ n27554 ;
  assign n30445 = n30307 ^ n29979 ;
  assign n30446 = n30445 ^ n27558 ;
  assign n30447 = n30304 ^ n29986 ;
  assign n30448 = n30447 ^ n27562 ;
  assign n30471 = n30301 ^ n29995 ;
  assign n30458 = n30292 ^ n30276 ;
  assign n30453 = n30290 ^ n30277 ;
  assign n30452 = n27412 & n30451 ;
  assign n30454 = n30453 ^ n30452 ;
  assign n30455 = n30453 ^ n27485 ;
  assign n30456 = ~n30454 & ~n30455 ;
  assign n30457 = n30456 ^ n27485 ;
  assign n30459 = n30458 ^ n30457 ;
  assign n30460 = n30458 ^ n27502 ;
  assign n30461 = n30459 & ~n30460 ;
  assign n30462 = n30461 ^ n27502 ;
  assign n30450 = n30295 ^ n30270 ;
  assign n30463 = n30462 ^ n30450 ;
  assign n30464 = n30462 ^ n27576 ;
  assign n30465 = ~n30463 & n30464 ;
  assign n30466 = n30465 ^ n27576 ;
  assign n30449 = n30299 ^ n30262 ;
  assign n30467 = n30466 ^ n30449 ;
  assign n30468 = n30466 ^ n27577 ;
  assign n30469 = ~n30467 & ~n30468 ;
  assign n30470 = n30469 ^ n27577 ;
  assign n30472 = n30471 ^ n30470 ;
  assign n30473 = n30471 ^ n27567 ;
  assign n30474 = n30472 & ~n30473 ;
  assign n30475 = n30474 ^ n27567 ;
  assign n30476 = n30475 ^ n30447 ;
  assign n30477 = ~n30448 & n30476 ;
  assign n30478 = n30477 ^ n27562 ;
  assign n30479 = n30478 ^ n30445 ;
  assign n30480 = ~n30446 & ~n30479 ;
  assign n30481 = n30480 ^ n27558 ;
  assign n30482 = n30481 ^ n30443 ;
  assign n30483 = n30444 & n30482 ;
  assign n30484 = n30483 ^ n27554 ;
  assign n30442 = n30312 ^ n29969 ;
  assign n30485 = n30484 ^ n30442 ;
  assign n30486 = n30440 ^ n27517 ;
  assign n30487 = n30486 ^ n30440 ;
  assign n30488 = n30487 ^ n30442 ;
  assign n30489 = ~n30485 & n30488 ;
  assign n30490 = n30489 ^ n30486 ;
  assign n30491 = n30441 & n30490 ;
  assign n30492 = n30491 ^ n27547 ;
  assign n30439 = n30318 ^ n29956 ;
  assign n30493 = n30492 ^ n30439 ;
  assign n30494 = n30437 ^ n27543 ;
  assign n30495 = n30494 ^ n30437 ;
  assign n30496 = n30495 ^ n30439 ;
  assign n30497 = ~n30493 & n30496 ;
  assign n30498 = n30497 ^ n30494 ;
  assign n30499 = ~n30438 & n30498 ;
  assign n30500 = n30499 ^ n27536 ;
  assign n30436 = n30332 ^ n30324 ;
  assign n30501 = n30500 ^ n30436 ;
  assign n30502 = n30500 ^ n27534 ;
  assign n30503 = ~n30501 & n30502 ;
  assign n30504 = n30503 ^ n27534 ;
  assign n30506 = n30505 ^ n30504 ;
  assign n30507 = n30434 ^ n27527 ;
  assign n30508 = n30507 ^ n30434 ;
  assign n30509 = n30508 ^ n30504 ;
  assign n30510 = n30506 & ~n30509 ;
  assign n30511 = n30510 ^ n30507 ;
  assign n30512 = ~n30435 & ~n30511 ;
  assign n30513 = n30512 ^ n27525 ;
  assign n30515 = n30514 ^ n30513 ;
  assign n30516 = n30514 ^ n27621 ;
  assign n30517 = n30515 & ~n30516 ;
  assign n30518 = n30517 ^ n27621 ;
  assign n30433 = n30365 ^ n30357 ;
  assign n30519 = n30518 ^ n30433 ;
  assign n30520 = n30518 ^ n27700 ;
  assign n30521 = n30519 & n30520 ;
  assign n30522 = n30521 ^ n27700 ;
  assign n30523 = n30522 ^ n30431 ;
  assign n30524 = ~n30432 & ~n30523 ;
  assign n30525 = n30524 ^ n27750 ;
  assign n30526 = n30525 ^ n27766 ;
  assign n30617 = n30527 ^ n30526 ;
  assign n30575 = n30522 ^ n30432 ;
  assign n30576 = n30433 ^ n27700 ;
  assign n30577 = n30576 ^ n30518 ;
  assign n30578 = n30516 ^ n30513 ;
  assign n30579 = n30511 ^ n27525 ;
  assign n30580 = n30439 ^ n27543 ;
  assign n30581 = n30580 ^ n30492 ;
  assign n30582 = n30490 ^ n27547 ;
  assign n30583 = n30470 ^ n27567 ;
  assign n30584 = n30583 ^ n30471 ;
  assign n30585 = n30449 ^ n27577 ;
  assign n30586 = n30585 ^ n30466 ;
  assign n30587 = n30457 ^ n27502 ;
  assign n30588 = n30587 ^ n30458 ;
  assign n30589 = n30464 ^ n30450 ;
  assign n30590 = ~n30588 & n30589 ;
  assign n30591 = ~n30586 & n30590 ;
  assign n30592 = ~n30584 & ~n30591 ;
  assign n30593 = n30475 ^ n30448 ;
  assign n30594 = ~n30592 & n30593 ;
  assign n30595 = n30478 ^ n30446 ;
  assign n30596 = n30594 & n30595 ;
  assign n30597 = n30481 ^ n27554 ;
  assign n30598 = n30597 ^ n30443 ;
  assign n30599 = ~n30596 & ~n30598 ;
  assign n30600 = n30442 ^ n27517 ;
  assign n30601 = n30600 ^ n30484 ;
  assign n30602 = n30599 & n30601 ;
  assign n30603 = ~n30582 & ~n30602 ;
  assign n30604 = n30581 & n30603 ;
  assign n30605 = n30498 ^ n27536 ;
  assign n30606 = n30604 & ~n30605 ;
  assign n30607 = n30436 ^ n27534 ;
  assign n30608 = n30607 ^ n30500 ;
  assign n30609 = n30606 & n30608 ;
  assign n30610 = n30505 ^ n27527 ;
  assign n30611 = n30610 ^ n30504 ;
  assign n30612 = ~n30609 & ~n30611 ;
  assign n30613 = n30579 & ~n30612 ;
  assign n30614 = ~n30578 & n30613 ;
  assign n30615 = ~n30577 & n30614 ;
  assign n30616 = n30575 & ~n30615 ;
  assign n30654 = n30617 ^ n30616 ;
  assign n1683 = n1666 ^ n1112 ;
  assign n1687 = n1686 ^ n1683 ;
  assign n1688 = n1687 ^ n915 ;
  assign n30655 = n30654 ^ n1688 ;
  assign n777 = n776 ^ n743 ;
  assign n787 = n786 ^ n777 ;
  assign n791 = n790 ^ n787 ;
  assign n30783 = n30654 ^ n791 ;
  assign n30656 = n30615 ^ n30575 ;
  assign n30657 = n30656 ^ n791 ;
  assign n30658 = n30614 ^ n30577 ;
  assign n2990 = n2983 ^ n1644 ;
  assign n2991 = n2990 ^ n721 ;
  assign n2992 = n2991 ^ n781 ;
  assign n30659 = n30658 ^ n2992 ;
  assign n30660 = n30613 ^ n30578 ;
  assign n30777 = n30660 ^ n2992 ;
  assign n30661 = n30660 ^ n714 ;
  assign n30774 = n30664 ^ n30660 ;
  assign n30665 = n30612 ^ n30579 ;
  assign n30666 = n30665 ^ n30664 ;
  assign n30767 = n30611 ^ n30609 ;
  assign n30667 = n30608 ^ n30606 ;
  assign n30671 = n30670 ^ n30667 ;
  assign n30675 = n30605 ^ n30604 ;
  assign n30672 = n28679 ^ n1494 ;
  assign n30673 = n30672 ^ n24981 ;
  assign n30674 = n30673 ^ n2933 ;
  assign n30676 = n30675 ^ n30674 ;
  assign n30680 = n30603 ^ n30581 ;
  assign n30677 = n28636 ^ n21159 ;
  assign n30678 = n30677 ^ n2921 ;
  assign n30679 = n30678 ^ n19827 ;
  assign n30681 = n30680 ^ n30679 ;
  assign n30682 = n30602 ^ n30582 ;
  assign n30686 = n30685 ^ n30682 ;
  assign n30689 = n30601 ^ n30599 ;
  assign n2364 = n2363 ^ n2297 ;
  assign n2374 = n2373 ^ n2364 ;
  assign n2378 = n2377 ^ n2374 ;
  assign n30690 = n30689 ^ n2378 ;
  assign n30693 = n28641 ^ n21174 ;
  assign n30694 = n30693 ^ n2233 ;
  assign n30695 = n30694 ^ n2368 ;
  assign n30752 = n30695 ^ n30689 ;
  assign n30691 = n30595 ^ n30594 ;
  assign n2218 = n2211 ^ n2160 ;
  assign n2225 = n2224 ^ n2218 ;
  assign n2229 = n2228 ^ n2225 ;
  assign n30692 = n30691 ^ n2229 ;
  assign n30698 = n30593 ^ n30592 ;
  assign n2126 = n2095 ^ n2071 ;
  assign n2127 = n2126 ^ n2123 ;
  assign n2131 = n2130 ^ n2127 ;
  assign n30699 = n30698 ^ n2131 ;
  assign n2099 = n2086 ^ n2056 ;
  assign n2112 = n2111 ^ n2099 ;
  assign n2116 = n2115 ^ n2112 ;
  assign n30742 = n30698 ^ n2116 ;
  assign n30700 = n30591 ^ n30584 ;
  assign n30701 = n30700 ^ n2116 ;
  assign n30703 = n28012 ^ n2006 ;
  assign n30704 = n30703 ^ n25009 ;
  assign n30705 = n30704 ^ n2108 ;
  assign n30702 = n30590 ^ n30586 ;
  assign n30706 = n30705 ^ n30702 ;
  assign n30710 = n30589 ^ n30588 ;
  assign n30707 = n3088 ^ n1997 ;
  assign n30708 = n30707 ^ n25018 ;
  assign n30709 = n30708 ^ n19844 ;
  assign n30711 = n30710 ^ n30709 ;
  assign n30712 = n21195 ^ n3076 ;
  assign n30713 = n30712 ^ n24700 ;
  assign n30714 = n30713 ^ n19851 ;
  assign n30715 = n30714 ^ n30588 ;
  assign n30723 = n30721 & n30722 ;
  assign n30716 = n28017 ^ n3044 ;
  assign n30717 = n30716 ^ n24696 ;
  assign n30718 = n30717 ^ n1793 ;
  assign n30724 = n30723 ^ n30718 ;
  assign n30726 = n30452 ^ n27485 ;
  assign n30727 = n30726 ^ n30453 ;
  assign n30725 = n30718 ^ n30714 ;
  assign n30728 = n30727 ^ n30725 ;
  assign n30729 = n30728 ^ n30714 ;
  assign n30730 = n30724 & ~n30729 ;
  assign n30731 = n30730 ^ n30725 ;
  assign n30732 = ~n30715 & n30731 ;
  assign n30733 = n30732 ^ n30714 ;
  assign n30734 = n30733 ^ n30709 ;
  assign n30735 = n30711 & ~n30734 ;
  assign n30736 = n30735 ^ n30710 ;
  assign n30737 = n30736 ^ n30702 ;
  assign n30738 = n30706 & ~n30737 ;
  assign n30739 = n30738 ^ n30705 ;
  assign n30740 = n30739 ^ n2116 ;
  assign n30741 = n30701 & n30740 ;
  assign n30743 = n30742 ^ n30741 ;
  assign n30744 = n30699 & n30743 ;
  assign n30745 = n30744 ^ n30698 ;
  assign n30746 = n30745 ^ n2229 ;
  assign n30747 = ~n30692 & n30746 ;
  assign n30696 = n30695 ^ n2229 ;
  assign n30748 = n30747 ^ n30696 ;
  assign n30749 = n30598 ^ n30596 ;
  assign n30750 = n30749 ^ n30695 ;
  assign n30751 = n30748 & n30750 ;
  assign n30753 = n30752 ^ n30751 ;
  assign n30754 = n30690 & n30753 ;
  assign n30755 = n30754 ^ n30689 ;
  assign n30756 = n30755 ^ n30685 ;
  assign n30757 = ~n30686 & n30756 ;
  assign n30687 = n30685 ^ n30679 ;
  assign n30758 = n30757 ^ n30687 ;
  assign n30759 = ~n30681 & ~n30758 ;
  assign n30760 = n30759 ^ n30680 ;
  assign n30761 = n30760 ^ n30674 ;
  assign n30762 = n30676 & n30761 ;
  assign n30763 = n30762 ^ n30675 ;
  assign n30764 = n30763 ^ n30667 ;
  assign n30765 = ~n30671 & n30764 ;
  assign n30766 = n30765 ^ n30670 ;
  assign n30768 = n30767 ^ n30766 ;
  assign n30769 = n30766 ^ n1535 ;
  assign n30770 = ~n30768 & n30769 ;
  assign n30771 = n30770 ^ n1535 ;
  assign n30772 = n30771 ^ n30664 ;
  assign n30773 = n30666 & n30772 ;
  assign n30775 = n30774 ^ n30773 ;
  assign n30776 = n30661 & n30775 ;
  assign n30778 = n30777 ^ n30776 ;
  assign n30779 = n30659 & ~n30778 ;
  assign n30780 = n30779 ^ n30658 ;
  assign n30781 = n30780 ^ n791 ;
  assign n30782 = ~n30657 & n30781 ;
  assign n30784 = n30783 ^ n30782 ;
  assign n30785 = ~n30655 & ~n30784 ;
  assign n30786 = n30785 ^ n30654 ;
  assign n30528 = n30527 ^ n30525 ;
  assign n30529 = n30526 & ~n30528 ;
  assign n30530 = n30529 ^ n27766 ;
  assign n29927 = n29868 ^ n29765 ;
  assign n30379 = n29931 ^ n29927 ;
  assign n30377 = n30376 ^ n29931 ;
  assign n30378 = ~n29936 & n30377 ;
  assign n30380 = n30379 ^ n30378 ;
  assign n29922 = n29178 ^ n28329 ;
  assign n29924 = n29923 ^ n29178 ;
  assign n29925 = n29922 & ~n29924 ;
  assign n29926 = n29925 ^ n28329 ;
  assign n30429 = n30380 ^ n29926 ;
  assign n30430 = n30429 ^ n27892 ;
  assign n30619 = n30530 ^ n30430 ;
  assign n30618 = ~n30616 & ~n30617 ;
  assign n30652 = n30619 ^ n30618 ;
  assign n1692 = n1673 ^ n1098 ;
  assign n1693 = n1692 ^ n928 ;
  assign n1694 = n1693 ^ n1295 ;
  assign n30653 = n30652 ^ n1694 ;
  assign n31286 = n30786 ^ n30653 ;
  assign n31287 = n31286 ^ n28754 ;
  assign n31288 = n31287 ^ n31024 ;
  assign n31289 = n31288 ^ n31286 ;
  assign n31290 = n31285 & ~n31289 ;
  assign n31291 = n31290 ^ n31287 ;
  assign n30850 = n30233 ^ n30232 ;
  assign n30909 = n30850 ^ n29904 ;
  assign n30910 = n30780 ^ n30657 ;
  assign n30911 = n30910 ^ n29206 ;
  assign n30912 = n30911 ^ n30850 ;
  assign n30913 = n30912 ^ n30910 ;
  assign n30914 = ~n30909 & n30913 ;
  assign n30915 = n30914 ^ n30911 ;
  assign n30926 = n30778 ^ n30658 ;
  assign n30922 = n30115 ^ n29029 ;
  assign n30569 = n30228 ^ n1183 ;
  assign n30923 = n30569 ^ n30115 ;
  assign n30924 = n30922 & ~n30923 ;
  assign n30925 = n30924 ^ n29029 ;
  assign n30927 = n30926 ^ n30925 ;
  assign n30929 = n30775 ^ n714 ;
  assign n31157 = n30929 ^ n30925 ;
  assign n30417 = n30225 ^ n30219 ;
  assign n30928 = n30417 ^ n29918 ;
  assign n30930 = n30929 ^ n29188 ;
  assign n30931 = n30930 ^ n30417 ;
  assign n30932 = n30931 ^ n30929 ;
  assign n30933 = ~n30928 & ~n30932 ;
  assign n30934 = n30933 ^ n30930 ;
  assign n29902 = n29901 ^ n29883 ;
  assign n30936 = n29909 ^ n29902 ;
  assign n30937 = n29909 ^ n29178 ;
  assign n30938 = n30936 & ~n30937 ;
  assign n30939 = n30938 ^ n29178 ;
  assign n30935 = n30771 ^ n30666 ;
  assign n30940 = n30939 ^ n30935 ;
  assign n30945 = n30768 ^ n1535 ;
  assign n30398 = n29880 ^ n29754 ;
  assign n30941 = n30398 ^ n30053 ;
  assign n30942 = n30053 ^ n29039 ;
  assign n30943 = n30941 & ~n30942 ;
  assign n30944 = n30943 ^ n29039 ;
  assign n30946 = n30945 ^ n30944 ;
  assign n30951 = n30763 ^ n30671 ;
  assign n31148 = n30951 ^ n30945 ;
  assign n30399 = n29878 ^ n29755 ;
  assign n30947 = n30399 ^ n29923 ;
  assign n30948 = n29923 ^ n29042 ;
  assign n30949 = ~n30947 & ~n30948 ;
  assign n30950 = n30949 ^ n29042 ;
  assign n30952 = n30951 ^ n30950 ;
  assign n29911 = n29874 ^ n29758 ;
  assign n30953 = n29929 ^ n29911 ;
  assign n30954 = n30760 ^ n30676 ;
  assign n30955 = n30954 ^ n29163 ;
  assign n30956 = n30955 ^ n29911 ;
  assign n30957 = n30956 ^ n30954 ;
  assign n30958 = n30953 & ~n30957 ;
  assign n30959 = n30958 ^ n30955 ;
  assign n31143 = n30954 ^ n30951 ;
  assign n30965 = n30755 ^ n30686 ;
  assign n30961 = n30028 ^ n29927 ;
  assign n30962 = n30028 ^ n29154 ;
  assign n30963 = ~n30961 & ~n30962 ;
  assign n30964 = n30963 ^ n29154 ;
  assign n30966 = n30965 ^ n30964 ;
  assign n30967 = n29931 ^ n28965 ;
  assign n30968 = n30753 ^ n2378 ;
  assign n30969 = n30968 ^ n30015 ;
  assign n30970 = n30969 ^ n29931 ;
  assign n30971 = n30970 ^ n30968 ;
  assign n30972 = ~n30967 & ~n30971 ;
  assign n30973 = n30972 ^ n30969 ;
  assign n31128 = n30968 ^ n30965 ;
  assign n30979 = n30745 ^ n30692 ;
  assign n30975 = n29709 ^ n28980 ;
  assign n30976 = n30358 ^ n28980 ;
  assign n30977 = n30975 & n30976 ;
  assign n30978 = n30977 ^ n29709 ;
  assign n30980 = n30979 ^ n30978 ;
  assign n30982 = n30743 ^ n2131 ;
  assign n31115 = n30982 ^ n30979 ;
  assign n30981 = n30348 ^ n29603 ;
  assign n30983 = n30982 ^ n28986 ;
  assign n30984 = n30983 ^ n30348 ;
  assign n30985 = n30984 ^ n30982 ;
  assign n30986 = ~n30981 & ~n30985 ;
  assign n30987 = n30986 ^ n30983 ;
  assign n30989 = n29593 ^ n28992 ;
  assign n30990 = n29939 ^ n29593 ;
  assign n30991 = n30989 & ~n30990 ;
  assign n30992 = n30991 ^ n28992 ;
  assign n30988 = n30739 ^ n30701 ;
  assign n30993 = n30992 ^ n30988 ;
  assign n30995 = n30736 ^ n30706 ;
  assign n31109 = n30995 ^ n30992 ;
  assign n30994 = n30335 ^ n28964 ;
  assign n30996 = n30995 ^ n29070 ;
  assign n30997 = n30996 ^ n30335 ;
  assign n30998 = n30997 ^ n30995 ;
  assign n30999 = n30994 & ~n30998 ;
  assign n31000 = n30999 ^ n30996 ;
  assign n31002 = n29945 ^ n28978 ;
  assign n31003 = n28998 ^ n28978 ;
  assign n31004 = ~n31002 & n31003 ;
  assign n31005 = n31004 ^ n28998 ;
  assign n30907 = n30731 ^ n30588 ;
  assign n31006 = n31005 ^ n30907 ;
  assign n31011 = n30727 ^ n30724 ;
  assign n31007 = n29951 ^ n28985 ;
  assign n31008 = n29004 ^ n28985 ;
  assign n31009 = n31007 & n31008 ;
  assign n31010 = n31009 ^ n29004 ;
  assign n31012 = n31011 ^ n31010 ;
  assign n31014 = n29577 ^ n29092 ;
  assign n31015 = n29958 ^ n29577 ;
  assign n31016 = n31014 & n31015 ;
  assign n31017 = n31016 ^ n29092 ;
  assign n31091 = n31017 ^ n31011 ;
  assign n31018 = n31017 ^ n31013 ;
  assign n31030 = n28217 ^ n28092 ;
  assign n31031 = n29528 ^ n28092 ;
  assign n31032 = ~n31030 & n31031 ;
  assign n31033 = n31032 ^ n28217 ;
  assign n30416 = n30177 ^ n28757 ;
  assign n30418 = n30417 ^ n27952 ;
  assign n30419 = n30418 ^ n30177 ;
  assign n30420 = n30419 ^ n30417 ;
  assign n30421 = ~n30416 & ~n30420 ;
  assign n30422 = n30421 ^ n30418 ;
  assign n30560 = n28766 ^ n27951 ;
  assign n30561 = n29507 ^ n28766 ;
  assign n30562 = ~n30560 & ~n30561 ;
  assign n30563 = n30562 ^ n27951 ;
  assign n30564 = n30563 ^ n30417 ;
  assign n30565 = n30564 ^ n30563 ;
  assign n29903 = n28754 ^ n27898 ;
  assign n29905 = n29904 ^ n28754 ;
  assign n29906 = n29903 & ~n29905 ;
  assign n29907 = n29906 ^ n27898 ;
  assign n29908 = n29907 ^ n29902 ;
  assign n29910 = n29909 ^ n29029 ;
  assign n29912 = n29911 ^ n28341 ;
  assign n29913 = n29912 ^ n29909 ;
  assign n29914 = n29913 ^ n29911 ;
  assign n29915 = ~n29910 & ~n29914 ;
  assign n29916 = n29915 ^ n29912 ;
  assign n29917 = n29206 ^ n28480 ;
  assign n29919 = n29918 ^ n29206 ;
  assign n29920 = ~n29917 & n29919 ;
  assign n29921 = n29920 ^ n28480 ;
  assign n30394 = n29921 ^ n29911 ;
  assign n30383 = n29871 ^ n29760 ;
  assign n29928 = n29927 ^ n29926 ;
  assign n30381 = n29928 & n30380 ;
  assign n30382 = n30381 ^ n29927 ;
  assign n30384 = n30383 ^ n30382 ;
  assign n30385 = n30053 ^ n29188 ;
  assign n30386 = n30383 ^ n28105 ;
  assign n30387 = n30386 ^ n30053 ;
  assign n30388 = n30387 ^ n30383 ;
  assign n30389 = n30385 & n30388 ;
  assign n30390 = n30389 ^ n30386 ;
  assign n30391 = ~n30384 & ~n30390 ;
  assign n30392 = n30391 ^ n30383 ;
  assign n30393 = n30392 ^ n29921 ;
  assign n30395 = n30394 ^ n30393 ;
  assign n30396 = n29916 & ~n30395 ;
  assign n30397 = n30396 ^ n30394 ;
  assign n30401 = n30398 ^ n29921 ;
  assign n30400 = n30399 ^ n30398 ;
  assign n30402 = n30401 ^ n30400 ;
  assign n30403 = n30397 & n30402 ;
  assign n30404 = n30403 ^ n30401 ;
  assign n30410 = n30398 ^ n29907 ;
  assign n30405 = n29359 ^ n28558 ;
  assign n30406 = n30115 ^ n29359 ;
  assign n30407 = n30405 & n30406 ;
  assign n30408 = n30407 ^ n28558 ;
  assign n30409 = n30408 ^ n29907 ;
  assign n30411 = n30410 ^ n30409 ;
  assign n30412 = ~n30404 & ~n30411 ;
  assign n30413 = n30412 ^ n30410 ;
  assign n30414 = ~n29908 & n30413 ;
  assign n30415 = n30414 ^ n29907 ;
  assign n30566 = n30565 ^ n30415 ;
  assign n30567 = n30422 & ~n30566 ;
  assign n30568 = n30567 ^ n30564 ;
  assign n30841 = n28744 ^ n28004 ;
  assign n30842 = n29514 ^ n28744 ;
  assign n30843 = ~n30841 & n30842 ;
  assign n30844 = n30843 ^ n28004 ;
  assign n30846 = n30844 ^ n30569 ;
  assign n30845 = n30844 ^ n30563 ;
  assign n30847 = n30846 ^ n30845 ;
  assign n30848 = n30568 & ~n30847 ;
  assign n30849 = n30848 ^ n30845 ;
  assign n30881 = n29497 ^ n28738 ;
  assign n30882 = n29497 ^ n28055 ;
  assign n30883 = n30881 & ~n30882 ;
  assign n30884 = n30883 ^ n28738 ;
  assign n30886 = n30884 ^ n30850 ;
  assign n30885 = n30884 ^ n30844 ;
  assign n30887 = n30886 ^ n30885 ;
  assign n30888 = n30849 & ~n30887 ;
  assign n30889 = n30888 ^ n30885 ;
  assign n30890 = n30238 ^ n30216 ;
  assign n31026 = n31024 ^ n30890 ;
  assign n31025 = n31024 ^ n30884 ;
  assign n31027 = n31026 ^ n31025 ;
  assign n31028 = n30889 & ~n31027 ;
  assign n31029 = n31028 ^ n31025 ;
  assign n31034 = n31033 ^ n31029 ;
  assign n31062 = n31034 ^ n26605 ;
  assign n30851 = n30850 ^ n30849 ;
  assign n30852 = n30851 ^ n27342 ;
  assign n30570 = n30569 ^ n30568 ;
  assign n30424 = n30413 ^ n29902 ;
  assign n30425 = n30424 ^ n27350 ;
  assign n30547 = n30408 ^ n30404 ;
  assign n30426 = n30399 ^ n30397 ;
  assign n30427 = n30426 ^ n27989 ;
  assign n30538 = n30392 ^ n29916 ;
  assign n30531 = n30530 ^ n30429 ;
  assign n30532 = ~n30430 & n30531 ;
  assign n30533 = n30532 ^ n27892 ;
  assign n30428 = n30390 ^ n30382 ;
  assign n30534 = n30533 ^ n30428 ;
  assign n30535 = n30533 ^ n27917 ;
  assign n30536 = ~n30534 & n30535 ;
  assign n30537 = n30536 ^ n27917 ;
  assign n30539 = n30538 ^ n30537 ;
  assign n30540 = n30426 ^ n27938 ;
  assign n30541 = n30540 ^ n30426 ;
  assign n30542 = n30541 ^ n30537 ;
  assign n30543 = ~n30539 & n30542 ;
  assign n30544 = n30543 ^ n30540 ;
  assign n30545 = n30427 & n30544 ;
  assign n30546 = n30545 ^ n27989 ;
  assign n30548 = n30547 ^ n30546 ;
  assign n30549 = n30547 ^ n28043 ;
  assign n30550 = n30548 & ~n30549 ;
  assign n30551 = n30550 ^ n28043 ;
  assign n30552 = n30551 ^ n30424 ;
  assign n30553 = n30425 & ~n30552 ;
  assign n30554 = n30553 ^ n27350 ;
  assign n30423 = n30422 ^ n30415 ;
  assign n30555 = n30554 ^ n30423 ;
  assign n30556 = n30554 ^ n27352 ;
  assign n30557 = n30555 & n30556 ;
  assign n30558 = n30557 ^ n27352 ;
  assign n30837 = n30570 ^ n30558 ;
  assign n30838 = n30570 ^ n27344 ;
  assign n30839 = n30837 & ~n30838 ;
  assign n30840 = n30839 ^ n27344 ;
  assign n30892 = n30851 ^ n30840 ;
  assign n30893 = n30852 & n30892 ;
  assign n30894 = n30893 ^ n27342 ;
  assign n30895 = n30894 ^ n27338 ;
  assign n30891 = n30890 ^ n30889 ;
  assign n31035 = n30894 ^ n30891 ;
  assign n31036 = ~n30895 & ~n31035 ;
  assign n31037 = n31036 ^ n27338 ;
  assign n31063 = n31062 ^ n31037 ;
  assign n30559 = n30558 ^ n27344 ;
  assign n30571 = n30570 ^ n30559 ;
  assign n30572 = n30544 ^ n27989 ;
  assign n30573 = n30537 ^ n27938 ;
  assign n30574 = n30573 ^ n30538 ;
  assign n30620 = n30618 & n30619 ;
  assign n30621 = n30428 ^ n27917 ;
  assign n30622 = n30621 ^ n30533 ;
  assign n30623 = ~n30620 & n30622 ;
  assign n30624 = n30574 & n30623 ;
  assign n30625 = n30572 & n30624 ;
  assign n30626 = n30546 ^ n28043 ;
  assign n30627 = n30626 ^ n30547 ;
  assign n30628 = ~n30625 & ~n30627 ;
  assign n30629 = n30551 ^ n30425 ;
  assign n30630 = n30628 & n30629 ;
  assign n30631 = n30423 ^ n27352 ;
  assign n30632 = n30631 ^ n30554 ;
  assign n30633 = n30630 & ~n30632 ;
  assign n30836 = ~n30571 & n30633 ;
  assign n30853 = n30852 ^ n30840 ;
  assign n30880 = ~n30836 & ~n30853 ;
  assign n30896 = n30895 ^ n30891 ;
  assign n31039 = n30880 & ~n30896 ;
  assign n31064 = n31063 ^ n31039 ;
  assign n31065 = n31064 ^ n3171 ;
  assign n30898 = n28582 ^ n3142 ;
  assign n30899 = n30898 ^ n2519 ;
  assign n30900 = n30899 ^ n3166 ;
  assign n30897 = n30896 ^ n30880 ;
  assign n30901 = n30900 ^ n30897 ;
  assign n30854 = n30853 ^ n30836 ;
  assign n30858 = n30857 ^ n30854 ;
  assign n30637 = n28598 ^ n3209 ;
  assign n30638 = n30637 ^ n25366 ;
  assign n30639 = n30638 ^ n2565 ;
  assign n30636 = n30632 ^ n30630 ;
  assign n30640 = n30639 ^ n30636 ;
  assign n30801 = n30643 ^ n2828 ;
  assign n30644 = n30627 ^ n30625 ;
  assign n30645 = n30644 ^ n30643 ;
  assign n30646 = n30624 ^ n30572 ;
  assign n30647 = n30646 ^ n1332 ;
  assign n30648 = n30623 ^ n30574 ;
  assign n1309 = n1269 ^ n1212 ;
  assign n1310 = n1309 ^ n1306 ;
  assign n1314 = n1313 ^ n1310 ;
  assign n30649 = n30648 ^ n1314 ;
  assign n30650 = n30622 ^ n30620 ;
  assign n1291 = n1197 ^ n1123 ;
  assign n1298 = n1297 ^ n1291 ;
  assign n1299 = n1298 ^ n1067 ;
  assign n30651 = n30650 ^ n1299 ;
  assign n30787 = n30786 ^ n1694 ;
  assign n30788 = ~n30653 & n30787 ;
  assign n30789 = n30788 ^ n30652 ;
  assign n30790 = n30789 ^ n1299 ;
  assign n30791 = ~n30651 & n30790 ;
  assign n30792 = n30791 ^ n30650 ;
  assign n30793 = n30792 ^ n1314 ;
  assign n30794 = n30649 & n30793 ;
  assign n30795 = n30794 ^ n30648 ;
  assign n30796 = n30795 ^ n1332 ;
  assign n30797 = n30647 & n30796 ;
  assign n30798 = n30797 ^ n1332 ;
  assign n30799 = n30798 ^ n30643 ;
  assign n30800 = ~n30645 & n30799 ;
  assign n30802 = n30801 ^ n30800 ;
  assign n30805 = n30629 ^ n30628 ;
  assign n30803 = n30636 ^ n2828 ;
  assign n30804 = n30803 ^ n30636 ;
  assign n30806 = n30805 ^ n30804 ;
  assign n30807 = n30802 & ~n30806 ;
  assign n30808 = n30807 ^ n30803 ;
  assign n30809 = n30640 & ~n30808 ;
  assign n30810 = n30809 ^ n30639 ;
  assign n2649 = n2648 ^ n2513 ;
  assign n2650 = n2649 ^ n2570 ;
  assign n2651 = n2650 ^ n2627 ;
  assign n30832 = n30810 ^ n2651 ;
  assign n30634 = n30633 ^ n30571 ;
  assign n30833 = n30810 ^ n30634 ;
  assign n30834 = n30832 & ~n30833 ;
  assign n30835 = n30834 ^ n2651 ;
  assign n30877 = n30854 ^ n30835 ;
  assign n30878 = n30858 & ~n30877 ;
  assign n30879 = n30878 ^ n30857 ;
  assign n31066 = n30897 ^ n30879 ;
  assign n31067 = ~n30901 & n31066 ;
  assign n31068 = n31067 ^ n30900 ;
  assign n31069 = n31068 ^ n3171 ;
  assign n31070 = n31065 & n31069 ;
  assign n31057 = n28571 ^ n2765 ;
  assign n31058 = n31057 ^ n3161 ;
  assign n31059 = n31058 ^ n1823 ;
  assign n31060 = n31059 ^ n3171 ;
  assign n31053 = n31033 ^ n31024 ;
  assign n31054 = ~n31029 & ~n31053 ;
  assign n31049 = n29489 ^ n28088 ;
  assign n31050 = n28226 ^ n28088 ;
  assign n31051 = n31049 & ~n31050 ;
  assign n31046 = n31033 ^ n27373 ;
  assign n31047 = n31046 ^ n28226 ;
  assign n31045 = n30243 ^ n30207 ;
  assign n31048 = n31047 ^ n31045 ;
  assign n31052 = n31051 ^ n31048 ;
  assign n31055 = n31054 ^ n31052 ;
  assign n31038 = n31037 ^ n31034 ;
  assign n31042 = n31039 ^ n31034 ;
  assign n31043 = n31038 & ~n31042 ;
  assign n31040 = n31039 ^ n31038 ;
  assign n31041 = n26605 & ~n31040 ;
  assign n31044 = n31043 ^ n31041 ;
  assign n31056 = n31055 ^ n31044 ;
  assign n31061 = n31060 ^ n31056 ;
  assign n31071 = n31070 ^ n31061 ;
  assign n31019 = n29968 ^ n29567 ;
  assign n31020 = n29567 ^ n28945 ;
  assign n31021 = n31019 & n31020 ;
  assign n31022 = n31021 ^ n28945 ;
  assign n31072 = n31071 ^ n31022 ;
  assign n31073 = n29974 ^ n29555 ;
  assign n31074 = n31068 ^ n31065 ;
  assign n31075 = n31074 ^ n28844 ;
  assign n31076 = n31075 ^ n29974 ;
  assign n31077 = n31076 ^ n31074 ;
  assign n31078 = ~n31073 & ~n31077 ;
  assign n31079 = n31078 ^ n31075 ;
  assign n30871 = n29981 ^ n28997 ;
  assign n30872 = n28997 ^ n28069 ;
  assign n30873 = ~n30871 & n30872 ;
  assign n30874 = n30873 ^ n28069 ;
  assign n30635 = n30634 ^ n2651 ;
  assign n30811 = n30810 ^ n30635 ;
  assign n30812 = n29018 ^ n28080 ;
  assign n30813 = n29990 ^ n29018 ;
  assign n30814 = ~n30812 & ~n30813 ;
  assign n30815 = n30814 ^ n28080 ;
  assign n30826 = n30811 & n30815 ;
  assign n30875 = n30874 ^ n30826 ;
  assign n30825 = n29987 ^ n29009 ;
  assign n30827 = n30826 ^ n28783 ;
  assign n30828 = n30827 ^ n29987 ;
  assign n30829 = n30828 ^ n30826 ;
  assign n30830 = ~n30825 & n30829 ;
  assign n30831 = n30830 ^ n30827 ;
  assign n30859 = n30858 ^ n30835 ;
  assign n30869 = n30859 ^ n30826 ;
  assign n30870 = ~n30831 & n30869 ;
  assign n30876 = n30875 ^ n30870 ;
  assign n30902 = n30901 ^ n30879 ;
  assign n31082 = n30902 ^ n30874 ;
  assign n31083 = ~n30876 & ~n31082 ;
  assign n31084 = n31083 ^ n30902 ;
  assign n31080 = n31074 ^ n31022 ;
  assign n31081 = n31080 ^ n31022 ;
  assign n31085 = n31084 ^ n31081 ;
  assign n31086 = n31079 & ~n31085 ;
  assign n31087 = n31086 ^ n31080 ;
  assign n31088 = n31072 & n31087 ;
  assign n31023 = n31022 ^ n31013 ;
  assign n31089 = n31088 ^ n31023 ;
  assign n31090 = ~n31018 & ~n31089 ;
  assign n31092 = n31091 ^ n31090 ;
  assign n31093 = n31012 & n31092 ;
  assign n31094 = n31093 ^ n31011 ;
  assign n31095 = n31094 ^ n31005 ;
  assign n31096 = n31006 & ~n31095 ;
  assign n31097 = n31096 ^ n30907 ;
  assign n31001 = n30733 ^ n30711 ;
  assign n31098 = n31097 ^ n31001 ;
  assign n31099 = n30325 ^ n28971 ;
  assign n31100 = n31001 ^ n29108 ;
  assign n31101 = n31100 ^ n30325 ;
  assign n31102 = n31101 ^ n31001 ;
  assign n31103 = ~n31099 & ~n31102 ;
  assign n31104 = n31103 ^ n31100 ;
  assign n31105 = ~n31098 & n31104 ;
  assign n31106 = n31105 ^ n31097 ;
  assign n31107 = n31106 ^ n30995 ;
  assign n31108 = ~n31000 & ~n31107 ;
  assign n31110 = n31109 ^ n31108 ;
  assign n31111 = ~n30993 & ~n31110 ;
  assign n31112 = n31111 ^ n30992 ;
  assign n31113 = n31112 ^ n30982 ;
  assign n31114 = ~n30987 & ~n31113 ;
  assign n31116 = n31115 ^ n31114 ;
  assign n31117 = ~n30980 & ~n31116 ;
  assign n31118 = n31117 ^ n30979 ;
  assign n30974 = n30749 ^ n30748 ;
  assign n31119 = n31118 ^ n30974 ;
  assign n31120 = n29890 ^ n28972 ;
  assign n31121 = n29937 ^ n28972 ;
  assign n31122 = ~n31120 & ~n31121 ;
  assign n31123 = n31122 ^ n29890 ;
  assign n31124 = n31123 ^ n30974 ;
  assign n31125 = ~n31119 & ~n31124 ;
  assign n31126 = n31125 ^ n31118 ;
  assign n31127 = n31126 ^ n30965 ;
  assign n31129 = n31128 ^ n31127 ;
  assign n31130 = n30973 & ~n31129 ;
  assign n31131 = n31130 ^ n31128 ;
  assign n31132 = ~n30966 & ~n31131 ;
  assign n31133 = n31132 ^ n30965 ;
  assign n30960 = n30758 ^ n30680 ;
  assign n31134 = n31133 ^ n30960 ;
  assign n31135 = n30008 ^ n29159 ;
  assign n31136 = n30383 ^ n29159 ;
  assign n31137 = ~n31135 & ~n31136 ;
  assign n31138 = n31137 ^ n30008 ;
  assign n31139 = n31138 ^ n30960 ;
  assign n31140 = n31134 & ~n31139 ;
  assign n31141 = n31140 ^ n31133 ;
  assign n31142 = n31141 ^ n30951 ;
  assign n31144 = n31143 ^ n31142 ;
  assign n31145 = ~n30959 & n31144 ;
  assign n31146 = n31145 ^ n31143 ;
  assign n31147 = ~n30952 & n31146 ;
  assign n31149 = n31148 ^ n31147 ;
  assign n31150 = n30946 & ~n31149 ;
  assign n31151 = n31150 ^ n30945 ;
  assign n31152 = n31151 ^ n30935 ;
  assign n31153 = ~n30940 & ~n31152 ;
  assign n31154 = n31153 ^ n30939 ;
  assign n31155 = n31154 ^ n30929 ;
  assign n31156 = n30934 & ~n31155 ;
  assign n31158 = n31157 ^ n31156 ;
  assign n31159 = n30927 & ~n31158 ;
  assign n31160 = n31159 ^ n30926 ;
  assign n30916 = n30177 ^ n29359 ;
  assign n30917 = n30890 ^ n30177 ;
  assign n30918 = ~n30916 & ~n30917 ;
  assign n30919 = n30918 ^ n29359 ;
  assign n30920 = n30919 ^ n30910 ;
  assign n30921 = n30920 ^ n30919 ;
  assign n31161 = n31160 ^ n30921 ;
  assign n31162 = ~n30915 & ~n31161 ;
  assign n31163 = n31162 ^ n30920 ;
  assign n31164 = n30784 ^ n1688 ;
  assign n31282 = n31164 ^ n30919 ;
  assign n31283 = n31163 & n31282 ;
  assign n31284 = n31283 ^ n30919 ;
  assign n31292 = n31291 ^ n31284 ;
  assign n31293 = n31292 ^ n27898 ;
  assign n31165 = n31164 ^ n31163 ;
  assign n31166 = n31165 ^ n28558 ;
  assign n31273 = n31160 ^ n30915 ;
  assign n31167 = n31158 ^ n30926 ;
  assign n31168 = n31167 ^ n28341 ;
  assign n31169 = n31154 ^ n30934 ;
  assign n31170 = n31169 ^ n28105 ;
  assign n31258 = n31149 ^ n30944 ;
  assign n31172 = n31146 ^ n30950 ;
  assign n31173 = n31172 ^ n28126 ;
  assign n31175 = n31139 ^ n31133 ;
  assign n31176 = n31175 ^ n28310 ;
  assign n31178 = n31126 ^ n30973 ;
  assign n31179 = n31178 ^ n28135 ;
  assign n31180 = n31124 ^ n31118 ;
  assign n31181 = n31180 ^ n28142 ;
  assign n31182 = n31116 ^ n30978 ;
  assign n31183 = n31182 ^ n28282 ;
  assign n31217 = n31106 ^ n31000 ;
  assign n31184 = n31104 ^ n31097 ;
  assign n31185 = n31184 ^ n28170 ;
  assign n31186 = n31094 ^ n31006 ;
  assign n31187 = n31186 ^ n27516 ;
  assign n31206 = n31092 ^ n31010 ;
  assign n31201 = n31089 ^ n31017 ;
  assign n31196 = n31087 ^ n31071 ;
  assign n30816 = n30815 ^ n30811 ;
  assign n30823 = n28211 & n30816 ;
  assign n30824 = n30823 ^ n28201 ;
  assign n30860 = n30859 ^ n30831 ;
  assign n30865 = n30860 ^ n30823 ;
  assign n30866 = ~n30824 & n30865 ;
  assign n30867 = n30866 ^ n28201 ;
  assign n30868 = n30867 ^ n28100 ;
  assign n30903 = n30902 ^ n30876 ;
  assign n31189 = n30903 ^ n30867 ;
  assign n31190 = n30868 & ~n31189 ;
  assign n31191 = n31190 ^ n28100 ;
  assign n31188 = n31084 ^ n31079 ;
  assign n31192 = n31191 ^ n31188 ;
  assign n31193 = n31191 ^ n28090 ;
  assign n31194 = ~n31192 & ~n31193 ;
  assign n31195 = n31194 ^ n28090 ;
  assign n31197 = n31196 ^ n31195 ;
  assign n31198 = n31196 ^ n28082 ;
  assign n31199 = ~n31197 & ~n31198 ;
  assign n31200 = n31199 ^ n28082 ;
  assign n31202 = n31201 ^ n31200 ;
  assign n31203 = n31201 ^ n28075 ;
  assign n31204 = ~n31202 & n31203 ;
  assign n31205 = n31204 ^ n28075 ;
  assign n31207 = n31206 ^ n31205 ;
  assign n31208 = n31206 ^ n28177 ;
  assign n31209 = ~n31207 & n31208 ;
  assign n31210 = n31209 ^ n28177 ;
  assign n31211 = n31210 ^ n31186 ;
  assign n31212 = n31187 & ~n31211 ;
  assign n31213 = n31212 ^ n27516 ;
  assign n31214 = n31213 ^ n31184 ;
  assign n31215 = ~n31185 & n31214 ;
  assign n31216 = n31215 ^ n28170 ;
  assign n31218 = n31217 ^ n31216 ;
  assign n31219 = n31110 ^ n30988 ;
  assign n31220 = n31219 ^ n28157 ;
  assign n31221 = n31220 ^ n31216 ;
  assign n31222 = n31221 ^ n31219 ;
  assign n31223 = n31218 & ~n31222 ;
  assign n31224 = n31223 ^ n31220 ;
  assign n31225 = n31112 ^ n30987 ;
  assign n31227 = n31225 ^ n28155 ;
  assign n31226 = n31225 ^ n31219 ;
  assign n31228 = n31227 ^ n31226 ;
  assign n31229 = n31224 & ~n31228 ;
  assign n31230 = n31229 ^ n31227 ;
  assign n31232 = n31182 ^ n28278 ;
  assign n31231 = n31225 ^ n31182 ;
  assign n31233 = n31232 ^ n31231 ;
  assign n31234 = ~n31230 & ~n31233 ;
  assign n31235 = n31234 ^ n31232 ;
  assign n31236 = ~n31183 & ~n31235 ;
  assign n31237 = n31236 ^ n28282 ;
  assign n31238 = n31237 ^ n31180 ;
  assign n31239 = n31181 & n31238 ;
  assign n31240 = n31239 ^ n28142 ;
  assign n31241 = n31240 ^ n31178 ;
  assign n31242 = ~n31179 & ~n31241 ;
  assign n31243 = n31242 ^ n28135 ;
  assign n31177 = n31131 ^ n30964 ;
  assign n31244 = n31243 ^ n31177 ;
  assign n31245 = n31243 ^ n28129 ;
  assign n31246 = n31244 & ~n31245 ;
  assign n31247 = n31246 ^ n28129 ;
  assign n31248 = n31247 ^ n31175 ;
  assign n31249 = n31176 & ~n31248 ;
  assign n31250 = n31249 ^ n28310 ;
  assign n31174 = n31141 ^ n30959 ;
  assign n31251 = n31250 ^ n31174 ;
  assign n31252 = n31250 ^ n28316 ;
  assign n31253 = n31251 & n31252 ;
  assign n31254 = n31253 ^ n28316 ;
  assign n31255 = n31254 ^ n31172 ;
  assign n31256 = ~n31173 & n31255 ;
  assign n31257 = n31256 ^ n28126 ;
  assign n31259 = n31258 ^ n31257 ;
  assign n31260 = n31258 ^ n28112 ;
  assign n31261 = ~n31259 & ~n31260 ;
  assign n31262 = n31261 ^ n28112 ;
  assign n31171 = n31151 ^ n30940 ;
  assign n31263 = n31262 ^ n31171 ;
  assign n31264 = n31262 ^ n28329 ;
  assign n31265 = n31263 & ~n31264 ;
  assign n31266 = n31265 ^ n28329 ;
  assign n31267 = n31266 ^ n31169 ;
  assign n31268 = n31170 & ~n31267 ;
  assign n31269 = n31268 ^ n28105 ;
  assign n31270 = n31269 ^ n31167 ;
  assign n31271 = ~n31168 & n31270 ;
  assign n31272 = n31271 ^ n28341 ;
  assign n31274 = n31273 ^ n31272 ;
  assign n31275 = n31165 ^ n28480 ;
  assign n31276 = n31275 ^ n31165 ;
  assign n31277 = n31276 ^ n31272 ;
  assign n31278 = ~n31274 & n31277 ;
  assign n31279 = n31278 ^ n31275 ;
  assign n31280 = n31166 & ~n31279 ;
  assign n31281 = n31280 ^ n28558 ;
  assign n31548 = n31292 ^ n31281 ;
  assign n31549 = ~n31293 & ~n31548 ;
  assign n31550 = n31549 ^ n27898 ;
  assign n31543 = n31286 ^ n31284 ;
  assign n31544 = n31291 & ~n31543 ;
  assign n31545 = n31544 ^ n31286 ;
  assign n31536 = n31045 ^ n29514 ;
  assign n31537 = n30789 ^ n30651 ;
  assign n31538 = n31537 ^ n28757 ;
  assign n31539 = n31538 ^ n31045 ;
  assign n31540 = n31539 ^ n31537 ;
  assign n31541 = n31536 & n31540 ;
  assign n31542 = n31541 ^ n31538 ;
  assign n31546 = n31545 ^ n31542 ;
  assign n31547 = n31546 ^ n27952 ;
  assign n31551 = n31550 ^ n31547 ;
  assign n31294 = n31293 ^ n31281 ;
  assign n31295 = n31272 ^ n28480 ;
  assign n31296 = n31295 ^ n31273 ;
  assign n31297 = n31269 ^ n31168 ;
  assign n31298 = n31266 ^ n31170 ;
  assign n31299 = n31171 ^ n28329 ;
  assign n31300 = n31299 ^ n31262 ;
  assign n31301 = n31260 ^ n31257 ;
  assign n31302 = n31174 ^ n28316 ;
  assign n31303 = n31302 ^ n31250 ;
  assign n31304 = n31247 ^ n31176 ;
  assign n31305 = n31177 ^ n28129 ;
  assign n31306 = n31305 ^ n31243 ;
  assign n31307 = n31230 ^ n28278 ;
  assign n31308 = n31217 ^ n28157 ;
  assign n31309 = n31308 ^ n31216 ;
  assign n31310 = n31210 ^ n31187 ;
  assign n31311 = n31205 ^ n28177 ;
  assign n31312 = n31311 ^ n31206 ;
  assign n30904 = n30903 ^ n30868 ;
  assign n31313 = n31188 ^ n28090 ;
  assign n31314 = n31313 ^ n31191 ;
  assign n31315 = n30904 & ~n31314 ;
  assign n31316 = n31195 ^ n28082 ;
  assign n31317 = n31316 ^ n31196 ;
  assign n31318 = n31315 & n31317 ;
  assign n31319 = n31200 ^ n28075 ;
  assign n31320 = n31319 ^ n31201 ;
  assign n31321 = ~n31318 & ~n31320 ;
  assign n31322 = n31312 & ~n31321 ;
  assign n31323 = n31310 & n31322 ;
  assign n31324 = n31213 ^ n31185 ;
  assign n31325 = ~n31323 & n31324 ;
  assign n31326 = ~n31309 & n31325 ;
  assign n31327 = n31224 ^ n28155 ;
  assign n31328 = ~n31326 & n31327 ;
  assign n31329 = n31307 & n31328 ;
  assign n31330 = n31235 ^ n28282 ;
  assign n31331 = n31329 & ~n31330 ;
  assign n31332 = n31237 ^ n31181 ;
  assign n31333 = n31331 & ~n31332 ;
  assign n31334 = n31240 ^ n31179 ;
  assign n31335 = ~n31333 & n31334 ;
  assign n31336 = ~n31306 & ~n31335 ;
  assign n31337 = n31304 & n31336 ;
  assign n31338 = ~n31303 & n31337 ;
  assign n31339 = n31254 ^ n31173 ;
  assign n31340 = ~n31338 & n31339 ;
  assign n31341 = ~n31301 & ~n31340 ;
  assign n31342 = ~n31300 & n31341 ;
  assign n31343 = ~n31298 & ~n31342 ;
  assign n31344 = n31297 & n31343 ;
  assign n31345 = ~n31296 & n31344 ;
  assign n31346 = n31279 ^ n28558 ;
  assign n31347 = ~n31345 & n31346 ;
  assign n31552 = ~n31294 & n31347 ;
  assign n31573 = n31551 & n31552 ;
  assign n31566 = n29497 ^ n28766 ;
  assign n31567 = n30278 ^ n29497 ;
  assign n31568 = ~n31566 & n31567 ;
  assign n31569 = n31568 ^ n28766 ;
  assign n31560 = n30792 ^ n30649 ;
  assign n31562 = n31560 ^ n31537 ;
  assign n31561 = n31560 ^ n31545 ;
  assign n31563 = n31562 ^ n31561 ;
  assign n31564 = n31542 & n31563 ;
  assign n31565 = n31564 ^ n31562 ;
  assign n31570 = n31569 ^ n31565 ;
  assign n31571 = n31570 ^ n27951 ;
  assign n31556 = n31550 ^ n31546 ;
  assign n31557 = n31550 ^ n27952 ;
  assign n31558 = ~n31556 & ~n31557 ;
  assign n31559 = n31558 ^ n27952 ;
  assign n31572 = n31571 ^ n31559 ;
  assign n31574 = n31573 ^ n31572 ;
  assign n31578 = n31577 ^ n31574 ;
  assign n31553 = n31552 ^ n31551 ;
  assign n31579 = n31578 ^ n31553 ;
  assign n31348 = n31347 ^ n31294 ;
  assign n2876 = n2861 ^ n2842 ;
  assign n2883 = n2882 ^ n2876 ;
  assign n2887 = n2886 ^ n2883 ;
  assign n31349 = n31344 ^ n31296 ;
  assign n1771 = n1746 ^ n1427 ;
  assign n1772 = n1771 ^ n1765 ;
  assign n1773 = n1772 ^ n1349 ;
  assign n31350 = n31349 ^ n1773 ;
  assign n31351 = n31336 ^ n31304 ;
  assign n31352 = ~n1590 & n31351 ;
  assign n31353 = n31337 ^ n31303 ;
  assign n31357 = ~n31353 & ~n31356 ;
  assign n31358 = ~n31352 & n31357 ;
  assign n31359 = n31358 ^ n31352 ;
  assign n887 = n856 ^ n826 ;
  assign n888 = n887 ^ n884 ;
  assign n892 = n891 ^ n888 ;
  assign n31360 = n31359 ^ n892 ;
  assign n31361 = n31340 ^ n31301 ;
  assign n31362 = n31339 ^ n31338 ;
  assign n31363 = ~n877 & n31362 ;
  assign n31364 = ~n31359 & n31363 ;
  assign n31365 = n31364 ^ n31359 ;
  assign n31366 = n31361 & ~n31365 ;
  assign n31367 = ~n31360 & n31366 ;
  assign n31368 = n31367 ^ n31365 ;
  assign n31369 = ~n31350 & ~n31368 ;
  assign n1158 = n1157 ^ n1070 ;
  assign n1159 = n1158 ^ n1151 ;
  assign n1160 = n1159 ^ n1142 ;
  assign n31370 = n31343 ^ n31297 ;
  assign n31371 = ~n1160 & ~n31370 ;
  assign n31372 = n31369 & ~n31371 ;
  assign n31373 = n31341 ^ n31300 ;
  assign n31375 = n996 & n31373 ;
  assign n31374 = n31373 ^ n996 ;
  assign n31376 = n31375 ^ n31374 ;
  assign n1753 = n1728 ^ n1416 ;
  assign n1754 = n1753 ^ n1003 ;
  assign n1755 = n1754 ^ n1145 ;
  assign n31377 = n31342 ^ n31298 ;
  assign n31378 = ~n1755 & ~n31377 ;
  assign n31379 = n31376 & n31378 ;
  assign n31380 = n31379 ^ n31376 ;
  assign n31381 = n31372 & n31380 ;
  assign n31385 = n31335 ^ n31306 ;
  assign n31386 = n31385 ^ n31384 ;
  assign n31387 = n31334 ^ n31333 ;
  assign n31391 = n31390 ^ n31387 ;
  assign n31392 = n31332 ^ n31331 ;
  assign n2943 = n2942 ^ n2939 ;
  assign n2944 = n2943 ^ n599 ;
  assign n2948 = n2947 ^ n2944 ;
  assign n31393 = n31392 ^ n2948 ;
  assign n31398 = n31330 ^ n31329 ;
  assign n31399 = n31398 ^ n31396 ;
  assign n31401 = n28875 ^ n593 ;
  assign n31402 = n31401 ^ n25827 ;
  assign n31403 = n31402 ^ n20760 ;
  assign n31400 = n31328 ^ n31307 ;
  assign n31404 = n31403 ^ n31400 ;
  assign n31459 = n21779 ^ n2395 ;
  assign n31460 = n31459 ^ n25832 ;
  assign n31461 = n31460 ^ n1469 ;
  assign n31462 = n31461 ^ n31400 ;
  assign n31457 = n31327 ^ n31326 ;
  assign n31408 = n31325 ^ n31309 ;
  assign n31405 = n21785 ^ n2386 ;
  assign n31406 = n31405 ^ n2356 ;
  assign n31407 = n31406 ^ n20768 ;
  assign n31409 = n31408 ^ n31407 ;
  assign n31411 = n31324 ^ n31323 ;
  assign n2343 = n2309 ^ n2267 ;
  assign n2344 = n2343 ^ n2340 ;
  assign n2348 = n2347 ^ n2344 ;
  assign n31412 = n31411 ^ n2348 ;
  assign n31413 = n31322 ^ n31310 ;
  assign n2331 = n2252 ^ n2199 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2333 = n2332 ^ n2321 ;
  assign n31414 = n31413 ^ n2333 ;
  assign n31416 = n28890 ^ n2184 ;
  assign n31417 = n31416 ^ n25842 ;
  assign n31418 = n31417 ^ n2328 ;
  assign n31415 = n31321 ^ n31312 ;
  assign n31419 = n31418 ^ n31415 ;
  assign n31421 = n28894 ^ n2177 ;
  assign n31422 = n31421 ^ n25868 ;
  assign n31423 = n31422 ^ n2021 ;
  assign n31420 = n31320 ^ n31318 ;
  assign n31424 = n31423 ^ n31420 ;
  assign n31426 = n28899 ^ n21801 ;
  assign n31427 = n31426 ^ n1943 ;
  assign n31428 = n31427 ^ n20390 ;
  assign n31425 = n31317 ^ n31315 ;
  assign n31429 = n31428 ^ n31425 ;
  assign n1878 = n1877 ^ n1868 ;
  assign n1891 = n1890 ^ n1878 ;
  assign n1895 = n1894 ^ n1891 ;
  assign n30905 = n30904 ^ n1895 ;
  assign n30819 = n28904 ^ n21810 ;
  assign n30820 = n30819 ^ n3002 ;
  assign n30821 = n30820 ^ n1885 ;
  assign n30817 = n30816 ^ n28211 ;
  assign n30818 = n3236 & n30817 ;
  assign n30822 = n30821 ^ n30818 ;
  assign n30861 = n30860 ^ n30824 ;
  assign n30862 = n30861 ^ n30818 ;
  assign n30863 = n30822 & ~n30862 ;
  assign n30864 = n30863 ^ n30821 ;
  assign n31430 = n30864 ^ n1895 ;
  assign n31431 = n30905 & ~n31430 ;
  assign n31432 = n31431 ^ n31314 ;
  assign n31436 = n31314 ^ n30904 ;
  assign n31433 = n28915 ^ n21805 ;
  assign n31434 = n31433 ^ n25850 ;
  assign n31435 = n31434 ^ n1938 ;
  assign n31437 = n31436 ^ n31435 ;
  assign n31438 = ~n31432 & n31437 ;
  assign n31439 = n31438 ^ n31435 ;
  assign n31440 = n31439 ^ n31425 ;
  assign n31441 = ~n31429 & n31440 ;
  assign n31442 = n31441 ^ n31428 ;
  assign n31443 = n31442 ^ n31423 ;
  assign n31444 = n31424 & n31443 ;
  assign n31445 = n31444 ^ n31423 ;
  assign n31446 = n31445 ^ n31415 ;
  assign n31447 = n31419 & ~n31446 ;
  assign n31448 = n31447 ^ n31418 ;
  assign n31449 = n31448 ^ n31413 ;
  assign n31450 = ~n31414 & n31449 ;
  assign n31451 = n31450 ^ n2333 ;
  assign n31452 = n31451 ^ n31411 ;
  assign n31453 = ~n31412 & n31452 ;
  assign n31410 = n31407 ^ n2348 ;
  assign n31454 = n31453 ^ n31410 ;
  assign n31455 = ~n31409 & ~n31454 ;
  assign n31456 = n31455 ^ n31408 ;
  assign n31458 = n31457 ^ n31456 ;
  assign n31463 = n31462 ^ n31458 ;
  assign n31464 = n31463 ^ n31462 ;
  assign n31465 = n31456 ^ n31400 ;
  assign n31466 = n31465 ^ n31462 ;
  assign n31467 = n31464 & ~n31466 ;
  assign n31468 = n31467 ^ n31462 ;
  assign n31469 = ~n31404 & n31468 ;
  assign n31470 = n31469 ^ n31403 ;
  assign n31471 = n31470 ^ n31398 ;
  assign n31472 = n31399 & ~n31471 ;
  assign n31397 = n31396 ^ n2948 ;
  assign n31473 = n31472 ^ n31397 ;
  assign n31474 = n31393 & ~n31473 ;
  assign n31475 = n31474 ^ n31392 ;
  assign n31476 = n31475 ^ n31387 ;
  assign n31477 = ~n31391 & n31476 ;
  assign n31478 = n31477 ^ n31390 ;
  assign n31479 = n31478 ^ n31384 ;
  assign n31480 = ~n31386 & ~n31479 ;
  assign n31481 = n31480 ^ n31385 ;
  assign n31482 = n31381 & ~n31481 ;
  assign n31483 = n31375 ^ n1755 ;
  assign n31484 = n31377 ^ n1755 ;
  assign n31485 = ~n31483 & n31484 ;
  assign n31486 = n31485 ^ n31377 ;
  assign n31488 = n31380 & ~n31486 ;
  assign n31487 = n31486 ^ n31370 ;
  assign n31489 = n31488 ^ n31487 ;
  assign n31490 = n31489 ^ n31487 ;
  assign n31491 = n31361 ^ n892 ;
  assign n31499 = n31361 ^ n877 ;
  assign n31492 = n31356 ^ n31353 ;
  assign n31493 = n31351 ^ n1590 ;
  assign n31494 = n31493 ^ n31356 ;
  assign n31495 = n31494 ^ n31352 ;
  assign n31496 = n31492 & ~n31495 ;
  assign n31497 = n31496 ^ n31353 ;
  assign n31498 = n31497 ^ n31361 ;
  assign n31500 = n31499 ^ n31498 ;
  assign n31501 = n31362 ^ n31361 ;
  assign n31502 = n31501 ^ n31499 ;
  assign n31503 = n31500 & ~n31502 ;
  assign n31504 = n31503 ^ n31499 ;
  assign n31505 = ~n31491 & n31504 ;
  assign n31506 = n31505 ^ n892 ;
  assign n31509 = n31490 & n31506 ;
  assign n31510 = n31509 ^ n31487 ;
  assign n31512 = n1773 ^ n1160 ;
  assign n31511 = n31370 ^ n1773 ;
  assign n31513 = n31512 ^ n31511 ;
  assign n31514 = ~n31510 & n31513 ;
  assign n31515 = n31514 ^ n31512 ;
  assign n31516 = ~n31350 & n31515 ;
  assign n31517 = n31516 ^ n1773 ;
  assign n31518 = ~n31482 & ~n31517 ;
  assign n31520 = n29387 ^ n1445 ;
  assign n31521 = n31520 ^ n1385 ;
  assign n31522 = n31521 ^ n2879 ;
  assign n31519 = n31346 ^ n31345 ;
  assign n31524 = n31522 ^ n31519 ;
  assign n31523 = n31519 & n31522 ;
  assign n31525 = n31524 ^ n31523 ;
  assign n31526 = ~n31518 & n31525 ;
  assign n31527 = ~n2887 & n31526 ;
  assign n31528 = ~n31348 & n31527 ;
  assign n31529 = n31528 ^ n31526 ;
  assign n31530 = n31348 ^ n2887 ;
  assign n31531 = n31523 ^ n2887 ;
  assign n31532 = ~n31530 & n31531 ;
  assign n31533 = n31532 ^ n31523 ;
  assign n31534 = ~n31529 & ~n31533 ;
  assign n2897 = n2872 ^ n2857 ;
  assign n2898 = n2897 ^ n2894 ;
  assign n2902 = n2901 ^ n2898 ;
  assign n31535 = n31534 ^ n2902 ;
  assign n31554 = n31553 ^ n2902 ;
  assign n31555 = n31535 & ~n31554 ;
  assign n31580 = n31579 ^ n31555 ;
  assign n31585 = n31584 ^ n31580 ;
  assign n31586 = n31585 ^ n28080 ;
  assign n32054 = n2782 & ~n31586 ;
  assign n3034 = n3030 ^ n3015 ;
  assign n3041 = n3040 ^ n3034 ;
  assign n3045 = n3044 ^ n3041 ;
  assign n32055 = n32054 ^ n3045 ;
  assign n31884 = n28080 & ~n31585 ;
  assign n32056 = n31884 ^ n28783 ;
  assign n31797 = n31011 ^ n29974 ;
  assign n31793 = n31580 & ~n31584 ;
  assign n31798 = n31793 ^ n29009 ;
  assign n31799 = n31798 ^ n31011 ;
  assign n31800 = n31799 ^ n31793 ;
  assign n31801 = ~n31797 & n31800 ;
  assign n31802 = n31801 ^ n31798 ;
  assign n31743 = n31572 & n31573 ;
  assign n31715 = n31570 ^ n31559 ;
  assign n31716 = n31571 & ~n31715 ;
  assign n31717 = n31716 ^ n27951 ;
  assign n31689 = n31569 ^ n31560 ;
  assign n31690 = ~n31565 & ~n31689 ;
  assign n31691 = n31690 ^ n31560 ;
  assign n31684 = n29528 ^ n28744 ;
  assign n31685 = n30277 ^ n29528 ;
  assign n31686 = n31684 & n31685 ;
  assign n31687 = n31686 ^ n28744 ;
  assign n31683 = n30795 ^ n30647 ;
  assign n31688 = n31687 ^ n31683 ;
  assign n31713 = n31691 ^ n31688 ;
  assign n31714 = n31713 ^ n28004 ;
  assign n31742 = n31717 ^ n31714 ;
  assign n31776 = n31743 ^ n31742 ;
  assign n31772 = n29378 ^ n2630 ;
  assign n31773 = n31772 ^ n25949 ;
  assign n31774 = n31773 ^ n2605 ;
  assign n31794 = n31776 ^ n31774 ;
  assign n31755 = n31574 ^ n31553 ;
  assign n31756 = n31755 ^ n2902 ;
  assign n31757 = n31756 ^ n31533 ;
  assign n31758 = n31757 ^ n31755 ;
  assign n31759 = n31574 ^ n2902 ;
  assign n31760 = n31759 ^ n31755 ;
  assign n31761 = ~n31758 & ~n31760 ;
  assign n31762 = n31761 ^ n31755 ;
  assign n31763 = ~n31578 & ~n31762 ;
  assign n31764 = n31763 ^ n31577 ;
  assign n31765 = n31529 & ~n31578 ;
  assign n31766 = ~n31764 & n31765 ;
  assign n31768 = ~n2902 & n31553 ;
  assign n31770 = n31766 & n31768 ;
  assign n31767 = n31766 ^ n31764 ;
  assign n31771 = n31770 ^ n31767 ;
  assign n31795 = n31794 ^ n31771 ;
  assign n31885 = n31802 ^ n31795 ;
  assign n32057 = n32056 ^ n31885 ;
  assign n32058 = n32057 ^ n32054 ;
  assign n32059 = n32055 & ~n32058 ;
  assign n32060 = n32059 ^ n3045 ;
  assign n32050 = n29816 ^ n1918 ;
  assign n32051 = n32050 ^ n3052 ;
  assign n32052 = n32051 ^ n21195 ;
  assign n31886 = n31885 ^ n31884 ;
  assign n31887 = n31885 ^ n28783 ;
  assign n31888 = n31886 & n31887 ;
  assign n31889 = n31888 ^ n28783 ;
  assign n31807 = n30907 ^ n29968 ;
  assign n31775 = n31774 ^ n31771 ;
  assign n31777 = n31776 ^ n31771 ;
  assign n31778 = n31775 & ~n31777 ;
  assign n31779 = n31778 ^ n31774 ;
  assign n31718 = n31717 ^ n31713 ;
  assign n31719 = n31714 & ~n31718 ;
  assign n31720 = n31719 ^ n28004 ;
  assign n31697 = n30271 ^ n29489 ;
  assign n31695 = n30798 ^ n30645 ;
  assign n31698 = n31695 ^ n28738 ;
  assign n31699 = n31698 ^ n30271 ;
  assign n31700 = n31699 ^ n31695 ;
  assign n31701 = ~n31697 & n31700 ;
  assign n31702 = n31701 ^ n31698 ;
  assign n31692 = n31691 ^ n31683 ;
  assign n31693 = n31688 & n31692 ;
  assign n31694 = n31693 ^ n31687 ;
  assign n31711 = n31702 ^ n31694 ;
  assign n31712 = n31711 ^ n28055 ;
  assign n31745 = n31720 ^ n31712 ;
  assign n31744 = ~n31742 & ~n31743 ;
  assign n31753 = n31745 ^ n31744 ;
  assign n2598 = n2597 ^ n2498 ;
  assign n2608 = n2607 ^ n2598 ;
  assign n2612 = n2611 ^ n2608 ;
  assign n31754 = n31753 ^ n2612 ;
  assign n31805 = n31779 ^ n31754 ;
  assign n31808 = n31805 ^ n28997 ;
  assign n31809 = n31808 ^ n29968 ;
  assign n31810 = n31809 ^ n31805 ;
  assign n31811 = ~n31807 & ~n31810 ;
  assign n31812 = n31811 ^ n31808 ;
  assign n31796 = n31795 ^ n31793 ;
  assign n31803 = n31796 & n31802 ;
  assign n31804 = n31803 ^ n31795 ;
  assign n31882 = n31812 ^ n31804 ;
  assign n31883 = n31882 ^ n28069 ;
  assign n31963 = n31889 ^ n31883 ;
  assign n32053 = n32052 ^ n31963 ;
  assign n32275 = n32060 ^ n32053 ;
  assign n2868 = n2828 ^ n2558 ;
  assign n2869 = n2868 ^ n2867 ;
  assign n2873 = n2872 ^ n2869 ;
  assign n35729 = n2873 ^ n2570 ;
  assign n35730 = n35729 ^ n29469 ;
  assign n35731 = n35730 ^ n24002 ;
  assign n1676 = n1673 ^ n1657 ;
  assign n1677 = n1676 ^ n1029 ;
  assign n1678 = n1677 ^ n1195 ;
  assign n1105 = n1022 ^ n963 ;
  assign n1115 = n1114 ^ n1105 ;
  assign n1116 = n1115 ^ n1098 ;
  assign n1188 = n1116 ^ n1047 ;
  assign n1198 = n1197 ^ n1188 ;
  assign n1205 = n1204 ^ n1198 ;
  assign n35456 = n1678 ^ n1205 ;
  assign n32022 = n29791 ^ n2428 ;
  assign n32023 = n32022 ^ n26486 ;
  assign n32024 = n32023 ^ n2363 ;
  assign n31667 = n30979 ^ n30335 ;
  assign n31668 = n30335 ^ n28978 ;
  assign n31669 = n31667 & ~n31668 ;
  assign n31670 = n31669 ^ n28978 ;
  assign n30906 = n30905 ^ n30864 ;
  assign n31671 = n31670 ^ n30906 ;
  assign n31824 = n30861 ^ n30822 ;
  assign n31676 = n30817 ^ n3236 ;
  assign n31672 = n29945 ^ n29577 ;
  assign n31673 = n30988 ^ n29945 ;
  assign n31674 = n31672 & n31673 ;
  assign n31675 = n31674 ^ n29577 ;
  assign n31677 = n31676 ^ n31675 ;
  assign n31682 = n30265 ^ n28092 ;
  assign n31696 = n31695 ^ n31694 ;
  assign n31703 = ~n31696 & n31702 ;
  assign n31704 = n31703 ^ n31695 ;
  assign n31705 = n31704 ^ n29021 ;
  assign n31706 = n31705 ^ n30265 ;
  assign n31707 = n31706 ^ n31704 ;
  assign n31708 = n31682 & n31707 ;
  assign n31709 = n31708 ^ n31705 ;
  assign n31591 = n30805 ^ n30802 ;
  assign n31710 = n31709 ^ n31591 ;
  assign n31747 = n31710 ^ n28217 ;
  assign n31721 = n31720 ^ n28055 ;
  assign n31722 = n31712 & n31721 ;
  assign n31723 = n31722 ^ n31720 ;
  assign n31748 = n31747 ^ n31723 ;
  assign n31746 = n31744 & n31745 ;
  assign n31751 = n31748 ^ n31746 ;
  assign n31752 = n31751 ^ n3224 ;
  assign n31780 = n31779 ^ n31753 ;
  assign n31781 = n31754 & ~n31780 ;
  assign n31782 = n31781 ^ n2612 ;
  assign n31783 = n31782 ^ n3224 ;
  assign n31784 = ~n31752 & n31783 ;
  assign n31749 = n31746 & ~n31748 ;
  assign n31738 = n30258 ^ n29012 ;
  assign n31739 = n29012 ^ n28088 ;
  assign n31740 = ~n31738 & n31739 ;
  assign n31734 = n31704 ^ n31591 ;
  assign n31735 = n31709 & n31734 ;
  assign n31729 = n31591 ^ n28088 ;
  assign n31728 = n30808 ^ n30639 ;
  assign n31730 = n31729 ^ n31728 ;
  assign n31727 = n28226 ^ n28217 ;
  assign n31731 = n31730 ^ n31727 ;
  assign n31732 = n31731 ^ n2705 ;
  assign n31733 = n31732 ^ n3224 ;
  assign n31736 = n31735 ^ n31733 ;
  assign n31724 = n31723 ^ n31710 ;
  assign n31725 = n31723 ^ n28217 ;
  assign n31726 = n31724 & ~n31725 ;
  assign n31737 = n31736 ^ n31726 ;
  assign n31741 = n31740 ^ n31737 ;
  assign n31750 = n31749 ^ n31741 ;
  assign n31785 = n31784 ^ n31750 ;
  assign n31678 = n29951 ^ n29567 ;
  assign n31679 = n30995 ^ n29951 ;
  assign n31680 = n31678 & ~n31679 ;
  assign n31681 = n31680 ^ n29567 ;
  assign n31786 = n31785 ^ n31681 ;
  assign n31791 = n31782 ^ n31752 ;
  assign n31787 = n31001 ^ n29958 ;
  assign n31788 = n29958 ^ n29555 ;
  assign n31789 = ~n31787 & ~n31788 ;
  assign n31790 = n31789 ^ n29555 ;
  assign n31792 = n31791 ^ n31790 ;
  assign n31806 = n31805 ^ n31804 ;
  assign n31813 = n31806 & n31812 ;
  assign n31814 = n31813 ^ n31805 ;
  assign n31815 = n31814 ^ n31790 ;
  assign n31816 = n31792 & n31815 ;
  assign n31817 = n31816 ^ n31791 ;
  assign n31818 = n31817 ^ n31681 ;
  assign n31819 = ~n31786 & n31818 ;
  assign n31820 = n31819 ^ n31785 ;
  assign n31821 = n31820 ^ n31675 ;
  assign n31822 = ~n31677 & ~n31821 ;
  assign n31823 = n31822 ^ n31676 ;
  assign n31825 = n31824 ^ n31823 ;
  assign n31826 = n30982 ^ n30325 ;
  assign n31827 = n31824 ^ n28985 ;
  assign n31828 = n31827 ^ n30982 ;
  assign n31829 = n31828 ^ n31824 ;
  assign n31830 = ~n31826 & ~n31829 ;
  assign n31831 = n31830 ^ n31827 ;
  assign n31832 = n31825 & ~n31831 ;
  assign n31833 = n31832 ^ n31824 ;
  assign n31834 = n31833 ^ n31670 ;
  assign n31835 = ~n31671 & n31834 ;
  assign n31836 = n31835 ^ n30906 ;
  assign n31665 = n31435 ^ n31432 ;
  assign n31661 = n30974 ^ n29939 ;
  assign n31662 = n29939 ^ n28971 ;
  assign n31663 = n31661 & ~n31662 ;
  assign n31664 = n31663 ^ n28971 ;
  assign n31666 = n31665 ^ n31664 ;
  assign n31911 = n31836 ^ n31666 ;
  assign n31876 = n31831 ^ n31823 ;
  assign n31877 = n31876 ^ n29004 ;
  assign n31878 = n31820 ^ n31677 ;
  assign n31879 = n31878 ^ n29092 ;
  assign n31896 = n31817 ^ n31786 ;
  assign n31880 = n31814 ^ n31792 ;
  assign n31881 = n31880 ^ n28844 ;
  assign n31890 = n31889 ^ n31882 ;
  assign n31891 = n31883 & n31890 ;
  assign n31892 = n31891 ^ n28069 ;
  assign n31893 = n31892 ^ n31880 ;
  assign n31894 = n31881 & ~n31893 ;
  assign n31895 = n31894 ^ n28844 ;
  assign n31897 = n31896 ^ n31895 ;
  assign n31898 = n31896 ^ n28945 ;
  assign n31899 = ~n31897 & n31898 ;
  assign n31900 = n31899 ^ n28945 ;
  assign n31901 = n31900 ^ n31878 ;
  assign n31902 = ~n31879 & ~n31901 ;
  assign n31903 = n31902 ^ n29092 ;
  assign n31904 = n31903 ^ n31876 ;
  assign n31905 = n31877 & ~n31904 ;
  assign n31906 = n31905 ^ n29004 ;
  assign n31875 = n31833 ^ n31671 ;
  assign n31907 = n31906 ^ n31875 ;
  assign n31908 = n31906 ^ n28998 ;
  assign n31909 = ~n31907 & n31908 ;
  assign n31910 = n31909 ^ n28998 ;
  assign n31912 = n31911 ^ n31910 ;
  assign n31913 = n31911 ^ n29108 ;
  assign n31914 = n31912 & ~n31913 ;
  assign n31915 = n31914 ^ n29108 ;
  assign n31837 = n31836 ^ n31664 ;
  assign n31838 = n31666 & ~n31837 ;
  assign n31839 = n31838 ^ n31665 ;
  assign n31659 = n31439 ^ n31429 ;
  assign n31655 = n30968 ^ n30348 ;
  assign n31656 = n30348 ^ n28964 ;
  assign n31657 = ~n31655 & ~n31656 ;
  assign n31658 = n31657 ^ n28964 ;
  assign n31660 = n31659 ^ n31658 ;
  assign n31873 = n31839 ^ n31660 ;
  assign n31874 = n31873 ^ n29070 ;
  assign n31974 = n31915 ^ n31874 ;
  assign n31960 = n31913 ^ n31910 ;
  assign n31961 = n31875 ^ n28998 ;
  assign n31962 = n31961 ^ n31906 ;
  assign n31964 = n31892 ^ n31881 ;
  assign n31965 = n31963 & ~n31964 ;
  assign n31966 = n31898 ^ n31895 ;
  assign n31967 = n31965 & ~n31966 ;
  assign n31968 = n31900 ^ n31879 ;
  assign n31969 = ~n31967 & ~n31968 ;
  assign n31970 = n31903 ^ n31877 ;
  assign n31971 = ~n31969 & n31970 ;
  assign n31972 = n31962 & n31971 ;
  assign n31973 = n31960 & ~n31972 ;
  assign n32021 = n31974 ^ n31973 ;
  assign n32025 = n32024 ^ n32021 ;
  assign n32027 = n29795 ^ n2402 ;
  assign n32028 = n32027 ^ n2216 ;
  assign n32029 = n32028 ^ n21174 ;
  assign n32026 = n31972 ^ n31960 ;
  assign n32030 = n32029 ^ n32026 ;
  assign n32034 = n31971 ^ n31962 ;
  assign n32031 = n29800 ^ n2409 ;
  assign n32032 = n32031 ^ n26497 ;
  assign n32033 = n32032 ^ n2211 ;
  assign n32035 = n32034 ^ n32033 ;
  assign n32036 = n31970 ^ n31969 ;
  assign n2082 = n2081 ^ n2036 ;
  assign n2092 = n2091 ^ n2082 ;
  assign n2096 = n2095 ^ n2092 ;
  assign n32037 = n32036 ^ n2096 ;
  assign n32041 = n31968 ^ n31967 ;
  assign n32038 = n29807 ^ n22319 ;
  assign n32039 = n32038 ^ n2014 ;
  assign n32040 = n32039 ^ n2086 ;
  assign n32042 = n32041 ^ n32040 ;
  assign n32043 = n31966 ^ n31965 ;
  assign n1990 = n1983 ^ n1962 ;
  assign n2003 = n2002 ^ n1990 ;
  assign n2007 = n2006 ^ n2003 ;
  assign n32044 = n32043 ^ n2007 ;
  assign n32046 = n3062 ^ n1927 ;
  assign n32047 = n32046 ^ n26112 ;
  assign n32048 = n32047 ^ n1997 ;
  assign n32045 = n31964 ^ n31963 ;
  assign n32049 = n32048 ^ n32045 ;
  assign n32061 = n32060 ^ n32052 ;
  assign n32062 = n32053 & ~n32061 ;
  assign n32063 = n32062 ^ n31963 ;
  assign n32064 = n32063 ^ n32045 ;
  assign n32065 = n32049 & ~n32064 ;
  assign n32066 = n32065 ^ n32048 ;
  assign n32067 = n32066 ^ n2007 ;
  assign n32068 = n32044 & n32067 ;
  assign n32069 = n32068 ^ n2007 ;
  assign n32070 = n32069 ^ n32040 ;
  assign n32071 = n32042 & ~n32070 ;
  assign n32072 = n32071 ^ n32041 ;
  assign n32073 = n32072 ^ n2096 ;
  assign n32074 = n32037 & ~n32073 ;
  assign n32075 = n32074 ^ n32036 ;
  assign n32076 = n32075 ^ n32033 ;
  assign n32077 = ~n32035 & ~n32076 ;
  assign n32078 = n32077 ^ n32034 ;
  assign n32079 = n32078 ^ n32026 ;
  assign n32080 = ~n32030 & ~n32079 ;
  assign n32081 = n32080 ^ n32029 ;
  assign n32082 = n32081 ^ n32021 ;
  assign n32083 = n32025 & ~n32082 ;
  assign n32084 = n32083 ^ n32024 ;
  assign n32017 = n29850 ^ n22373 ;
  assign n32018 = n32017 ^ n26481 ;
  assign n32019 = n32018 ^ n21165 ;
  assign n31916 = n31915 ^ n31873 ;
  assign n31917 = ~n31874 & n31916 ;
  assign n31918 = n31917 ^ n29070 ;
  assign n31840 = n31839 ^ n31658 ;
  assign n31841 = n31660 & n31840 ;
  assign n31842 = n31841 ^ n31659 ;
  assign n31653 = n31442 ^ n31424 ;
  assign n31649 = n30965 ^ n30358 ;
  assign n31650 = n30358 ^ n29593 ;
  assign n31651 = ~n31649 & n31650 ;
  assign n31652 = n31651 ^ n29593 ;
  assign n31654 = n31653 ^ n31652 ;
  assign n31871 = n31842 ^ n31654 ;
  assign n31872 = n31871 ^ n28992 ;
  assign n31976 = n31918 ^ n31872 ;
  assign n31975 = n31973 & n31974 ;
  assign n32016 = n31976 ^ n31975 ;
  assign n32020 = n32019 ^ n32016 ;
  assign n32667 = n32084 ^ n32020 ;
  assign n32234 = n31475 ^ n31391 ;
  assign n32235 = n32234 ^ n30929 ;
  assign n32236 = n32234 ^ n30383 ;
  assign n32237 = n32235 & ~n32236 ;
  assign n32238 = n32237 ^ n30383 ;
  assign n32233 = n32081 ^ n32025 ;
  assign n32239 = n32238 ^ n32233 ;
  assign n32113 = n31396 ^ n31393 ;
  assign n32114 = n32113 ^ n31472 ;
  assign n32241 = n32114 ^ n30935 ;
  assign n32242 = n32114 ^ n29927 ;
  assign n32243 = ~n32241 & ~n32242 ;
  assign n32244 = n32243 ^ n29927 ;
  assign n32240 = n32078 ^ n32030 ;
  assign n32245 = n32244 ^ n32240 ;
  assign n31943 = n31470 ^ n31399 ;
  assign n32247 = n31943 ^ n30945 ;
  assign n32248 = n31943 ^ n29931 ;
  assign n32249 = ~n32247 & ~n32248 ;
  assign n32250 = n32249 ^ n29931 ;
  assign n32246 = n32075 ^ n32035 ;
  assign n32251 = n32250 ^ n32246 ;
  assign n32256 = n32072 ^ n32037 ;
  assign n32252 = n30951 ^ n29937 ;
  assign n31610 = n31461 ^ n31404 ;
  assign n31608 = n31461 ^ n31457 ;
  assign n31609 = n31458 & n31608 ;
  assign n31611 = n31610 ^ n31609 ;
  assign n32253 = n31611 ^ n30951 ;
  assign n32254 = n32252 & ~n32253 ;
  assign n32255 = n32254 ^ n29937 ;
  assign n32257 = n32256 ^ n32255 ;
  assign n31618 = n31608 ^ n31456 ;
  assign n32258 = n31618 ^ n30954 ;
  assign n32259 = n32069 ^ n32042 ;
  assign n32260 = n32259 ^ n30358 ;
  assign n32261 = n32260 ^ n31618 ;
  assign n32262 = n32261 ^ n32259 ;
  assign n32263 = ~n32258 & n32262 ;
  assign n32264 = n32263 ^ n32260 ;
  assign n32266 = n30960 ^ n30348 ;
  assign n31624 = n31409 ^ n2348 ;
  assign n31625 = n31624 ^ n31453 ;
  assign n32267 = n31625 ^ n30960 ;
  assign n32268 = ~n32266 & ~n32267 ;
  assign n32269 = n32268 ^ n30348 ;
  assign n32265 = n32066 ^ n32044 ;
  assign n32270 = n32269 ^ n32265 ;
  assign n32639 = n32063 ^ n32049 ;
  assign n31641 = n31448 ^ n31414 ;
  assign n32271 = n31641 ^ n30968 ;
  assign n32272 = n30968 ^ n30335 ;
  assign n32273 = n32271 & n32272 ;
  assign n32274 = n32273 ^ n30335 ;
  assign n32276 = n32275 ^ n32274 ;
  assign n32626 = n32057 ^ n32055 ;
  assign n32277 = n31653 ^ n30979 ;
  assign n32278 = n30979 ^ n29945 ;
  assign n32279 = n32277 & n32278 ;
  assign n32280 = n32279 ^ n29945 ;
  assign n31587 = n31586 ^ n2782 ;
  assign n32281 = n32280 ^ n31587 ;
  assign n32386 = n31530 ^ n31518 ;
  assign n32387 = n32386 ^ n31522 ;
  assign n32388 = n32387 ^ n31530 ;
  assign n32389 = ~n31524 & ~n32388 ;
  assign n32390 = n32389 ^ n32386 ;
  assign n32381 = n29990 ^ n29021 ;
  assign n32382 = n31074 ^ n29990 ;
  assign n32383 = ~n32381 & n32382 ;
  assign n32384 = n32383 ^ n29021 ;
  assign n32481 = n32390 ^ n32384 ;
  assign n32287 = n30902 ^ n30258 ;
  assign n32288 = n30258 ^ n29489 ;
  assign n32289 = n32287 & ~n32288 ;
  assign n32290 = n32289 ^ n29489 ;
  assign n32286 = n31524 ^ n31518 ;
  assign n32291 = n32290 ^ n32286 ;
  assign n32370 = n30265 ^ n29528 ;
  assign n32371 = n30859 ^ n30265 ;
  assign n32372 = n32370 & ~n32371 ;
  assign n32373 = n32372 ^ n29528 ;
  assign n32292 = n30271 ^ n29497 ;
  assign n32293 = n30811 ^ n30271 ;
  assign n32294 = n32292 & n32293 ;
  assign n32295 = n32294 ^ n29497 ;
  assign n31593 = ~n31368 & ~n31506 ;
  assign n31594 = ~n31481 & n31593 ;
  assign n31595 = n31594 ^ n31506 ;
  assign n31596 = n31488 & n31595 ;
  assign n31597 = n31596 ^ n31486 ;
  assign n32132 = n31597 ^ n1160 ;
  assign n32133 = n32132 ^ n31370 ;
  assign n32296 = n32295 ^ n32133 ;
  assign n32297 = n30278 ^ n29507 ;
  assign n32298 = n31591 ^ n30278 ;
  assign n32299 = n32297 & n32298 ;
  assign n32300 = n32299 ^ n29507 ;
  assign n32140 = n31595 ^ n31374 ;
  assign n32301 = n32300 ^ n32140 ;
  assign n32348 = n31045 ^ n30177 ;
  assign n32349 = n31695 ^ n31045 ;
  assign n32350 = n32348 & n32349 ;
  assign n32351 = n32350 ^ n30177 ;
  assign n32302 = n31537 ^ n30850 ;
  assign n32303 = n30850 ^ n29918 ;
  assign n32304 = ~n32302 & ~n32303 ;
  assign n32305 = n32304 ^ n29918 ;
  assign n32197 = n31493 ^ n31481 ;
  assign n32306 = n32305 ^ n32197 ;
  assign n32311 = n31478 ^ n31386 ;
  assign n32307 = n31286 ^ n30569 ;
  assign n32308 = n30569 ^ n29909 ;
  assign n32309 = ~n32307 & n32308 ;
  assign n32310 = n32309 ^ n29909 ;
  assign n32312 = n32311 ^ n32310 ;
  assign n32112 = n30910 ^ n29902 ;
  assign n32115 = n32114 ^ n29923 ;
  assign n32116 = n32115 ^ n30910 ;
  assign n32117 = n32116 ^ n32114 ;
  assign n32118 = ~n32112 & n32117 ;
  assign n32119 = n32118 ^ n32115 ;
  assign n31942 = n30926 ^ n30398 ;
  assign n31944 = n31943 ^ n29929 ;
  assign n31945 = n31944 ^ n30926 ;
  assign n31946 = n31945 ^ n31943 ;
  assign n31947 = ~n31942 & n31946 ;
  assign n31948 = n31947 ^ n31944 ;
  assign n31607 = n30929 ^ n30399 ;
  assign n31612 = n31611 ^ n30008 ;
  assign n31613 = n31612 ^ n30929 ;
  assign n31614 = n31613 ^ n31611 ;
  assign n31615 = n31607 & ~n31614 ;
  assign n31616 = n31615 ^ n31612 ;
  assign n31617 = n30935 ^ n29911 ;
  assign n31619 = n31618 ^ n30028 ;
  assign n31620 = n31619 ^ n30935 ;
  assign n31621 = n31620 ^ n31618 ;
  assign n31622 = n31617 & ~n31621 ;
  assign n31623 = n31622 ^ n31619 ;
  assign n31626 = n30945 ^ n30383 ;
  assign n31627 = n30383 ^ n30015 ;
  assign n31628 = ~n31626 & n31627 ;
  assign n31629 = n31628 ^ n30015 ;
  assign n31630 = n31629 ^ n31625 ;
  assign n31635 = n31451 ^ n31412 ;
  assign n31631 = n30951 ^ n29927 ;
  assign n31632 = n29927 ^ n29890 ;
  assign n31633 = ~n31631 & ~n31632 ;
  assign n31634 = n31633 ^ n29890 ;
  assign n31636 = n31635 ^ n31634 ;
  assign n31637 = n30954 ^ n29931 ;
  assign n31638 = n29931 ^ n29709 ;
  assign n31639 = ~n31637 & ~n31638 ;
  assign n31640 = n31639 ^ n29709 ;
  assign n31642 = n31641 ^ n31640 ;
  assign n31647 = n31445 ^ n31419 ;
  assign n31643 = n30960 ^ n29937 ;
  assign n31644 = n29937 ^ n29603 ;
  assign n31645 = ~n31643 & ~n31644 ;
  assign n31646 = n31645 ^ n29603 ;
  assign n31648 = n31647 ^ n31646 ;
  assign n31843 = n31842 ^ n31652 ;
  assign n31844 = ~n31654 & ~n31843 ;
  assign n31845 = n31844 ^ n31653 ;
  assign n31846 = n31845 ^ n31646 ;
  assign n31847 = n31648 & ~n31846 ;
  assign n31848 = n31847 ^ n31647 ;
  assign n31849 = n31848 ^ n31640 ;
  assign n31850 = ~n31642 & ~n31849 ;
  assign n31851 = n31850 ^ n31641 ;
  assign n31852 = n31851 ^ n31634 ;
  assign n31853 = ~n31636 & n31852 ;
  assign n31854 = n31853 ^ n31635 ;
  assign n31855 = n31854 ^ n31625 ;
  assign n31856 = ~n31630 & ~n31855 ;
  assign n31857 = n31856 ^ n31629 ;
  assign n31858 = n31857 ^ n31618 ;
  assign n31859 = n31623 & ~n31858 ;
  assign n31860 = n31859 ^ n31618 ;
  assign n31949 = n31860 ^ n31611 ;
  assign n31950 = ~n31616 & n31949 ;
  assign n31951 = n31950 ^ n31860 ;
  assign n32120 = n31951 ^ n31943 ;
  assign n32121 = n31948 & ~n32120 ;
  assign n32122 = n32121 ^ n31943 ;
  assign n32313 = n32122 ^ n32114 ;
  assign n32314 = ~n32119 & n32313 ;
  assign n32315 = n32314 ^ n32114 ;
  assign n32316 = n32315 ^ n32234 ;
  assign n32317 = n31164 ^ n30417 ;
  assign n32318 = n32234 ^ n30053 ;
  assign n32319 = n32318 ^ n32234 ;
  assign n32320 = n32319 ^ n31164 ;
  assign n32321 = ~n32317 & n32320 ;
  assign n32322 = n32321 ^ n32318 ;
  assign n32323 = ~n32316 & n32322 ;
  assign n32324 = n32323 ^ n32234 ;
  assign n32325 = n32324 ^ n32310 ;
  assign n32326 = ~n32312 & n32325 ;
  assign n32327 = n32326 ^ n32311 ;
  assign n32328 = n32327 ^ n32197 ;
  assign n32329 = ~n32306 & n32328 ;
  assign n32330 = n32329 ^ n32305 ;
  assign n32207 = n31481 ^ n1590 ;
  assign n32208 = n31492 ^ n31351 ;
  assign n32209 = n32208 ^ n31492 ;
  assign n32210 = n32209 ^ n31481 ;
  assign n32211 = n32207 & n32210 ;
  assign n32212 = n32211 ^ n32208 ;
  assign n32331 = n32330 ^ n32212 ;
  assign n32332 = n31560 ^ n30890 ;
  assign n32333 = n30890 ^ n30115 ;
  assign n32334 = n32332 & n32333 ;
  assign n32335 = n32334 ^ n30115 ;
  assign n32336 = n32335 ^ n32212 ;
  assign n32337 = ~n32331 & ~n32336 ;
  assign n32338 = n32337 ^ n32335 ;
  assign n32192 = n31362 ^ n877 ;
  assign n32177 = ~n31359 & ~n31481 ;
  assign n32178 = ~n31497 & n32177 ;
  assign n32179 = n32178 ^ n31497 ;
  assign n32193 = n32192 ^ n32179 ;
  assign n32339 = n32338 ^ n32193 ;
  assign n32340 = n31683 ^ n31024 ;
  assign n32341 = n32193 ^ n29904 ;
  assign n32342 = n32341 ^ n31683 ;
  assign n32343 = n32342 ^ n32193 ;
  assign n32344 = n32340 & n32343 ;
  assign n32345 = n32344 ^ n32341 ;
  assign n32346 = ~n32339 & n32345 ;
  assign n32347 = n32346 ^ n32338 ;
  assign n32352 = n32351 ^ n32347 ;
  assign n32180 = n32179 ^ n31362 ;
  assign n32181 = n31491 ^ n877 ;
  assign n32182 = n32181 ^ n31491 ;
  assign n32183 = n32182 ^ n32179 ;
  assign n32184 = n32180 & n32183 ;
  assign n32185 = n32184 ^ n32181 ;
  assign n32353 = n32347 ^ n32185 ;
  assign n32354 = n32352 & n32353 ;
  assign n32355 = n32354 ^ n32351 ;
  assign n32356 = n32355 ^ n32140 ;
  assign n32357 = ~n32301 & n32356 ;
  assign n32358 = n32357 ^ n32355 ;
  assign n32149 = n31595 ^ n31373 ;
  assign n32150 = n31374 & ~n32149 ;
  assign n32148 = n31484 ^ n996 ;
  assign n32151 = n32150 ^ n32148 ;
  assign n32359 = n32358 ^ n32151 ;
  assign n32360 = n30277 ^ n29514 ;
  assign n32361 = n31728 ^ n30277 ;
  assign n32362 = n32360 & n32361 ;
  assign n32363 = n32362 ^ n29514 ;
  assign n32364 = n32363 ^ n32358 ;
  assign n32365 = ~n32359 & ~n32364 ;
  assign n32366 = n32365 ^ n32363 ;
  assign n32367 = n32366 ^ n32133 ;
  assign n32368 = n32296 & ~n32367 ;
  assign n32369 = n32368 ^ n32366 ;
  assign n32374 = n32373 ^ n32369 ;
  assign n31598 = n31597 ^ n31370 ;
  assign n31599 = n31350 ^ n1160 ;
  assign n31600 = n31599 ^ n31350 ;
  assign n31601 = n31600 ^ n31597 ;
  assign n31602 = ~n31598 & n31601 ;
  assign n31603 = n31602 ^ n31599 ;
  assign n32375 = n32369 ^ n31603 ;
  assign n32376 = ~n32374 & ~n32375 ;
  assign n32377 = n32376 ^ n32373 ;
  assign n32378 = n32377 ^ n32286 ;
  assign n32379 = n32291 & n32378 ;
  assign n32380 = n32379 ^ n32290 ;
  assign n32482 = n32481 ^ n32380 ;
  assign n32504 = n32482 ^ n28092 ;
  assign n32394 = n32373 ^ n31603 ;
  assign n32395 = n32394 ^ n32369 ;
  assign n32396 = n32395 ^ n28744 ;
  assign n32397 = n32366 ^ n32296 ;
  assign n32398 = n32397 ^ n28766 ;
  assign n32401 = n32355 ^ n32301 ;
  assign n32402 = n32401 ^ n28754 ;
  assign n32403 = n32351 ^ n32185 ;
  assign n32404 = n32403 ^ n32347 ;
  assign n32405 = n32404 ^ n29359 ;
  assign n32406 = n32345 ^ n32338 ;
  assign n32407 = n32406 ^ n29206 ;
  assign n32409 = n32327 ^ n32306 ;
  assign n32410 = n32409 ^ n29188 ;
  assign n32412 = n32322 ^ n32315 ;
  assign n32413 = n32412 ^ n29039 ;
  assign n32123 = n32122 ^ n32119 ;
  assign n32124 = n32123 ^ n29042 ;
  assign n31952 = n31951 ^ n31948 ;
  assign n31953 = n31952 ^ n29163 ;
  assign n31862 = n31857 ^ n31623 ;
  assign n31863 = n31862 ^ n29154 ;
  assign n31864 = n31854 ^ n31630 ;
  assign n31865 = n31864 ^ n28965 ;
  assign n31867 = n31848 ^ n31642 ;
  assign n31868 = n31867 ^ n28980 ;
  assign n31869 = n31845 ^ n31648 ;
  assign n31870 = n31869 ^ n28986 ;
  assign n31919 = n31918 ^ n31871 ;
  assign n31920 = ~n31872 & n31919 ;
  assign n31921 = n31920 ^ n28992 ;
  assign n31922 = n31921 ^ n31869 ;
  assign n31923 = ~n31870 & n31922 ;
  assign n31924 = n31923 ^ n28986 ;
  assign n31925 = n31924 ^ n31867 ;
  assign n31926 = ~n31868 & ~n31925 ;
  assign n31927 = n31926 ^ n28980 ;
  assign n31866 = n31851 ^ n31636 ;
  assign n31928 = n31927 ^ n31866 ;
  assign n31929 = n31927 ^ n28972 ;
  assign n31930 = ~n31928 & ~n31929 ;
  assign n31931 = n31930 ^ n28972 ;
  assign n31932 = n31931 ^ n31864 ;
  assign n31933 = ~n31865 & n31932 ;
  assign n31934 = n31933 ^ n28965 ;
  assign n31935 = n31934 ^ n31862 ;
  assign n31936 = n31863 & n31935 ;
  assign n31937 = n31936 ^ n29154 ;
  assign n31861 = n31860 ^ n31616 ;
  assign n31938 = n31937 ^ n31861 ;
  assign n31939 = n31937 ^ n29159 ;
  assign n31940 = n31938 & n31939 ;
  assign n31941 = n31940 ^ n29159 ;
  assign n32109 = n31952 ^ n31941 ;
  assign n32110 = ~n31953 & n32109 ;
  assign n32111 = n32110 ^ n29163 ;
  assign n32414 = n32123 ^ n32111 ;
  assign n32415 = ~n32124 & n32414 ;
  assign n32416 = n32415 ^ n29042 ;
  assign n32417 = n32416 ^ n32412 ;
  assign n32418 = n32413 & ~n32417 ;
  assign n32419 = n32418 ^ n29039 ;
  assign n32411 = n32324 ^ n32312 ;
  assign n32420 = n32419 ^ n32411 ;
  assign n32421 = n32419 ^ n29178 ;
  assign n32422 = ~n32420 & ~n32421 ;
  assign n32423 = n32422 ^ n29178 ;
  assign n32424 = n32423 ^ n32409 ;
  assign n32425 = n32410 & n32424 ;
  assign n32426 = n32425 ^ n29188 ;
  assign n32408 = n32336 ^ n32330 ;
  assign n32427 = n32426 ^ n32408 ;
  assign n32428 = n32426 ^ n29029 ;
  assign n32429 = ~n32427 & n32428 ;
  assign n32430 = n32429 ^ n29029 ;
  assign n32431 = n32430 ^ n32406 ;
  assign n32432 = ~n32407 & n32431 ;
  assign n32433 = n32432 ^ n29206 ;
  assign n32434 = n32433 ^ n32404 ;
  assign n32435 = n32405 & n32434 ;
  assign n32436 = n32435 ^ n29359 ;
  assign n32437 = n32436 ^ n32401 ;
  assign n32438 = n32402 & n32437 ;
  assign n32439 = n32438 ^ n28754 ;
  assign n32399 = n32363 ^ n32151 ;
  assign n32400 = n32399 ^ n32358 ;
  assign n32440 = n32439 ^ n32400 ;
  assign n32441 = n32439 ^ n28757 ;
  assign n32442 = n32440 & n32441 ;
  assign n32443 = n32442 ^ n28757 ;
  assign n32444 = n32443 ^ n32397 ;
  assign n32445 = n32398 & ~n32444 ;
  assign n32446 = n32445 ^ n28766 ;
  assign n32447 = n32446 ^ n32395 ;
  assign n32448 = n32396 & ~n32447 ;
  assign n32449 = n32448 ^ n28744 ;
  assign n32393 = n32377 ^ n32291 ;
  assign n32450 = n32449 ^ n32393 ;
  assign n32451 = n32449 ^ n28738 ;
  assign n32452 = ~n32450 & ~n32451 ;
  assign n32453 = n32452 ^ n28738 ;
  assign n32505 = n32504 ^ n32453 ;
  assign n32454 = n32393 ^ n28738 ;
  assign n32455 = n32454 ^ n32449 ;
  assign n32456 = n32436 ^ n32402 ;
  assign n32457 = n32433 ^ n32405 ;
  assign n32458 = n32411 ^ n29178 ;
  assign n32459 = n32458 ^ n32419 ;
  assign n32125 = n32124 ^ n32111 ;
  assign n31954 = n31953 ^ n31941 ;
  assign n31955 = n31861 ^ n29159 ;
  assign n31956 = n31955 ^ n31937 ;
  assign n31957 = n31934 ^ n31863 ;
  assign n31958 = n31866 ^ n28972 ;
  assign n31959 = n31958 ^ n31927 ;
  assign n31977 = ~n31975 & ~n31976 ;
  assign n31978 = n31921 ^ n31870 ;
  assign n31979 = n31977 & ~n31978 ;
  assign n31980 = n31924 ^ n31868 ;
  assign n31981 = n31979 & ~n31980 ;
  assign n31982 = n31959 & n31981 ;
  assign n31983 = n31931 ^ n31865 ;
  assign n31984 = ~n31982 & n31983 ;
  assign n31985 = n31957 & ~n31984 ;
  assign n31986 = n31956 & n31985 ;
  assign n32126 = n31954 & n31986 ;
  assign n32460 = ~n32125 & ~n32126 ;
  assign n32461 = n32416 ^ n32413 ;
  assign n32462 = ~n32460 & ~n32461 ;
  assign n32463 = n32459 & n32462 ;
  assign n32464 = n32423 ^ n32410 ;
  assign n32465 = ~n32463 & ~n32464 ;
  assign n32466 = n32408 ^ n29029 ;
  assign n32467 = n32466 ^ n32426 ;
  assign n32468 = n32465 & n32467 ;
  assign n32469 = n32430 ^ n32407 ;
  assign n32470 = n32468 & ~n32469 ;
  assign n32471 = ~n32457 & ~n32470 ;
  assign n32472 = n32456 & n32471 ;
  assign n32473 = n32400 ^ n28757 ;
  assign n32474 = n32473 ^ n32439 ;
  assign n32475 = n32472 & n32474 ;
  assign n32476 = n32443 ^ n32398 ;
  assign n32477 = n32475 & ~n32476 ;
  assign n32478 = n32446 ^ n32396 ;
  assign n32479 = ~n32477 & n32478 ;
  assign n32480 = ~n32455 & n32479 ;
  assign n32506 = n32505 ^ n32480 ;
  assign n32499 = n30193 ^ n2675 ;
  assign n32500 = n32499 ^ n26755 ;
  assign n32501 = n32500 ^ n1841 ;
  assign n32507 = n32506 ^ n32501 ;
  assign n32508 = n32479 ^ n32455 ;
  assign n3129 = n3128 ^ n2669 ;
  assign n3139 = n3138 ^ n3129 ;
  assign n3143 = n3142 ^ n3139 ;
  assign n32509 = n32508 ^ n3143 ;
  assign n32513 = n32478 ^ n32477 ;
  assign n32510 = n30200 ^ n22733 ;
  assign n32511 = n32510 ^ n26581 ;
  assign n32512 = n32511 ^ n3135 ;
  assign n32514 = n32513 ^ n32512 ;
  assign n32515 = n32476 ^ n32475 ;
  assign n32519 = n32518 ^ n32515 ;
  assign n32521 = n30211 ^ n22741 ;
  assign n32522 = n32521 ^ n2645 ;
  assign n32523 = n32522 ^ n3209 ;
  assign n32520 = n32474 ^ n32472 ;
  assign n32524 = n32523 ^ n32520 ;
  assign n32528 = n32471 ^ n32456 ;
  assign n32525 = n30215 ^ n22748 ;
  assign n32526 = n32525 ^ n26450 ;
  assign n32527 = n32526 ^ n2546 ;
  assign n32529 = n32528 ^ n32527 ;
  assign n32530 = n32470 ^ n32457 ;
  assign n32534 = n32533 ^ n32530 ;
  assign n32535 = n32469 ^ n32468 ;
  assign n1280 = n1241 ^ n1183 ;
  assign n1281 = n1280 ^ n1277 ;
  assign n1285 = n1284 ^ n1281 ;
  assign n32536 = n32535 ^ n1285 ;
  assign n32537 = n32467 ^ n32465 ;
  assign n32538 = n32537 ^ n1270 ;
  assign n32539 = n32464 ^ n32463 ;
  assign n1119 = n1082 ^ n1037 ;
  assign n1120 = n1119 ^ n1103 ;
  assign n1124 = n1123 ^ n1120 ;
  assign n32540 = n32539 ^ n1124 ;
  assign n32541 = n32462 ^ n32459 ;
  assign n32542 = n32541 ^ n1116 ;
  assign n32543 = n32461 ^ n32460 ;
  assign n32544 = n32543 ^ n1657 ;
  assign n32127 = n32126 ^ n32125 ;
  assign n32128 = n32127 ^ n1648 ;
  assign n31987 = n31986 ^ n31954 ;
  assign n31988 = n31987 ^ n2987 ;
  assign n31992 = n31985 ^ n31956 ;
  assign n31993 = n31992 ^ n31991 ;
  assign n31994 = n31984 ^ n31957 ;
  assign n31995 = n31994 ^ n638 ;
  assign n31999 = n31983 ^ n31982 ;
  assign n32000 = n31999 ^ n31998 ;
  assign n32004 = n31981 ^ n31959 ;
  assign n32005 = n32004 ^ n32003 ;
  assign n32009 = n31980 ^ n31979 ;
  assign n32010 = n32009 ^ n32008 ;
  assign n32012 = n29786 ^ n1475 ;
  assign n32013 = n32012 ^ n26472 ;
  assign n32014 = n32013 ^ n21159 ;
  assign n32011 = n31978 ^ n31977 ;
  assign n32015 = n32014 ^ n32011 ;
  assign n32085 = n32084 ^ n32016 ;
  assign n32086 = ~n32020 & n32085 ;
  assign n32087 = n32086 ^ n32019 ;
  assign n32088 = n32087 ^ n32011 ;
  assign n32089 = n32015 & ~n32088 ;
  assign n32090 = n32089 ^ n32014 ;
  assign n32091 = n32090 ^ n32008 ;
  assign n32092 = n32010 & ~n32091 ;
  assign n32093 = n32092 ^ n32009 ;
  assign n32094 = n32093 ^ n32003 ;
  assign n32095 = ~n32005 & ~n32094 ;
  assign n32096 = n32095 ^ n32004 ;
  assign n32097 = n32096 ^ n31998 ;
  assign n32098 = ~n32000 & n32097 ;
  assign n32099 = n32098 ^ n31999 ;
  assign n32100 = n32099 ^ n638 ;
  assign n32101 = n31995 & n32100 ;
  assign n32102 = n32101 ^ n31994 ;
  assign n32103 = n32102 ^ n31991 ;
  assign n32104 = ~n31993 & ~n32103 ;
  assign n32105 = n32104 ^ n31992 ;
  assign n32106 = n32105 ^ n2987 ;
  assign n32107 = ~n31988 & n32106 ;
  assign n32108 = n32107 ^ n31987 ;
  assign n32545 = n32127 ^ n32108 ;
  assign n32546 = n32128 & n32545 ;
  assign n32547 = n32546 ^ n1648 ;
  assign n32548 = n32547 ^ n1657 ;
  assign n32549 = ~n32544 & ~n32548 ;
  assign n32550 = n32549 ^ n32543 ;
  assign n32551 = n32550 ^ n1116 ;
  assign n32552 = ~n32542 & n32551 ;
  assign n32553 = n32552 ^ n32541 ;
  assign n32554 = n32553 ^ n1124 ;
  assign n32555 = n32540 & n32554 ;
  assign n32556 = n32555 ^ n32539 ;
  assign n32557 = n32556 ^ n1270 ;
  assign n32558 = n32538 & ~n32557 ;
  assign n32559 = n32558 ^ n32537 ;
  assign n32560 = n32559 ^ n1285 ;
  assign n32561 = ~n32536 & ~n32560 ;
  assign n32562 = n32561 ^ n32535 ;
  assign n32563 = n32562 ^ n32530 ;
  assign n32564 = ~n32534 & ~n32563 ;
  assign n32565 = n32564 ^ n32533 ;
  assign n32566 = n32565 ^ n32527 ;
  assign n32567 = ~n32529 & ~n32566 ;
  assign n32568 = n32567 ^ n32528 ;
  assign n32569 = n32568 ^ n32520 ;
  assign n32570 = ~n32524 & ~n32569 ;
  assign n32571 = n32570 ^ n32523 ;
  assign n32572 = n32571 ^ n32515 ;
  assign n32573 = n32519 & ~n32572 ;
  assign n32574 = n32573 ^ n32518 ;
  assign n32575 = n32574 ^ n32512 ;
  assign n32576 = ~n32514 & ~n32575 ;
  assign n32577 = n32576 ^ n32513 ;
  assign n32578 = n32577 ^ n3143 ;
  assign n32579 = ~n32509 & n32578 ;
  assign n32580 = n32579 ^ n32508 ;
  assign n32581 = n32580 ^ n32501 ;
  assign n32582 = n32507 & ~n32581 ;
  assign n32494 = n31553 ^ n31535 ;
  assign n32492 = n32384 ^ n28088 ;
  assign n32493 = n32492 ^ n29012 ;
  assign n32495 = n32494 ^ n32493 ;
  assign n2769 = n2748 ^ n2719 ;
  assign n2773 = n2772 ^ n2769 ;
  assign n2774 = n2773 ^ n2765 ;
  assign n32496 = n32495 ^ n2774 ;
  assign n32489 = n31071 ^ n29987 ;
  assign n32490 = n29987 ^ n29012 ;
  assign n32491 = n32489 & ~n32490 ;
  assign n32497 = n32496 ^ n32491 ;
  assign n32483 = n32482 ^ n32480 ;
  assign n32486 = n32480 ^ n32453 ;
  assign n32487 = ~n32483 & n32486 ;
  assign n32484 = n32483 ^ n32453 ;
  assign n32485 = n28092 & ~n32484 ;
  assign n32488 = n32487 ^ n32485 ;
  assign n32498 = n32497 ^ n32488 ;
  assign n32502 = n32501 ^ n32498 ;
  assign n32385 = n32384 ^ n32380 ;
  assign n32391 = n32390 ^ n32380 ;
  assign n32392 = ~n32385 & ~n32391 ;
  assign n32503 = n32502 ^ n32392 ;
  assign n32583 = n32582 ^ n32503 ;
  assign n32282 = n31659 ^ n30982 ;
  assign n32283 = n30982 ^ n29951 ;
  assign n32284 = n32282 & n32283 ;
  assign n32285 = n32284 ^ n29951 ;
  assign n32584 = n32583 ^ n32285 ;
  assign n32589 = n32580 ^ n32507 ;
  assign n32585 = n30988 ^ n29958 ;
  assign n32586 = n31665 ^ n30988 ;
  assign n32587 = n32585 & ~n32586 ;
  assign n32588 = n32587 ^ n29958 ;
  assign n32590 = n32589 ^ n32588 ;
  assign n32593 = n32571 ^ n32519 ;
  assign n32594 = n30907 ^ n29981 ;
  assign n32595 = n31676 ^ n29981 ;
  assign n32596 = ~n32594 & ~n32595 ;
  assign n32597 = n32596 ^ n30907 ;
  assign n32598 = n32593 & ~n32597 ;
  assign n32592 = n32574 ^ n32514 ;
  assign n32599 = n32598 ^ n32592 ;
  assign n32600 = n31824 ^ n31001 ;
  assign n32601 = n32598 ^ n29974 ;
  assign n32602 = n32601 ^ n31824 ;
  assign n32603 = n32602 ^ n32598 ;
  assign n32604 = ~n32600 & ~n32603 ;
  assign n32605 = n32604 ^ n32601 ;
  assign n32606 = ~n32599 & ~n32605 ;
  assign n32607 = n32606 ^ n32598 ;
  assign n32591 = n32577 ^ n32509 ;
  assign n32608 = n32607 ^ n32591 ;
  assign n32609 = n30995 ^ n30906 ;
  assign n32610 = n32591 ^ n29968 ;
  assign n32611 = n32610 ^ n30906 ;
  assign n32612 = n32611 ^ n32591 ;
  assign n32613 = ~n32609 & ~n32612 ;
  assign n32614 = n32613 ^ n32610 ;
  assign n32615 = n32608 & n32614 ;
  assign n32616 = n32615 ^ n32607 ;
  assign n32617 = n32616 ^ n32588 ;
  assign n32618 = ~n32590 & ~n32617 ;
  assign n32619 = n32618 ^ n32589 ;
  assign n32620 = n32619 ^ n32285 ;
  assign n32621 = n32584 & n32620 ;
  assign n32622 = n32621 ^ n32583 ;
  assign n32623 = n32622 ^ n32280 ;
  assign n32624 = n32281 & n32623 ;
  assign n32625 = n32624 ^ n31587 ;
  assign n32627 = n32626 ^ n32625 ;
  assign n32628 = n31647 ^ n30974 ;
  assign n32629 = n32626 ^ n30325 ;
  assign n32630 = n32629 ^ n31647 ;
  assign n32631 = n32630 ^ n32626 ;
  assign n32632 = ~n32628 & n32631 ;
  assign n32633 = n32632 ^ n32629 ;
  assign n32634 = ~n32627 & n32633 ;
  assign n32635 = n32634 ^ n32626 ;
  assign n32636 = n32635 ^ n32274 ;
  assign n32637 = n32276 & ~n32636 ;
  assign n32638 = n32637 ^ n32275 ;
  assign n32640 = n32639 ^ n32638 ;
  assign n32641 = n31635 ^ n30965 ;
  assign n32642 = n32639 ^ n29939 ;
  assign n32643 = n32642 ^ n31635 ;
  assign n32644 = n32643 ^ n32639 ;
  assign n32645 = ~n32641 & n32644 ;
  assign n32646 = n32645 ^ n32642 ;
  assign n32647 = n32640 & ~n32646 ;
  assign n32648 = n32647 ^ n32639 ;
  assign n32649 = n32648 ^ n32265 ;
  assign n32650 = n32270 & ~n32649 ;
  assign n32651 = n32650 ^ n32269 ;
  assign n32652 = n32651 ^ n32259 ;
  assign n32653 = ~n32264 & n32652 ;
  assign n32654 = n32653 ^ n32259 ;
  assign n32655 = n32654 ^ n32255 ;
  assign n32656 = ~n32257 & n32655 ;
  assign n32657 = n32656 ^ n32256 ;
  assign n32658 = n32657 ^ n32246 ;
  assign n32659 = n32251 & n32658 ;
  assign n32660 = n32659 ^ n32250 ;
  assign n32661 = n32660 ^ n32240 ;
  assign n32662 = ~n32245 & n32661 ;
  assign n32663 = n32662 ^ n32244 ;
  assign n32664 = n32663 ^ n32233 ;
  assign n32665 = n32239 & n32664 ;
  assign n32666 = n32665 ^ n32238 ;
  assign n32668 = n32667 ^ n32666 ;
  assign n32669 = n32311 ^ n30926 ;
  assign n32670 = n32667 ^ n29911 ;
  assign n32671 = n32670 ^ n30926 ;
  assign n32672 = n32671 ^ n32667 ;
  assign n32673 = n32669 & ~n32672 ;
  assign n32674 = n32673 ^ n32670 ;
  assign n32675 = ~n32668 & n32674 ;
  assign n32676 = n32675 ^ n32667 ;
  assign n32202 = n32087 ^ n32015 ;
  assign n32198 = n32197 ^ n30910 ;
  assign n32199 = n32197 ^ n30399 ;
  assign n32200 = n32198 & ~n32199 ;
  assign n32201 = n32200 ^ n30399 ;
  assign n32228 = n32202 ^ n32201 ;
  assign n32800 = n32676 ^ n32228 ;
  assign n32802 = n32800 ^ n30008 ;
  assign n32801 = ~n30008 & n32800 ;
  assign n32803 = n32802 ^ n32801 ;
  assign n32804 = ~n29929 & ~n32803 ;
  assign n32805 = n32676 ^ n32202 ;
  assign n32204 = n32090 ^ n32010 ;
  assign n32806 = n32204 ^ n32201 ;
  assign n32206 = n31164 ^ n30398 ;
  assign n32213 = n32212 ^ n31164 ;
  assign n32214 = ~n32206 & ~n32213 ;
  assign n32215 = n32214 ^ n30398 ;
  assign n32807 = n32806 ^ n32215 ;
  assign n32808 = n32807 ^ n32204 ;
  assign n32809 = n32808 ^ n32676 ;
  assign n32810 = n32809 ^ n32215 ;
  assign n32811 = n32805 & n32810 ;
  assign n32812 = n32811 ^ n32807 ;
  assign n32813 = n32804 & n32812 ;
  assign n32814 = n32813 ^ n32803 ;
  assign n32718 = n32674 ^ n32666 ;
  assign n32719 = n32718 ^ n30028 ;
  assign n32720 = n32663 ^ n32239 ;
  assign n32721 = n32720 ^ n30015 ;
  assign n32722 = n32660 ^ n32245 ;
  assign n32723 = n32722 ^ n29890 ;
  assign n32724 = n32657 ^ n32251 ;
  assign n32725 = n32724 ^ n29709 ;
  assign n32726 = n32654 ^ n32257 ;
  assign n32727 = n32726 ^ n29603 ;
  assign n32728 = n32651 ^ n32264 ;
  assign n32729 = n32728 ^ n29593 ;
  assign n32730 = n32648 ^ n32270 ;
  assign n32731 = n32730 ^ n28964 ;
  assign n32732 = n32646 ^ n32638 ;
  assign n32733 = n32732 ^ n28971 ;
  assign n32734 = n32635 ^ n32276 ;
  assign n32735 = n32734 ^ n28978 ;
  assign n32763 = n32633 ^ n32625 ;
  assign n32736 = n32622 ^ n32281 ;
  assign n32737 = n32736 ^ n29577 ;
  assign n32738 = n32619 ^ n32584 ;
  assign n32739 = n32738 ^ n29567 ;
  assign n32752 = n32616 ^ n32590 ;
  assign n32741 = n32597 ^ n32593 ;
  assign n32742 = ~n29018 & ~n32741 ;
  assign n32743 = n32742 ^ n29009 ;
  assign n32744 = n32605 ^ n32592 ;
  assign n32745 = n32744 ^ n32742 ;
  assign n32746 = ~n32743 & ~n32745 ;
  assign n32747 = n32746 ^ n29009 ;
  assign n32740 = n32614 ^ n32607 ;
  assign n32748 = n32747 ^ n32740 ;
  assign n32749 = n32747 ^ n28997 ;
  assign n32750 = ~n32748 & ~n32749 ;
  assign n32751 = n32750 ^ n28997 ;
  assign n32753 = n32752 ^ n32751 ;
  assign n32754 = n32752 ^ n29555 ;
  assign n32755 = n32753 & n32754 ;
  assign n32756 = n32755 ^ n29555 ;
  assign n32757 = n32756 ^ n32738 ;
  assign n32758 = ~n32739 & ~n32757 ;
  assign n32759 = n32758 ^ n29567 ;
  assign n32760 = n32759 ^ n32736 ;
  assign n32761 = ~n32737 & ~n32760 ;
  assign n32762 = n32761 ^ n29577 ;
  assign n32764 = n32763 ^ n32762 ;
  assign n32765 = n32763 ^ n28985 ;
  assign n32766 = ~n32764 & n32765 ;
  assign n32767 = n32766 ^ n28985 ;
  assign n32768 = n32767 ^ n32734 ;
  assign n32769 = ~n32735 & n32768 ;
  assign n32770 = n32769 ^ n28978 ;
  assign n32771 = n32770 ^ n32732 ;
  assign n32772 = ~n32733 & ~n32771 ;
  assign n32773 = n32772 ^ n28971 ;
  assign n32774 = n32773 ^ n32730 ;
  assign n32775 = ~n32731 & ~n32774 ;
  assign n32776 = n32775 ^ n28964 ;
  assign n32777 = n32776 ^ n32728 ;
  assign n32778 = n32729 & ~n32777 ;
  assign n32779 = n32778 ^ n29593 ;
  assign n32780 = n32779 ^ n32726 ;
  assign n32781 = ~n32727 & ~n32780 ;
  assign n32782 = n32781 ^ n29603 ;
  assign n32783 = n32782 ^ n32724 ;
  assign n32784 = n32725 & ~n32783 ;
  assign n32785 = n32784 ^ n29709 ;
  assign n32786 = n32785 ^ n32722 ;
  assign n32787 = n32723 & ~n32786 ;
  assign n32788 = n32787 ^ n29890 ;
  assign n32789 = n32788 ^ n32720 ;
  assign n32790 = ~n32721 & n32789 ;
  assign n32791 = n32790 ^ n30015 ;
  assign n32792 = n32791 ^ n32718 ;
  assign n32793 = ~n32719 & ~n32792 ;
  assign n32794 = n32793 ^ n30028 ;
  assign n32827 = n32801 ^ n29929 ;
  assign n32828 = n32812 ^ n32801 ;
  assign n32829 = n32827 & n32828 ;
  assign n32830 = n32829 ^ n29929 ;
  assign n32868 = ~n32794 & ~n32830 ;
  assign n32869 = ~n32814 & n32868 ;
  assign n32870 = n32869 ^ n32830 ;
  assign n32220 = n32093 ^ n32005 ;
  assign n32191 = n31286 ^ n29902 ;
  assign n32194 = n32193 ^ n31286 ;
  assign n32195 = ~n32191 & n32194 ;
  assign n32196 = n32195 ^ n29902 ;
  assign n32797 = n32220 ^ n32196 ;
  assign n32203 = ~n32201 & n32202 ;
  assign n32205 = n32204 ^ n32203 ;
  assign n32216 = n32215 ^ n32203 ;
  assign n32217 = n32205 & ~n32216 ;
  assign n32218 = n32217 ^ n32204 ;
  assign n32229 = n32228 ^ n32203 ;
  assign n32230 = ~n32204 & ~n32229 ;
  assign n32231 = ~n32215 & n32230 ;
  assign n32232 = n32231 ^ n32229 ;
  assign n32677 = ~n32232 & ~n32676 ;
  assign n32795 = ~n32218 & n32677 ;
  assign n32796 = n32795 ^ n32218 ;
  assign n32798 = n32797 ^ n32796 ;
  assign n32799 = n32798 ^ n29923 ;
  assign n32871 = n32870 ^ n32799 ;
  assign n32879 = n32800 ^ n32794 ;
  assign n32880 = n30008 ^ n29929 ;
  assign n32881 = n32880 ^ n32812 ;
  assign n32882 = n32881 ^ n29929 ;
  assign n32883 = n32882 ^ n32794 ;
  assign n32884 = n32883 ^ n32812 ;
  assign n32885 = n32879 & n32884 ;
  assign n32886 = n32885 ^ n32881 ;
  assign n32867 = n32802 ^ n32794 ;
  assign n32893 = n32767 ^ n32735 ;
  assign n32894 = n32765 ^ n32762 ;
  assign n32895 = n32740 ^ n28997 ;
  assign n32896 = n32895 ^ n32747 ;
  assign n32897 = n32754 ^ n32751 ;
  assign n32898 = ~n32896 & ~n32897 ;
  assign n32899 = n32756 ^ n32739 ;
  assign n32900 = n32898 & ~n32899 ;
  assign n32901 = n32759 ^ n32737 ;
  assign n32902 = ~n32900 & ~n32901 ;
  assign n32903 = n32894 & ~n32902 ;
  assign n32904 = ~n32893 & n32903 ;
  assign n32905 = n32770 ^ n32733 ;
  assign n32906 = ~n32904 & n32905 ;
  assign n32907 = n32773 ^ n32731 ;
  assign n32908 = n32906 & ~n32907 ;
  assign n32909 = n32776 ^ n32729 ;
  assign n32910 = ~n32908 & n32909 ;
  assign n32911 = n32779 ^ n32727 ;
  assign n32912 = n32910 & ~n32911 ;
  assign n32913 = n32782 ^ n32725 ;
  assign n32914 = n32912 & ~n32913 ;
  assign n32915 = n32785 ^ n32723 ;
  assign n32916 = n32914 & ~n32915 ;
  assign n32917 = n32788 ^ n32721 ;
  assign n32918 = ~n32916 & ~n32917 ;
  assign n32919 = n32791 ^ n32719 ;
  assign n32920 = ~n32918 & n32919 ;
  assign n33011 = ~n32867 & n32920 ;
  assign n33012 = ~n32886 & n33011 ;
  assign n33013 = ~n32871 & ~n33012 ;
  assign n32872 = n32870 ^ n32798 ;
  assign n32815 = n32796 ^ n32196 ;
  assign n32189 = n32096 ^ n32000 ;
  assign n32816 = n32220 ^ n32189 ;
  assign n32176 = n31537 ^ n30417 ;
  assign n32186 = n32185 ^ n31537 ;
  assign n32187 = ~n32176 & n32186 ;
  assign n32188 = n32187 ^ n30417 ;
  assign n32817 = n32816 ^ n32188 ;
  assign n32818 = n32817 ^ n32189 ;
  assign n32819 = n32818 ^ n32196 ;
  assign n32820 = n32819 ^ n32188 ;
  assign n32821 = n32815 & n32820 ;
  assign n32822 = n32821 ^ n32817 ;
  assign n32823 = n32822 ^ n30053 ;
  assign n32873 = n32823 ^ n29923 ;
  assign n32874 = n32873 ^ n32823 ;
  assign n32875 = n32874 ^ n32870 ;
  assign n32876 = ~n32872 & ~n32875 ;
  assign n32877 = n32876 ^ n32873 ;
  assign n33047 = n33013 ^ n32877 ;
  assign n33048 = n33012 ^ n32871 ;
  assign n33049 = n2992 ^ n1664 ;
  assign n33050 = n33049 ^ n769 ;
  assign n33051 = n33050 ^ n847 ;
  assign n33052 = n32920 ^ n32867 ;
  assign n33057 = n33052 & n33055 ;
  assign n33056 = n33055 ^ n33052 ;
  assign n33058 = n33057 ^ n33056 ;
  assign n33059 = n33011 ^ n32886 ;
  assign n33060 = ~n762 & ~n33059 ;
  assign n33061 = n33058 & n33060 ;
  assign n33062 = n33061 ^ n33058 ;
  assign n33063 = ~n33051 & n33062 ;
  assign n33064 = ~n33048 & n33063 ;
  assign n843 = n842 ^ n791 ;
  assign n853 = n852 ^ n843 ;
  assign n857 = n856 ^ n853 ;
  assign n33065 = n33064 ^ n857 ;
  assign n33066 = n33047 & ~n33065 ;
  assign n33082 = n33064 ^ n33062 ;
  assign n33067 = n33047 ^ n857 ;
  assign n33069 = n33057 ^ n762 ;
  assign n33070 = n33059 ^ n33057 ;
  assign n33071 = n33069 & ~n33070 ;
  assign n33072 = n33071 ^ n762 ;
  assign n33068 = n33051 ^ n33047 ;
  assign n33073 = n33072 ^ n33068 ;
  assign n33074 = n33073 ^ n33048 ;
  assign n33075 = n33074 ^ n33068 ;
  assign n33076 = n33072 ^ n857 ;
  assign n33077 = n33076 ^ n33068 ;
  assign n33078 = ~n33075 & n33077 ;
  assign n33079 = n33078 ^ n33068 ;
  assign n33080 = ~n33067 & ~n33079 ;
  assign n33081 = n33080 ^ n33047 ;
  assign n33083 = n32919 ^ n32918 ;
  assign n33084 = n33083 ^ n1553 ;
  assign n33088 = n32917 ^ n32916 ;
  assign n33089 = n33088 ^ n33087 ;
  assign n33093 = n32915 ^ n32914 ;
  assign n33090 = n27201 ^ n1512 ;
  assign n33091 = n33090 ^ n30674 ;
  assign n33092 = n33091 ^ n2942 ;
  assign n33094 = n33093 ^ n33092 ;
  assign n33098 = n32913 ^ n32912 ;
  assign n33095 = n30679 ^ n23072 ;
  assign n33096 = n33095 ^ n2930 ;
  assign n33097 = n33096 ^ n21772 ;
  assign n33099 = n33098 ^ n33097 ;
  assign n33100 = n32911 ^ n32910 ;
  assign n33104 = n33103 ^ n33100 ;
  assign n33108 = n32909 ^ n32908 ;
  assign n33105 = n2915 ^ n2378 ;
  assign n33106 = n33105 ^ n27212 ;
  assign n33107 = n33106 ^ n21779 ;
  assign n33109 = n33108 ^ n33107 ;
  assign n33113 = n32907 ^ n32906 ;
  assign n33110 = n30695 ^ n23080 ;
  assign n33111 = n33110 ^ n2314 ;
  assign n33112 = n33111 ^ n21785 ;
  assign n33114 = n33113 ^ n33112 ;
  assign n33115 = n32905 ^ n32904 ;
  assign n2299 = n2292 ^ n2229 ;
  assign n2306 = n2305 ^ n2299 ;
  assign n2310 = n2309 ^ n2306 ;
  assign n33116 = n33115 ^ n2310 ;
  assign n33117 = n32903 ^ n32893 ;
  assign n2195 = n2164 ^ n2131 ;
  assign n2196 = n2195 ^ n2192 ;
  assign n2200 = n2199 ^ n2196 ;
  assign n33118 = n33117 ^ n2200 ;
  assign n33119 = n32902 ^ n32894 ;
  assign n2168 = n2155 ^ n2116 ;
  assign n2181 = n2180 ^ n2168 ;
  assign n2185 = n2184 ^ n2181 ;
  assign n33120 = n33119 ^ n2185 ;
  assign n33122 = n30705 ^ n2063 ;
  assign n33123 = n33122 ^ n27222 ;
  assign n33124 = n33123 ^ n2177 ;
  assign n33121 = n32901 ^ n32900 ;
  assign n33125 = n33124 ^ n33121 ;
  assign n33129 = n32899 ^ n32898 ;
  assign n33126 = n30709 ^ n2051 ;
  assign n33127 = n33126 ^ n27226 ;
  assign n33128 = n33127 ^ n21801 ;
  assign n33130 = n33129 ^ n33128 ;
  assign n33132 = n30714 ^ n23096 ;
  assign n33133 = n33132 ^ n27240 ;
  assign n33134 = n33133 ^ n21805 ;
  assign n33131 = n32897 ^ n32896 ;
  assign n33135 = n33134 ^ n33131 ;
  assign n33136 = n30718 ^ n3080 ;
  assign n33137 = n33136 ^ n27230 ;
  assign n33138 = n33137 ^ n1877 ;
  assign n33139 = n33138 ^ n32896 ;
  assign n33145 = n30721 ^ n3074 ;
  assign n33146 = n33145 ^ n1850 ;
  assign n33147 = n33146 ^ n21810 ;
  assign n33140 = n31059 ^ n3183 ;
  assign n33141 = n33140 ^ n23528 ;
  assign n33142 = n33141 ^ n1826 ;
  assign n33143 = n32741 ^ n29018 ;
  assign n33144 = n33142 & n33143 ;
  assign n33148 = n33147 ^ n33144 ;
  assign n33149 = n32744 ^ n32743 ;
  assign n33150 = n33149 ^ n33144 ;
  assign n33151 = n33148 & n33150 ;
  assign n33152 = n33151 ^ n33147 ;
  assign n33153 = n33152 ^ n32896 ;
  assign n33154 = ~n33139 & n33153 ;
  assign n33155 = n33154 ^ n33138 ;
  assign n33156 = n33155 ^ n33134 ;
  assign n33157 = ~n33135 & n33156 ;
  assign n33158 = n33157 ^ n33134 ;
  assign n33159 = n33158 ^ n33128 ;
  assign n33160 = n33130 & n33159 ;
  assign n33161 = n33160 ^ n33128 ;
  assign n33162 = n33161 ^ n33121 ;
  assign n33163 = n33125 & ~n33162 ;
  assign n33164 = n33163 ^ n33124 ;
  assign n33165 = n33164 ^ n33119 ;
  assign n33166 = n33120 & ~n33165 ;
  assign n33167 = n33166 ^ n2185 ;
  assign n33168 = n33167 ^ n2200 ;
  assign n33169 = n33118 & ~n33168 ;
  assign n33170 = n33169 ^ n33117 ;
  assign n33171 = n33170 ^ n2310 ;
  assign n33172 = ~n33116 & ~n33171 ;
  assign n33173 = n33172 ^ n33115 ;
  assign n33174 = n33173 ^ n33112 ;
  assign n33175 = ~n33114 & n33174 ;
  assign n33176 = n33175 ^ n33113 ;
  assign n33177 = n33176 ^ n33107 ;
  assign n33178 = n33109 & n33177 ;
  assign n33179 = n33178 ^ n33108 ;
  assign n33180 = n33179 ^ n33100 ;
  assign n33181 = n33104 & ~n33180 ;
  assign n33182 = n33181 ^ n33103 ;
  assign n33183 = n33182 ^ n33097 ;
  assign n33184 = n33099 & ~n33183 ;
  assign n33185 = n33184 ^ n33098 ;
  assign n33186 = n33185 ^ n33092 ;
  assign n33187 = n33094 & ~n33186 ;
  assign n33188 = n33187 ^ n33093 ;
  assign n33189 = n33188 ^ n33087 ;
  assign n33190 = n33089 & ~n33189 ;
  assign n33191 = n33190 ^ n33088 ;
  assign n33192 = n33191 ^ n1553 ;
  assign n33193 = n33084 & ~n33192 ;
  assign n33194 = n33193 ^ n33083 ;
  assign n33195 = n33081 & n33194 ;
  assign n33196 = n33082 & n33195 ;
  assign n33199 = n33066 & n33196 ;
  assign n33197 = n33196 ^ n33081 ;
  assign n33200 = n33199 ^ n33197 ;
  assign n33014 = ~n32877 & ~n33013 ;
  assign n32219 = n32218 ^ n32196 ;
  assign n32221 = n32220 ^ n32188 ;
  assign n32222 = n32221 ^ n32196 ;
  assign n32223 = n32222 ^ n32188 ;
  assign n32224 = n32219 & n32223 ;
  assign n32225 = n32224 ^ n32221 ;
  assign n32227 = n32225 ^ n32188 ;
  assign n32190 = n32189 ^ n32188 ;
  assign n32678 = ~n32190 & n32677 ;
  assign n32679 = n32227 & n32678 ;
  assign n32680 = n32220 & n32679 ;
  assign n32681 = n32232 ^ n32196 ;
  assign n32682 = n32680 & n32681 ;
  assign n32683 = n32682 ^ n32679 ;
  assign n32684 = n32683 ^ n32189 ;
  assign n32226 = ~n32190 & ~n32225 ;
  assign n32685 = n32684 ^ n32226 ;
  assign n32139 = n31560 ^ n30569 ;
  assign n32141 = n32140 ^ n31560 ;
  assign n32142 = ~n32139 & n32141 ;
  assign n32143 = n32142 ^ n30569 ;
  assign n32138 = n32099 ^ n31995 ;
  assign n32169 = n32143 ^ n32138 ;
  assign n32841 = n32685 ^ n32169 ;
  assign n32843 = n32841 ^ n29909 ;
  assign n32824 = ~n32814 & ~n32823 ;
  assign n32825 = ~n32799 & n32824 ;
  assign n32826 = ~n32794 & n32825 ;
  assign n32832 = n32822 ^ n29923 ;
  assign n32831 = n32830 ^ n32822 ;
  assign n32833 = n32832 ^ n32831 ;
  assign n32834 = n32822 ^ n32798 ;
  assign n32835 = n32834 ^ n32831 ;
  assign n32836 = ~n32833 & n32835 ;
  assign n32837 = n32836 ^ n32831 ;
  assign n32838 = ~n32823 & ~n32837 ;
  assign n32839 = n32838 ^ n30053 ;
  assign n32840 = ~n32826 & n32839 ;
  assign n32857 = n32843 ^ n32840 ;
  assign n33023 = n33014 ^ n32857 ;
  assign n1704 = n1688 ^ n1195 ;
  assign n1708 = n1707 ^ n1704 ;
  assign n1709 = n1708 ^ n977 ;
  assign n33039 = n33023 ^ n1709 ;
  assign n33793 = n33200 ^ n33039 ;
  assign n32989 = n32556 ^ n32538 ;
  assign n34681 = n33793 ^ n32989 ;
  assign n34682 = n32989 ^ n32133 ;
  assign n34683 = n34681 & n34682 ;
  assign n34684 = n34683 ^ n32133 ;
  assign n33348 = n32234 ^ n30945 ;
  assign n33349 = n32204 ^ n30945 ;
  assign n33350 = ~n33348 & ~n33349 ;
  assign n33351 = n33350 ^ n32234 ;
  assign n33352 = n33167 ^ n33118 ;
  assign n33354 = n33351 & ~n33352 ;
  assign n33379 = n32114 ^ n30951 ;
  assign n33380 = n32202 ^ n30951 ;
  assign n33381 = ~n33379 & n33380 ;
  assign n33382 = n33381 ^ n32114 ;
  assign n33383 = n33164 ^ n33120 ;
  assign n33397 = n32240 ^ n31618 ;
  assign n33398 = n31618 ^ n30965 ;
  assign n33399 = n33397 & n33398 ;
  assign n33400 = n33399 ^ n30965 ;
  assign n33401 = n33155 ^ n33135 ;
  assign n33404 = n33400 & n33401 ;
  assign n33418 = n33149 ^ n33148 ;
  assign n33414 = n31635 ^ n30974 ;
  assign n33415 = n32256 ^ n31635 ;
  assign n33416 = ~n33414 & n33415 ;
  assign n33417 = n33416 ^ n30974 ;
  assign n33419 = n33418 ^ n33417 ;
  assign n33424 = n33143 ^ n33142 ;
  assign n33420 = n31641 ^ n30979 ;
  assign n33421 = n32259 ^ n31641 ;
  assign n33422 = n33420 & n33421 ;
  assign n33423 = n33422 ^ n30979 ;
  assign n33425 = n33424 ^ n33423 ;
  assign n33473 = n31647 ^ n30982 ;
  assign n33474 = n32265 ^ n31647 ;
  assign n33475 = n33473 & ~n33474 ;
  assign n33476 = n33475 ^ n30982 ;
  assign n33465 = n31011 ^ n29987 ;
  assign n33466 = n31785 ^ n31011 ;
  assign n33467 = n33465 & ~n33466 ;
  assign n33462 = n32568 ^ n32524 ;
  assign n33427 = n31013 ^ n29990 ;
  assign n33428 = n31791 ^ n31013 ;
  assign n33429 = ~n33427 & n33428 ;
  assign n33430 = n33429 ^ n29990 ;
  assign n33460 = n33430 ^ n29012 ;
  assign n33461 = n33460 ^ n29987 ;
  assign n33463 = n33462 ^ n33461 ;
  assign n33464 = n33463 ^ n3193 ;
  assign n33468 = n33467 ^ n33464 ;
  assign n32129 = n32128 ^ n32108 ;
  assign n31592 = n31591 ^ n31024 ;
  assign n31604 = n31603 ^ n31591 ;
  assign n31605 = n31592 & ~n31604 ;
  assign n31606 = n31605 ^ n31024 ;
  assign n32130 = n32129 ^ n31606 ;
  assign n32145 = n32102 ^ n31993 ;
  assign n32144 = ~n32138 & n32143 ;
  assign n32146 = n32145 ^ n32144 ;
  assign n32147 = n31683 ^ n30850 ;
  assign n32152 = n32151 ^ n31683 ;
  assign n32153 = n32147 & ~n32152 ;
  assign n32154 = n32153 ^ n30850 ;
  assign n32155 = n32154 ^ n32144 ;
  assign n32156 = ~n32146 & ~n32155 ;
  assign n32157 = n32156 ^ n32145 ;
  assign n32158 = n32157 ^ n31606 ;
  assign n32131 = n31695 ^ n30890 ;
  assign n32134 = n32133 ^ n31695 ;
  assign n32135 = ~n32131 & n32134 ;
  assign n32136 = n32135 ^ n30890 ;
  assign n32137 = n32136 ^ n32129 ;
  assign n32159 = n32158 ^ n32137 ;
  assign n32161 = n32105 ^ n31988 ;
  assign n32160 = n32157 ^ n32137 ;
  assign n32162 = n32161 ^ n32160 ;
  assign n32163 = n32162 ^ n32137 ;
  assign n32164 = n32159 & n32163 ;
  assign n32165 = n32164 ^ n32137 ;
  assign n32166 = n32130 & ~n32165 ;
  assign n32167 = n32166 ^ n32129 ;
  assign n32168 = n32145 & ~n32154 ;
  assign n32170 = n32169 ^ n32144 ;
  assign n32171 = ~n32168 & ~n32170 ;
  assign n32172 = n31606 & n32171 ;
  assign n32173 = n32129 & n32172 ;
  assign n32174 = n32173 ^ n32171 ;
  assign n32175 = n32167 & n32174 ;
  assign n32686 = n32175 & n32685 ;
  assign n32687 = n32686 ^ n32167 ;
  assign n32688 = n32687 ^ n32167 ;
  assign n32689 = n32173 ^ n32136 ;
  assign n32690 = ~n32161 & ~n32689 ;
  assign n32691 = n32688 & n32690 ;
  assign n32692 = n32691 ^ n32687 ;
  assign n32693 = n31728 ^ n31045 ;
  assign n32694 = n32286 ^ n31728 ;
  assign n32695 = n32693 & n32694 ;
  assign n32696 = n32695 ^ n31045 ;
  assign n32697 = n32547 ^ n32544 ;
  assign n32935 = n32696 & ~n32697 ;
  assign n32698 = n32697 ^ n32696 ;
  assign n32936 = n32935 ^ n32698 ;
  assign n32937 = ~n32692 & ~n32936 ;
  assign n32929 = n30811 ^ n30278 ;
  assign n32930 = n32390 ^ n30811 ;
  assign n32931 = n32929 & n32930 ;
  assign n32932 = n32931 ^ n30278 ;
  assign n32933 = n32550 ^ n32542 ;
  assign n32953 = ~n32932 & ~n32933 ;
  assign n32985 = n30902 ^ n30271 ;
  assign n32986 = n31580 ^ n30902 ;
  assign n32987 = n32985 & n32986 ;
  assign n32988 = n32987 ^ n30271 ;
  assign n32990 = n32989 ^ n32988 ;
  assign n33226 = ~n32953 & ~n32990 ;
  assign n33227 = ~n32936 & n33226 ;
  assign n32943 = n30859 ^ n30277 ;
  assign n32944 = n32494 ^ n30859 ;
  assign n32945 = ~n32943 & ~n32944 ;
  assign n32946 = n32945 ^ n30277 ;
  assign n32947 = n32553 ^ n32540 ;
  assign n33228 = n32946 & n32947 ;
  assign n33229 = n33227 & ~n33228 ;
  assign n33230 = n32937 & n33229 ;
  assign n33231 = n32988 ^ n32946 ;
  assign n33232 = n33231 ^ n32947 ;
  assign n32949 = n32935 ^ n32932 ;
  assign n32950 = n32935 ^ n32933 ;
  assign n32951 = ~n32949 & n32950 ;
  assign n32952 = n32951 ^ n32933 ;
  assign n33233 = n33232 ^ n32952 ;
  assign n33234 = n33233 ^ n33231 ;
  assign n33235 = n32988 ^ n32947 ;
  assign n33236 = n33235 ^ n33231 ;
  assign n33237 = n33234 & n33236 ;
  assign n33238 = n33237 ^ n33231 ;
  assign n33239 = ~n32990 & ~n33238 ;
  assign n33240 = n33239 ^ n32989 ;
  assign n33241 = ~n33230 & ~n33240 ;
  assign n33225 = n32559 ^ n32536 ;
  assign n33242 = n33241 ^ n33225 ;
  assign n33243 = n31074 ^ n30265 ;
  assign n33244 = n31795 ^ n31074 ;
  assign n33245 = n33243 & ~n33244 ;
  assign n33246 = n33245 ^ n30265 ;
  assign n33300 = n33246 ^ n33225 ;
  assign n33301 = ~n33242 & ~n33300 ;
  assign n33302 = n33301 ^ n33246 ;
  assign n33293 = n31805 ^ n31071 ;
  assign n33294 = n32562 ^ n32534 ;
  assign n33295 = n33294 ^ n30258 ;
  assign n33296 = n33295 ^ n31805 ;
  assign n33297 = n33296 ^ n33294 ;
  assign n33298 = ~n33293 & n33297 ;
  assign n33299 = n33298 ^ n33295 ;
  assign n33303 = n33302 ^ n33299 ;
  assign n33304 = n33303 ^ n29489 ;
  assign n32701 = ~n32170 & n32685 ;
  assign n32702 = n32157 & ~n32168 ;
  assign n32703 = n32701 & n32702 ;
  assign n32704 = n32703 ^ n32157 ;
  assign n32705 = n32704 ^ n32136 ;
  assign n32708 = n32704 ^ n32161 ;
  assign n32709 = n32705 & ~n32708 ;
  assign n32706 = n32161 ^ n32130 ;
  assign n32710 = n32709 ^ n32706 ;
  assign n32711 = n32710 ^ n29904 ;
  assign n32712 = n32161 ^ n32136 ;
  assign n32713 = n32712 ^ n32704 ;
  assign n32714 = n32713 ^ n30115 ;
  assign n32842 = n32841 ^ n32840 ;
  assign n32844 = ~n32842 & ~n32843 ;
  assign n32845 = n32844 ^ n29909 ;
  assign n32716 = n32154 ^ n32145 ;
  assign n32715 = ~n32144 & ~n32701 ;
  assign n32717 = n32716 ^ n32715 ;
  assign n32846 = n32845 ^ n32717 ;
  assign n32847 = n32845 ^ n29918 ;
  assign n32848 = ~n32846 & ~n32847 ;
  assign n32849 = n32848 ^ n29918 ;
  assign n32850 = n32849 ^ n32713 ;
  assign n32851 = ~n32714 & ~n32850 ;
  assign n32852 = n32851 ^ n30115 ;
  assign n32853 = n32852 ^ n32710 ;
  assign n32854 = n32711 & ~n32853 ;
  assign n32855 = n32854 ^ n29904 ;
  assign n32699 = n32698 ^ n32692 ;
  assign n32925 = n30177 & n32699 ;
  assign n32700 = n32699 ^ n30177 ;
  assign n32926 = n32925 ^ n32700 ;
  assign n32927 = n32855 & n32926 ;
  assign n32938 = ~n32935 & ~n32937 ;
  assign n32934 = n32933 ^ n32932 ;
  assign n32939 = n32938 ^ n32934 ;
  assign n32963 = ~n29507 & n32939 ;
  assign n32954 = n32937 & ~n32953 ;
  assign n32955 = ~n32952 & n32954 ;
  assign n32956 = n32955 ^ n32952 ;
  assign n32948 = n32947 ^ n32946 ;
  assign n32957 = n32956 ^ n32948 ;
  assign n32958 = n32957 ^ n29514 ;
  assign n32984 = n32956 ^ n32946 ;
  assign n32991 = n32990 ^ n32947 ;
  assign n32992 = n32991 ^ n32946 ;
  assign n32993 = n32992 ^ n32990 ;
  assign n32994 = n32984 & n32993 ;
  assign n32995 = n32994 ^ n32991 ;
  assign n32996 = n32995 ^ n29497 ;
  assign n33249 = ~n32958 & ~n32996 ;
  assign n33250 = ~n32963 & n33249 ;
  assign n33251 = n32927 & n33250 ;
  assign n33253 = n32995 ^ n32957 ;
  assign n32959 = n32939 ^ n32925 ;
  assign n32960 = n32925 ^ n29507 ;
  assign n32961 = n32959 & n32960 ;
  assign n32962 = n32961 ^ n29507 ;
  assign n33252 = n32995 ^ n32962 ;
  assign n33254 = n33253 ^ n33252 ;
  assign n33255 = n32995 ^ n29514 ;
  assign n33256 = n33255 ^ n33253 ;
  assign n33257 = n33254 & ~n33256 ;
  assign n33258 = n33257 ^ n33253 ;
  assign n33259 = ~n32996 & ~n33258 ;
  assign n33260 = n33259 ^ n29497 ;
  assign n33261 = ~n33251 & n33260 ;
  assign n33247 = n33246 ^ n33242 ;
  assign n33289 = n33261 ^ n33247 ;
  assign n33290 = n33261 ^ n29528 ;
  assign n33291 = n33289 & ~n33290 ;
  assign n33292 = n33291 ^ n29528 ;
  assign n33305 = n33304 ^ n33292 ;
  assign n33248 = n33247 ^ n29528 ;
  assign n33262 = n33261 ^ n33248 ;
  assign n32964 = n32927 & ~n32963 ;
  assign n32965 = ~n32962 & n32964 ;
  assign n32966 = n32965 ^ n32962 ;
  assign n32983 = n32966 ^ n32957 ;
  assign n32997 = n32996 ^ n29514 ;
  assign n32998 = n32997 ^ n32957 ;
  assign n32999 = n32998 ^ n32996 ;
  assign n33000 = ~n32983 & ~n32999 ;
  assign n33001 = n33000 ^ n32997 ;
  assign n32856 = n32855 ^ n32700 ;
  assign n32858 = n32849 ^ n32714 ;
  assign n32859 = n32717 ^ n29918 ;
  assign n32860 = n32859 ^ n32845 ;
  assign n32861 = n30115 ^ n29904 ;
  assign n32862 = n32861 ^ n32710 ;
  assign n32863 = n32862 ^ n32851 ;
  assign n32864 = ~n32860 & n32863 ;
  assign n32865 = n32858 & n32864 ;
  assign n32866 = ~n32857 & n32865 ;
  assign n32878 = ~n32871 & ~n32877 ;
  assign n32887 = n32878 & ~n32886 ;
  assign n32888 = ~n32867 & n32887 ;
  assign n32889 = n32888 ^ n32878 ;
  assign n32890 = n32889 ^ n32877 ;
  assign n32891 = n32866 & ~n32890 ;
  assign n32921 = ~n32871 & ~n32920 ;
  assign n32922 = n32891 & n32921 ;
  assign n32892 = n32891 ^ n32865 ;
  assign n32923 = n32922 ^ n32892 ;
  assign n32924 = ~n32856 & ~n32923 ;
  assign n32940 = n32939 ^ n29507 ;
  assign n32928 = ~n32925 & ~n32927 ;
  assign n32941 = n32940 ^ n32928 ;
  assign n32942 = n32924 & ~n32941 ;
  assign n32967 = n32966 ^ n32958 ;
  assign n33002 = n32942 & n32967 ;
  assign n33003 = n33002 ^ n33001 ;
  assign n33263 = ~n33001 & n33003 ;
  assign n33306 = ~n33262 & ~n33263 ;
  assign n33441 = ~n33305 & n33306 ;
  assign n33432 = n33302 ^ n33294 ;
  assign n33433 = n33299 & n33432 ;
  assign n33434 = n33433 ^ n33294 ;
  assign n33426 = n32565 ^ n32529 ;
  assign n33431 = n33430 ^ n33426 ;
  assign n33435 = n33434 ^ n33431 ;
  assign n33454 = n33441 ^ n33435 ;
  assign n33437 = n33303 ^ n33292 ;
  assign n33438 = ~n33304 & ~n33437 ;
  assign n33439 = n33438 ^ n29489 ;
  assign n33457 = n33454 ^ n33439 ;
  assign n33458 = ~n29021 & ~n33457 ;
  assign n33455 = n33439 ^ n33435 ;
  assign n33456 = ~n33454 & n33455 ;
  assign n33459 = n33458 ^ n33456 ;
  assign n33469 = n33468 ^ n33459 ;
  assign n33443 = n30900 ^ n3157 ;
  assign n33444 = n33443 ^ n2522 ;
  assign n33445 = n33444 ^ n3188 ;
  assign n33470 = n33469 ^ n33445 ;
  assign n33452 = n33434 ^ n33430 ;
  assign n33453 = n33431 & ~n33452 ;
  assign n33471 = n33470 ^ n33453 ;
  assign n33436 = n33435 ^ n29021 ;
  assign n33440 = n33439 ^ n33436 ;
  assign n33442 = n33441 ^ n33440 ;
  assign n33446 = n33445 ^ n33442 ;
  assign n33307 = n33306 ^ n33305 ;
  assign n33311 = n33310 ^ n33307 ;
  assign n33015 = ~n32857 & n33014 ;
  assign n33016 = ~n32860 & ~n33015 ;
  assign n33017 = n32858 & n33016 ;
  assign n33018 = n33017 ^ n32863 ;
  assign n1423 = n1360 ^ n1314 ;
  assign n1424 = n1423 ^ n1410 ;
  assign n1428 = n1427 ^ n1424 ;
  assign n33019 = n33018 ^ n1428 ;
  assign n33024 = n1709 & n33023 ;
  assign n1713 = n1694 ^ n1204 ;
  assign n1714 = n1713 ^ n983 ;
  assign n1715 = n1714 ^ n1416 ;
  assign n33025 = n33024 ^ n1715 ;
  assign n33026 = n33015 ^ n32860 ;
  assign n33027 = n33026 ^ n1715 ;
  assign n33028 = n33025 & ~n33027 ;
  assign n33029 = n33028 ^ n33024 ;
  assign n1412 = n1299 ^ n1219 ;
  assign n1419 = n1418 ^ n1412 ;
  assign n1420 = n1419 ^ n1157 ;
  assign n33021 = n33018 ^ n1420 ;
  assign n33020 = n33016 ^ n32858 ;
  assign n33022 = n33021 ^ n33020 ;
  assign n33030 = n33029 ^ n33022 ;
  assign n33031 = n33030 ^ n33021 ;
  assign n33032 = n33020 ^ n33018 ;
  assign n33033 = n33032 ^ n33021 ;
  assign n33034 = ~n33031 & n33033 ;
  assign n33035 = n33034 ^ n33021 ;
  assign n33036 = n33019 & ~n33035 ;
  assign n33037 = n33036 ^ n1428 ;
  assign n33038 = n33020 ^ n1420 ;
  assign n33040 = n33039 ^ n33024 ;
  assign n33041 = ~n1715 & ~n33026 ;
  assign n33042 = n33040 & n33041 ;
  assign n33043 = n33042 ^ n33040 ;
  assign n33044 = n33019 & n33043 ;
  assign n33045 = n33038 & n33044 ;
  assign n33046 = ~n33037 & n33045 ;
  assign n33201 = n33046 & ~n33200 ;
  assign n33202 = n33201 ^ n33037 ;
  assign n32968 = n32967 ^ n32942 ;
  assign n33010 = ~n2873 & n32968 ;
  assign n33004 = n30639 ^ n3212 ;
  assign n33005 = n33004 ^ n27168 ;
  assign n33006 = n33005 ^ n2577 ;
  assign n33007 = n33006 ^ n33003 ;
  assign n32970 = n32941 ^ n32924 ;
  assign n33203 = ~n32970 & ~n32973 ;
  assign n32975 = n32923 ^ n32856 ;
  assign n33204 = n32975 ^ n1446 ;
  assign n32976 = n1446 & ~n32975 ;
  assign n33205 = n33204 ^ n32976 ;
  assign n33206 = n33203 & ~n33205 ;
  assign n33207 = n33206 ^ n33205 ;
  assign n33265 = n33007 & ~n33207 ;
  assign n33266 = ~n33010 & n33265 ;
  assign n33267 = n33202 & n33266 ;
  assign n32969 = n32968 ^ n2873 ;
  assign n32974 = n32973 ^ n32970 ;
  assign n32977 = n32976 ^ n32970 ;
  assign n32978 = n32974 & ~n32977 ;
  assign n32979 = n32978 ^ n32973 ;
  assign n32980 = n32979 ^ n32968 ;
  assign n32981 = ~n32969 & n32980 ;
  assign n32982 = n32981 ^ n2873 ;
  assign n33268 = n33003 ^ n32982 ;
  assign n33269 = n33007 & ~n33268 ;
  assign n33270 = n33269 ^ n33006 ;
  assign n33271 = ~n33267 & ~n33270 ;
  assign n2652 = n2651 ^ n2516 ;
  assign n2653 = n2652 ^ n2582 ;
  assign n2654 = n2653 ^ n2630 ;
  assign n33272 = n33271 ^ n2654 ;
  assign n33264 = n33263 ^ n33262 ;
  assign n33286 = n33264 ^ n2654 ;
  assign n33287 = ~n33272 & n33286 ;
  assign n33288 = n33287 ^ n2654 ;
  assign n33447 = n33307 ^ n33288 ;
  assign n33448 = ~n33311 & n33447 ;
  assign n33449 = n33448 ^ n33310 ;
  assign n33450 = n33449 ^ n33445 ;
  assign n33451 = ~n33446 & n33450 ;
  assign n33472 = n33471 ^ n33451 ;
  assign n33477 = n33476 ^ n33472 ;
  assign n33285 = n32275 ^ n31659 ;
  assign n33312 = n33311 ^ n33288 ;
  assign n33313 = n33312 ^ n30995 ;
  assign n33314 = n33313 ^ n32275 ;
  assign n33315 = n33314 ^ n33312 ;
  assign n33316 = n33285 & n33315 ;
  assign n33317 = n33316 ^ n33313 ;
  assign n33218 = n32626 ^ n31665 ;
  assign n30908 = n30907 ^ n30906 ;
  assign n31588 = n31587 ^ n30906 ;
  assign n31589 = ~n30908 & n31588 ;
  assign n31590 = n31589 ^ n30907 ;
  assign n33008 = n33007 ^ n32982 ;
  assign n33009 = n33008 ^ n33007 ;
  assign n33208 = n33202 & ~n33207 ;
  assign n33209 = ~n33010 & n33208 ;
  assign n33210 = ~n33009 & n33209 ;
  assign n33211 = n33210 ^ n33008 ;
  assign n33219 = ~n31590 & n33211 ;
  assign n33220 = n33219 ^ n31001 ;
  assign n33221 = n33220 ^ n32626 ;
  assign n33222 = n33221 ^ n33219 ;
  assign n33223 = ~n33218 & n33222 ;
  assign n33224 = n33223 ^ n33220 ;
  assign n33273 = n33272 ^ n33264 ;
  assign n33318 = n33273 ^ n33219 ;
  assign n33319 = ~n33224 & ~n33318 ;
  assign n33320 = n33319 ^ n33273 ;
  assign n33479 = n33320 ^ n33312 ;
  assign n33480 = ~n33317 & n33479 ;
  assign n33481 = n33480 ^ n33312 ;
  assign n33478 = n33449 ^ n33446 ;
  assign n33482 = n33481 ^ n33478 ;
  assign n33483 = n32639 ^ n31653 ;
  assign n33484 = n33478 ^ n30988 ;
  assign n33485 = n33484 ^ n32639 ;
  assign n33486 = n33485 ^ n33478 ;
  assign n33487 = ~n33483 & n33486 ;
  assign n33488 = n33487 ^ n33484 ;
  assign n33489 = n33482 & n33488 ;
  assign n33490 = n33489 ^ n33481 ;
  assign n33491 = n33490 ^ n33472 ;
  assign n33492 = n33477 & n33491 ;
  assign n33493 = n33492 ^ n33476 ;
  assign n33494 = n33493 ^ n33423 ;
  assign n33495 = ~n33425 & n33494 ;
  assign n33496 = n33495 ^ n33424 ;
  assign n33497 = n33496 ^ n33417 ;
  assign n33498 = ~n33419 & ~n33497 ;
  assign n33499 = n33498 ^ n33418 ;
  assign n33326 = n33152 ^ n33139 ;
  assign n33500 = n33499 ^ n33326 ;
  assign n33501 = n32246 ^ n31625 ;
  assign n33502 = n33326 ^ n30968 ;
  assign n33503 = n33502 ^ n33326 ;
  assign n33504 = n33503 ^ n32246 ;
  assign n33505 = ~n33501 & ~n33504 ;
  assign n33506 = n33505 ^ n33502 ;
  assign n33507 = n33500 & ~n33506 ;
  assign n33508 = n33507 ^ n33326 ;
  assign n33509 = ~n33404 & ~n33508 ;
  assign n33391 = n33158 ^ n33130 ;
  assign n33392 = n32233 ^ n31611 ;
  assign n33393 = n32233 ^ n30960 ;
  assign n33394 = n33392 & ~n33393 ;
  assign n33395 = n33394 ^ n30960 ;
  assign n33510 = ~n33391 & n33395 ;
  assign n33511 = n33509 & n33510 ;
  assign n33512 = n33511 ^ n33509 ;
  assign n33385 = n33161 ^ n33125 ;
  assign n33386 = n32667 ^ n31943 ;
  assign n33387 = n31943 ^ n30954 ;
  assign n33388 = n33386 & ~n33387 ;
  assign n33389 = n33388 ^ n30954 ;
  assign n33513 = ~n33385 & n33389 ;
  assign n33514 = n33512 & n33513 ;
  assign n33515 = n33514 ^ n33512 ;
  assign n33516 = ~n33383 & n33515 ;
  assign n33517 = ~n33382 & n33516 ;
  assign n33518 = n33517 ^ n33515 ;
  assign n33553 = ~n33354 & n33518 ;
  assign n33353 = n33352 ^ n33351 ;
  assign n33355 = n33354 ^ n33353 ;
  assign n33384 = n33383 ^ n33382 ;
  assign n33390 = n33389 ^ n33385 ;
  assign n33396 = n33395 ^ n33391 ;
  assign n33402 = n33401 ^ n33400 ;
  assign n33403 = n33402 ^ n33391 ;
  assign n33405 = n33404 ^ n33403 ;
  assign n33406 = ~n33396 & n33405 ;
  assign n33407 = n33406 ^ n33395 ;
  assign n33408 = n33407 ^ n33385 ;
  assign n33409 = ~n33390 & n33408 ;
  assign n33410 = n33409 ^ n33389 ;
  assign n33411 = n33410 ^ n33382 ;
  assign n33412 = n33384 & n33411 ;
  assign n33413 = n33412 ^ n33383 ;
  assign n33552 = ~n33354 & n33413 ;
  assign n33619 = ~n33355 & ~n33552 ;
  assign n33620 = ~n33553 & n33619 ;
  assign n33357 = n32311 ^ n30935 ;
  assign n33358 = n32220 ^ n30935 ;
  assign n33359 = ~n33357 & n33358 ;
  assign n33360 = n33359 ^ n32311 ;
  assign n33347 = n33170 ^ n33116 ;
  assign n33361 = n33360 ^ n33347 ;
  assign n33621 = n33620 ^ n33361 ;
  assign n33519 = ~n33413 & ~n33518 ;
  assign n33561 = n33519 ^ n33353 ;
  assign n33562 = n33561 ^ n29931 ;
  assign n33610 = n33410 & ~n33515 ;
  assign n33611 = n33610 ^ n33384 ;
  assign n33565 = n33508 ^ n33402 ;
  assign n33566 = n33565 ^ n29939 ;
  assign n33567 = n33506 ^ n33499 ;
  assign n33568 = n33567 ^ n30335 ;
  assign n33569 = n33496 ^ n33419 ;
  assign n33570 = n33569 ^ n30325 ;
  assign n33571 = n33493 ^ n33425 ;
  assign n33572 = n33571 ^ n29945 ;
  assign n33573 = n33490 ^ n33477 ;
  assign n33574 = n33573 ^ n29951 ;
  assign n33575 = n33488 ^ n33481 ;
  assign n33576 = n33575 ^ n29958 ;
  assign n33321 = n33320 ^ n33317 ;
  assign n33322 = n33321 ^ n29968 ;
  assign n33212 = n33211 ^ n31590 ;
  assign n33216 = n29981 & ~n33212 ;
  assign n33217 = n33216 ^ n29974 ;
  assign n33274 = n33273 ^ n33224 ;
  assign n33282 = n33274 ^ n33216 ;
  assign n33283 = ~n33217 & n33282 ;
  assign n33284 = n33283 ^ n29974 ;
  assign n33577 = n33321 ^ n33284 ;
  assign n33578 = ~n33322 & n33577 ;
  assign n33579 = n33578 ^ n29968 ;
  assign n33580 = n33579 ^ n33575 ;
  assign n33581 = n33576 & n33580 ;
  assign n33582 = n33581 ^ n29958 ;
  assign n33583 = n33582 ^ n33573 ;
  assign n33584 = ~n33574 & n33583 ;
  assign n33585 = n33584 ^ n29951 ;
  assign n33586 = n33585 ^ n33571 ;
  assign n33587 = n33572 & n33586 ;
  assign n33588 = n33587 ^ n29945 ;
  assign n33589 = n33588 ^ n33569 ;
  assign n33590 = ~n33570 & ~n33589 ;
  assign n33591 = n33590 ^ n30325 ;
  assign n33592 = n33591 ^ n33567 ;
  assign n33593 = n33568 & ~n33592 ;
  assign n33594 = n33593 ^ n30335 ;
  assign n33595 = n33594 ^ n33565 ;
  assign n33596 = n33566 & n33595 ;
  assign n33597 = n33596 ^ n29939 ;
  assign n33598 = n33597 ^ n30348 ;
  assign n33601 = n33401 ^ n33396 ;
  assign n33599 = n33508 ^ n33400 ;
  assign n33600 = n33402 & ~n33599 ;
  assign n33602 = n33601 ^ n33600 ;
  assign n33603 = n33602 ^ n33597 ;
  assign n33604 = ~n33598 & n33603 ;
  assign n33605 = n33604 ^ n30348 ;
  assign n33563 = n33407 & ~n33512 ;
  assign n33564 = n33563 ^ n33390 ;
  assign n33606 = n33605 ^ n33564 ;
  assign n33607 = n33605 ^ n30358 ;
  assign n33608 = ~n33606 & ~n33607 ;
  assign n33609 = n33608 ^ n30358 ;
  assign n33612 = n33611 ^ n33609 ;
  assign n33613 = n33611 ^ n29937 ;
  assign n33614 = ~n33612 & n33613 ;
  assign n33615 = n33614 ^ n29937 ;
  assign n33616 = n33615 ^ n33561 ;
  assign n33617 = ~n33562 & n33616 ;
  assign n33618 = n33617 ^ n29931 ;
  assign n33622 = n33621 ^ n33618 ;
  assign n33623 = n33621 ^ n29927 ;
  assign n33624 = ~n33622 & n33623 ;
  assign n33625 = n33624 ^ n29927 ;
  assign n33356 = n33355 ^ n33347 ;
  assign n33362 = ~n33356 & ~n33361 ;
  assign n33363 = n33362 ^ n33355 ;
  assign n33520 = n33347 & n33360 ;
  assign n33554 = ~n33363 & ~n33520 ;
  assign n33555 = ~n33553 & n33554 ;
  assign n33556 = ~n33552 & n33555 ;
  assign n33557 = n33556 ^ n33554 ;
  assign n33558 = n33557 ^ n33363 ;
  assign n33367 = n32197 ^ n30929 ;
  assign n33368 = n32189 ^ n30929 ;
  assign n33369 = n33367 & ~n33368 ;
  assign n33370 = n33369 ^ n32197 ;
  assign n33364 = n33173 ^ n33114 ;
  assign n33521 = n33370 ^ n33364 ;
  assign n33559 = n33558 ^ n33521 ;
  assign n33560 = n33559 ^ n30383 ;
  assign n33692 = n33625 ^ n33560 ;
  assign n33668 = n33615 ^ n33562 ;
  assign n33669 = n33613 ^ n33609 ;
  assign n33670 = n33564 ^ n30358 ;
  assign n33671 = n33670 ^ n33605 ;
  assign n33672 = n33588 ^ n33570 ;
  assign n33673 = n33585 ^ n33572 ;
  assign n33323 = n33322 ^ n33284 ;
  assign n33674 = n33579 ^ n33576 ;
  assign n33675 = ~n33323 & n33674 ;
  assign n33676 = n33582 ^ n33574 ;
  assign n33677 = n33675 & n33676 ;
  assign n33678 = n33673 & ~n33677 ;
  assign n33679 = ~n33672 & ~n33678 ;
  assign n33680 = n33591 ^ n33568 ;
  assign n33681 = n33679 & ~n33680 ;
  assign n33682 = n33594 ^ n33566 ;
  assign n33683 = ~n33681 & n33682 ;
  assign n33684 = n33602 ^ n30348 ;
  assign n33685 = n33684 ^ n33597 ;
  assign n33686 = n33683 & ~n33685 ;
  assign n33687 = n33671 & ~n33686 ;
  assign n33688 = n33669 & n33687 ;
  assign n33689 = ~n33668 & n33688 ;
  assign n33690 = n33623 ^ n33618 ;
  assign n33691 = n33689 & n33690 ;
  assign n33912 = n33692 ^ n33691 ;
  assign n2952 = n2951 ^ n2948 ;
  assign n2953 = n2952 ^ n608 ;
  assign n2957 = n2956 ^ n2953 ;
  assign n33913 = n33912 ^ n2957 ;
  assign n33914 = n33690 ^ n33689 ;
  assign n33918 = n33917 ^ n33914 ;
  assign n33920 = n31403 ^ n596 ;
  assign n33921 = n33920 ^ n27799 ;
  assign n33922 = n33921 ^ n22776 ;
  assign n33919 = n33688 ^ n33668 ;
  assign n33923 = n33922 ^ n33919 ;
  assign n33927 = n33687 ^ n33669 ;
  assign n33924 = n31461 ^ n23944 ;
  assign n33925 = n33924 ^ n27803 ;
  assign n33926 = n33925 ^ n1475 ;
  assign n33928 = n33927 ^ n33926 ;
  assign n33932 = n33686 ^ n33671 ;
  assign n33929 = n31407 ^ n23884 ;
  assign n33930 = n33929 ^ n2439 ;
  assign n33931 = n33930 ^ n22373 ;
  assign n33933 = n33932 ^ n33931 ;
  assign n33934 = n33685 ^ n33683 ;
  assign n2424 = n2421 ^ n2390 ;
  assign n2425 = n2424 ^ n2348 ;
  assign n2429 = n2428 ^ n2425 ;
  assign n33935 = n33934 ^ n2429 ;
  assign n33936 = n33682 ^ n33681 ;
  assign n2412 = n2333 ^ n2277 ;
  assign n2413 = n2412 ^ n2411 ;
  assign n2414 = n2413 ^ n2402 ;
  assign n33937 = n33936 ^ n2414 ;
  assign n33939 = n31418 ^ n2259 ;
  assign n33940 = n33939 ^ n27436 ;
  assign n33941 = n33940 ^ n2409 ;
  assign n33938 = n33680 ^ n33679 ;
  assign n33942 = n33941 ^ n33938 ;
  assign n33944 = n31423 ^ n2249 ;
  assign n33945 = n33944 ^ n27469 ;
  assign n33946 = n33945 ^ n2081 ;
  assign n33943 = n33678 ^ n33672 ;
  assign n33947 = n33946 ^ n33943 ;
  assign n33949 = n31428 ^ n23898 ;
  assign n33950 = n33949 ^ n1988 ;
  assign n33951 = n33950 ^ n22319 ;
  assign n33948 = n33677 ^ n33673 ;
  assign n33952 = n33951 ^ n33948 ;
  assign n33956 = n33676 ^ n33675 ;
  assign n33953 = n31435 ^ n23902 ;
  assign n33954 = n33953 ^ n27448 ;
  assign n33955 = n33954 ^ n1983 ;
  assign n33957 = n33956 ^ n33955 ;
  assign n33958 = n33674 ^ n33323 ;
  assign n1911 = n1910 ^ n1895 ;
  assign n1924 = n1923 ^ n1911 ;
  assign n1928 = n1927 ^ n1924 ;
  assign n33959 = n33958 ^ n1928 ;
  assign n33279 = n30821 ^ n23907 ;
  assign n33280 = n33279 ^ n3032 ;
  assign n33281 = n33280 ^ n1918 ;
  assign n33324 = n33323 ^ n33281 ;
  assign n33213 = n33212 ^ n29981 ;
  assign n33214 = n2756 & ~n33213 ;
  assign n33215 = n33214 ^ n3242 ;
  assign n33275 = n33274 ^ n33217 ;
  assign n33276 = n33275 ^ n3242 ;
  assign n33277 = n33215 & ~n33276 ;
  assign n33278 = n33277 ^ n33214 ;
  assign n33960 = n33281 ^ n33278 ;
  assign n33961 = ~n33324 & ~n33960 ;
  assign n33962 = n33961 ^ n33323 ;
  assign n33963 = n33962 ^ n1928 ;
  assign n33964 = n33959 & ~n33963 ;
  assign n33965 = n33964 ^ n1928 ;
  assign n33966 = n33965 ^ n33955 ;
  assign n33967 = ~n33957 & ~n33966 ;
  assign n33968 = n33967 ^ n33956 ;
  assign n33969 = n33968 ^ n33948 ;
  assign n33970 = ~n33952 & ~n33969 ;
  assign n33971 = n33970 ^ n33951 ;
  assign n33972 = n33971 ^ n33943 ;
  assign n33973 = ~n33947 & n33972 ;
  assign n33974 = n33973 ^ n33946 ;
  assign n33975 = n33974 ^ n33938 ;
  assign n33976 = n33942 & ~n33975 ;
  assign n33977 = n33976 ^ n33941 ;
  assign n33978 = n33977 ^ n33936 ;
  assign n33979 = ~n33937 & n33978 ;
  assign n33980 = n33979 ^ n2414 ;
  assign n33981 = n33980 ^ n2429 ;
  assign n33982 = ~n33935 & ~n33981 ;
  assign n33983 = n33982 ^ n33934 ;
  assign n33984 = n33983 ^ n33931 ;
  assign n33985 = n33933 & n33984 ;
  assign n33986 = n33985 ^ n33932 ;
  assign n33987 = n33986 ^ n33926 ;
  assign n33988 = ~n33928 & ~n33987 ;
  assign n33989 = n33988 ^ n33927 ;
  assign n33990 = n33989 ^ n33919 ;
  assign n33991 = n33923 & n33990 ;
  assign n33992 = n33991 ^ n33922 ;
  assign n33993 = n33992 ^ n33914 ;
  assign n33994 = ~n33918 & n33993 ;
  assign n33995 = n33994 ^ n33917 ;
  assign n33996 = n33995 ^ n2957 ;
  assign n33997 = n33913 & ~n33996 ;
  assign n33998 = n33997 ^ n33912 ;
  assign n33342 = n32212 ^ n32138 ;
  assign n33343 = n32138 ^ n30926 ;
  assign n33344 = ~n33342 & ~n33343 ;
  assign n33345 = n33344 ^ n30926 ;
  assign n33341 = n33176 ^ n33109 ;
  assign n33346 = n33345 ^ n33341 ;
  assign n33632 = n33364 ^ n33346 ;
  assign n33630 = n33558 ^ n33370 ;
  assign n33631 = n33521 & ~n33630 ;
  assign n33633 = n33632 ^ n33631 ;
  assign n33694 = n33633 ^ n29911 ;
  assign n33626 = n33625 ^ n33559 ;
  assign n33627 = n33560 & n33626 ;
  assign n33628 = n33627 ^ n30383 ;
  assign n33695 = n33694 ^ n33628 ;
  assign n33693 = ~n33691 & ~n33692 ;
  assign n33910 = n33695 ^ n33693 ;
  assign n33911 = n33910 ^ n33909 ;
  assign n34680 = n33998 ^ n33911 ;
  assign n34685 = n34684 ^ n34680 ;
  assign n33999 = n33998 ^ n33909 ;
  assign n34000 = ~n33911 & ~n33999 ;
  assign n34001 = n34000 ^ n33910 ;
  assign n33529 = n32193 ^ n32145 ;
  assign n33340 = n33179 ^ n33104 ;
  assign n33530 = n33340 ^ n30910 ;
  assign n33531 = n33530 ^ n32145 ;
  assign n33532 = n33531 ^ n33340 ;
  assign n33533 = ~n33529 & n33532 ;
  assign n33534 = n33533 ^ n33530 ;
  assign n33365 = n33364 ^ n33341 ;
  assign n33366 = n33365 ^ n33363 ;
  assign n33371 = n33370 ^ n33366 ;
  assign n33372 = n33371 ^ n33365 ;
  assign n33373 = n33363 ^ n33341 ;
  assign n33374 = n33373 ^ n33365 ;
  assign n33375 = ~n33372 & n33374 ;
  assign n33376 = n33375 ^ n33365 ;
  assign n33377 = ~n33346 & n33376 ;
  assign n33378 = n33377 ^ n33345 ;
  assign n33522 = ~n33346 & ~n33354 ;
  assign n33523 = n33521 & n33522 ;
  assign n33524 = ~n33520 & n33523 ;
  assign n33525 = ~n33519 & n33524 ;
  assign n33526 = ~n33378 & n33525 ;
  assign n33527 = n33526 ^ n33378 ;
  assign n33637 = n33534 ^ n33527 ;
  assign n33639 = n33637 ^ n30399 ;
  assign n33629 = n33628 ^ n29911 ;
  assign n33634 = n33633 ^ n33628 ;
  assign n33635 = ~n33629 & n33634 ;
  assign n33636 = n33635 ^ n29911 ;
  assign n33697 = n33639 ^ n33636 ;
  assign n33696 = ~n33693 & ~n33695 ;
  assign n33877 = n33697 ^ n33696 ;
  assign n33881 = n33880 ^ n33877 ;
  assign n34882 = n34001 ^ n33881 ;
  assign n34503 = n33995 ^ n33913 ;
  assign n34499 = n32947 ^ n32151 ;
  assign n33743 = n33051 ^ n33048 ;
  assign n33744 = n33062 & ~n33072 ;
  assign n33745 = n33194 & n33744 ;
  assign n33746 = n33745 ^ n33072 ;
  assign n33771 = n33746 ^ n33067 ;
  assign n33772 = n33771 ^ n33051 ;
  assign n33773 = n33772 ^ n33067 ;
  assign n33774 = ~n33743 & n33773 ;
  assign n33775 = n33774 ^ n33771 ;
  assign n34500 = n33775 ^ n32151 ;
  assign n34501 = ~n34499 & n34500 ;
  assign n34502 = n34501 ^ n32947 ;
  assign n34504 = n34503 ^ n34502 ;
  assign n33747 = n33746 ^ n33743 ;
  assign n34485 = n33747 ^ n32933 ;
  assign n34486 = n33747 ^ n32140 ;
  assign n34487 = ~n34485 & n34486 ;
  assign n34488 = n34487 ^ n32140 ;
  assign n34686 = n34503 ^ n34488 ;
  assign n34064 = n33986 ^ n33928 ;
  assign n33712 = n33194 ^ n33056 ;
  assign n34065 = n33712 ^ n32129 ;
  assign n34066 = n33712 ^ n32193 ;
  assign n34067 = n34065 & ~n34066 ;
  assign n34068 = n34067 ^ n32193 ;
  assign n34473 = ~n34064 & ~n34068 ;
  assign n34070 = n32697 ^ n32185 ;
  assign n33730 = n33194 ^ n33052 ;
  assign n33731 = n33056 & ~n33730 ;
  assign n33728 = n33055 ^ n762 ;
  assign n33729 = n33728 ^ n33059 ;
  assign n33732 = n33731 ^ n33729 ;
  assign n34071 = n33732 ^ n32185 ;
  assign n34072 = n34070 & n34071 ;
  assign n34073 = n34072 ^ n32697 ;
  assign n34474 = n34473 ^ n34073 ;
  assign n34329 = n33989 ^ n33923 ;
  assign n34475 = n34473 ^ n34329 ;
  assign n34476 = ~n34474 & n34475 ;
  assign n34477 = n34476 ^ n34073 ;
  assign n34687 = n34686 ^ n34477 ;
  assign n34489 = n33992 ^ n33918 ;
  assign n34688 = n34687 ^ n34489 ;
  assign n34689 = n34688 ^ n34686 ;
  assign n34690 = n34502 ^ n34477 ;
  assign n34691 = n34690 ^ n34686 ;
  assign n34692 = ~n34689 & ~n34691 ;
  assign n34693 = n34692 ^ n34686 ;
  assign n34694 = ~n34504 & n34693 ;
  assign n34695 = n34694 ^ n34503 ;
  assign n34074 = n32212 ^ n32161 ;
  assign n34075 = n33983 ^ n33933 ;
  assign n33661 = n33191 ^ n33084 ;
  assign n34076 = n34075 ^ n33661 ;
  assign n34077 = n34076 ^ n34075 ;
  assign n34078 = n34077 ^ n32212 ;
  assign n34079 = n34074 & ~n34078 ;
  assign n34080 = n34079 ^ n34076 ;
  assign n33543 = n33188 ^ n33089 ;
  assign n34082 = n33543 ^ n32145 ;
  assign n34083 = n33543 ^ n32197 ;
  assign n34084 = n34082 & n34083 ;
  assign n34085 = n34084 ^ n32197 ;
  assign n34081 = n33980 ^ n33935 ;
  assign n34086 = n34085 ^ n34081 ;
  assign n33328 = n33185 ^ n33094 ;
  assign n34087 = n33328 ^ n32138 ;
  assign n34088 = n33977 ^ n33937 ;
  assign n34089 = n34088 ^ n32311 ;
  assign n34090 = n34089 ^ n32138 ;
  assign n34091 = n34090 ^ n34088 ;
  assign n34092 = n34087 & n34091 ;
  assign n34093 = n34092 ^ n34089 ;
  assign n34096 = n32204 ^ n31943 ;
  assign n34097 = n33341 ^ n32204 ;
  assign n34098 = n34096 & n34097 ;
  assign n34099 = n34098 ^ n31943 ;
  assign n34095 = n33968 ^ n33952 ;
  assign n34100 = n34099 ^ n34095 ;
  assign n34101 = n33364 ^ n31611 ;
  assign n34102 = n33364 ^ n32202 ;
  assign n34103 = n34101 & n34102 ;
  assign n34104 = n34103 ^ n32202 ;
  assign n34105 = n32667 ^ n31618 ;
  assign n34106 = n33347 ^ n32667 ;
  assign n34107 = n34105 & ~n34106 ;
  assign n34108 = n34107 ^ n31618 ;
  assign n34109 = n33962 ^ n33959 ;
  assign n34111 = ~n34108 & ~n34109 ;
  assign n34110 = n34109 ^ n34108 ;
  assign n34112 = n34111 ^ n34110 ;
  assign n34113 = n33965 ^ n33957 ;
  assign n34114 = n34112 & n34113 ;
  assign n34115 = ~n34104 & n34114 ;
  assign n34116 = n34115 ^ n34112 ;
  assign n34117 = n34100 & n34116 ;
  assign n34119 = n32220 ^ n32114 ;
  assign n34120 = n33340 ^ n32220 ;
  assign n34121 = ~n34119 & n34120 ;
  assign n34122 = n34121 ^ n32114 ;
  assign n34118 = n33971 ^ n33947 ;
  assign n34123 = n34122 ^ n34118 ;
  assign n34124 = n34117 & ~n34123 ;
  assign n34280 = n33275 ^ n33215 ;
  assign n34129 = n33385 ^ n32246 ;
  assign n34130 = n33213 ^ n2756 ;
  assign n34131 = n34130 ^ n31641 ;
  assign n34132 = n34131 ^ n33385 ;
  assign n34133 = n34132 ^ n34130 ;
  assign n34134 = n34129 & ~n34133 ;
  assign n34135 = n34134 ^ n34131 ;
  assign n34170 = n33202 ^ n32974 ;
  assign n34171 = n34170 ^ n1446 ;
  assign n34172 = n34171 ^ n32974 ;
  assign n34173 = n33204 & n34172 ;
  assign n34174 = n34173 ^ n34170 ;
  assign n34166 = n31676 ^ n31013 ;
  assign n34167 = n32589 ^ n31013 ;
  assign n34168 = n34166 & n34167 ;
  assign n34169 = n34168 ^ n31676 ;
  assign n34175 = n34174 ^ n34169 ;
  assign n34155 = n33202 ^ n1446 ;
  assign n34156 = n34155 ^ n32975 ;
  assign n34024 = ~n33029 & n33043 ;
  assign n34025 = ~n33200 & n34024 ;
  assign n34026 = n34025 ^ n33029 ;
  assign n34145 = n34026 ^ n33020 ;
  assign n34146 = n33038 & ~n34145 ;
  assign n34144 = n33019 ^ n1420 ;
  assign n34147 = n34146 ^ n34144 ;
  assign n34140 = n31791 ^ n31074 ;
  assign n34141 = n32592 ^ n31791 ;
  assign n34142 = ~n34140 & ~n34141 ;
  assign n34143 = n34142 ^ n31074 ;
  assign n34148 = n34147 ^ n34143 ;
  assign n34023 = n32593 ^ n31805 ;
  assign n34027 = n34026 ^ n33038 ;
  assign n34028 = n34027 ^ n30902 ;
  assign n34029 = n34028 ^ n32593 ;
  assign n34030 = n34029 ^ n34027 ;
  assign n34031 = ~n34023 & ~n34030 ;
  assign n34032 = n34031 ^ n34028 ;
  assign n33817 = n31795 ^ n30859 ;
  assign n33818 = n33462 ^ n31795 ;
  assign n33819 = n33817 & ~n33818 ;
  assign n33820 = n33819 ^ n30859 ;
  assign n33789 = n33426 ^ n30811 ;
  assign n33790 = n33426 ^ n31580 ;
  assign n33791 = ~n33789 & n33790 ;
  assign n33792 = n33791 ^ n30811 ;
  assign n33794 = n33793 ^ n33792 ;
  assign n33742 = n33225 ^ n32390 ;
  assign n33748 = n33747 ^ n31591 ;
  assign n33749 = n33748 ^ n33747 ;
  assign n33750 = n33749 ^ n32390 ;
  assign n33751 = ~n33742 & n33750 ;
  assign n33752 = n33751 ^ n33748 ;
  assign n33733 = n32286 ^ n31695 ;
  assign n33734 = n32989 ^ n32286 ;
  assign n33735 = n33733 & n33734 ;
  assign n33736 = n33735 ^ n31695 ;
  assign n33708 = n32947 ^ n31603 ;
  assign n33709 = n32947 ^ n31683 ;
  assign n33710 = ~n33708 & ~n33709 ;
  assign n33711 = n33710 ^ n31683 ;
  assign n33713 = n33712 ^ n33711 ;
  assign n33657 = n32933 ^ n32133 ;
  assign n33658 = n32133 ^ n31560 ;
  assign n33659 = ~n33657 & ~n33658 ;
  assign n33660 = n33659 ^ n31560 ;
  assign n33662 = n33661 ^ n33660 ;
  assign n33544 = n32697 ^ n31537 ;
  assign n33545 = n32697 ^ n32151 ;
  assign n33546 = ~n33544 & n33545 ;
  assign n33547 = n33546 ^ n31537 ;
  assign n33548 = n33547 ^ n33543 ;
  assign n33329 = n32140 ^ n32129 ;
  assign n33330 = n32140 ^ n31286 ;
  assign n33331 = n33329 & n33330 ;
  assign n33332 = n33331 ^ n31286 ;
  assign n33333 = n33332 ^ n33328 ;
  assign n33338 = n33182 ^ n33099 ;
  assign n33334 = n32161 ^ n31164 ;
  assign n33335 = n32185 ^ n32161 ;
  assign n33336 = ~n33334 & n33335 ;
  assign n33337 = n33336 ^ n31164 ;
  assign n33339 = n33338 ^ n33337 ;
  assign n33528 = n33527 ^ n33340 ;
  assign n33535 = n33528 & n33534 ;
  assign n33536 = n33535 ^ n33527 ;
  assign n33537 = n33536 ^ n33337 ;
  assign n33538 = ~n33339 & n33537 ;
  assign n33539 = n33538 ^ n33338 ;
  assign n33540 = n33539 ^ n33328 ;
  assign n33541 = n33333 & ~n33540 ;
  assign n33542 = n33541 ^ n33332 ;
  assign n33654 = n33543 ^ n33542 ;
  assign n33655 = n33548 & ~n33654 ;
  assign n33656 = n33655 ^ n33547 ;
  assign n33705 = n33660 ^ n33656 ;
  assign n33706 = ~n33662 & n33705 ;
  assign n33707 = n33706 ^ n33661 ;
  assign n33725 = n33711 ^ n33707 ;
  assign n33726 = n33713 & ~n33725 ;
  assign n33727 = n33726 ^ n33712 ;
  assign n33753 = n33736 ^ n33727 ;
  assign n33754 = n33732 ^ n33727 ;
  assign n33755 = ~n33753 & ~n33754 ;
  assign n33756 = n33755 ^ n33736 ;
  assign n33768 = n33756 ^ n33747 ;
  assign n33769 = ~n33752 & ~n33768 ;
  assign n33770 = n33769 ^ n33747 ;
  assign n33785 = n33775 ^ n33770 ;
  assign n33776 = n32494 ^ n31728 ;
  assign n33777 = n33294 ^ n32494 ;
  assign n33778 = n33776 & ~n33777 ;
  assign n33779 = n33778 ^ n31728 ;
  assign n33786 = n33779 ^ n33770 ;
  assign n33787 = n33785 & n33786 ;
  assign n33788 = n33787 ^ n33779 ;
  assign n33806 = n33792 ^ n33788 ;
  assign n33807 = ~n33794 & ~n33806 ;
  assign n33808 = n33807 ^ n33793 ;
  assign n34033 = n33820 ^ n33808 ;
  assign n33809 = n33200 ^ n33023 ;
  assign n33810 = n1715 ^ n1709 ;
  assign n33811 = n33810 ^ n33026 ;
  assign n33812 = n33811 ^ n1715 ;
  assign n33813 = n33812 ^ n33026 ;
  assign n33814 = n33813 ^ n33200 ;
  assign n33815 = n33809 & ~n33814 ;
  assign n33816 = n33815 ^ n33811 ;
  assign n34034 = n33816 ^ n33808 ;
  assign n34035 = ~n34033 & n34034 ;
  assign n34036 = n34035 ^ n33820 ;
  assign n34149 = n34036 ^ n34027 ;
  assign n34150 = ~n34032 & n34149 ;
  assign n34151 = n34150 ^ n34027 ;
  assign n34152 = n34151 ^ n34147 ;
  assign n34153 = ~n34148 & n34152 ;
  assign n34154 = n34153 ^ n34151 ;
  assign n34157 = n34156 ^ n34154 ;
  assign n34158 = n32591 ^ n31785 ;
  assign n34159 = n34156 ^ n31071 ;
  assign n34160 = n34159 ^ n32591 ;
  assign n34161 = n34160 ^ n34156 ;
  assign n34162 = n34158 & n34161 ;
  assign n34163 = n34162 ^ n34159 ;
  assign n34164 = ~n34157 & ~n34163 ;
  assign n34165 = n34164 ^ n34156 ;
  assign n34239 = n34174 ^ n34165 ;
  assign n34240 = n34175 & n34239 ;
  assign n33663 = n33662 ^ n33656 ;
  assign n33664 = n33663 ^ n30569 ;
  assign n33645 = n33539 ^ n33333 ;
  assign n33550 = n33536 ^ n33339 ;
  assign n33551 = n33550 ^ n30398 ;
  assign n33638 = n33637 ^ n33636 ;
  assign n33640 = ~n33638 & n33639 ;
  assign n33641 = n33640 ^ n30399 ;
  assign n33642 = n33641 ^ n33550 ;
  assign n33643 = ~n33551 & ~n33642 ;
  assign n33644 = n33643 ^ n30398 ;
  assign n33646 = n33645 ^ n33644 ;
  assign n33647 = n33645 ^ n29902 ;
  assign n33648 = ~n33646 & ~n33647 ;
  assign n33649 = n33648 ^ n29902 ;
  assign n33549 = n33548 ^ n33542 ;
  assign n33650 = n33649 ^ n33549 ;
  assign n33651 = n33649 ^ n30417 ;
  assign n33652 = n33650 & n33651 ;
  assign n33653 = n33652 ^ n30417 ;
  assign n33665 = n33664 ^ n33653 ;
  assign n33666 = n33549 ^ n30417 ;
  assign n33667 = n33666 ^ n33649 ;
  assign n33698 = n33696 & n33697 ;
  assign n33699 = n33641 ^ n33551 ;
  assign n33700 = n33698 & ~n33699 ;
  assign n33701 = n33647 ^ n33644 ;
  assign n33702 = ~n33700 & ~n33701 ;
  assign n33703 = ~n33667 & ~n33702 ;
  assign n33704 = ~n33665 & n33703 ;
  assign n33716 = n33663 ^ n33653 ;
  assign n33717 = ~n33664 & ~n33716 ;
  assign n33718 = n33717 ^ n30569 ;
  assign n33714 = n33713 ^ n33707 ;
  assign n33715 = n33714 ^ n30850 ;
  assign n33719 = n33718 ^ n33715 ;
  assign n33720 = ~n33704 & n33719 ;
  assign n33737 = n33736 ^ n33732 ;
  assign n33738 = n33737 ^ n33727 ;
  assign n33739 = n33738 ^ n30890 ;
  assign n33721 = n33718 ^ n33714 ;
  assign n33722 = n33718 ^ n30850 ;
  assign n33723 = ~n33721 & n33722 ;
  assign n33724 = n33723 ^ n30850 ;
  assign n33740 = n33739 ^ n33724 ;
  assign n33741 = n33720 & ~n33740 ;
  assign n33759 = n33738 ^ n33724 ;
  assign n33760 = ~n33739 & n33759 ;
  assign n33761 = n33760 ^ n30890 ;
  assign n33757 = n33756 ^ n33752 ;
  assign n33758 = n33757 ^ n31024 ;
  assign n33762 = n33761 ^ n33758 ;
  assign n33763 = n33741 & ~n33762 ;
  assign n33780 = n33779 ^ n33775 ;
  assign n33781 = n33780 ^ n33770 ;
  assign n33782 = n33781 ^ n31045 ;
  assign n33764 = n33761 ^ n33757 ;
  assign n33765 = n33761 ^ n31024 ;
  assign n33766 = ~n33764 & ~n33765 ;
  assign n33767 = n33766 ^ n31024 ;
  assign n33783 = n33782 ^ n33767 ;
  assign n33784 = ~n33763 & ~n33783 ;
  assign n33797 = n33781 ^ n33767 ;
  assign n33798 = ~n33782 & ~n33797 ;
  assign n33799 = n33798 ^ n31045 ;
  assign n33795 = n33794 ^ n33788 ;
  assign n33796 = n33795 ^ n30278 ;
  assign n33800 = n33799 ^ n33796 ;
  assign n33801 = n33784 & n33800 ;
  assign n33821 = n33820 ^ n33816 ;
  assign n33822 = n33821 ^ n33808 ;
  assign n33823 = n33822 ^ n30277 ;
  assign n33802 = n33799 ^ n33795 ;
  assign n33803 = n33799 ^ n30278 ;
  assign n33804 = n33802 & n33803 ;
  assign n33805 = n33804 ^ n30278 ;
  assign n33824 = n33823 ^ n33805 ;
  assign n34022 = n33801 & ~n33824 ;
  assign n34039 = n33822 ^ n33805 ;
  assign n34040 = n33823 & n34039 ;
  assign n34041 = n34040 ^ n30277 ;
  assign n34037 = n34036 ^ n34032 ;
  assign n34038 = n34037 ^ n30271 ;
  assign n34042 = n34041 ^ n34038 ;
  assign n34193 = n34022 & n34042 ;
  assign n34182 = n34041 ^ n34037 ;
  assign n34183 = n34041 ^ n30271 ;
  assign n34184 = ~n34182 & n34183 ;
  assign n34185 = n34184 ^ n30271 ;
  assign n34180 = n34151 ^ n34148 ;
  assign n34181 = n34180 ^ n30265 ;
  assign n34194 = n34185 ^ n34181 ;
  assign n34195 = ~n34193 & ~n34194 ;
  assign n34186 = n34185 ^ n34180 ;
  assign n34187 = n34181 & n34186 ;
  assign n34188 = n34187 ^ n30265 ;
  assign n34178 = n34163 ^ n34154 ;
  assign n34179 = n34178 ^ n30258 ;
  assign n34196 = n34188 ^ n34179 ;
  assign n34197 = n34195 & ~n34196 ;
  assign n34189 = n34188 ^ n34178 ;
  assign n34190 = ~n34179 & n34189 ;
  assign n34191 = n34190 ^ n30258 ;
  assign n34232 = n34197 ^ n34191 ;
  assign n34176 = n34175 ^ n34165 ;
  assign n34236 = n34232 ^ n34176 ;
  assign n34237 = n29990 & ~n34236 ;
  assign n34231 = n34197 ^ n34176 ;
  assign n34233 = n34231 & ~n34232 ;
  assign n34226 = ~n32979 & ~n33208 ;
  assign n34227 = n34226 ^ n32969 ;
  assign n34224 = n34169 ^ n29987 ;
  assign n34225 = n34224 ^ n31011 ;
  assign n34228 = n34227 ^ n34225 ;
  assign n34229 = n34228 ^ n3227 ;
  assign n34221 = n32583 ^ n31824 ;
  assign n34222 = n31824 ^ n31011 ;
  assign n34223 = ~n34221 & ~n34222 ;
  assign n34230 = n34229 ^ n34223 ;
  assign n34234 = n34233 ^ n34230 ;
  assign n2662 = n2612 ^ n2532 ;
  assign n2672 = n2671 ^ n2662 ;
  assign n2676 = n2675 ^ n2672 ;
  assign n34235 = n34234 ^ n2676 ;
  assign n34238 = n34237 ^ n34235 ;
  assign n34241 = n34240 ^ n34238 ;
  assign n34177 = n34176 ^ n29990 ;
  assign n34192 = n34191 ^ n34177 ;
  assign n34198 = n34197 ^ n34192 ;
  assign n34199 = n34198 ^ n2676 ;
  assign n34202 = n31577 ^ n2592 ;
  assign n34203 = n34202 ^ n3122 ;
  assign n34204 = n34203 ^ n22733 ;
  assign n34201 = n34194 ^ n34193 ;
  assign n34205 = n34204 ^ n34201 ;
  assign n34043 = n34042 ^ n34022 ;
  assign n34019 = n24002 ^ n2902 ;
  assign n34020 = n34019 ^ n27522 ;
  assign n34021 = n34020 ^ n3101 ;
  assign n34044 = n34043 ^ n34021 ;
  assign n33826 = n3110 ^ n2887 ;
  assign n33827 = n33826 ^ n27867 ;
  assign n33828 = n33827 ^ n22741 ;
  assign n33825 = n33824 ^ n33801 ;
  assign n33829 = n33828 ^ n33825 ;
  assign n33831 = n31522 ^ n2849 ;
  assign n33832 = n33831 ^ n27861 ;
  assign n33833 = n33832 ^ n22748 ;
  assign n33830 = n33800 ^ n33784 ;
  assign n33834 = n33833 ^ n33830 ;
  assign n33836 = n2837 ^ n1773 ;
  assign n33837 = n33836 ^ n27856 ;
  assign n33838 = n33837 ^ n2639 ;
  assign n33835 = n33783 ^ n33763 ;
  assign n33839 = n33838 ^ n33835 ;
  assign n33840 = n33762 ^ n33741 ;
  assign n1260 = n1259 ^ n1160 ;
  assign n1261 = n1260 ^ n1253 ;
  assign n1262 = n1261 ^ n1241 ;
  assign n33841 = n33840 ^ n1262 ;
  assign n33850 = n33719 ^ n33704 ;
  assign n959 = n908 ^ n892 ;
  assign n960 = n959 ^ n956 ;
  assign n964 = n963 ^ n960 ;
  assign n33848 = n33703 ^ n33665 ;
  assign n33849 = n964 & n33848 ;
  assign n33851 = n33850 ^ n33849 ;
  assign n33852 = n33849 ^ n1083 ;
  assign n33853 = ~n33851 & ~n33852 ;
  assign n33854 = n33853 ^ n33850 ;
  assign n33843 = n1755 ^ n1738 ;
  assign n33844 = n33843 ^ n1090 ;
  assign n33845 = n33844 ^ n1247 ;
  assign n33846 = n33845 ^ n33840 ;
  assign n33842 = n33740 ^ n33720 ;
  assign n33847 = n33846 ^ n33842 ;
  assign n33855 = n33854 ^ n33847 ;
  assign n33856 = n33855 ^ n33846 ;
  assign n33857 = n33842 ^ n33840 ;
  assign n33858 = n33857 ^ n33846 ;
  assign n33859 = ~n33856 & ~n33858 ;
  assign n33860 = n33859 ^ n33846 ;
  assign n33861 = ~n33841 & n33860 ;
  assign n33862 = n33861 ^ n1262 ;
  assign n33863 = n33845 ^ n33842 ;
  assign n33864 = n33848 ^ n964 ;
  assign n33865 = n33864 ^ n33849 ;
  assign n33866 = ~n1083 & n33850 ;
  assign n33867 = n33865 & n33866 ;
  assign n33868 = n33867 ^ n33865 ;
  assign n33869 = ~n33841 & n33868 ;
  assign n33870 = ~n33863 & n33869 ;
  assign n33871 = ~n33862 & n33870 ;
  assign n33872 = n33702 ^ n33667 ;
  assign n33873 = n33701 ^ n33700 ;
  assign n33882 = ~n33877 & n33880 ;
  assign n33883 = n33882 ^ n33881 ;
  assign n33884 = n33699 ^ n33698 ;
  assign n33885 = ~n1611 & ~n33884 ;
  assign n33886 = ~n33883 & ~n33885 ;
  assign n33887 = ~n33876 & n33886 ;
  assign n33888 = ~n33873 & n33887 ;
  assign n33889 = n33888 ^ n949 ;
  assign n33890 = n33872 & ~n33889 ;
  assign n33906 = n33888 ^ n33886 ;
  assign n33891 = n33872 ^ n949 ;
  assign n33894 = n33882 ^ n1611 ;
  assign n33895 = n33884 ^ n1611 ;
  assign n33896 = n33894 & ~n33895 ;
  assign n33897 = n33896 ^ n33882 ;
  assign n33892 = n33873 ^ n33872 ;
  assign n33893 = n33892 ^ n33876 ;
  assign n33898 = n33897 ^ n33893 ;
  assign n33899 = n33898 ^ n33892 ;
  assign n33900 = n33876 ^ n949 ;
  assign n33901 = n33900 ^ n33892 ;
  assign n33902 = ~n33899 & n33901 ;
  assign n33903 = n33902 ^ n33892 ;
  assign n33904 = ~n33891 & ~n33903 ;
  assign n33905 = n33904 ^ n33872 ;
  assign n34002 = n33905 & ~n34001 ;
  assign n34003 = n33906 & n34002 ;
  assign n34006 = n33890 & n34003 ;
  assign n34004 = n34003 ^ n33905 ;
  assign n34007 = n34006 ^ n34004 ;
  assign n34008 = n33871 & ~n34007 ;
  assign n34009 = n34008 ^ n33862 ;
  assign n34010 = n34009 ^ n33838 ;
  assign n34011 = ~n33839 & n34010 ;
  assign n34012 = n34011 ^ n33838 ;
  assign n34013 = n34012 ^ n33830 ;
  assign n34014 = ~n33834 & n34013 ;
  assign n34015 = n34014 ^ n33833 ;
  assign n34016 = n34015 ^ n33825 ;
  assign n34017 = n33829 & ~n34016 ;
  assign n34018 = n34017 ^ n33828 ;
  assign n34206 = n34021 ^ n34018 ;
  assign n34207 = ~n34044 & ~n34206 ;
  assign n34208 = n34207 ^ n34043 ;
  assign n34209 = n34208 ^ n34201 ;
  assign n34210 = n34205 & n34209 ;
  assign n34211 = n34210 ^ n34204 ;
  assign n34200 = n34196 ^ n34195 ;
  assign n34212 = n34211 ^ n34200 ;
  assign n34213 = n31774 ^ n2633 ;
  assign n34214 = n34213 ^ n27927 ;
  assign n34215 = n34214 ^ n2669 ;
  assign n34216 = n34215 ^ n34211 ;
  assign n34217 = n34212 & n34216 ;
  assign n34218 = n34217 ^ n34215 ;
  assign n34219 = n34218 ^ n2676 ;
  assign n34220 = n34199 & n34219 ;
  assign n34242 = n34241 ^ n34220 ;
  assign n34136 = n33391 ^ n32256 ;
  assign n34137 = n32256 ^ n31647 ;
  assign n34138 = ~n34136 & n34137 ;
  assign n34139 = n34138 ^ n31647 ;
  assign n34243 = n34242 ^ n34139 ;
  assign n34248 = n34218 ^ n34199 ;
  assign n34244 = n33401 ^ n32259 ;
  assign n34245 = n32259 ^ n31653 ;
  assign n34246 = n34244 & n34245 ;
  assign n34247 = n34246 ^ n31653 ;
  assign n34249 = n34248 ^ n34247 ;
  assign n34254 = n34215 ^ n34200 ;
  assign n34255 = n34254 ^ n34211 ;
  assign n34250 = n33326 ^ n32265 ;
  assign n34251 = n33326 ^ n31659 ;
  assign n34252 = n34250 & n34251 ;
  assign n34253 = n34252 ^ n31659 ;
  assign n34256 = n34255 ^ n34253 ;
  assign n34045 = n34044 ^ n34018 ;
  assign n34046 = n32275 ^ n30906 ;
  assign n34047 = n33424 ^ n32275 ;
  assign n34048 = n34046 & ~n34047 ;
  assign n34049 = n34048 ^ n30906 ;
  assign n34258 = ~n34045 & n34049 ;
  assign n34257 = n34208 ^ n34205 ;
  assign n34259 = n34258 ^ n34257 ;
  assign n34260 = n33418 ^ n32639 ;
  assign n34261 = n34258 ^ n31665 ;
  assign n34262 = n34261 ^ n33418 ;
  assign n34263 = n34262 ^ n34258 ;
  assign n34264 = n34260 & ~n34263 ;
  assign n34265 = n34264 ^ n34261 ;
  assign n34266 = ~n34259 & n34265 ;
  assign n34267 = n34266 ^ n34258 ;
  assign n34268 = n34267 ^ n34255 ;
  assign n34269 = ~n34256 & ~n34268 ;
  assign n34270 = n34269 ^ n34267 ;
  assign n34271 = n34270 ^ n34247 ;
  assign n34272 = n34249 & ~n34271 ;
  assign n34273 = n34272 ^ n34248 ;
  assign n34274 = n34273 ^ n34139 ;
  assign n34275 = n34243 & ~n34274 ;
  assign n34276 = n34275 ^ n34242 ;
  assign n34277 = n34276 ^ n34130 ;
  assign n34278 = n34135 & ~n34277 ;
  assign n34279 = n34278 ^ n34130 ;
  assign n34281 = n34280 ^ n34279 ;
  assign n34282 = n33383 ^ n32240 ;
  assign n34283 = n34280 ^ n31635 ;
  assign n34284 = n34283 ^ n33383 ;
  assign n34285 = n34284 ^ n34280 ;
  assign n34286 = ~n34282 & ~n34285 ;
  assign n34287 = n34286 ^ n34283 ;
  assign n34288 = ~n34281 & ~n34287 ;
  assign n34289 = n34288 ^ n34280 ;
  assign n34125 = n32233 ^ n31625 ;
  assign n34126 = n33352 ^ n32233 ;
  assign n34127 = ~n34125 & ~n34126 ;
  assign n34128 = n34127 ^ n31625 ;
  assign n34290 = n34289 ^ n34128 ;
  assign n33325 = n33324 ^ n33278 ;
  assign n34291 = n34289 ^ n33325 ;
  assign n34292 = n34290 & ~n34291 ;
  assign n34293 = n34292 ^ n33325 ;
  assign n34294 = n34124 & ~n34293 ;
  assign n34296 = n34113 ^ n34104 ;
  assign n34297 = n34113 ^ n34111 ;
  assign n34298 = n34296 & ~n34297 ;
  assign n34299 = n34298 ^ n34111 ;
  assign n34295 = n34122 ^ n34095 ;
  assign n34300 = n34299 ^ n34295 ;
  assign n34301 = n34300 ^ n34099 ;
  assign n34302 = n34301 ^ n34295 ;
  assign n34303 = n34299 ^ n34118 ;
  assign n34304 = n34303 ^ n34295 ;
  assign n34305 = ~n34302 & n34304 ;
  assign n34306 = n34305 ^ n34295 ;
  assign n34307 = ~n34123 & n34306 ;
  assign n34308 = n34307 ^ n34122 ;
  assign n34309 = ~n34294 & ~n34308 ;
  assign n34094 = n33974 ^ n33942 ;
  assign n34310 = n34309 ^ n34094 ;
  assign n34311 = n33338 ^ n32189 ;
  assign n34312 = n34094 ^ n32234 ;
  assign n34313 = n34312 ^ n32189 ;
  assign n34314 = n34313 ^ n34094 ;
  assign n34315 = ~n34311 & ~n34314 ;
  assign n34316 = n34315 ^ n34312 ;
  assign n34317 = ~n34310 & n34316 ;
  assign n34318 = n34317 ^ n34309 ;
  assign n34319 = n34318 ^ n34088 ;
  assign n34320 = n34093 & n34319 ;
  assign n34321 = n34320 ^ n34088 ;
  assign n34322 = n34321 ^ n34081 ;
  assign n34323 = ~n34086 & ~n34322 ;
  assign n34324 = n34323 ^ n34085 ;
  assign n34325 = n34324 ^ n34075 ;
  assign n34326 = ~n34080 & ~n34325 ;
  assign n34327 = n34326 ^ n34075 ;
  assign n34069 = n34068 ^ n34064 ;
  assign n34478 = n34473 ^ n34069 ;
  assign n34479 = n34073 & n34329 ;
  assign n34480 = n34478 & n34479 ;
  assign n34481 = n34480 ^ n34478 ;
  assign n34696 = n34503 ^ n34481 ;
  assign n34697 = ~n34488 & n34489 ;
  assign n34698 = n34481 & n34697 ;
  assign n34699 = n34698 ^ n34481 ;
  assign n34700 = n34502 & n34699 ;
  assign n34701 = n34696 & n34700 ;
  assign n34702 = n34701 ^ n34699 ;
  assign n34703 = ~n34327 & n34702 ;
  assign n34704 = ~n34695 & n34703 ;
  assign n34705 = n34704 ^ n34695 ;
  assign n34967 = n34882 ^ n34705 ;
  assign n34884 = n33225 ^ n31603 ;
  assign n34885 = n33816 ^ n31603 ;
  assign n34886 = n34884 & n34885 ;
  assign n34887 = n34886 ^ n33225 ;
  assign n34968 = n34967 ^ n34887 ;
  assign n34969 = n34968 ^ n34680 ;
  assign n34970 = n34969 ^ n34882 ;
  assign n34971 = n34970 ^ n34887 ;
  assign n34972 = n34685 & ~n34971 ;
  assign n34973 = n34972 ^ n34968 ;
  assign n35006 = n34973 ^ n31683 ;
  assign n34706 = n34705 ^ n34685 ;
  assign n34707 = n34706 ^ n31560 ;
  assign n34490 = n34489 ^ n34488 ;
  assign n34482 = ~n34327 & n34481 ;
  assign n34483 = n34477 & n34482 ;
  assign n34484 = n34483 ^ n34477 ;
  assign n34491 = n34490 ^ n34484 ;
  assign n34492 = n34491 ^ n31286 ;
  assign n34337 = n34327 ^ n34069 ;
  assign n34338 = n34337 ^ n30910 ;
  assign n34339 = n34324 ^ n34080 ;
  assign n34340 = n34339 ^ n30926 ;
  assign n34423 = n34321 ^ n34086 ;
  assign n34342 = n34316 ^ n34309 ;
  assign n34343 = n34342 ^ n30945 ;
  assign n34398 = n34116 & ~n34293 ;
  assign n34399 = ~n34299 & n34398 ;
  assign n34400 = n34399 ^ n34299 ;
  assign n34401 = n34400 ^ n34100 ;
  assign n34352 = n34293 ^ n34110 ;
  assign n34353 = n34352 ^ n30965 ;
  assign n34354 = n34128 ^ n33325 ;
  assign n34355 = n34354 ^ n34289 ;
  assign n34356 = n34355 ^ n30968 ;
  assign n34383 = n34287 ^ n34279 ;
  assign n34357 = n34276 ^ n34135 ;
  assign n34358 = n34357 ^ n30979 ;
  assign n34359 = n34273 ^ n34243 ;
  assign n34360 = n34359 ^ n30982 ;
  assign n34361 = n34270 ^ n34249 ;
  assign n34362 = n34361 ^ n30988 ;
  assign n34050 = n34049 ^ n34045 ;
  assign n34364 = ~n30907 & ~n34050 ;
  assign n34365 = n34364 ^ n31001 ;
  assign n34366 = n34265 ^ n34257 ;
  assign n34367 = n34366 ^ n34364 ;
  assign n34368 = n34365 & n34367 ;
  assign n34369 = n34368 ^ n31001 ;
  assign n34363 = n34267 ^ n34256 ;
  assign n34370 = n34369 ^ n34363 ;
  assign n34371 = n34369 ^ n30995 ;
  assign n34372 = ~n34370 & n34371 ;
  assign n34373 = n34372 ^ n30995 ;
  assign n34374 = n34373 ^ n34361 ;
  assign n34375 = n34362 & ~n34374 ;
  assign n34376 = n34375 ^ n30988 ;
  assign n34377 = n34376 ^ n34359 ;
  assign n34378 = n34360 & ~n34377 ;
  assign n34379 = n34378 ^ n30982 ;
  assign n34380 = n34379 ^ n34357 ;
  assign n34381 = ~n34358 & ~n34380 ;
  assign n34382 = n34381 ^ n30979 ;
  assign n34384 = n34383 ^ n34382 ;
  assign n34385 = n34383 ^ n30974 ;
  assign n34386 = n34384 & n34385 ;
  assign n34387 = n34386 ^ n30974 ;
  assign n34388 = n34387 ^ n34355 ;
  assign n34389 = n34356 & ~n34388 ;
  assign n34390 = n34389 ^ n30968 ;
  assign n34391 = n34390 ^ n34352 ;
  assign n34392 = n34353 & n34391 ;
  assign n34393 = n34392 ^ n30965 ;
  assign n34344 = n34293 ^ n34108 ;
  assign n34345 = n34113 ^ n34109 ;
  assign n34346 = n34345 ^ n34104 ;
  assign n34347 = n34346 ^ n34113 ;
  assign n34348 = n34347 ^ n34104 ;
  assign n34349 = n34348 ^ n34293 ;
  assign n34350 = ~n34344 & n34349 ;
  assign n34351 = n34350 ^ n34346 ;
  assign n34394 = n34393 ^ n34351 ;
  assign n34395 = n34393 ^ n30960 ;
  assign n34396 = n34394 & n34395 ;
  assign n34397 = n34396 ^ n30960 ;
  assign n34402 = n34401 ^ n34397 ;
  assign n34403 = n34401 ^ n30954 ;
  assign n34404 = n34402 & ~n34403 ;
  assign n34405 = n34404 ^ n30954 ;
  assign n34406 = n34405 ^ n30951 ;
  assign n34407 = n34400 ^ n34095 ;
  assign n34408 = n34123 ^ n34099 ;
  assign n34409 = n34408 ^ n34123 ;
  assign n34410 = n34409 ^ n34400 ;
  assign n34411 = ~n34407 & n34410 ;
  assign n34412 = n34411 ^ n34408 ;
  assign n34413 = n34412 ^ n34405 ;
  assign n34414 = n34406 & ~n34413 ;
  assign n34415 = n34414 ^ n30951 ;
  assign n34416 = n34415 ^ n34342 ;
  assign n34417 = n34343 & n34416 ;
  assign n34418 = n34417 ^ n30945 ;
  assign n34341 = n34318 ^ n34093 ;
  assign n34419 = n34418 ^ n34341 ;
  assign n34420 = n34418 ^ n30935 ;
  assign n34421 = n34419 & n34420 ;
  assign n34422 = n34421 ^ n30935 ;
  assign n34424 = n34423 ^ n34422 ;
  assign n34425 = n34423 ^ n30929 ;
  assign n34426 = ~n34424 & n34425 ;
  assign n34427 = n34426 ^ n30929 ;
  assign n34428 = n34427 ^ n34339 ;
  assign n34429 = ~n34340 & n34428 ;
  assign n34430 = n34429 ^ n30926 ;
  assign n34431 = n34430 ^ n34337 ;
  assign n34432 = n34338 & n34431 ;
  assign n34433 = n34432 ^ n30910 ;
  assign n34328 = n34327 ^ n34073 ;
  assign n34330 = n34329 ^ n34328 ;
  assign n34331 = n34330 ^ n34073 ;
  assign n34332 = n34331 ^ n34064 ;
  assign n34333 = n34332 ^ n34329 ;
  assign n34334 = ~n34069 & n34333 ;
  assign n34335 = n34334 ^ n34330 ;
  assign n34469 = n34433 ^ n34335 ;
  assign n34470 = n34433 ^ n31164 ;
  assign n34471 = ~n34469 & n34470 ;
  assign n34472 = n34471 ^ n31164 ;
  assign n34495 = n34491 ^ n34472 ;
  assign n34496 = n34492 & n34495 ;
  assign n34497 = n34496 ^ n31286 ;
  assign n34676 = n34497 ^ n31537 ;
  assign n34498 = n34488 ^ n34484 ;
  assign n34505 = n34504 ^ n34489 ;
  assign n34506 = n34505 ^ n34504 ;
  assign n34507 = n34506 ^ n34484 ;
  assign n34508 = n34498 & n34507 ;
  assign n34509 = n34508 ^ n34505 ;
  assign n34677 = n34509 ^ n34497 ;
  assign n34678 = n34676 & ~n34677 ;
  assign n34679 = n34678 ^ n31537 ;
  assign n34963 = n34706 ^ n34679 ;
  assign n34964 = n34707 & n34963 ;
  assign n34965 = n34964 ^ n31560 ;
  assign n35007 = n35006 ^ n34965 ;
  assign n34708 = n34707 ^ n34679 ;
  assign n34336 = n34335 ^ n31164 ;
  assign n34434 = n34433 ^ n34336 ;
  assign n34435 = n34430 ^ n34338 ;
  assign n34436 = n34425 ^ n34422 ;
  assign n34437 = n34341 ^ n30935 ;
  assign n34438 = n34437 ^ n34418 ;
  assign n34439 = n34403 ^ n34397 ;
  assign n34440 = n34351 ^ n30960 ;
  assign n34441 = n34440 ^ n34393 ;
  assign n34442 = n34387 ^ n34356 ;
  assign n34443 = n34385 ^ n34382 ;
  assign n34444 = n34363 ^ n30995 ;
  assign n34445 = n34444 ^ n34369 ;
  assign n34446 = n34373 ^ n34362 ;
  assign n34447 = ~n34445 & ~n34446 ;
  assign n34448 = n34376 ^ n34360 ;
  assign n34449 = n34447 & ~n34448 ;
  assign n34450 = n34379 ^ n34358 ;
  assign n34451 = ~n34449 & ~n34450 ;
  assign n34452 = n34443 & ~n34451 ;
  assign n34453 = ~n34442 & n34452 ;
  assign n34454 = n34390 ^ n34353 ;
  assign n34455 = ~n34453 & n34454 ;
  assign n34456 = n34441 & n34455 ;
  assign n34457 = ~n34439 & ~n34456 ;
  assign n34458 = n34412 ^ n30951 ;
  assign n34459 = n34458 ^ n34405 ;
  assign n34460 = n34457 & n34459 ;
  assign n34461 = n34415 ^ n34343 ;
  assign n34462 = n34460 & n34461 ;
  assign n34463 = n34438 & n34462 ;
  assign n34464 = n34436 & ~n34463 ;
  assign n34465 = n34427 ^ n34340 ;
  assign n34466 = ~n34464 & n34465 ;
  assign n34467 = ~n34435 & n34466 ;
  assign n34468 = n34434 & n34467 ;
  assign n34493 = n34492 ^ n34472 ;
  assign n34494 = ~n34468 & ~n34493 ;
  assign n34510 = n34509 ^ n31537 ;
  assign n34511 = n34510 ^ n34497 ;
  assign n34709 = ~n34494 & ~n34511 ;
  assign n35005 = ~n34708 & n34709 ;
  assign n35067 = n35007 ^ n35005 ;
  assign n35457 = n35456 ^ n35067 ;
  assign n34710 = n34709 ^ n34708 ;
  assign n34711 = n34710 ^ n1678 ;
  assign n34512 = n34511 ^ n34494 ;
  assign n1667 = n1666 ^ n1648 ;
  assign n1668 = n1667 ^ n842 ;
  assign n1669 = n1668 ^ n1017 ;
  assign n34513 = n34512 ^ n1669 ;
  assign n34523 = n34466 ^ n34435 ;
  assign n34524 = n680 & n34523 ;
  assign n34520 = n31991 ^ n1625 ;
  assign n34521 = n34520 ^ n2983 ;
  assign n34522 = n34521 ^ n738 ;
  assign n34525 = n34524 ^ n34522 ;
  assign n34526 = n34467 ^ n34434 ;
  assign n34527 = n34526 ^ n34522 ;
  assign n34528 = n34525 & n34527 ;
  assign n34529 = n34528 ^ n34524 ;
  assign n34515 = n2987 ^ n1664 ;
  assign n34516 = n34515 ^ n743 ;
  assign n34517 = n34516 ^ n1631 ;
  assign n34518 = n34517 ^ n34512 ;
  assign n34514 = n34493 ^ n34468 ;
  assign n34519 = n34518 ^ n34514 ;
  assign n34530 = n34529 ^ n34519 ;
  assign n34531 = n34530 ^ n34518 ;
  assign n34532 = n34514 ^ n34512 ;
  assign n34533 = n34532 ^ n34518 ;
  assign n34534 = ~n34531 & n34533 ;
  assign n34535 = n34534 ^ n34518 ;
  assign n34536 = ~n34513 & n34535 ;
  assign n34537 = n34536 ^ n1669 ;
  assign n34538 = n34523 ^ n680 ;
  assign n34539 = n34538 ^ n34524 ;
  assign n34540 = ~n34522 & n34526 ;
  assign n34541 = n34539 & n34540 ;
  assign n34542 = n34541 ^ n34539 ;
  assign n34543 = ~n34514 & n34542 ;
  assign n34544 = ~n34517 & n34543 ;
  assign n34545 = n34544 ^ n34513 ;
  assign n34546 = n34544 ^ n34542 ;
  assign n34547 = n34512 & n34546 ;
  assign n34548 = n34545 & n34547 ;
  assign n34549 = n34548 ^ n34546 ;
  assign n34550 = ~n34537 & n34549 ;
  assign n34554 = n34465 ^ n34464 ;
  assign n34555 = n34554 ^ n34553 ;
  assign n34559 = n34463 ^ n34436 ;
  assign n34560 = n34559 ^ n34558 ;
  assign n34564 = n34462 ^ n34438 ;
  assign n34565 = n34564 ^ n34563 ;
  assign n34567 = n32014 ^ n1487 ;
  assign n34568 = n34567 ^ n28679 ;
  assign n34569 = n34568 ^ n23072 ;
  assign n34566 = n34461 ^ n34460 ;
  assign n34570 = n34569 ^ n34566 ;
  assign n34572 = n32019 ^ n28636 ;
  assign n34573 = n34572 ^ n23133 ;
  assign n34574 = n34573 ^ n24544 ;
  assign n34571 = n34459 ^ n34457 ;
  assign n34575 = n34574 ^ n34571 ;
  assign n34583 = n34454 ^ n34453 ;
  assign n34584 = n32033 ^ n24557 ;
  assign n34585 = n34584 ^ n28641 ;
  assign n34586 = n34585 ^ n2292 ;
  assign n34587 = ~n34583 & n34586 ;
  assign n34582 = n34455 ^ n34441 ;
  assign n34588 = n34587 ^ n34582 ;
  assign n34589 = n32029 ^ n24549 ;
  assign n34590 = n34589 ^ n2297 ;
  assign n34591 = n34590 ^ n23080 ;
  assign n34592 = n34591 ^ n34582 ;
  assign n34593 = n34588 & ~n34592 ;
  assign n34594 = n34593 ^ n34587 ;
  assign n34578 = n32024 ^ n24589 ;
  assign n34579 = n34578 ^ n28665 ;
  assign n34580 = n34579 ^ n2915 ;
  assign n34576 = n34456 ^ n34439 ;
  assign n34577 = n34576 ^ n34571 ;
  assign n34581 = n34580 ^ n34577 ;
  assign n34595 = n34594 ^ n34581 ;
  assign n34596 = n34595 ^ n34577 ;
  assign n34597 = n34580 ^ n34571 ;
  assign n34598 = n34597 ^ n34577 ;
  assign n34599 = ~n34596 & ~n34598 ;
  assign n34600 = n34599 ^ n34577 ;
  assign n34601 = ~n34575 & ~n34600 ;
  assign n34602 = n34601 ^ n34574 ;
  assign n34603 = n34586 ^ n34583 ;
  assign n34604 = n34603 ^ n34587 ;
  assign n34605 = ~n34582 & ~n34591 ;
  assign n34606 = ~n34604 & n34605 ;
  assign n34607 = n34606 ^ n34604 ;
  assign n34608 = ~n34575 & ~n34607 ;
  assign n34609 = n34452 ^ n34442 ;
  assign n2148 = n2147 ^ n2096 ;
  assign n2161 = n2160 ^ n2148 ;
  assign n2165 = n2164 ^ n2161 ;
  assign n34610 = n34609 ^ n2165 ;
  assign n34614 = n34451 ^ n34443 ;
  assign n34611 = n32040 ^ n24562 ;
  assign n34612 = n34611 ^ n2071 ;
  assign n34613 = n34612 ^ n2155 ;
  assign n34615 = n34614 ^ n34613 ;
  assign n34616 = n34450 ^ n34449 ;
  assign n2038 = n2031 ^ n2007 ;
  assign n2057 = n2056 ^ n2038 ;
  assign n2064 = n2063 ^ n2057 ;
  assign n34617 = n34616 ^ n2064 ;
  assign n34619 = n32048 ^ n1969 ;
  assign n34620 = n34619 ^ n28012 ;
  assign n34621 = n34620 ^ n2051 ;
  assign n34618 = n34448 ^ n34447 ;
  assign n34622 = n34621 ^ n34618 ;
  assign n34626 = n34446 ^ n34445 ;
  assign n34623 = n32052 ^ n1957 ;
  assign n34624 = n34623 ^ n3088 ;
  assign n34625 = n34624 ^ n23096 ;
  assign n34627 = n34626 ^ n34625 ;
  assign n3064 = n3060 ^ n3045 ;
  assign n3077 = n3076 ^ n3064 ;
  assign n3081 = n3080 ^ n3077 ;
  assign n34628 = n34445 ^ n3081 ;
  assign n34630 = n28017 ^ n2782 ;
  assign n34631 = n34630 ^ n3022 ;
  assign n34632 = n34631 ^ n3074 ;
  assign n34051 = n34050 ^ n30907 ;
  assign n34052 = n3010 ^ n2774 ;
  assign n34053 = n34052 ^ n3179 ;
  assign n34054 = n34053 ^ n23528 ;
  assign n34629 = n34051 & n34054 ;
  assign n34633 = n34632 ^ n34629 ;
  assign n34634 = n34366 ^ n34365 ;
  assign n34635 = n34634 ^ n34629 ;
  assign n34636 = n34633 & n34635 ;
  assign n34637 = n34636 ^ n34632 ;
  assign n34638 = n34637 ^ n34445 ;
  assign n34639 = ~n34628 & n34638 ;
  assign n34640 = n34639 ^ n3081 ;
  assign n34641 = n34640 ^ n34625 ;
  assign n34642 = ~n34627 & n34641 ;
  assign n34643 = n34642 ^ n34625 ;
  assign n34644 = n34643 ^ n34618 ;
  assign n34645 = n34622 & ~n34644 ;
  assign n34646 = n34645 ^ n34621 ;
  assign n34647 = n34646 ^ n2064 ;
  assign n34648 = n34617 & ~n34647 ;
  assign n34649 = n34648 ^ n34616 ;
  assign n34650 = n34649 ^ n34613 ;
  assign n34651 = n34615 & ~n34650 ;
  assign n34652 = n34651 ^ n34614 ;
  assign n34653 = n34652 ^ n2165 ;
  assign n34654 = n34610 & ~n34653 ;
  assign n34655 = n34654 ^ n34609 ;
  assign n34656 = n34608 & n34655 ;
  assign n34657 = ~n34602 & n34656 ;
  assign n34660 = n34576 & ~n34580 ;
  assign n34661 = n34657 & n34660 ;
  assign n34658 = n34657 ^ n34569 ;
  assign n34659 = n34658 ^ n34602 ;
  assign n34662 = n34661 ^ n34659 ;
  assign n34663 = ~n34570 & n34662 ;
  assign n34664 = n34663 ^ n34569 ;
  assign n34665 = n34664 ^ n34563 ;
  assign n34666 = ~n34565 & ~n34665 ;
  assign n34667 = n34666 ^ n34564 ;
  assign n34668 = n34667 ^ n34558 ;
  assign n34669 = ~n34560 & n34668 ;
  assign n34670 = n34669 ^ n34559 ;
  assign n34671 = n34670 ^ n34553 ;
  assign n34672 = n34555 & n34671 ;
  assign n34673 = n34672 ^ n34554 ;
  assign n34674 = n34550 & n34673 ;
  assign n34675 = n34674 ^ n34537 ;
  assign n35454 = n34710 ^ n34675 ;
  assign n35455 = n34711 & ~n35454 ;
  assign n35458 = n35457 ^ n35455 ;
  assign n35450 = n33273 ^ n32592 ;
  assign n35192 = n34015 ^ n33829 ;
  assign n35451 = n35192 ^ n33273 ;
  assign n35452 = n35450 & n35451 ;
  assign n35453 = n35452 ^ n32592 ;
  assign n35459 = n35458 ^ n35453 ;
  assign n34062 = n34012 ^ n33834 ;
  assign n34063 = n34062 ^ n33211 ;
  assign n34712 = n34711 ^ n34675 ;
  assign n34713 = n34712 ^ n32593 ;
  assign n34714 = n34713 ^ n34062 ;
  assign n34715 = n34714 ^ n34712 ;
  assign n34716 = n34063 & ~n34715 ;
  assign n34717 = n34716 ^ n34713 ;
  assign n34737 = n34673 ^ n34523 ;
  assign n34742 = n34673 ^ n680 ;
  assign n34743 = ~n34737 & n34742 ;
  assign n34738 = n34522 ^ n680 ;
  assign n34739 = n34738 ^ n34526 ;
  assign n34744 = n34743 ^ n34739 ;
  assign n34723 = n34156 ^ n33294 ;
  assign n34724 = n33854 & n33868 ;
  assign n34725 = ~n34007 & n34724 ;
  assign n34726 = n34725 ^ n33854 ;
  assign n34727 = n34726 ^ n33863 ;
  assign n34728 = n34727 ^ n34156 ;
  assign n34729 = ~n34723 & n34728 ;
  assign n34730 = n34729 ^ n33294 ;
  assign n34745 = n34744 ^ n34730 ;
  assign n34748 = n34007 ^ n33848 ;
  assign n34749 = n33864 & n34748 ;
  assign n34746 = n33850 ^ n964 ;
  assign n34747 = n34746 ^ n1083 ;
  assign n34750 = n34749 ^ n34747 ;
  assign n34751 = n34750 ^ n34147 ;
  assign n34752 = n34673 ^ n34538 ;
  assign n34753 = n34752 ^ n33225 ;
  assign n34754 = n34753 ^ n34752 ;
  assign n34755 = n34754 ^ n34750 ;
  assign n34756 = n34751 & n34755 ;
  assign n34757 = n34756 ^ n34753 ;
  assign n34761 = n34007 ^ n33864 ;
  assign n34762 = n34761 ^ n34027 ;
  assign n34763 = n34027 ^ n32989 ;
  assign n34764 = n34762 & n34763 ;
  assign n34765 = n34764 ^ n32989 ;
  assign n34760 = n34670 ^ n34555 ;
  assign n34766 = n34765 ^ n34760 ;
  assign n34781 = n34667 ^ n34560 ;
  assign n34767 = n33816 ^ n32947 ;
  assign n34768 = ~n33883 & ~n34001 ;
  assign n34769 = ~n33885 & n34768 ;
  assign n34770 = ~n33897 & n34769 ;
  assign n34771 = n34770 ^ n33897 ;
  assign n34772 = n34771 ^ n33876 ;
  assign n34773 = n33891 ^ n33873 ;
  assign n34774 = n34773 ^ n33891 ;
  assign n34775 = n34774 ^ n34771 ;
  assign n34776 = ~n34772 & n34775 ;
  assign n34777 = n34776 ^ n34773 ;
  assign n34778 = n34777 ^ n33816 ;
  assign n34779 = ~n34767 & n34778 ;
  assign n34780 = n34779 ^ n32947 ;
  assign n34782 = n34781 ^ n34780 ;
  assign n35276 = n34664 ^ n34565 ;
  assign n34789 = n34662 ^ n34566 ;
  assign n34783 = ~n33882 & ~n34768 ;
  assign n34784 = n34783 ^ n33895 ;
  assign n34785 = n34784 ^ n32697 ;
  assign n34786 = n34784 ^ n33775 ;
  assign n34787 = n34785 & ~n34786 ;
  assign n34788 = n34787 ^ n32697 ;
  assign n34790 = n34789 ^ n34788 ;
  assign n35256 = ~n34594 & ~n34607 ;
  assign n35257 = n34655 & n35256 ;
  assign n35258 = n35257 ^ n34594 ;
  assign n35264 = n35258 ^ n34576 ;
  assign n35267 = n35258 ^ n34580 ;
  assign n35268 = n35264 & n35267 ;
  assign n35265 = n34580 ^ n34575 ;
  assign n35269 = n35268 ^ n35265 ;
  assign n35272 = n35269 ^ n34789 ;
  assign n35244 = n34680 ^ n32161 ;
  assign n35245 = n34680 ^ n33732 ;
  assign n35246 = ~n35244 & n35245 ;
  assign n35247 = n35246 ^ n32161 ;
  assign n34808 = n34655 ^ n34603 ;
  assign n34804 = n33661 ^ n32138 ;
  assign n34805 = n34489 ^ n32138 ;
  assign n34806 = ~n34804 & ~n34805 ;
  assign n34807 = n34806 ^ n33661 ;
  assign n34809 = n34808 ^ n34807 ;
  assign n34810 = n34329 ^ n32189 ;
  assign n34811 = n34652 ^ n34610 ;
  assign n34812 = n34811 ^ n33543 ;
  assign n34813 = n34812 ^ n34329 ;
  assign n34814 = n34813 ^ n34811 ;
  assign n34815 = n34810 & ~n34814 ;
  assign n34816 = n34815 ^ n34812 ;
  assign n34821 = n34649 ^ n34615 ;
  assign n34817 = n34064 ^ n33328 ;
  assign n34818 = n33328 ^ n32220 ;
  assign n34819 = n34817 & ~n34818 ;
  assign n34820 = n34819 ^ n32220 ;
  assign n34822 = n34821 ^ n34820 ;
  assign n34827 = n34646 ^ n34617 ;
  assign n34823 = n33338 ^ n32204 ;
  assign n34824 = n34075 ^ n33338 ;
  assign n34825 = n34823 & n34824 ;
  assign n34826 = n34825 ^ n32204 ;
  assign n34828 = n34827 ^ n34826 ;
  assign n34833 = n34643 ^ n34622 ;
  assign n34829 = n33340 ^ n32202 ;
  assign n34830 = n34081 ^ n33340 ;
  assign n34831 = n34829 & n34830 ;
  assign n34832 = n34831 ^ n32202 ;
  assign n34834 = n34833 ^ n34832 ;
  assign n35218 = n34640 ^ n34627 ;
  assign n34839 = n34637 ^ n34628 ;
  assign n34835 = n34094 ^ n33364 ;
  assign n34836 = n33364 ^ n32233 ;
  assign n34837 = ~n34835 & n34836 ;
  assign n34838 = n34837 ^ n32233 ;
  assign n34840 = n34839 ^ n34838 ;
  assign n34845 = n34634 ^ n34633 ;
  assign n34841 = n33347 ^ n32240 ;
  assign n34842 = n34118 ^ n33347 ;
  assign n34843 = ~n34841 & ~n34842 ;
  assign n34844 = n34843 ^ n32240 ;
  assign n34846 = n34845 ^ n34844 ;
  assign n34847 = n34095 ^ n33352 ;
  assign n34055 = n34054 ^ n34051 ;
  assign n34848 = n34055 ^ n32246 ;
  assign n34849 = n34848 ^ n34095 ;
  assign n34850 = n34849 ^ n34055 ;
  assign n34851 = ~n34847 & ~n34850 ;
  assign n34852 = n34851 ^ n34848 ;
  assign n35172 = n34113 ^ n33383 ;
  assign n35173 = n33383 ^ n32256 ;
  assign n35174 = n35172 & n35173 ;
  assign n35175 = n35174 ^ n32256 ;
  assign n35030 = n33312 ^ n32583 ;
  assign n34719 = n34010 ^ n33835 ;
  assign n35031 = n34719 ^ n31785 ;
  assign n35032 = n35031 ^ n33312 ;
  assign n35033 = n35032 ^ n34719 ;
  assign n35034 = n35030 & n35033 ;
  assign n35035 = n35034 ^ n35031 ;
  assign n34863 = n33845 ^ n33841 ;
  assign n34861 = n34726 ^ n33842 ;
  assign n34862 = ~n33863 & ~n34861 ;
  assign n34864 = n34863 ^ n34862 ;
  assign n34857 = n32589 ^ n31791 ;
  assign n34858 = n33273 ^ n32589 ;
  assign n34859 = n34857 & ~n34858 ;
  assign n34860 = n34859 ^ n31791 ;
  assign n34865 = n34864 ^ n34860 ;
  assign n34866 = n34174 ^ n31580 ;
  assign n34867 = n32593 ^ n31580 ;
  assign n34868 = ~n34866 & n34867 ;
  assign n34869 = n34868 ^ n32593 ;
  assign n34870 = n34869 ^ n34761 ;
  assign n34871 = n34156 ^ n33462 ;
  assign n34872 = n33462 ^ n32494 ;
  assign n34873 = n34871 & n34872 ;
  assign n34874 = n34873 ^ n32494 ;
  assign n34875 = n34874 ^ n34777 ;
  assign n34876 = n33294 ^ n32286 ;
  assign n34877 = n34027 ^ n33294 ;
  assign n34878 = ~n34876 & ~n34877 ;
  assign n34879 = n34878 ^ n32286 ;
  assign n34880 = n34784 & n34879 ;
  assign n34881 = ~n34680 & n34684 ;
  assign n34883 = n34882 ^ n34881 ;
  assign n34888 = n34887 ^ n34881 ;
  assign n34889 = n34883 & n34888 ;
  assign n34890 = n34889 ^ n34882 ;
  assign n34891 = n34890 ^ n34784 ;
  assign n34892 = n34891 ^ n34695 ;
  assign n34893 = n34892 ^ n34891 ;
  assign n34894 = n34881 ^ n34685 ;
  assign n34895 = ~n34882 & ~n34894 ;
  assign n34896 = n34887 & n34895 ;
  assign n34897 = n34896 ^ n34894 ;
  assign n34898 = ~n34890 & ~n34897 ;
  assign n34901 = n34893 & n34898 ;
  assign n34902 = n34901 ^ n34891 ;
  assign n34903 = n34147 ^ n33426 ;
  assign n34904 = n34147 ^ n32390 ;
  assign n34905 = ~n34903 & n34904 ;
  assign n34906 = n34905 ^ n33426 ;
  assign n34908 = n34906 ^ n34879 ;
  assign n34907 = n34906 ^ n34784 ;
  assign n34909 = n34908 ^ n34907 ;
  assign n34910 = n34902 & n34909 ;
  assign n34911 = n34910 ^ n34908 ;
  assign n34912 = n33876 ^ n33873 ;
  assign n34913 = n34912 ^ n34771 ;
  assign n34914 = n34913 ^ n34906 ;
  assign n34915 = ~n34911 & ~n34914 ;
  assign n34916 = n34915 ^ n34913 ;
  assign n34917 = ~n34897 & ~n34914 ;
  assign n34918 = n34702 & n34917 ;
  assign n34919 = ~n34327 & n34918 ;
  assign n34920 = ~n34916 & n34919 ;
  assign n34923 = n34880 & n34920 ;
  assign n34921 = n34920 ^ n34916 ;
  assign n34924 = n34923 ^ n34921 ;
  assign n34925 = n34924 ^ n34874 ;
  assign n34926 = n34875 & n34925 ;
  assign n34927 = n34926 ^ n34924 ;
  assign n34928 = n34927 ^ n34869 ;
  assign n34929 = ~n34870 & ~n34928 ;
  assign n34930 = n34929 ^ n34761 ;
  assign n34931 = n34930 ^ n34750 ;
  assign n34932 = n32592 ^ n31795 ;
  assign n34933 = n34227 ^ n32592 ;
  assign n34934 = ~n34932 & n34933 ;
  assign n34935 = n34934 ^ n31795 ;
  assign n34936 = n34935 ^ n34930 ;
  assign n34937 = ~n34931 & ~n34936 ;
  assign n34938 = n34937 ^ n34935 ;
  assign n34939 = n34938 ^ n34727 ;
  assign n34940 = n33211 ^ n32591 ;
  assign n34941 = n34727 ^ n31805 ;
  assign n34942 = n34941 ^ n33211 ;
  assign n34943 = n34942 ^ n34727 ;
  assign n34944 = ~n34940 & n34943 ;
  assign n34945 = n34944 ^ n34941 ;
  assign n34946 = n34939 & n34945 ;
  assign n34947 = n34946 ^ n34727 ;
  assign n35027 = n34947 ^ n34864 ;
  assign n35028 = ~n34865 & ~n35027 ;
  assign n35029 = n35028 ^ n34947 ;
  assign n35133 = n35029 ^ n34719 ;
  assign n35134 = n35035 & ~n35133 ;
  assign n35135 = n35134 ^ n34719 ;
  assign n35128 = n31676 ^ n31587 ;
  assign n35129 = n33478 ^ n31587 ;
  assign n35130 = ~n35128 & ~n35129 ;
  assign n35131 = n35130 ^ n31676 ;
  assign n35132 = n35131 ^ n34062 ;
  assign n35136 = n35135 ^ n35132 ;
  assign n35137 = n35136 ^ n31013 ;
  assign n35036 = n35035 ^ n35029 ;
  assign n35037 = n35036 ^ n31071 ;
  assign n34950 = n34945 ^ n34938 ;
  assign n34951 = n34950 ^ n30902 ;
  assign n34952 = n34935 ^ n34750 ;
  assign n34953 = n34952 ^ n34930 ;
  assign n34954 = n34953 ^ n30859 ;
  assign n34956 = n34924 ^ n34875 ;
  assign n34957 = n34956 ^ n31728 ;
  assign n34960 = n34879 ^ n34784 ;
  assign n34958 = n34705 & n34898 ;
  assign n34959 = n34958 ^ n34890 ;
  assign n34961 = n34960 ^ n34959 ;
  assign n34962 = n34961 ^ n31695 ;
  assign n34966 = n34965 ^ n31683 ;
  assign n34974 = n34973 ^ n34965 ;
  assign n34975 = ~n34966 & ~n34974 ;
  assign n34976 = n34975 ^ n31683 ;
  assign n34977 = n34976 ^ n34961 ;
  assign n34978 = ~n34962 & ~n34977 ;
  assign n34979 = n34978 ^ n31695 ;
  assign n34980 = n34979 ^ n31591 ;
  assign n34981 = n34959 ^ n34784 ;
  assign n34982 = n34914 ^ n34879 ;
  assign n34983 = n34982 ^ n34914 ;
  assign n34984 = n34983 ^ n34959 ;
  assign n34985 = n34981 & ~n34984 ;
  assign n34986 = n34985 ^ n34982 ;
  assign n34987 = n34986 ^ n34979 ;
  assign n34988 = n34980 & n34987 ;
  assign n34989 = n34988 ^ n31591 ;
  assign n34990 = n34989 ^ n34956 ;
  assign n34991 = ~n34957 & ~n34990 ;
  assign n34992 = n34991 ^ n31728 ;
  assign n34955 = n34927 ^ n34870 ;
  assign n34993 = n34992 ^ n34955 ;
  assign n34994 = n34992 ^ n30811 ;
  assign n34995 = n34993 & n34994 ;
  assign n34996 = n34995 ^ n30811 ;
  assign n34997 = n34996 ^ n34953 ;
  assign n34998 = n34954 & ~n34997 ;
  assign n34999 = n34998 ^ n30859 ;
  assign n35000 = n34999 ^ n34950 ;
  assign n35001 = ~n34951 & ~n35000 ;
  assign n35002 = n35001 ^ n30902 ;
  assign n34948 = n34947 ^ n34865 ;
  assign n35023 = n35002 ^ n34948 ;
  assign n35024 = n35002 ^ n31074 ;
  assign n35025 = n35023 & ~n35024 ;
  assign n35026 = n35025 ^ n31074 ;
  assign n35125 = n35026 ^ n31071 ;
  assign n35126 = n35037 & n35125 ;
  assign n35127 = n35126 ^ n31071 ;
  assign n35138 = n35137 ^ n35127 ;
  assign n34949 = n34948 ^ n31074 ;
  assign n35003 = n35002 ^ n34949 ;
  assign n35004 = n34999 ^ n34951 ;
  assign n35008 = ~n35005 & n35007 ;
  assign n35009 = n34976 ^ n34962 ;
  assign n35010 = n35008 & ~n35009 ;
  assign n35011 = n34986 ^ n31591 ;
  assign n35012 = n35011 ^ n34979 ;
  assign n35013 = n35010 & n35012 ;
  assign n35014 = n34989 ^ n34957 ;
  assign n35015 = ~n35013 & ~n35014 ;
  assign n35016 = n34955 ^ n30811 ;
  assign n35017 = n35016 ^ n34992 ;
  assign n35018 = n35015 & n35017 ;
  assign n35019 = n34996 ^ n34954 ;
  assign n35020 = n35018 & ~n35019 ;
  assign n35021 = n35004 & n35020 ;
  assign n35022 = ~n35003 & ~n35021 ;
  assign n35038 = n35037 ^ n35026 ;
  assign n35124 = n35022 & n35038 ;
  assign n35139 = n35138 ^ n35124 ;
  assign n3144 = n3143 ^ n2717 ;
  assign n3154 = n3153 ^ n3144 ;
  assign n3158 = n3157 ^ n3154 ;
  assign n35140 = n35139 ^ n3158 ;
  assign n35040 = n32512 ^ n24677 ;
  assign n35041 = n35040 ^ n28582 ;
  assign n35042 = n35041 ^ n3150 ;
  assign n35039 = n35038 ^ n35022 ;
  assign n35043 = n35042 ^ n35039 ;
  assign n35045 = n32523 ^ n24649 ;
  assign n35046 = n35045 ^ n2648 ;
  assign n35047 = n35046 ^ n3212 ;
  assign n35044 = n35020 ^ n35004 ;
  assign n35048 = n35047 ^ n35044 ;
  assign n35052 = n35019 ^ n35018 ;
  assign n35049 = n32527 ^ n24512 ;
  assign n35050 = n35049 ^ n28598 ;
  assign n35051 = n35050 ^ n2558 ;
  assign n35053 = n35052 ^ n35051 ;
  assign n35054 = n35017 ^ n35015 ;
  assign n35058 = n35057 ^ n35054 ;
  assign n35059 = n35014 ^ n35013 ;
  assign n1397 = n1396 ^ n1285 ;
  assign n1398 = n1397 ^ n1369 ;
  assign n1399 = n1398 ^ n1379 ;
  assign n35060 = n35059 ^ n1399 ;
  assign n35061 = n35012 ^ n35010 ;
  assign n35062 = n35061 ^ n1362 ;
  assign n1215 = n1175 ^ n1124 ;
  assign n1216 = n1215 ^ n1212 ;
  assign n1220 = n1219 ^ n1216 ;
  assign n35087 = n35061 ^ n1220 ;
  assign n35063 = n35009 ^ n35008 ;
  assign n35064 = n35063 ^ n1220 ;
  assign n35065 = n1678 & n34710 ;
  assign n35066 = n35065 ^ n1205 ;
  assign n35068 = n35067 ^ n35065 ;
  assign n35069 = n35066 & n35068 ;
  assign n35070 = n35069 ^ n1205 ;
  assign n35074 = n35065 ^ n34711 ;
  assign n35075 = ~n1205 & n35067 ;
  assign n35076 = n35074 & n35075 ;
  assign n35077 = n35076 ^ n35074 ;
  assign n35071 = n35070 ^ n35063 ;
  assign n35080 = n35071 ^ n34537 ;
  assign n35081 = n35080 ^ n35071 ;
  assign n35082 = n35077 & n35081 ;
  assign n35083 = ~n35070 & n35082 ;
  assign n35084 = n35083 ^ n35070 ;
  assign n35072 = n35071 ^ n35070 ;
  assign n35085 = n35084 ^ n35072 ;
  assign n35086 = ~n35064 & n35085 ;
  assign n35088 = n35087 ^ n35086 ;
  assign n35089 = n35062 & n35088 ;
  assign n35090 = n35089 ^ n35061 ;
  assign n35091 = n34675 & n35077 ;
  assign n35092 = n34549 & n35062 ;
  assign n35093 = n35091 & n35092 ;
  assign n35094 = n34673 & n35093 ;
  assign n35095 = ~n35090 & n35094 ;
  assign n35098 = ~n1220 & n35063 ;
  assign n35100 = n35095 & n35098 ;
  assign n35096 = n35095 ^ n35090 ;
  assign n35097 = n35096 ^ n1399 ;
  assign n35101 = n35100 ^ n35097 ;
  assign n35102 = ~n35060 & ~n35101 ;
  assign n35103 = n35102 ^ n35059 ;
  assign n35104 = n35103 ^ n35054 ;
  assign n35105 = ~n35058 & ~n35104 ;
  assign n35106 = n35105 ^ n35057 ;
  assign n35107 = n35106 ^ n35051 ;
  assign n35108 = n35053 & ~n35107 ;
  assign n35109 = n35108 ^ n35052 ;
  assign n35110 = n35109 ^ n35047 ;
  assign n35111 = ~n35048 & n35110 ;
  assign n35112 = n35111 ^ n35047 ;
  assign n35116 = n35115 ^ n35112 ;
  assign n35117 = n35021 ^ n35003 ;
  assign n35118 = n35117 ^ n35115 ;
  assign n35119 = n35116 & n35118 ;
  assign n35120 = n35119 ^ n35115 ;
  assign n35121 = n35120 ^ n35039 ;
  assign n35122 = n35043 & ~n35121 ;
  assign n35123 = n35122 ^ n35042 ;
  assign n35141 = n35140 ^ n35123 ;
  assign n34853 = n34109 ^ n33385 ;
  assign n34854 = n33385 ^ n32259 ;
  assign n34855 = n34853 & n34854 ;
  assign n34856 = n34855 ^ n32259 ;
  assign n35142 = n35141 ^ n34856 ;
  assign n35144 = n33391 ^ n33325 ;
  assign n35145 = n33391 ^ n32265 ;
  assign n35146 = n35144 & n35145 ;
  assign n35147 = n35146 ^ n32265 ;
  assign n35143 = n35120 ^ n35043 ;
  assign n35148 = n35147 ^ n35143 ;
  assign n35155 = n35118 ^ n35112 ;
  assign n35149 = n35109 ^ n35048 ;
  assign n35150 = n33326 ^ n32275 ;
  assign n35151 = n34130 ^ n32275 ;
  assign n35152 = ~n35150 & n35151 ;
  assign n35153 = n35152 ^ n33326 ;
  assign n35154 = ~n35149 & ~n35153 ;
  assign n35156 = n35155 ^ n35154 ;
  assign n35157 = n34280 ^ n33401 ;
  assign n35158 = n35154 ^ n32639 ;
  assign n35159 = n35158 ^ n34280 ;
  assign n35160 = n35159 ^ n35154 ;
  assign n35161 = n35157 & n35160 ;
  assign n35162 = n35161 ^ n35158 ;
  assign n35163 = n35156 & ~n35162 ;
  assign n35164 = n35163 ^ n35155 ;
  assign n35165 = n35164 ^ n35143 ;
  assign n35166 = n35148 & ~n35165 ;
  assign n35167 = n35166 ^ n35147 ;
  assign n35168 = n35167 ^ n34856 ;
  assign n35169 = n35142 & ~n35168 ;
  assign n35170 = n35169 ^ n35141 ;
  assign n35176 = n35175 ^ n35170 ;
  assign n35196 = n32501 ^ n2723 ;
  assign n35197 = n35196 ^ n28571 ;
  assign n35198 = n35197 ^ n1844 ;
  assign n35193 = n35131 ^ n31011 ;
  assign n35194 = n35193 ^ n31824 ;
  assign n35195 = n35194 ^ n35192 ;
  assign n35199 = n35198 ^ n35195 ;
  assign n35189 = n33472 ^ n32626 ;
  assign n35190 = n32626 ^ n31824 ;
  assign n35191 = ~n35189 & n35190 ;
  assign n35200 = n35199 ^ n35191 ;
  assign n35183 = n35136 ^ n35127 ;
  assign n35186 = n35127 ^ n35124 ;
  assign n35187 = ~n35183 & ~n35186 ;
  assign n35184 = n35183 ^ n35124 ;
  assign n35185 = ~n31013 & n35184 ;
  assign n35188 = n35187 ^ n35185 ;
  assign n35201 = n35200 ^ n35188 ;
  assign n35202 = n35201 ^ n3158 ;
  assign n35181 = n35135 ^ n35131 ;
  assign n35182 = ~n35132 & ~n35181 ;
  assign n35203 = n35202 ^ n35182 ;
  assign n35179 = n35123 ^ n3158 ;
  assign n35180 = n35140 & n35179 ;
  assign n35204 = n35203 ^ n35180 ;
  assign n35205 = n35204 ^ n34055 ;
  assign n35171 = n35170 ^ n34055 ;
  assign n35206 = n35205 ^ n35171 ;
  assign n35207 = n35176 & ~n35206 ;
  assign n35208 = n35207 ^ n35171 ;
  assign n35209 = ~n34852 & n35208 ;
  assign n35210 = n35209 ^ n34055 ;
  assign n35211 = n35210 ^ n34844 ;
  assign n35212 = ~n34846 & ~n35211 ;
  assign n35213 = n35212 ^ n34845 ;
  assign n35214 = n35213 ^ n34838 ;
  assign n35215 = ~n34840 & n35214 ;
  assign n35216 = n35215 ^ n34839 ;
  assign n35219 = n35218 ^ n35216 ;
  assign n35220 = n34088 ^ n33341 ;
  assign n35221 = n35218 ^ n32667 ;
  assign n35222 = n35221 ^ n34088 ;
  assign n35223 = n35222 ^ n35218 ;
  assign n35224 = ~n35220 & n35223 ;
  assign n35225 = n35224 ^ n35221 ;
  assign n35226 = n35219 & ~n35225 ;
  assign n35217 = n35216 ^ n34832 ;
  assign n35227 = n35226 ^ n35217 ;
  assign n35228 = n34834 & n35227 ;
  assign n35229 = n35228 ^ n34833 ;
  assign n35230 = n35229 ^ n34826 ;
  assign n35231 = n34828 & ~n35230 ;
  assign n35232 = n35231 ^ n34827 ;
  assign n35233 = n35232 ^ n34820 ;
  assign n35234 = ~n34822 & n35233 ;
  assign n35235 = n35234 ^ n34821 ;
  assign n35236 = n35235 ^ n34811 ;
  assign n35237 = n34816 & n35236 ;
  assign n35238 = n35237 ^ n34811 ;
  assign n35239 = n35238 ^ n34808 ;
  assign n35240 = n34809 & ~n35239 ;
  assign n35241 = n35240 ^ n35238 ;
  assign n35248 = n35247 ^ n35241 ;
  assign n34795 = n34655 ^ n34586 ;
  assign n34800 = n34655 ^ n34583 ;
  assign n34801 = ~n34795 & ~n34800 ;
  assign n34796 = n34583 ^ n34582 ;
  assign n34797 = n34796 ^ n34591 ;
  assign n34802 = n34801 ^ n34797 ;
  assign n34791 = n33712 ^ n32145 ;
  assign n34792 = n34503 ^ n32145 ;
  assign n34793 = ~n34791 & n34792 ;
  assign n34794 = n34793 ^ n33712 ;
  assign n34803 = n34802 ^ n34794 ;
  assign n35242 = n35241 ^ n34802 ;
  assign n35243 = n34803 & ~n35242 ;
  assign n35249 = n35248 ^ n35243 ;
  assign n35255 = n34580 ^ n34576 ;
  assign n35259 = n35258 ^ n35255 ;
  assign n35250 = n33747 ^ n32129 ;
  assign n35251 = n34882 ^ n32129 ;
  assign n35252 = ~n35250 & n35251 ;
  assign n35253 = n35252 ^ n33747 ;
  assign n35254 = n35253 ^ n35247 ;
  assign n35260 = n35259 ^ n35254 ;
  assign n35261 = n35260 ^ n35253 ;
  assign n35262 = n35249 & ~n35261 ;
  assign n35263 = n35262 ^ n35254 ;
  assign n35270 = n35269 ^ n35253 ;
  assign n35271 = ~n35263 & ~n35270 ;
  assign n35273 = n35272 ^ n35271 ;
  assign n35274 = n34790 & n35273 ;
  assign n35275 = n35274 ^ n34789 ;
  assign n35277 = n35276 ^ n35275 ;
  assign n35278 = n34913 ^ n33793 ;
  assign n35279 = n35276 ^ n32933 ;
  assign n35280 = n35279 ^ n34913 ;
  assign n35281 = n35280 ^ n35276 ;
  assign n35282 = n35278 & n35281 ;
  assign n35283 = n35282 ^ n35279 ;
  assign n35284 = n35277 & ~n35283 ;
  assign n35285 = n35284 ^ n35276 ;
  assign n35286 = n35285 ^ n34780 ;
  assign n35287 = ~n34782 & ~n35286 ;
  assign n35288 = n35287 ^ n34781 ;
  assign n35289 = n35288 ^ n34760 ;
  assign n35290 = ~n34766 & n35289 ;
  assign n35291 = n35290 ^ n34765 ;
  assign n35292 = n35291 ^ n34752 ;
  assign n35293 = ~n34757 & n35292 ;
  assign n34758 = n34752 ^ n34730 ;
  assign n35294 = n35293 ^ n34758 ;
  assign n35295 = ~n34745 & n35294 ;
  assign n34732 = ~n34529 & n34542 ;
  assign n34733 = n34673 & n34732 ;
  assign n34734 = n34733 ^ n34529 ;
  assign n34731 = n34517 ^ n34514 ;
  assign n34735 = n34734 ^ n34731 ;
  assign n34736 = n34735 ^ n34730 ;
  assign n35296 = n35295 ^ n34736 ;
  assign n35297 = n34864 ^ n33426 ;
  assign n35298 = n34864 ^ n34174 ;
  assign n35299 = n35297 & n35298 ;
  assign n35300 = n35299 ^ n33426 ;
  assign n35301 = n35300 ^ n34735 ;
  assign n35302 = n35296 & ~n35301 ;
  assign n35303 = n35302 ^ n34735 ;
  assign n34718 = n34227 ^ n33462 ;
  assign n34720 = n34719 ^ n34227 ;
  assign n34721 = n34718 & n34720 ;
  assign n34722 = n34721 ^ n33462 ;
  assign n35304 = n35303 ^ n34722 ;
  assign n35307 = n34517 ^ n34513 ;
  assign n35305 = n34734 ^ n34514 ;
  assign n35306 = n34731 & ~n35305 ;
  assign n35308 = n35307 ^ n35306 ;
  assign n35309 = n35308 ^ n34722 ;
  assign n35310 = n35304 & n35309 ;
  assign n35311 = n35310 ^ n35303 ;
  assign n35447 = n35311 ^ n34712 ;
  assign n35448 = n34717 & n35447 ;
  assign n35449 = n35448 ^ n34712 ;
  assign n35460 = n35459 ^ n35449 ;
  assign n35461 = n35460 ^ n31795 ;
  assign n35313 = n35309 ^ n35303 ;
  assign n35314 = n35313 ^ n32494 ;
  assign n35316 = n35294 ^ n34744 ;
  assign n35317 = n35316 ^ n32286 ;
  assign n35319 = n35288 ^ n34766 ;
  assign n35320 = n35319 ^ n32133 ;
  assign n35421 = n35285 ^ n34782 ;
  assign n35321 = n35283 ^ n35275 ;
  assign n35322 = n35321 ^ n32140 ;
  assign n35324 = n35269 ^ n35263 ;
  assign n35325 = n35324 ^ n32193 ;
  assign n35401 = n35241 ^ n34803 ;
  assign n35326 = n35238 ^ n34809 ;
  assign n35327 = n35326 ^ n32311 ;
  assign n35389 = n35232 ^ n34822 ;
  assign n35330 = n35216 ^ n34834 ;
  assign n35331 = n35330 ^ n35226 ;
  assign n35332 = n35331 ^ n31611 ;
  assign n35376 = n35225 ^ n35216 ;
  assign n35333 = n35213 ^ n34840 ;
  assign n35334 = n35333 ^ n31625 ;
  assign n35367 = n35210 ^ n34846 ;
  assign n35342 = n35167 ^ n35142 ;
  assign n35343 = n35342 ^ n31653 ;
  assign n35351 = n35164 ^ n35148 ;
  assign n35344 = n35153 ^ n35149 ;
  assign n35345 = n30906 & n35344 ;
  assign n35346 = n35345 ^ n31665 ;
  assign n35347 = n35162 ^ n35155 ;
  assign n35348 = n35347 ^ n35345 ;
  assign n35349 = n35346 & ~n35348 ;
  assign n35350 = n35349 ^ n31665 ;
  assign n35352 = n35351 ^ n35350 ;
  assign n35353 = n35351 ^ n31659 ;
  assign n35354 = ~n35352 & ~n35353 ;
  assign n35355 = n35354 ^ n31659 ;
  assign n35356 = n35355 ^ n35342 ;
  assign n35357 = n35343 & n35356 ;
  assign n35358 = n35357 ^ n31653 ;
  assign n35340 = n35204 ^ n35175 ;
  assign n35341 = n35340 ^ n35170 ;
  assign n35359 = n35358 ^ n35341 ;
  assign n35360 = n35358 ^ n31647 ;
  assign n35361 = n35359 & n35360 ;
  assign n35362 = n35361 ^ n31647 ;
  assign n35335 = n35204 ^ n34852 ;
  assign n35336 = n35335 ^ n35170 ;
  assign n35337 = n35336 ^ n34852 ;
  assign n35338 = ~n35176 & ~n35337 ;
  assign n35339 = n35338 ^ n35335 ;
  assign n35363 = n35362 ^ n35339 ;
  assign n35364 = n35362 ^ n31641 ;
  assign n35365 = ~n35363 & ~n35364 ;
  assign n35366 = n35365 ^ n31641 ;
  assign n35368 = n35367 ^ n35366 ;
  assign n35369 = n35333 ^ n31635 ;
  assign n35370 = n35369 ^ n35333 ;
  assign n35371 = n35370 ^ n35366 ;
  assign n35372 = ~n35368 & n35371 ;
  assign n35373 = n35372 ^ n35369 ;
  assign n35374 = ~n35334 & n35373 ;
  assign n35375 = n35374 ^ n31625 ;
  assign n35377 = n35376 ^ n35375 ;
  assign n35378 = n31618 ^ n31611 ;
  assign n35379 = n35378 ^ n35375 ;
  assign n35380 = n35379 ^ n31611 ;
  assign n35381 = ~n35377 & n35380 ;
  assign n35382 = n35381 ^ n35378 ;
  assign n35383 = n35332 & ~n35382 ;
  assign n35384 = n35383 ^ n35331 ;
  assign n35329 = n35229 ^ n34828 ;
  assign n35385 = n35384 ^ n35329 ;
  assign n35386 = n35384 ^ n31943 ;
  assign n35387 = n35385 & ~n35386 ;
  assign n35388 = n35387 ^ n31943 ;
  assign n35390 = n35389 ^ n35388 ;
  assign n35391 = n35389 ^ n32114 ;
  assign n35392 = n35390 & ~n35391 ;
  assign n35393 = n35392 ^ n32114 ;
  assign n35328 = n35235 ^ n34816 ;
  assign n35394 = n35393 ^ n35328 ;
  assign n35395 = n35393 ^ n32234 ;
  assign n35396 = ~n35394 & ~n35395 ;
  assign n35397 = n35396 ^ n32234 ;
  assign n35398 = n35397 ^ n35326 ;
  assign n35399 = n35327 & ~n35398 ;
  assign n35400 = n35399 ^ n32311 ;
  assign n35402 = n35401 ^ n35400 ;
  assign n35403 = n35401 ^ n32197 ;
  assign n35404 = ~n35402 & ~n35403 ;
  assign n35405 = n35404 ^ n32197 ;
  assign n35406 = n35405 ^ n32212 ;
  assign n35407 = n35259 ^ n35249 ;
  assign n35408 = n35407 ^ n32212 ;
  assign n35409 = n35406 & n35408 ;
  assign n35410 = n35409 ^ n35407 ;
  assign n35411 = n35410 ^ n35324 ;
  assign n35412 = n35325 & ~n35411 ;
  assign n35413 = n35412 ^ n32193 ;
  assign n35323 = n35273 ^ n34788 ;
  assign n35414 = n35413 ^ n35323 ;
  assign n35415 = n35323 ^ n32185 ;
  assign n35416 = n35414 & ~n35415 ;
  assign n35417 = n35416 ^ n35413 ;
  assign n35418 = n35417 ^ n35321 ;
  assign n35419 = n35322 & n35418 ;
  assign n35420 = n35419 ^ n32140 ;
  assign n35422 = n35421 ^ n35420 ;
  assign n35423 = n35420 ^ n32151 ;
  assign n35424 = n35422 & ~n35423 ;
  assign n35425 = n35424 ^ n35421 ;
  assign n35426 = n35425 ^ n35319 ;
  assign n35427 = ~n35320 & n35426 ;
  assign n35428 = n35427 ^ n32133 ;
  assign n35318 = n35291 ^ n34757 ;
  assign n35429 = n35428 ^ n35318 ;
  assign n35430 = n35318 ^ n31603 ;
  assign n35431 = ~n35429 & ~n35430 ;
  assign n35432 = n35431 ^ n35428 ;
  assign n35433 = n35432 ^ n35316 ;
  assign n35434 = n35317 & n35433 ;
  assign n35435 = n35434 ^ n32286 ;
  assign n35315 = n35300 ^ n35296 ;
  assign n35436 = n35435 ^ n35315 ;
  assign n35437 = n35315 ^ n32390 ;
  assign n35438 = n35436 & ~n35437 ;
  assign n35439 = n35438 ^ n35435 ;
  assign n35440 = n35439 ^ n35313 ;
  assign n35441 = ~n35314 & ~n35440 ;
  assign n35442 = n35441 ^ n32494 ;
  assign n35312 = n35311 ^ n34717 ;
  assign n35443 = n35442 ^ n35312 ;
  assign n35444 = n35312 ^ n31580 ;
  assign n35445 = n35443 & ~n35444 ;
  assign n35446 = n35445 ^ n35442 ;
  assign n35462 = n35461 ^ n35446 ;
  assign n35463 = n35442 ^ n31580 ;
  assign n35464 = n35463 ^ n35312 ;
  assign n35465 = n35428 ^ n31603 ;
  assign n35466 = n35465 ^ n35318 ;
  assign n35467 = n35423 ^ n35421 ;
  assign n35468 = n35417 ^ n35322 ;
  assign n35469 = n35339 ^ n31641 ;
  assign n35470 = n35469 ^ n35362 ;
  assign n35471 = n35360 ^ n35341 ;
  assign n35472 = n35353 ^ n35350 ;
  assign n35473 = n35355 ^ n35343 ;
  assign n35474 = n35472 & n35473 ;
  assign n35475 = n35471 & n35474 ;
  assign n35476 = ~n35470 & ~n35475 ;
  assign n35477 = n35367 ^ n31635 ;
  assign n35478 = n35477 ^ n35366 ;
  assign n35479 = ~n35476 & n35478 ;
  assign n35480 = n35373 ^ n31625 ;
  assign n35481 = n35479 & ~n35480 ;
  assign n35482 = n35376 ^ n31618 ;
  assign n35483 = n35482 ^ n35375 ;
  assign n35484 = ~n35481 & ~n35483 ;
  assign n35485 = n35382 ^ n35331 ;
  assign n35486 = n35484 & ~n35485 ;
  assign n35487 = n35329 ^ n31943 ;
  assign n35488 = n35487 ^ n35384 ;
  assign n35489 = ~n35486 & n35488 ;
  assign n35490 = n35388 ^ n32114 ;
  assign n35491 = n35490 ^ n35389 ;
  assign n35492 = n35489 & n35491 ;
  assign n35493 = n35328 ^ n32234 ;
  assign n35494 = n35493 ^ n35393 ;
  assign n35495 = n35492 & n35494 ;
  assign n35496 = n35397 ^ n32311 ;
  assign n35497 = n35496 ^ n35326 ;
  assign n35498 = n35495 & n35497 ;
  assign n35499 = n35400 ^ n32197 ;
  assign n35500 = n35499 ^ n35401 ;
  assign n35501 = ~n35498 & n35500 ;
  assign n35502 = n35407 ^ n35406 ;
  assign n35503 = ~n35501 & ~n35502 ;
  assign n35504 = n35410 ^ n35325 ;
  assign n35505 = n35503 & n35504 ;
  assign n35506 = n35413 ^ n32185 ;
  assign n35507 = n35506 ^ n35323 ;
  assign n35508 = n35505 & n35507 ;
  assign n35509 = ~n35468 & ~n35508 ;
  assign n35510 = ~n35467 & ~n35509 ;
  assign n35511 = n35425 ^ n35320 ;
  assign n35512 = n35510 & n35511 ;
  assign n35513 = n35466 & ~n35512 ;
  assign n35514 = n35432 ^ n35317 ;
  assign n35515 = n35513 & n35514 ;
  assign n35516 = n35435 ^ n32390 ;
  assign n35517 = n35516 ^ n35315 ;
  assign n35518 = n35515 & ~n35517 ;
  assign n35519 = n35439 ^ n35314 ;
  assign n35520 = ~n35518 & ~n35519 ;
  assign n35521 = ~n35464 & n35520 ;
  assign n35725 = ~n35462 & n35521 ;
  assign n35715 = n34045 ^ n33312 ;
  assign n35716 = ~n35070 & ~n35091 ;
  assign n35717 = n35716 ^ n35064 ;
  assign n35718 = n35717 ^ n32591 ;
  assign n35719 = n35718 ^ n34045 ;
  assign n35720 = n35719 ^ n35717 ;
  assign n35721 = ~n35715 & ~n35720 ;
  assign n35722 = n35721 ^ n35718 ;
  assign n35712 = n35453 ^ n35449 ;
  assign n35713 = n35459 & n35712 ;
  assign n35714 = n35713 ^ n35458 ;
  assign n35723 = n35722 ^ n35714 ;
  assign n35708 = n35460 ^ n35446 ;
  assign n35709 = n35461 & ~n35708 ;
  assign n35710 = n35709 ^ n31795 ;
  assign n35711 = n35710 ^ n31805 ;
  assign n35724 = n35723 ^ n35711 ;
  assign n35726 = n35725 ^ n35724 ;
  assign n35727 = n35726 ^ n34061 ;
  assign n35522 = n35521 ^ n35462 ;
  assign n35523 = n35522 ^ n34061 ;
  assign n35524 = n35520 ^ n35464 ;
  assign n35525 = n35524 ^ n2850 ;
  assign n35527 = n2797 ^ n1428 ;
  assign n35528 = n35527 ^ n29387 ;
  assign n35529 = n35528 ^ n2837 ;
  assign n35526 = n35519 ^ n35518 ;
  assign n35530 = n35529 ^ n35526 ;
  assign n35532 = n1420 ^ n1321 ;
  assign n35533 = n35532 ^ n1746 ;
  assign n35534 = n35533 ^ n1259 ;
  assign n35699 = n35534 ^ n35529 ;
  assign n35531 = n35517 ^ n35515 ;
  assign n35535 = n35534 ^ n35531 ;
  assign n35536 = n35514 ^ n35513 ;
  assign n1734 = n1715 ^ n1306 ;
  assign n1735 = n1734 ^ n1070 ;
  assign n1739 = n1738 ^ n1735 ;
  assign n35537 = n35536 ^ n1739 ;
  assign n1725 = n1709 ^ n1297 ;
  assign n1729 = n1728 ^ n1725 ;
  assign n1730 = n1729 ^ n1064 ;
  assign n35693 = n1739 ^ n1730 ;
  assign n35538 = n35512 ^ n35466 ;
  assign n35539 = n35538 ^ n1730 ;
  assign n35540 = n35511 ^ n35510 ;
  assign n909 = n908 ^ n857 ;
  assign n922 = n921 ^ n909 ;
  assign n929 = n928 ^ n922 ;
  assign n35541 = n35540 ^ n929 ;
  assign n35543 = n33051 ^ n1686 ;
  assign n35544 = n35543 ^ n826 ;
  assign n35545 = n35544 ^ n919 ;
  assign n35687 = n35545 ^ n929 ;
  assign n35542 = n35509 ^ n35467 ;
  assign n35546 = n35545 ^ n35542 ;
  assign n35684 = n35545 ^ n819 ;
  assign n35547 = n35508 ^ n35468 ;
  assign n35548 = n35547 ^ n819 ;
  assign n35552 = n35507 ^ n35505 ;
  assign n35553 = n35552 ^ n35551 ;
  assign n35554 = n35504 ^ n35503 ;
  assign n35555 = n35554 ^ n1574 ;
  assign n35559 = n35500 ^ n35498 ;
  assign n35556 = n33092 ^ n29416 ;
  assign n35557 = n35556 ^ n1530 ;
  assign n35558 = n35557 ^ n2951 ;
  assign n35560 = n35559 ^ n35558 ;
  assign n35569 = n35497 ^ n35495 ;
  assign n35566 = n33097 ^ n25051 ;
  assign n35567 = n35566 ^ n2939 ;
  assign n35568 = n35567 ^ n23877 ;
  assign n35570 = n35569 ^ n35568 ;
  assign n35574 = n35491 ^ n35489 ;
  assign n35658 = n35657 ^ n35574 ;
  assign n35571 = n33107 ^ n2921 ;
  assign n35572 = n35571 ^ n28875 ;
  assign n35573 = n35572 ^ n23944 ;
  assign n35575 = n35574 ^ n35573 ;
  assign n35576 = n33112 ^ n24991 ;
  assign n35577 = n35576 ^ n2395 ;
  assign n35578 = n35577 ^ n23884 ;
  assign n35652 = n35578 ^ n35573 ;
  assign n35579 = n35488 ^ n35486 ;
  assign n35580 = n35579 ^ n35578 ;
  assign n35581 = n35485 ^ n35484 ;
  assign n2380 = n2373 ^ n2310 ;
  assign n2387 = n2386 ^ n2380 ;
  assign n2391 = n2390 ^ n2387 ;
  assign n35582 = n35581 ^ n2391 ;
  assign n2270 = n2233 ^ n2200 ;
  assign n2271 = n2270 ^ n2267 ;
  assign n2278 = n2277 ^ n2271 ;
  assign n35646 = n2391 ^ n2278 ;
  assign n35583 = n35483 ^ n35481 ;
  assign n35584 = n35583 ^ n2278 ;
  assign n35585 = n35480 ^ n35479 ;
  assign n2237 = n2224 ^ n2185 ;
  assign n2253 = n2252 ^ n2237 ;
  assign n2260 = n2259 ^ n2253 ;
  assign n35586 = n35585 ^ n2260 ;
  assign n35588 = n33124 ^ n2123 ;
  assign n35589 = n35588 ^ n28890 ;
  assign n35590 = n35589 ^ n2249 ;
  assign n35640 = n35590 ^ n2260 ;
  assign n35587 = n35478 ^ n35476 ;
  assign n35591 = n35590 ^ n35587 ;
  assign n35595 = n35475 ^ n35470 ;
  assign n35592 = n33128 ^ n2111 ;
  assign n35593 = n35592 ^ n28894 ;
  assign n35594 = n35593 ^ n23898 ;
  assign n35596 = n35595 ^ n35594 ;
  assign n35622 = n28899 ^ n25009 ;
  assign n35623 = n35622 ^ n33134 ;
  assign n35624 = n35623 ^ n23902 ;
  assign n35634 = n35624 ^ n35594 ;
  assign n35610 = n33147 ^ n24700 ;
  assign n35611 = n35610 ^ n1868 ;
  assign n35612 = n35611 ^ n23907 ;
  assign n35600 = n35347 ^ n35346 ;
  assign n35597 = n33142 ^ n24696 ;
  assign n35598 = n35597 ^ n28904 ;
  assign n35599 = n35598 ^ n1863 ;
  assign n35601 = n35600 ^ n35599 ;
  assign n35605 = n35344 ^ n30906 ;
  assign n35606 = n35604 & n35605 ;
  assign n35607 = n35606 ^ n35599 ;
  assign n35608 = n35601 & ~n35607 ;
  assign n35609 = n35608 ^ n35600 ;
  assign n35613 = n35612 ^ n35609 ;
  assign n35619 = n35609 ^ n35472 ;
  assign n35620 = ~n35613 & n35619 ;
  assign n35614 = n33138 ^ n25018 ;
  assign n35615 = n35614 ^ n28915 ;
  assign n35616 = n35615 ^ n1910 ;
  assign n35617 = n35616 ^ n35472 ;
  assign n35621 = n35620 ^ n35617 ;
  assign n35627 = n35624 ^ n35616 ;
  assign n35625 = n35473 ^ n35472 ;
  assign n35626 = n35625 ^ n35624 ;
  assign n35628 = n35627 ^ n35626 ;
  assign n35629 = n35621 & ~n35628 ;
  assign n35630 = n35629 ^ n35627 ;
  assign n35631 = n35474 ^ n35471 ;
  assign n35632 = n35631 ^ n35624 ;
  assign n35633 = n35630 & ~n35632 ;
  assign n35635 = n35634 ^ n35633 ;
  assign n35636 = n35596 & ~n35635 ;
  assign n35637 = n35636 ^ n35595 ;
  assign n35638 = n35637 ^ n35590 ;
  assign n35639 = n35591 & n35638 ;
  assign n35641 = n35640 ^ n35639 ;
  assign n35642 = n35586 & n35641 ;
  assign n35643 = n35642 ^ n2260 ;
  assign n35644 = n35643 ^ n2278 ;
  assign n35645 = n35584 & n35644 ;
  assign n35647 = n35646 ^ n35645 ;
  assign n35648 = ~n35582 & ~n35647 ;
  assign n35649 = n35648 ^ n35581 ;
  assign n35650 = n35649 ^ n35578 ;
  assign n35651 = n35580 & ~n35650 ;
  assign n35653 = n35652 ^ n35651 ;
  assign n35654 = ~n35575 & ~n35653 ;
  assign n35659 = n35658 ^ n35654 ;
  assign n35662 = n35657 ^ n35568 ;
  assign n35660 = n35494 ^ n35492 ;
  assign n35661 = n35660 ^ n35568 ;
  assign n35663 = n35662 ^ n35661 ;
  assign n35664 = ~n35659 & ~n35663 ;
  assign n35665 = n35664 ^ n35662 ;
  assign n35666 = ~n35570 & ~n35665 ;
  assign n35667 = n35666 ^ n35569 ;
  assign n35668 = n35667 ^ n35558 ;
  assign n35669 = ~n35560 & ~n35668 ;
  assign n35564 = n35563 ^ n35558 ;
  assign n35670 = n35669 ^ n35564 ;
  assign n35672 = n35502 ^ n35501 ;
  assign n35673 = n35672 ^ n35554 ;
  assign n35671 = n35563 ^ n35554 ;
  assign n35674 = n35673 ^ n35671 ;
  assign n35675 = n35670 & ~n35674 ;
  assign n35676 = n35675 ^ n35671 ;
  assign n35677 = ~n35555 & ~n35676 ;
  assign n35678 = n35677 ^ n35554 ;
  assign n35679 = n35678 ^ n35551 ;
  assign n35680 = ~n35553 & n35679 ;
  assign n35681 = n35680 ^ n35552 ;
  assign n35682 = n35681 ^ n819 ;
  assign n35683 = n35548 & ~n35682 ;
  assign n35685 = n35684 ^ n35683 ;
  assign n35686 = ~n35546 & n35685 ;
  assign n35688 = n35687 ^ n35686 ;
  assign n35689 = ~n35541 & ~n35688 ;
  assign n35690 = n35689 ^ n35540 ;
  assign n35691 = n35690 ^ n1730 ;
  assign n35692 = ~n35539 & ~n35691 ;
  assign n35694 = n35693 ^ n35692 ;
  assign n35695 = n35537 & ~n35694 ;
  assign n35696 = n35695 ^ n35536 ;
  assign n35697 = n35696 ^ n35534 ;
  assign n35698 = ~n35535 & n35697 ;
  assign n35700 = n35699 ^ n35698 ;
  assign n35701 = ~n35530 & n35700 ;
  assign n35702 = n35701 ^ n35529 ;
  assign n35703 = n35702 ^ n2850 ;
  assign n35704 = n35525 & ~n35703 ;
  assign n35705 = n35704 ^ n35524 ;
  assign n35706 = n35705 ^ n34061 ;
  assign n35707 = n35523 & n35706 ;
  assign n35728 = n35727 ^ n35707 ;
  assign n35732 = n35731 ^ n35728 ;
  assign n33327 = n33326 ^ n33325 ;
  assign n34056 = n34055 ^ n33325 ;
  assign n34057 = n33327 & n34056 ;
  assign n34058 = n34057 ^ n33326 ;
  assign n35733 = n35732 ^ n34058 ;
  assign n35777 = n32275 & n35733 ;
  assign n35778 = n35777 ^ n32639 ;
  assign n35771 = n33006 ^ n3215 ;
  assign n35772 = n35771 ^ n29378 ;
  assign n35773 = n35772 ^ n2592 ;
  assign n35758 = n33478 ^ n32589 ;
  assign n35759 = n34257 ^ n33478 ;
  assign n35760 = n35758 & ~n35759 ;
  assign n35761 = n35760 ^ n32589 ;
  assign n35762 = n35761 ^ n35717 ;
  assign n35763 = n35762 ^ n35761 ;
  assign n35764 = n35763 ^ n35714 ;
  assign n35765 = n35722 & ~n35764 ;
  assign n35766 = n35765 ^ n35762 ;
  assign n35752 = n35716 ^ n1220 ;
  assign n35755 = n35716 ^ n35063 ;
  assign n35756 = n35752 & n35755 ;
  assign n35753 = n35063 ^ n35062 ;
  assign n35757 = n35756 ^ n35753 ;
  assign n35767 = n35766 ^ n35757 ;
  assign n35768 = n35767 ^ n31791 ;
  assign n35748 = n35723 ^ n35710 ;
  assign n35749 = n35723 ^ n31805 ;
  assign n35750 = n35748 & ~n35749 ;
  assign n35751 = n35750 ^ n31805 ;
  assign n35769 = n35768 ^ n35751 ;
  assign n35747 = n35724 & n35725 ;
  assign n35770 = n35769 ^ n35747 ;
  assign n35774 = n35773 ^ n35770 ;
  assign n35744 = n35731 ^ n35726 ;
  assign n35745 = n35728 & ~n35744 ;
  assign n35746 = n35745 ^ n35731 ;
  assign n35775 = n35774 ^ n35746 ;
  assign n35737 = n34845 ^ n34109 ;
  assign n35738 = ~n34058 & ~n35732 ;
  assign n35739 = n35738 ^ n33401 ;
  assign n35740 = n35739 ^ n34845 ;
  assign n35741 = n35740 ^ n35738 ;
  assign n35742 = ~n35737 & n35741 ;
  assign n35743 = n35742 ^ n35739 ;
  assign n35776 = n35775 ^ n35743 ;
  assign n35819 = n35777 ^ n35776 ;
  assign n35820 = n35778 & n35819 ;
  assign n35821 = n35820 ^ n32639 ;
  assign n35822 = n35821 ^ n32265 ;
  assign n35813 = n34839 ^ n34113 ;
  assign n35814 = n34839 ^ n33391 ;
  assign n35815 = ~n35813 & ~n35814 ;
  assign n35816 = n35815 ^ n33391 ;
  assign n35810 = ~n35747 & ~n35769 ;
  assign n35807 = n35101 ^ n35059 ;
  assign n35798 = n34255 ^ n33472 ;
  assign n35799 = n35761 ^ n35757 ;
  assign n35800 = ~n35766 & n35799 ;
  assign n35801 = n35800 ^ n35761 ;
  assign n35802 = n35801 ^ n32583 ;
  assign n35803 = n35802 ^ n34255 ;
  assign n35804 = n35803 ^ n35801 ;
  assign n35805 = n35798 & ~n35804 ;
  assign n35806 = n35805 ^ n35802 ;
  assign n35808 = n35807 ^ n35806 ;
  assign n35794 = n35767 ^ n35751 ;
  assign n35795 = ~n35768 & ~n35794 ;
  assign n35796 = n35795 ^ n31791 ;
  assign n35797 = n35796 ^ n31785 ;
  assign n35809 = n35808 ^ n35797 ;
  assign n35811 = n35810 ^ n35809 ;
  assign n35791 = n35773 ^ n35746 ;
  assign n35792 = n35774 & n35791 ;
  assign n2655 = n2654 ^ n2519 ;
  assign n2656 = n2655 ^ n2597 ;
  assign n2657 = n2656 ^ n2633 ;
  assign n35789 = n35773 ^ n2657 ;
  assign n35793 = n35792 ^ n35789 ;
  assign n35812 = n35811 ^ n35793 ;
  assign n35817 = n35816 ^ n35812 ;
  assign n35786 = n35775 ^ n35738 ;
  assign n35787 = ~n35743 & n35786 ;
  assign n35788 = n35787 ^ n35738 ;
  assign n35818 = n35817 ^ n35788 ;
  assign n35823 = n35822 ^ n35818 ;
  assign n35783 = n3242 ^ n1890 ;
  assign n35784 = n35783 ^ n29816 ;
  assign n35785 = n35784 ^ n3060 ;
  assign n35824 = n35823 ^ n35785 ;
  assign n35734 = n35733 ^ n32275 ;
  assign n35735 = n3230 & n35734 ;
  assign n35736 = n35735 ^ n3023 ;
  assign n35779 = n35778 ^ n35776 ;
  assign n35780 = n35779 ^ n35735 ;
  assign n35781 = n35736 & n35780 ;
  assign n35782 = n35781 ^ n3023 ;
  assign n35825 = n35824 ^ n35782 ;
  assign n36096 = n35688 ^ n35540 ;
  assign n35924 = n35103 ^ n35058 ;
  assign n36092 = n35924 ^ n34045 ;
  assign n36093 = n34045 ^ n33211 ;
  assign n36094 = n36092 & ~n36093 ;
  assign n36095 = n36094 ^ n33211 ;
  assign n36097 = n36096 ^ n36095 ;
  assign n35838 = n35685 ^ n35542 ;
  assign n35834 = n35192 ^ n34227 ;
  assign n35835 = n35807 ^ n35192 ;
  assign n35836 = n35834 & n35835 ;
  assign n35837 = n35836 ^ n34227 ;
  assign n35839 = n35838 ^ n35837 ;
  assign n36080 = n35681 ^ n35548 ;
  assign n35844 = n35678 ^ n35553 ;
  assign n35840 = n34719 ^ n34156 ;
  assign n35841 = n35717 ^ n34719 ;
  assign n35842 = n35840 & n35841 ;
  assign n35843 = n35842 ^ n34156 ;
  assign n35845 = n35844 ^ n35843 ;
  assign n35847 = n34864 ^ n34147 ;
  assign n35848 = n35458 ^ n34864 ;
  assign n35849 = ~n35847 & ~n35848 ;
  assign n35850 = n35849 ^ n34147 ;
  assign n35846 = n35676 ^ n1574 ;
  assign n35851 = n35850 ^ n35846 ;
  assign n35856 = n35672 ^ n35670 ;
  assign n35852 = n34727 ^ n34027 ;
  assign n35853 = n34727 ^ n34712 ;
  assign n35854 = n35852 & ~n35853 ;
  assign n35855 = n35854 ^ n34027 ;
  assign n35857 = n35856 ^ n35855 ;
  assign n36061 = n35667 ^ n35560 ;
  assign n36052 = n34761 ^ n34735 ;
  assign n36053 = n34761 ^ n33793 ;
  assign n36054 = n36052 & n36053 ;
  assign n36055 = n36054 ^ n33793 ;
  assign n36043 = n35660 ^ n35659 ;
  assign n35859 = n34913 ^ n34752 ;
  assign n35860 = n34913 ^ n33747 ;
  assign n35861 = ~n35859 & n35860 ;
  assign n35862 = n35861 ^ n33747 ;
  assign n35858 = n35653 ^ n35574 ;
  assign n35863 = n35862 ^ n35858 ;
  assign n35868 = n35649 ^ n35580 ;
  assign n35864 = n34784 ^ n34760 ;
  assign n35865 = n34760 ^ n33732 ;
  assign n35866 = n35864 & n35865 ;
  assign n35867 = n35866 ^ n34784 ;
  assign n35869 = n35868 ^ n35867 ;
  assign n35874 = n35647 ^ n35581 ;
  assign n35870 = n34882 ^ n34781 ;
  assign n35871 = n34882 ^ n33712 ;
  assign n35872 = ~n35870 & n35871 ;
  assign n35873 = n35872 ^ n33712 ;
  assign n35875 = n35874 ^ n35873 ;
  assign n35877 = n35276 ^ n34680 ;
  assign n35878 = n34680 ^ n33661 ;
  assign n35879 = ~n35877 & ~n35878 ;
  assign n35880 = n35879 ^ n33661 ;
  assign n35876 = n35643 ^ n35584 ;
  assign n35881 = n35880 ^ n35876 ;
  assign n35883 = n35641 ^ n35585 ;
  assign n36030 = n35883 ^ n35880 ;
  assign n35882 = n34789 ^ n34503 ;
  assign n35884 = n35883 ^ n33543 ;
  assign n35885 = n35884 ^ n34789 ;
  assign n35886 = n35885 ^ n35883 ;
  assign n35887 = n35882 & ~n35886 ;
  assign n35888 = n35887 ^ n35884 ;
  assign n35893 = n35637 ^ n35591 ;
  assign n35889 = n34489 ^ n33328 ;
  assign n35890 = n35269 ^ n34489 ;
  assign n35891 = ~n35889 & ~n35890 ;
  assign n35892 = n35891 ^ n33328 ;
  assign n35894 = n35893 ^ n35892 ;
  assign n35895 = n35259 ^ n34329 ;
  assign n35896 = n35635 ^ n35595 ;
  assign n35897 = n35896 ^ n33338 ;
  assign n35898 = n35897 ^ n35259 ;
  assign n35899 = n35898 ^ n35896 ;
  assign n35900 = ~n35895 & ~n35899 ;
  assign n35901 = n35900 ^ n35897 ;
  assign n35903 = n34064 ^ n33340 ;
  assign n35904 = n34802 ^ n34064 ;
  assign n35905 = ~n35903 & ~n35904 ;
  assign n35906 = n35905 ^ n33340 ;
  assign n35902 = n35631 ^ n35630 ;
  assign n35907 = n35906 ^ n35902 ;
  assign n35909 = n34808 ^ n34075 ;
  assign n35910 = n34075 ^ n33341 ;
  assign n35911 = ~n35909 & n35910 ;
  assign n35912 = n35911 ^ n33341 ;
  assign n36018 = n35912 ^ n35902 ;
  assign n35908 = n35625 ^ n35621 ;
  assign n35913 = n35912 ^ n35908 ;
  assign n36002 = n34811 ^ n34081 ;
  assign n36003 = n34081 ^ n33364 ;
  assign n36004 = n36002 & ~n36003 ;
  assign n36005 = n36004 ^ n33364 ;
  assign n36015 = n36005 ^ n35912 ;
  assign n35914 = n34833 ^ n34118 ;
  assign n35956 = n33445 ^ n3161 ;
  assign n35957 = n35956 ^ n2534 ;
  assign n35958 = n35957 ^ n3197 ;
  assign n35959 = n35958 ^ n35936 ;
  assign n35952 = n35106 ^ n35053 ;
  assign n35953 = n35952 ^ n32626 ;
  assign n35954 = n35953 ^ n35924 ;
  assign n35951 = n31824 ^ n31676 ;
  assign n35955 = n35954 ^ n35951 ;
  assign n35960 = n35959 ^ n35955 ;
  assign n35915 = n33424 ^ n31587 ;
  assign n35916 = n34248 ^ n31587 ;
  assign n35917 = ~n35915 & n35916 ;
  assign n35918 = n35917 ^ n33424 ;
  assign n35919 = n35918 ^ n35801 ;
  assign n35920 = n35919 ^ n35807 ;
  assign n35921 = n35920 ^ n35918 ;
  assign n35922 = ~n35806 & n35921 ;
  assign n35923 = n35922 ^ n35919 ;
  assign n35949 = n35924 ^ n35918 ;
  assign n35950 = n35923 & n35949 ;
  assign n35961 = n35960 ^ n35950 ;
  assign n35926 = n35808 ^ n35796 ;
  assign n35927 = n35808 ^ n31785 ;
  assign n35928 = n35926 & ~n35927 ;
  assign n35929 = n35928 ^ n31785 ;
  assign n35930 = n35929 ^ n31676 ;
  assign n35925 = n35924 ^ n35923 ;
  assign n35947 = n35929 ^ n35925 ;
  assign n35948 = ~n35930 & ~n35947 ;
  assign n35962 = n35961 ^ n35948 ;
  assign n35944 = n33418 ^ n32626 ;
  assign n35945 = n34242 ^ n33418 ;
  assign n35946 = ~n35944 & n35945 ;
  assign n35963 = n35962 ^ n35946 ;
  assign n35931 = n35930 ^ n35925 ;
  assign n35932 = n35809 & n35810 ;
  assign n35943 = n35931 & n35932 ;
  assign n35964 = n35963 ^ n35943 ;
  assign n35933 = n35932 ^ n35931 ;
  assign n35937 = n35936 ^ n35933 ;
  assign n35938 = n35811 ^ n2657 ;
  assign n35939 = n35793 & n35938 ;
  assign n35940 = n35939 ^ n2657 ;
  assign n35941 = n35940 ^ n35933 ;
  assign n35942 = n35937 & ~n35941 ;
  assign n35965 = n35964 ^ n35942 ;
  assign n35966 = n35965 ^ n33383 ;
  assign n35967 = n35966 ^ n34833 ;
  assign n35968 = n35967 ^ n35965 ;
  assign n35969 = n35914 & n35968 ;
  assign n35970 = n35969 ^ n35966 ;
  assign n35978 = n35218 ^ n34095 ;
  assign n35979 = n34095 ^ n33385 ;
  assign n35980 = n35978 & n35979 ;
  assign n35981 = n35980 ^ n33385 ;
  assign n35977 = n35940 ^ n35937 ;
  assign n35982 = n35981 ^ n35977 ;
  assign n35983 = n35812 ^ n35788 ;
  assign n35984 = n35817 & ~n35983 ;
  assign n35985 = n35984 ^ n35816 ;
  assign n35986 = n35985 ^ n35977 ;
  assign n35987 = n35982 & ~n35986 ;
  assign n35988 = n35987 ^ n35981 ;
  assign n35971 = n34827 ^ n34094 ;
  assign n35972 = n34094 ^ n33352 ;
  assign n35973 = ~n35971 & n35972 ;
  assign n35974 = n35973 ^ n33352 ;
  assign n35975 = n35974 ^ n35965 ;
  assign n35976 = n35975 ^ n35974 ;
  assign n35989 = n35988 ^ n35976 ;
  assign n35990 = ~n35970 & ~n35989 ;
  assign n35991 = n35990 ^ n35975 ;
  assign n35992 = n34088 ^ n33347 ;
  assign n35993 = n34821 ^ n34088 ;
  assign n35994 = n35992 & n35993 ;
  assign n35995 = n35994 ^ n33347 ;
  assign n35997 = n35995 ^ n35974 ;
  assign n35830 = n35605 ^ n35604 ;
  assign n35996 = n35995 ^ n35830 ;
  assign n35998 = n35997 ^ n35996 ;
  assign n35999 = n35991 & n35998 ;
  assign n36000 = n35999 ^ n35996 ;
  assign n36007 = n36005 ^ n35995 ;
  assign n36001 = n35607 ^ n35600 ;
  assign n36006 = n36005 ^ n36001 ;
  assign n36008 = n36007 ^ n36006 ;
  assign n36009 = ~n36000 & ~n36008 ;
  assign n36010 = n36009 ^ n36007 ;
  assign n36011 = n35612 ^ n35472 ;
  assign n36012 = n36011 ^ n35609 ;
  assign n36013 = n36012 ^ n36005 ;
  assign n36014 = ~n36010 & n36013 ;
  assign n36016 = n36015 ^ n36014 ;
  assign n36017 = n35913 & ~n36016 ;
  assign n36019 = n36018 ^ n36017 ;
  assign n36020 = ~n35907 & ~n36019 ;
  assign n36021 = n36020 ^ n35906 ;
  assign n36022 = n36021 ^ n35896 ;
  assign n36023 = n35901 & n36022 ;
  assign n36024 = n36023 ^ n35896 ;
  assign n36025 = n36024 ^ n35892 ;
  assign n36026 = n35894 & ~n36025 ;
  assign n36027 = n36026 ^ n35893 ;
  assign n36028 = n36027 ^ n35883 ;
  assign n36029 = n35888 & n36028 ;
  assign n36031 = n36030 ^ n36029 ;
  assign n36032 = n35881 & n36031 ;
  assign n36033 = n36032 ^ n35880 ;
  assign n36034 = n36033 ^ n35873 ;
  assign n36035 = ~n35875 & ~n36034 ;
  assign n36036 = n36035 ^ n35874 ;
  assign n36037 = n36036 ^ n35867 ;
  assign n36038 = n35869 & ~n36037 ;
  assign n36039 = n36038 ^ n35868 ;
  assign n36040 = n36039 ^ n35858 ;
  assign n36041 = ~n35863 & ~n36040 ;
  assign n36042 = n36041 ^ n35862 ;
  assign n36044 = n36043 ^ n36042 ;
  assign n36048 = n36043 ^ n33775 ;
  assign n36045 = n34777 ^ n33775 ;
  assign n36046 = n34777 ^ n34744 ;
  assign n36047 = n36045 & ~n36046 ;
  assign n36049 = n36048 ^ n36047 ;
  assign n36050 = n36044 & ~n36049 ;
  assign n36051 = n36050 ^ n36043 ;
  assign n36056 = n36055 ^ n36051 ;
  assign n36057 = n35665 ^ n35569 ;
  assign n36058 = n36057 ^ n36051 ;
  assign n36059 = ~n36056 & n36058 ;
  assign n36060 = n36059 ^ n36055 ;
  assign n36062 = n36061 ^ n36060 ;
  assign n36063 = n34750 ^ n33816 ;
  assign n36064 = n36061 ^ n35308 ;
  assign n36065 = n36064 ^ n36061 ;
  assign n36066 = n36065 ^ n34750 ;
  assign n36067 = n36063 & n36066 ;
  assign n36068 = n36067 ^ n36064 ;
  assign n36069 = ~n36062 & ~n36068 ;
  assign n36070 = n36069 ^ n36061 ;
  assign n36071 = n36070 ^ n35855 ;
  assign n36072 = ~n35857 & ~n36071 ;
  assign n36073 = n36072 ^ n35856 ;
  assign n36074 = n36073 ^ n35846 ;
  assign n36075 = ~n35851 & ~n36074 ;
  assign n36076 = n36075 ^ n35850 ;
  assign n36077 = n36076 ^ n35843 ;
  assign n36078 = ~n35845 & n36077 ;
  assign n36079 = n36078 ^ n35844 ;
  assign n36081 = n36080 ^ n36079 ;
  assign n36082 = n34174 ^ n34062 ;
  assign n36083 = n35757 ^ n34174 ;
  assign n36084 = ~n36082 & n36083 ;
  assign n36085 = n36084 ^ n34062 ;
  assign n36086 = n36085 ^ n36079 ;
  assign n36087 = ~n36081 & n36086 ;
  assign n36088 = n36087 ^ n36080 ;
  assign n36089 = n36088 ^ n35837 ;
  assign n36090 = ~n35839 & n36089 ;
  assign n36091 = n36090 ^ n35838 ;
  assign n36226 = n36095 ^ n36091 ;
  assign n36227 = ~n36097 & n36226 ;
  assign n36228 = n36227 ^ n36096 ;
  assign n36219 = n35952 ^ n34257 ;
  assign n36220 = n35690 ^ n35539 ;
  assign n36221 = n36220 ^ n33273 ;
  assign n36222 = n36221 ^ n35952 ;
  assign n36223 = n36222 ^ n36220 ;
  assign n36224 = n36219 & ~n36223 ;
  assign n36225 = n36224 ^ n36221 ;
  assign n36229 = n36228 ^ n36225 ;
  assign n36099 = n36088 ^ n35839 ;
  assign n36100 = n36099 ^ n33462 ;
  assign n36103 = n36073 ^ n35851 ;
  assign n36104 = n36103 ^ n33225 ;
  assign n36105 = n36068 ^ n36060 ;
  assign n36106 = n36105 ^ n32947 ;
  assign n36107 = n36057 ^ n36055 ;
  assign n36108 = n36107 ^ n36051 ;
  assign n36109 = n36108 ^ n32933 ;
  assign n36111 = n36039 ^ n35863 ;
  assign n36112 = n36111 ^ n32129 ;
  assign n36113 = n36036 ^ n35869 ;
  assign n36114 = n36113 ^ n32161 ;
  assign n36115 = n36033 ^ n35875 ;
  assign n36116 = n36115 ^ n32145 ;
  assign n36117 = n36031 ^ n35876 ;
  assign n36118 = n36117 ^ n32138 ;
  assign n36167 = n36027 ^ n35888 ;
  assign n36119 = n36024 ^ n35894 ;
  assign n36120 = n36119 ^ n32220 ;
  assign n36122 = n35991 ^ n35830 ;
  assign n36123 = n36122 ^ n32246 ;
  assign n36132 = n35988 ^ n35970 ;
  assign n36125 = n35821 ^ n35818 ;
  assign n36126 = n35822 & ~n36125 ;
  assign n36127 = n36126 ^ n32265 ;
  assign n36124 = n35985 ^ n35982 ;
  assign n36128 = n36127 ^ n36124 ;
  assign n36129 = n36127 ^ n32259 ;
  assign n36130 = ~n36128 & n36129 ;
  assign n36131 = n36130 ^ n32259 ;
  assign n36133 = n36132 ^ n36131 ;
  assign n36134 = n36132 ^ n32256 ;
  assign n36135 = n36133 & ~n36134 ;
  assign n36136 = n36135 ^ n32256 ;
  assign n36137 = n36136 ^ n36122 ;
  assign n36138 = n36123 & n36137 ;
  assign n36139 = n36138 ^ n32246 ;
  assign n36140 = n36139 ^ n32240 ;
  assign n36141 = n36001 ^ n36000 ;
  assign n36142 = n36141 ^ n36139 ;
  assign n36143 = ~n36140 & ~n36142 ;
  assign n36144 = n36143 ^ n32240 ;
  assign n36145 = n36144 ^ n32233 ;
  assign n36146 = n36012 ^ n36010 ;
  assign n36147 = n36146 ^ n36144 ;
  assign n36148 = n36145 & n36147 ;
  assign n36149 = n36148 ^ n32233 ;
  assign n36150 = n36149 ^ n32667 ;
  assign n36151 = n36016 ^ n35908 ;
  assign n36152 = n36151 ^ n36149 ;
  assign n36153 = ~n36150 & ~n36152 ;
  assign n36154 = n36153 ^ n32667 ;
  assign n36155 = n36154 ^ n32202 ;
  assign n36156 = n36019 ^ n35906 ;
  assign n36157 = n36156 ^ n36154 ;
  assign n36158 = ~n36155 & n36157 ;
  assign n36159 = n36158 ^ n32202 ;
  assign n36121 = n36021 ^ n35901 ;
  assign n36160 = n36159 ^ n36121 ;
  assign n36161 = n36159 ^ n32204 ;
  assign n36162 = ~n36160 & n36161 ;
  assign n36163 = n36162 ^ n32204 ;
  assign n36164 = n36163 ^ n36119 ;
  assign n36165 = ~n36120 & ~n36164 ;
  assign n36166 = n36165 ^ n32220 ;
  assign n36168 = n36167 ^ n36166 ;
  assign n36169 = n36167 ^ n32189 ;
  assign n36170 = n36168 & n36169 ;
  assign n36171 = n36170 ^ n32189 ;
  assign n36172 = n36171 ^ n36117 ;
  assign n36173 = ~n36118 & ~n36172 ;
  assign n36174 = n36173 ^ n32138 ;
  assign n36175 = n36174 ^ n36115 ;
  assign n36176 = n36116 & ~n36175 ;
  assign n36177 = n36176 ^ n32145 ;
  assign n36178 = n36177 ^ n36113 ;
  assign n36179 = ~n36114 & ~n36178 ;
  assign n36180 = n36179 ^ n32161 ;
  assign n36181 = n36180 ^ n36111 ;
  assign n36182 = ~n36112 & ~n36181 ;
  assign n36183 = n36182 ^ n32129 ;
  assign n36110 = n36049 ^ n36042 ;
  assign n36184 = n36183 ^ n36110 ;
  assign n36185 = n36183 ^ n32697 ;
  assign n36186 = ~n36184 & n36185 ;
  assign n36187 = n36186 ^ n32697 ;
  assign n36188 = n36187 ^ n36108 ;
  assign n36189 = n36109 & n36188 ;
  assign n36190 = n36189 ^ n32933 ;
  assign n36191 = n36190 ^ n36105 ;
  assign n36192 = ~n36106 & ~n36191 ;
  assign n36193 = n36192 ^ n32947 ;
  assign n36194 = n36193 ^ n32989 ;
  assign n36195 = n36070 ^ n35857 ;
  assign n36196 = n36195 ^ n36193 ;
  assign n36197 = ~n36194 & ~n36196 ;
  assign n36198 = n36197 ^ n32989 ;
  assign n36199 = n36198 ^ n36103 ;
  assign n36200 = ~n36104 & ~n36199 ;
  assign n36201 = n36200 ^ n33225 ;
  assign n36202 = n36201 ^ n33294 ;
  assign n36203 = n36076 ^ n35845 ;
  assign n36204 = n36203 ^ n36201 ;
  assign n36205 = ~n36202 & ~n36204 ;
  assign n36206 = n36205 ^ n33294 ;
  assign n36101 = n36085 ^ n36080 ;
  assign n36102 = n36101 ^ n36079 ;
  assign n36207 = n36206 ^ n36102 ;
  assign n36208 = n36206 ^ n33426 ;
  assign n36209 = ~n36207 & ~n36208 ;
  assign n36210 = n36209 ^ n33426 ;
  assign n36211 = n36210 ^ n36099 ;
  assign n36212 = n36100 & n36211 ;
  assign n36213 = n36212 ^ n33462 ;
  assign n36098 = n36097 ^ n36091 ;
  assign n36214 = n36213 ^ n36098 ;
  assign n36215 = n36213 ^ n32593 ;
  assign n36216 = ~n36214 & n36215 ;
  assign n36217 = n36216 ^ n32593 ;
  assign n36218 = n36217 ^ n32592 ;
  assign n36230 = n36229 ^ n36218 ;
  assign n36231 = n36198 ^ n36104 ;
  assign n36232 = n36195 ^ n36194 ;
  assign n36233 = n36187 ^ n32933 ;
  assign n36234 = n36233 ^ n36108 ;
  assign n36235 = n36110 ^ n32697 ;
  assign n36236 = n36235 ^ n36183 ;
  assign n36237 = n36163 ^ n36120 ;
  assign n36238 = n36161 ^ n36121 ;
  assign n36239 = n36124 ^ n32259 ;
  assign n36240 = n36239 ^ n36127 ;
  assign n36241 = ~n35823 & ~n36240 ;
  assign n36242 = n36131 ^ n32256 ;
  assign n36243 = n36242 ^ n36132 ;
  assign n36244 = n36241 & n36243 ;
  assign n36245 = n36136 ^ n36123 ;
  assign n36246 = ~n36244 & n36245 ;
  assign n36247 = n36141 ^ n36140 ;
  assign n36248 = ~n36246 & ~n36247 ;
  assign n36249 = n36146 ^ n36145 ;
  assign n36250 = n36248 & n36249 ;
  assign n36251 = n36151 ^ n36150 ;
  assign n36252 = ~n36250 & ~n36251 ;
  assign n36253 = n36156 ^ n36155 ;
  assign n36254 = n36252 & ~n36253 ;
  assign n36255 = ~n36238 & ~n36254 ;
  assign n36256 = n36237 & n36255 ;
  assign n36257 = n36166 ^ n32189 ;
  assign n36258 = n36257 ^ n36167 ;
  assign n36259 = n36256 & n36258 ;
  assign n36260 = n36171 ^ n36118 ;
  assign n36261 = n36259 & n36260 ;
  assign n36262 = n36174 ^ n32145 ;
  assign n36263 = n36262 ^ n36115 ;
  assign n36264 = ~n36261 & ~n36263 ;
  assign n36265 = n36177 ^ n36114 ;
  assign n36266 = ~n36264 & ~n36265 ;
  assign n36267 = n36180 ^ n36112 ;
  assign n36268 = n36266 & n36267 ;
  assign n36269 = n36236 & n36268 ;
  assign n36270 = ~n36234 & ~n36269 ;
  assign n36271 = n36190 ^ n36106 ;
  assign n36272 = ~n36270 & n36271 ;
  assign n36273 = ~n36232 & n36272 ;
  assign n36274 = ~n36231 & ~n36273 ;
  assign n36275 = n36203 ^ n36202 ;
  assign n36276 = n36274 & n36275 ;
  assign n36277 = n36102 ^ n33426 ;
  assign n36278 = n36277 ^ n36206 ;
  assign n36279 = n36276 & ~n36278 ;
  assign n36280 = n36210 ^ n36100 ;
  assign n36281 = ~n36279 & n36280 ;
  assign n36282 = n36098 ^ n32593 ;
  assign n36283 = n36282 ^ n36213 ;
  assign n36284 = n36281 & ~n36283 ;
  assign n36483 = n36230 & n36284 ;
  assign n36479 = n35694 ^ n35536 ;
  assign n36470 = n34255 ^ n33312 ;
  assign n36471 = n35149 ^ n34255 ;
  assign n36472 = n36470 & ~n36471 ;
  assign n36473 = n36472 ^ n33312 ;
  assign n36475 = n36473 ^ n36220 ;
  assign n36474 = n36473 ^ n36228 ;
  assign n36476 = n36475 ^ n36474 ;
  assign n36477 = ~n36225 & ~n36476 ;
  assign n36478 = n36477 ^ n36475 ;
  assign n36480 = n36479 ^ n36478 ;
  assign n36481 = n36480 ^ n32591 ;
  assign n36466 = n36229 ^ n36217 ;
  assign n36467 = n36229 ^ n32592 ;
  assign n36468 = ~n36466 & ~n36467 ;
  assign n36469 = n36468 ^ n32592 ;
  assign n36482 = n36481 ^ n36469 ;
  assign n36484 = n36483 ^ n36482 ;
  assign n36286 = n33833 ^ n2894 ;
  assign n36287 = n36286 ^ n30211 ;
  assign n36288 = n36287 ^ n24512 ;
  assign n36285 = n36284 ^ n36230 ;
  assign n36289 = n36288 ^ n36285 ;
  assign n36296 = n33838 ^ n2882 ;
  assign n36297 = n36296 ^ n30215 ;
  assign n36298 = n36297 ^ n2642 ;
  assign n36295 = n36283 ^ n36281 ;
  assign n36299 = n36298 ^ n36295 ;
  assign n36300 = n36280 ^ n36279 ;
  assign n1386 = n1385 ^ n1262 ;
  assign n1387 = n1386 ^ n1352 ;
  assign n1388 = n1387 ^ n1379 ;
  assign n36301 = n36300 ^ n1388 ;
  assign n36302 = n33845 ^ n1765 ;
  assign n36303 = n36302 ^ n1183 ;
  assign n36304 = n36303 ^ n1346 ;
  assign n36456 = n36304 ^ n1388 ;
  assign n36305 = n36278 ^ n36276 ;
  assign n36306 = n36305 ^ n36304 ;
  assign n36307 = n36275 ^ n36274 ;
  assign n36308 = n36307 ^ n1176 ;
  assign n36309 = n36273 ^ n36231 ;
  assign n1040 = n1003 ^ n964 ;
  assign n1041 = n1040 ^ n1037 ;
  assign n1048 = n1047 ^ n1041 ;
  assign n36310 = n36309 ^ n1048 ;
  assign n36311 = n36272 ^ n36232 ;
  assign n1007 = n991 ^ n949 ;
  assign n1023 = n1022 ^ n1007 ;
  assign n1030 = n1029 ^ n1023 ;
  assign n36312 = n36311 ^ n1030 ;
  assign n36444 = n36317 ^ n1030 ;
  assign n36313 = n36269 ^ n36234 ;
  assign n36314 = n36313 ^ n1632 ;
  assign n36323 = n36268 ^ n36236 ;
  assign n36324 = n36323 ^ n36322 ;
  assign n36328 = n36267 ^ n36266 ;
  assign n36329 = n36328 ^ n36327 ;
  assign n36330 = n36265 ^ n36264 ;
  assign n2961 = n2960 ^ n2957 ;
  assign n2962 = n2961 ^ n620 ;
  assign n2966 = n2965 ^ n2962 ;
  assign n36331 = n36330 ^ n2966 ;
  assign n36332 = n36263 ^ n36261 ;
  assign n36336 = n36335 ^ n36332 ;
  assign n36340 = n33922 ^ n599 ;
  assign n36341 = n36340 ^ n29775 ;
  assign n36342 = n36341 ^ n24537 ;
  assign n36339 = n36260 ^ n36259 ;
  assign n36343 = n36342 ^ n36339 ;
  assign n36345 = n33926 ^ n25823 ;
  assign n36346 = n36345 ^ n29780 ;
  assign n36347 = n36346 ^ n1487 ;
  assign n36423 = n36347 ^ n36342 ;
  assign n36344 = n36258 ^ n36256 ;
  assign n36348 = n36347 ^ n36344 ;
  assign n36352 = n36255 ^ n36237 ;
  assign n36349 = n33931 ^ n25827 ;
  assign n36350 = n36349 ^ n29786 ;
  assign n36351 = n36350 ^ n24544 ;
  assign n36353 = n36352 ^ n36351 ;
  assign n36355 = n25832 ^ n2429 ;
  assign n36356 = n36355 ^ n29850 ;
  assign n36357 = n36356 ^ n24589 ;
  assign n36417 = n36357 ^ n36351 ;
  assign n36354 = n36254 ^ n36238 ;
  assign n36358 = n36357 ^ n36354 ;
  assign n36360 = n2414 ^ n2356 ;
  assign n36361 = n36360 ^ n29791 ;
  assign n36362 = n36361 ^ n24549 ;
  assign n36359 = n36253 ^ n36252 ;
  assign n36363 = n36362 ^ n36359 ;
  assign n36365 = n33941 ^ n2340 ;
  assign n36366 = n36365 ^ n29795 ;
  assign n36367 = n36366 ^ n24557 ;
  assign n36411 = n36367 ^ n36362 ;
  assign n36364 = n36251 ^ n36250 ;
  assign n36368 = n36367 ^ n36364 ;
  assign n36370 = n33946 ^ n2330 ;
  assign n36371 = n36370 ^ n29800 ;
  assign n36372 = n36371 ^ n2147 ;
  assign n36369 = n36249 ^ n36248 ;
  assign n36373 = n36372 ^ n36369 ;
  assign n36378 = n36245 ^ n36244 ;
  assign n36375 = n33955 ^ n25868 ;
  assign n36376 = n36375 ^ n29807 ;
  assign n36377 = n36376 ^ n2031 ;
  assign n36379 = n36378 ^ n36377 ;
  assign n36380 = n36243 ^ n36241 ;
  assign n1944 = n1943 ^ n1928 ;
  assign n1963 = n1962 ^ n1944 ;
  assign n1970 = n1969 ^ n1963 ;
  assign n36381 = n36380 ^ n1970 ;
  assign n36386 = n36240 ^ n35823 ;
  assign n36382 = n33281 ^ n25850 ;
  assign n36383 = n36382 ^ n3062 ;
  assign n36384 = n36383 ^ n1957 ;
  assign n36387 = n36386 ^ n36384 ;
  assign n36388 = n35785 ^ n35782 ;
  assign n36389 = ~n35824 & ~n36388 ;
  assign n36390 = n36389 ^ n35823 ;
  assign n36391 = n36390 ^ n36384 ;
  assign n36392 = ~n36387 & ~n36391 ;
  assign n36385 = n36384 ^ n1970 ;
  assign n36393 = n36392 ^ n36385 ;
  assign n36394 = ~n36381 & ~n36393 ;
  assign n36395 = n36394 ^ n36380 ;
  assign n36396 = n36395 ^ n36377 ;
  assign n36397 = ~n36379 & ~n36396 ;
  assign n36398 = n36397 ^ n36377 ;
  assign n36405 = n36398 ^ n36372 ;
  assign n36374 = n36247 ^ n36246 ;
  assign n36399 = n36398 ^ n36374 ;
  assign n36400 = n33951 ^ n25842 ;
  assign n36401 = n36400 ^ n2036 ;
  assign n36402 = n36401 ^ n24562 ;
  assign n36403 = n36402 ^ n36374 ;
  assign n36404 = ~n36399 & n36403 ;
  assign n36406 = n36405 ^ n36404 ;
  assign n36407 = ~n36373 & n36406 ;
  assign n36408 = n36407 ^ n36372 ;
  assign n36409 = n36408 ^ n36367 ;
  assign n36410 = n36368 & n36409 ;
  assign n36412 = n36411 ^ n36410 ;
  assign n36413 = ~n36363 & n36412 ;
  assign n36414 = n36413 ^ n36362 ;
  assign n36415 = n36414 ^ n36354 ;
  assign n36416 = ~n36358 & n36415 ;
  assign n36418 = n36417 ^ n36416 ;
  assign n36419 = ~n36353 & ~n36418 ;
  assign n36420 = n36419 ^ n36352 ;
  assign n36421 = n36420 ^ n36347 ;
  assign n36422 = ~n36348 & ~n36421 ;
  assign n36424 = n36423 ^ n36422 ;
  assign n36425 = ~n36343 & n36424 ;
  assign n36426 = n36425 ^ n36342 ;
  assign n36427 = n36426 ^ n36335 ;
  assign n36428 = n36336 & n36427 ;
  assign n36337 = n36335 ^ n2966 ;
  assign n36429 = n36428 ^ n36337 ;
  assign n36430 = ~n36331 & ~n36429 ;
  assign n36431 = n36430 ^ n36330 ;
  assign n36432 = n36431 ^ n36327 ;
  assign n36433 = ~n36329 & n36432 ;
  assign n36434 = n36433 ^ n36328 ;
  assign n36435 = n36434 ^ n36322 ;
  assign n36436 = ~n36324 & n36435 ;
  assign n36437 = n36436 ^ n36323 ;
  assign n36438 = n36437 ^ n1632 ;
  assign n36439 = n36314 & ~n36438 ;
  assign n36318 = n36317 ^ n1632 ;
  assign n36440 = n36439 ^ n36318 ;
  assign n36441 = n36271 ^ n36270 ;
  assign n36442 = n36441 ^ n36317 ;
  assign n36443 = n36440 & n36442 ;
  assign n36445 = n36444 ^ n36443 ;
  assign n36446 = n36312 & ~n36445 ;
  assign n36447 = n36446 ^ n36311 ;
  assign n36448 = n36447 ^ n1048 ;
  assign n36449 = n36310 & ~n36448 ;
  assign n36450 = n36449 ^ n36309 ;
  assign n36451 = n36450 ^ n1176 ;
  assign n36452 = n36308 & ~n36451 ;
  assign n36453 = n36452 ^ n36307 ;
  assign n36454 = n36453 ^ n36304 ;
  assign n36455 = ~n36306 & n36454 ;
  assign n36457 = n36456 ^ n36455 ;
  assign n36458 = n36301 & n36457 ;
  assign n36459 = n36458 ^ n1388 ;
  assign n36460 = n36459 ^ n36295 ;
  assign n36461 = n36299 & ~n36460 ;
  assign n36462 = n36461 ^ n36298 ;
  assign n36463 = n36462 ^ n36288 ;
  assign n36464 = ~n36289 & n36463 ;
  assign n36290 = n33828 ^ n3116 ;
  assign n36291 = n36290 ^ n30206 ;
  assign n36292 = n36291 ^ n24649 ;
  assign n36293 = n36292 ^ n36288 ;
  assign n36465 = n36464 ^ n36293 ;
  assign n36485 = n36484 ^ n36465 ;
  assign n35829 = n34839 ^ n33325 ;
  assign n35831 = n35830 ^ n33325 ;
  assign n35832 = n35829 & n35831 ;
  assign n35833 = n35832 ^ n34839 ;
  assign n36486 = n36485 ^ n35833 ;
  assign n36487 = n36486 ^ n33326 ;
  assign n35826 = n35198 ^ n2767 ;
  assign n35827 = n35826 ^ n31059 ;
  assign n35828 = n35827 ^ n1847 ;
  assign n37309 = n36487 ^ n35828 ;
  assign n38168 = n37309 ^ n36012 ;
  assign n38169 = n37309 ^ n35825 ;
  assign n38170 = n38168 & n38169 ;
  assign n38171 = n38170 ^ n36012 ;
  assign n37255 = n36459 ^ n36299 ;
  assign n37948 = n37255 ^ n35732 ;
  assign n36592 = n35844 ^ n34777 ;
  assign n36597 = n36418 ^ n36352 ;
  assign n36593 = n34913 ^ n34735 ;
  assign n36594 = n35846 ^ n34735 ;
  assign n36595 = n36593 & n36594 ;
  assign n36596 = n36595 ^ n34913 ;
  assign n36598 = n36597 ^ n36596 ;
  assign n36599 = n36061 ^ n34752 ;
  assign n36600 = n36412 ^ n36359 ;
  assign n36601 = n36600 ^ n34882 ;
  assign n36602 = n36601 ^ n36061 ;
  assign n36603 = n36602 ^ n36600 ;
  assign n36604 = ~n36599 & n36603 ;
  assign n36605 = n36604 ^ n36601 ;
  assign n36606 = n36414 ^ n36358 ;
  assign n36761 = n36606 ^ n36600 ;
  assign n36611 = n36408 ^ n36368 ;
  assign n36607 = n34760 ^ n34680 ;
  assign n36608 = n36057 ^ n34760 ;
  assign n36609 = n36607 & ~n36608 ;
  assign n36610 = n36609 ^ n34680 ;
  assign n36612 = n36611 ^ n36610 ;
  assign n36614 = n36406 ^ n36369 ;
  assign n36756 = n36614 ^ n36610 ;
  assign n36613 = n36043 ^ n34781 ;
  assign n36615 = n36614 ^ n34503 ;
  assign n36616 = n36615 ^ n34781 ;
  assign n36617 = n36616 ^ n36614 ;
  assign n36618 = ~n36613 & n36617 ;
  assign n36619 = n36618 ^ n36615 ;
  assign n36624 = n36403 ^ n36398 ;
  assign n36620 = n35858 ^ n35276 ;
  assign n36621 = n35858 ^ n34489 ;
  assign n36622 = ~n36620 & n36621 ;
  assign n36623 = n36622 ^ n34489 ;
  assign n36625 = n36624 ^ n36623 ;
  assign n36741 = n36395 ^ n36379 ;
  assign n36627 = n35874 ^ n34064 ;
  assign n36628 = n35874 ^ n35269 ;
  assign n36629 = n36627 & ~n36628 ;
  assign n36630 = n36629 ^ n34064 ;
  assign n36626 = n36393 ^ n36380 ;
  assign n36631 = n36630 ^ n36626 ;
  assign n36632 = n35876 ^ n35259 ;
  assign n36633 = n36390 ^ n36387 ;
  assign n36634 = n36633 ^ n34075 ;
  assign n36635 = n36634 ^ n35876 ;
  assign n36636 = n36635 ^ n36633 ;
  assign n36637 = n36632 & ~n36636 ;
  assign n36638 = n36637 ^ n36634 ;
  assign n36641 = n35883 ^ n34802 ;
  assign n36642 = n35883 ^ n34081 ;
  assign n36643 = n36641 & ~n36642 ;
  assign n36644 = n36643 ^ n34081 ;
  assign n36645 = n36644 ^ n35825 ;
  assign n36723 = n35779 ^ n35736 ;
  assign n36580 = n35734 ^ n3230 ;
  assign n36724 = n36723 ^ n36580 ;
  assign n36561 = n35700 ^ n35526 ;
  assign n36504 = n34248 ^ n33478 ;
  assign n36505 = n35155 ^ n34248 ;
  assign n36506 = ~n36504 & ~n36505 ;
  assign n36507 = n36506 ^ n33478 ;
  assign n36509 = n36507 ^ n36473 ;
  assign n36508 = n36507 ^ n36479 ;
  assign n36510 = n36509 ^ n36508 ;
  assign n36511 = ~n36478 & ~n36510 ;
  assign n36512 = n36511 ^ n36509 ;
  assign n36552 = n35143 ^ n34242 ;
  assign n36553 = n34242 ^ n33472 ;
  assign n36554 = ~n36552 & n36553 ;
  assign n36555 = n36554 ^ n33472 ;
  assign n36557 = n36555 ^ n36507 ;
  assign n36513 = n35696 ^ n35535 ;
  assign n36556 = n36555 ^ n36513 ;
  assign n36558 = n36557 ^ n36556 ;
  assign n36559 = n36512 & n36558 ;
  assign n36560 = n36559 ^ n36557 ;
  assign n36562 = n36561 ^ n36560 ;
  assign n36515 = n36480 ^ n36469 ;
  assign n36516 = ~n36481 & ~n36515 ;
  assign n36517 = n36516 ^ n32591 ;
  assign n36518 = n36517 ^ n32589 ;
  assign n36514 = n36513 ^ n36512 ;
  assign n36548 = n36517 ^ n36514 ;
  assign n36549 = ~n36518 & n36548 ;
  assign n36550 = n36549 ^ n32589 ;
  assign n36551 = n36550 ^ n32583 ;
  assign n36563 = n36562 ^ n36551 ;
  assign n36503 = ~n36482 & n36483 ;
  assign n36519 = n36518 ^ n36514 ;
  assign n36564 = ~n36503 & n36519 ;
  assign n36667 = ~n36563 & n36564 ;
  assign n36661 = n36562 ^ n36550 ;
  assign n36662 = n36562 ^ n32583 ;
  assign n36663 = n36661 & n36662 ;
  assign n36664 = n36663 ^ n32583 ;
  assign n36665 = n36664 ^ n31587 ;
  assign n36656 = n34130 ^ n33424 ;
  assign n36657 = n35141 ^ n34130 ;
  assign n36658 = ~n36656 & n36657 ;
  assign n36659 = n36658 ^ n33424 ;
  assign n36650 = n35702 ^ n35525 ;
  assign n36652 = n36650 ^ n36555 ;
  assign n36651 = n36650 ^ n36561 ;
  assign n36653 = n36652 ^ n36651 ;
  assign n36654 = ~n36560 & ~n36653 ;
  assign n36655 = n36654 ^ n36652 ;
  assign n36660 = n36659 ^ n36655 ;
  assign n36666 = n36665 ^ n36660 ;
  assign n36690 = n36667 ^ n36666 ;
  assign n36681 = n34215 ^ n2636 ;
  assign n36682 = n36681 ^ n30193 ;
  assign n36683 = n36682 ^ n2717 ;
  assign n36691 = n36690 ^ n36683 ;
  assign n36543 = n34204 ^ n2607 ;
  assign n36544 = n36543 ^ n3128 ;
  assign n36545 = n36544 ^ n24677 ;
  assign n36522 = n36484 ^ n36292 ;
  assign n36523 = n36465 & n36522 ;
  assign n36524 = n36523 ^ n36292 ;
  assign n36546 = n36545 ^ n36524 ;
  assign n36520 = n36519 ^ n36503 ;
  assign n36500 = n34021 ^ n25949 ;
  assign n36501 = n36500 ^ n30200 ;
  assign n36502 = n36501 ^ n3104 ;
  assign n36521 = n36520 ^ n36502 ;
  assign n36541 = n36524 ^ n36502 ;
  assign n36542 = n36521 & n36541 ;
  assign n36547 = n36546 ^ n36542 ;
  assign n36565 = n36564 ^ n36563 ;
  assign n36692 = n36565 ^ n36545 ;
  assign n36693 = n36547 & ~n36692 ;
  assign n36694 = n36693 ^ n36545 ;
  assign n36695 = n36694 ^ n36683 ;
  assign n36696 = ~n36691 & n36695 ;
  assign n2707 = n2703 ^ n2676 ;
  assign n2720 = n2719 ^ n2707 ;
  assign n2724 = n2723 ^ n2720 ;
  assign n36684 = n36683 ^ n2724 ;
  assign n36679 = n32626 ^ n31587 ;
  assign n36677 = n36650 ^ n33418 ;
  assign n36676 = n35705 ^ n35523 ;
  assign n36678 = n36677 ^ n36676 ;
  assign n36680 = n36679 ^ n36678 ;
  assign n36685 = n36684 ^ n36680 ;
  assign n36674 = n36659 ^ n36650 ;
  assign n36675 = n36655 & n36674 ;
  assign n36686 = n36685 ^ n36675 ;
  assign n36672 = n36664 ^ n36660 ;
  assign n36673 = ~n36665 & ~n36672 ;
  assign n36687 = n36686 ^ n36673 ;
  assign n36669 = n34280 ^ n33418 ;
  assign n36670 = n35204 ^ n34280 ;
  assign n36671 = ~n36669 & n36670 ;
  assign n36688 = n36687 ^ n36671 ;
  assign n36668 = ~n36666 & n36667 ;
  assign n36689 = n36688 ^ n36668 ;
  assign n36697 = n36696 ^ n36689 ;
  assign n36646 = n35902 ^ n34821 ;
  assign n36647 = n34821 ^ n34118 ;
  assign n36648 = n36646 & ~n36647 ;
  assign n36649 = n36648 ^ n34118 ;
  assign n36698 = n36697 ^ n36649 ;
  assign n36540 = n36012 ^ n34833 ;
  assign n36566 = n36565 ^ n36547 ;
  assign n36567 = n36566 ^ n34113 ;
  assign n36568 = n36567 ^ n36012 ;
  assign n36569 = n36568 ^ n36566 ;
  assign n36570 = ~n36540 & ~n36569 ;
  assign n36571 = n36570 ^ n36567 ;
  assign n36493 = n36001 ^ n35218 ;
  assign n36494 = ~n35833 & n36485 ;
  assign n36495 = n36494 ^ n34109 ;
  assign n36496 = n36495 ^ n36001 ;
  assign n36497 = n36496 ^ n36494 ;
  assign n36498 = n36493 & ~n36497 ;
  assign n36499 = n36498 ^ n36495 ;
  assign n36525 = n36524 ^ n36521 ;
  assign n36572 = n36525 ^ n36494 ;
  assign n36573 = ~n36499 & ~n36572 ;
  assign n36574 = n36573 ^ n36494 ;
  assign n36700 = n36574 ^ n36566 ;
  assign n36701 = n36571 & ~n36700 ;
  assign n36702 = n36701 ^ n36566 ;
  assign n36699 = n36694 ^ n36691 ;
  assign n36703 = n36702 ^ n36699 ;
  assign n36704 = n35908 ^ n34827 ;
  assign n36705 = n36699 ^ n34095 ;
  assign n36706 = n36705 ^ n35908 ;
  assign n36707 = n36706 ^ n36699 ;
  assign n36708 = n36704 & ~n36707 ;
  assign n36709 = n36708 ^ n36705 ;
  assign n36710 = n36703 & n36709 ;
  assign n36711 = n36710 ^ n36702 ;
  assign n36712 = n36711 ^ n36649 ;
  assign n36713 = n36698 & ~n36712 ;
  assign n36714 = n36713 ^ n36697 ;
  assign n36715 = n36714 ^ n36580 ;
  assign n36716 = n35896 ^ n34811 ;
  assign n36717 = n36580 ^ n34094 ;
  assign n36718 = n36717 ^ n35896 ;
  assign n36719 = n36718 ^ n36580 ;
  assign n36720 = ~n36716 & n36719 ;
  assign n36721 = n36720 ^ n36717 ;
  assign n36722 = ~n36715 & n36721 ;
  assign n36725 = n36724 ^ n36722 ;
  assign n36726 = n34808 ^ n34088 ;
  assign n36727 = n35893 ^ n34808 ;
  assign n36728 = n36726 & n36727 ;
  assign n36729 = n36728 ^ n34088 ;
  assign n36730 = n36729 ^ n36723 ;
  assign n36731 = n36725 & n36730 ;
  assign n36732 = n36731 ^ n36729 ;
  assign n36733 = n36732 ^ n35825 ;
  assign n36734 = n36645 & ~n36733 ;
  assign n36735 = n36734 ^ n36644 ;
  assign n36736 = n36735 ^ n36633 ;
  assign n36737 = ~n36638 & ~n36736 ;
  assign n36639 = n36633 ^ n36630 ;
  assign n36738 = n36737 ^ n36639 ;
  assign n36739 = n36631 & ~n36738 ;
  assign n36740 = n36739 ^ n36630 ;
  assign n36742 = n36741 ^ n36740 ;
  assign n36743 = n35868 ^ n34789 ;
  assign n36744 = n36741 ^ n34329 ;
  assign n36745 = n36744 ^ n35868 ;
  assign n36746 = n36745 ^ n36741 ;
  assign n36747 = ~n36743 & n36746 ;
  assign n36748 = n36747 ^ n36744 ;
  assign n36749 = ~n36742 & ~n36748 ;
  assign n36750 = n36749 ^ n36741 ;
  assign n36751 = n36750 ^ n36623 ;
  assign n36752 = n36625 & n36751 ;
  assign n36753 = n36752 ^ n36624 ;
  assign n36754 = n36753 ^ n36614 ;
  assign n36755 = ~n36619 & n36754 ;
  assign n36757 = n36756 ^ n36755 ;
  assign n36758 = ~n36612 & ~n36757 ;
  assign n36759 = n36758 ^ n36611 ;
  assign n36760 = n36759 ^ n36606 ;
  assign n36762 = n36761 ^ n36760 ;
  assign n36763 = ~n36605 & ~n36762 ;
  assign n36764 = n36763 ^ n36761 ;
  assign n36770 = n36606 ^ n36596 ;
  assign n36765 = n35856 ^ n34744 ;
  assign n36766 = n35856 ^ n34784 ;
  assign n36767 = ~n36765 & n36766 ;
  assign n36768 = n36767 ^ n34784 ;
  assign n36769 = n36768 ^ n36596 ;
  assign n36771 = n36770 ^ n36769 ;
  assign n36772 = n36764 & n36771 ;
  assign n36773 = n36772 ^ n36770 ;
  assign n36774 = ~n36598 & n36773 ;
  assign n36775 = n36774 ^ n36597 ;
  assign n36776 = n36775 ^ n35308 ;
  assign n36777 = n36776 ^ n36775 ;
  assign n36778 = n36777 ^ n34777 ;
  assign n36779 = n36592 & n36778 ;
  assign n36780 = n36779 ^ n36776 ;
  assign n36782 = n36420 ^ n36348 ;
  assign n36586 = n36080 ^ n34712 ;
  assign n36587 = n34761 ^ n34712 ;
  assign n36588 = n36586 & ~n36587 ;
  assign n36589 = n36588 ^ n34761 ;
  assign n36783 = n36782 ^ n36589 ;
  assign n36781 = n36775 ^ n36589 ;
  assign n36784 = n36783 ^ n36781 ;
  assign n36785 = ~n36780 & ~n36784 ;
  assign n36786 = n36785 ^ n36783 ;
  assign n36590 = n36424 ^ n36339 ;
  assign n36875 = n36786 ^ n36590 ;
  assign n36798 = n36773 ^ n36597 ;
  assign n36799 = n36798 ^ n33747 ;
  assign n36801 = n36759 ^ n36605 ;
  assign n36802 = n36801 ^ n33712 ;
  assign n36803 = n36757 ^ n36611 ;
  assign n36804 = n36803 ^ n33661 ;
  assign n36805 = n36753 ^ n36619 ;
  assign n36806 = n36805 ^ n33543 ;
  assign n36808 = n36738 ^ n36626 ;
  assign n36809 = n36808 ^ n33340 ;
  assign n36810 = n36735 ^ n36638 ;
  assign n36811 = n36810 ^ n33341 ;
  assign n36831 = n36729 ^ n36725 ;
  assign n36814 = n36711 ^ n36698 ;
  assign n36815 = n36814 ^ n33383 ;
  assign n36816 = n36709 ^ n36702 ;
  assign n36817 = n36816 ^ n33385 ;
  assign n36527 = ~n33326 & ~n36486 ;
  assign n36528 = n36527 ^ n33401 ;
  assign n36526 = n36525 ^ n36499 ;
  assign n36536 = n36527 ^ n36526 ;
  assign n36537 = ~n36528 & ~n36536 ;
  assign n36538 = n36537 ^ n33401 ;
  assign n36539 = n36538 ^ n33391 ;
  assign n36575 = n36574 ^ n36571 ;
  assign n36818 = n36575 ^ n36538 ;
  assign n36819 = ~n36539 & n36818 ;
  assign n36820 = n36819 ^ n33391 ;
  assign n36821 = n36820 ^ n36816 ;
  assign n36822 = n36817 & ~n36821 ;
  assign n36823 = n36822 ^ n33385 ;
  assign n36824 = n36823 ^ n36814 ;
  assign n36825 = ~n36815 & n36824 ;
  assign n36826 = n36825 ^ n33383 ;
  assign n36813 = n36721 ^ n36714 ;
  assign n36827 = n36826 ^ n36813 ;
  assign n36828 = n36826 ^ n33352 ;
  assign n36829 = n36827 & n36828 ;
  assign n36830 = n36829 ^ n33352 ;
  assign n36832 = n36831 ^ n36830 ;
  assign n36833 = n36831 ^ n33347 ;
  assign n36834 = ~n36832 & ~n36833 ;
  assign n36835 = n36834 ^ n33347 ;
  assign n36812 = n36732 ^ n36645 ;
  assign n36836 = n36835 ^ n36812 ;
  assign n36837 = n36835 ^ n33364 ;
  assign n36838 = ~n36836 & ~n36837 ;
  assign n36839 = n36838 ^ n33364 ;
  assign n36840 = n36839 ^ n36810 ;
  assign n36841 = ~n36811 & ~n36840 ;
  assign n36842 = n36841 ^ n33341 ;
  assign n36843 = n36842 ^ n36808 ;
  assign n36844 = n36809 & n36843 ;
  assign n36845 = n36844 ^ n33340 ;
  assign n36846 = n36845 ^ n33338 ;
  assign n36847 = n36748 ^ n36740 ;
  assign n36848 = n36847 ^ n36845 ;
  assign n36849 = n36846 & ~n36848 ;
  assign n36850 = n36849 ^ n33338 ;
  assign n36807 = n36750 ^ n36625 ;
  assign n36851 = n36850 ^ n36807 ;
  assign n36852 = n36850 ^ n33328 ;
  assign n36853 = ~n36851 & n36852 ;
  assign n36854 = n36853 ^ n33328 ;
  assign n36855 = n36854 ^ n36805 ;
  assign n36856 = n36806 & ~n36855 ;
  assign n36857 = n36856 ^ n33543 ;
  assign n36858 = n36857 ^ n36803 ;
  assign n36859 = n36804 & ~n36858 ;
  assign n36860 = n36859 ^ n33661 ;
  assign n36861 = n36860 ^ n36801 ;
  assign n36862 = ~n36802 & n36861 ;
  assign n36863 = n36862 ^ n33712 ;
  assign n36800 = n36768 ^ n36764 ;
  assign n36864 = n36863 ^ n36800 ;
  assign n36865 = n36800 ^ n33732 ;
  assign n36866 = ~n36864 & n36865 ;
  assign n36867 = n36866 ^ n36863 ;
  assign n36868 = n36867 ^ n36798 ;
  assign n36869 = n36799 & ~n36868 ;
  assign n36870 = n36869 ^ n33747 ;
  assign n36797 = n36782 ^ n36780 ;
  assign n36871 = n36870 ^ n36797 ;
  assign n36872 = n36797 ^ n33775 ;
  assign n36873 = n36871 & n36872 ;
  assign n36874 = n36873 ^ n36870 ;
  assign n36876 = n36875 ^ n36874 ;
  assign n36794 = n36426 ^ n36336 ;
  assign n36585 = n35838 ^ n34750 ;
  assign n36591 = n36590 ^ n36589 ;
  assign n36787 = n36591 & n36786 ;
  assign n36788 = n36787 ^ n36590 ;
  assign n36789 = n36788 ^ n35458 ;
  assign n36790 = n36789 ^ n34750 ;
  assign n36791 = n36790 ^ n36788 ;
  assign n36792 = ~n36585 & n36791 ;
  assign n36793 = n36792 ^ n36789 ;
  assign n36795 = n36794 ^ n36793 ;
  assign n36877 = n36795 ^ n33793 ;
  assign n36878 = n36877 ^ n36795 ;
  assign n36879 = n36878 ^ n36874 ;
  assign n36880 = ~n36876 & ~n36879 ;
  assign n36881 = n36880 ^ n36877 ;
  assign n36897 = n36881 ^ n33816 ;
  assign n36898 = n36807 ^ n33328 ;
  assign n36899 = n36898 ^ n36850 ;
  assign n36900 = n36847 ^ n36846 ;
  assign n36901 = n36839 ^ n33341 ;
  assign n36902 = n36901 ^ n36810 ;
  assign n36903 = n36812 ^ n33364 ;
  assign n36904 = n36903 ^ n36835 ;
  assign n36905 = n36813 ^ n33352 ;
  assign n36906 = n36905 ^ n36826 ;
  assign n36576 = n36575 ^ n36539 ;
  assign n36907 = n36820 ^ n36817 ;
  assign n36908 = n36576 & ~n36907 ;
  assign n36909 = n36823 ^ n33383 ;
  assign n36910 = n36909 ^ n36814 ;
  assign n36911 = n36908 & n36910 ;
  assign n36912 = ~n36906 & ~n36911 ;
  assign n36913 = n36830 ^ n33347 ;
  assign n36914 = n36913 ^ n36831 ;
  assign n36915 = ~n36912 & n36914 ;
  assign n36916 = ~n36904 & n36915 ;
  assign n36917 = ~n36902 & ~n36916 ;
  assign n36918 = n36842 ^ n36809 ;
  assign n36919 = n36917 & ~n36918 ;
  assign n36920 = ~n36900 & ~n36919 ;
  assign n36921 = ~n36899 & n36920 ;
  assign n36922 = n36854 ^ n33543 ;
  assign n36923 = n36922 ^ n36805 ;
  assign n36924 = n36921 & ~n36923 ;
  assign n36925 = n36857 ^ n36804 ;
  assign n36926 = n36924 & ~n36925 ;
  assign n36927 = n36860 ^ n33712 ;
  assign n36928 = n36927 ^ n36801 ;
  assign n36929 = ~n36926 & ~n36928 ;
  assign n36930 = n36865 ^ n36863 ;
  assign n36931 = ~n36929 & n36930 ;
  assign n36932 = n36867 ^ n36799 ;
  assign n36933 = n36931 & ~n36932 ;
  assign n36934 = n36870 ^ n33775 ;
  assign n36935 = n36934 ^ n36797 ;
  assign n36936 = n36933 & n36935 ;
  assign n36937 = n36874 ^ n33793 ;
  assign n36938 = n36937 ^ n36875 ;
  assign n36939 = ~n36936 & ~n36938 ;
  assign n36940 = n36897 & ~n36939 ;
  assign n36894 = n36429 ^ n36330 ;
  assign n36885 = n35717 ^ n34727 ;
  assign n36886 = n36096 ^ n35717 ;
  assign n36887 = n36885 & n36886 ;
  assign n36888 = n36887 ^ n34727 ;
  assign n36890 = n36888 ^ n36794 ;
  assign n36889 = n36888 ^ n36788 ;
  assign n36891 = n36890 ^ n36889 ;
  assign n36892 = ~n36793 & ~n36891 ;
  assign n36893 = n36892 ^ n36890 ;
  assign n36895 = n36894 ^ n36893 ;
  assign n36796 = n36795 ^ n33816 ;
  assign n36882 = n36796 & ~n36881 ;
  assign n36883 = n36882 ^ n36795 ;
  assign n36884 = n36883 ^ n34027 ;
  assign n36896 = n36895 ^ n36884 ;
  assign n37199 = n36940 ^ n36896 ;
  assign n37069 = n34517 ^ n1652 ;
  assign n37070 = n37069 ^ n791 ;
  assign n37071 = n37070 ^ n1686 ;
  assign n1682 = n1669 ^ n1114 ;
  assign n1689 = n1688 ^ n1682 ;
  assign n1690 = n1689 ^ n928 ;
  assign n37197 = n37071 ^ n1690 ;
  assign n37065 = n34522 ^ n1646 ;
  assign n37066 = n37065 ^ n2992 ;
  assign n37067 = n37066 ^ n786 ;
  assign n37064 = n36938 ^ n36936 ;
  assign n37068 = n37067 ^ n37064 ;
  assign n37074 = n36935 ^ n36933 ;
  assign n37075 = n37074 ^ n722 ;
  assign n37079 = n36932 ^ n36931 ;
  assign n37080 = n37079 ^ n37078 ;
  assign n37084 = n36930 ^ n36929 ;
  assign n37184 = n37084 ^ n37079 ;
  assign n37085 = n37084 ^ n37083 ;
  assign n37181 = n37089 ^ n37083 ;
  assign n37086 = n36928 ^ n36926 ;
  assign n37090 = n37089 ^ n37086 ;
  assign n37092 = n34569 ^ n1499 ;
  assign n37093 = n37092 ^ n30674 ;
  assign n37094 = n37093 ^ n25051 ;
  assign n37091 = n36925 ^ n36924 ;
  assign n37095 = n37094 ^ n37091 ;
  assign n37100 = n36923 ^ n36921 ;
  assign n37096 = n34574 ^ n26517 ;
  assign n37097 = n37096 ^ n30679 ;
  assign n37098 = n37097 ^ n24981 ;
  assign n37101 = n37100 ^ n37098 ;
  assign n37103 = n34580 ^ n26472 ;
  assign n37104 = n37103 ^ n30685 ;
  assign n37105 = n37104 ^ n2921 ;
  assign n37102 = n36920 ^ n36899 ;
  assign n37106 = n37105 ^ n37102 ;
  assign n37111 = n36919 ^ n36900 ;
  assign n37107 = n34591 ^ n26481 ;
  assign n37108 = n37107 ^ n2378 ;
  assign n37109 = n37108 ^ n24991 ;
  assign n37112 = n37111 ^ n37109 ;
  assign n37116 = n36918 ^ n36917 ;
  assign n37113 = n34586 ^ n26486 ;
  assign n37114 = n37113 ^ n30695 ;
  assign n37115 = n37114 ^ n2373 ;
  assign n37117 = n37116 ^ n37115 ;
  assign n2217 = n2216 ^ n2165 ;
  assign n2230 = n2229 ^ n2217 ;
  assign n2234 = n2233 ^ n2230 ;
  assign n37165 = n37115 ^ n2234 ;
  assign n37118 = n36916 ^ n36902 ;
  assign n37119 = n37118 ^ n2234 ;
  assign n37123 = n36915 ^ n36904 ;
  assign n37120 = n34613 ^ n26497 ;
  assign n37121 = n37120 ^ n2131 ;
  assign n37122 = n37121 ^ n2224 ;
  assign n37124 = n37123 ^ n37122 ;
  assign n37126 = n34621 ^ n2014 ;
  assign n37127 = n37126 ^ n30705 ;
  assign n37128 = n37127 ^ n2111 ;
  assign n37125 = n36911 ^ n36906 ;
  assign n37129 = n37128 ^ n37125 ;
  assign n37133 = n36910 ^ n36908 ;
  assign n37150 = n37133 ^ n37128 ;
  assign n37130 = n34625 ^ n2002 ;
  assign n37131 = n37130 ^ n30709 ;
  assign n37132 = n37131 ^ n25009 ;
  assign n37134 = n37133 ^ n37132 ;
  assign n37138 = n36907 ^ n36576 ;
  assign n37147 = n37138 ^ n37132 ;
  assign n37135 = n25018 ^ n3081 ;
  assign n37136 = n37135 ^ n30714 ;
  assign n37137 = n37136 ^ n26112 ;
  assign n37139 = n37138 ^ n37137 ;
  assign n36533 = n34632 ^ n3052 ;
  assign n36534 = n36533 ^ n30718 ;
  assign n36535 = n36534 ^ n24700 ;
  assign n36489 = n34054 ^ n3040 ;
  assign n36490 = n36489 ^ n30721 ;
  assign n36491 = n36490 ^ n24696 ;
  assign n36488 = n35828 & n36487 ;
  assign n36492 = n36491 ^ n36488 ;
  assign n36529 = n36528 ^ n36526 ;
  assign n36530 = n36529 ^ n36491 ;
  assign n36531 = ~n36492 & ~n36530 ;
  assign n36532 = n36531 ^ n36529 ;
  assign n37140 = n36535 ^ n36532 ;
  assign n37141 = n37137 ^ n36576 ;
  assign n37142 = n37141 ^ n37137 ;
  assign n37143 = n37142 ^ n36532 ;
  assign n37144 = n37140 & ~n37143 ;
  assign n37145 = n37144 ^ n37141 ;
  assign n37146 = n37139 & ~n37145 ;
  assign n37148 = n37147 ^ n37146 ;
  assign n37149 = ~n37134 & ~n37148 ;
  assign n37151 = n37150 ^ n37149 ;
  assign n37152 = n37129 & ~n37151 ;
  assign n37153 = n37152 ^ n37128 ;
  assign n2098 = n2091 ^ n2064 ;
  assign n2117 = n2116 ^ n2098 ;
  assign n2124 = n2123 ^ n2117 ;
  assign n37154 = n37153 ^ n2124 ;
  assign n37155 = n36914 ^ n36912 ;
  assign n37158 = n37155 ^ n37153 ;
  assign n37159 = ~n37154 & n37158 ;
  assign n37156 = n37155 ^ n37122 ;
  assign n37160 = n37159 ^ n37156 ;
  assign n37161 = n37124 & ~n37160 ;
  assign n37162 = n37161 ^ n37123 ;
  assign n37163 = n37162 ^ n2234 ;
  assign n37164 = n37119 & n37163 ;
  assign n37166 = n37165 ^ n37164 ;
  assign n37167 = ~n37117 & ~n37166 ;
  assign n37168 = n37167 ^ n37116 ;
  assign n37169 = n37168 ^ n37109 ;
  assign n37170 = ~n37112 & ~n37169 ;
  assign n37110 = n37109 ^ n37105 ;
  assign n37171 = n37170 ^ n37110 ;
  assign n37172 = n37106 & n37171 ;
  assign n37173 = n37172 ^ n37105 ;
  assign n37174 = n37173 ^ n37098 ;
  assign n37175 = n37101 & n37174 ;
  assign n37099 = n37098 ^ n37094 ;
  assign n37176 = n37175 ^ n37099 ;
  assign n37177 = n37095 & n37176 ;
  assign n37178 = n37177 ^ n37094 ;
  assign n37179 = n37178 ^ n37086 ;
  assign n37180 = n37090 & ~n37179 ;
  assign n37182 = n37181 ^ n37180 ;
  assign n37183 = n37085 & ~n37182 ;
  assign n37185 = n37184 ^ n37183 ;
  assign n37186 = n37080 & n37185 ;
  assign n37187 = n37186 ^ n37079 ;
  assign n37188 = n37187 ^ n722 ;
  assign n37189 = ~n37075 & ~n37188 ;
  assign n37190 = n37189 ^ n37074 ;
  assign n37072 = n37071 ^ n37067 ;
  assign n37073 = n37072 ^ n37071 ;
  assign n37191 = n37190 ^ n37073 ;
  assign n37192 = n37068 & ~n37191 ;
  assign n37193 = n37192 ^ n37072 ;
  assign n37194 = n36939 ^ n36897 ;
  assign n37195 = n37194 ^ n37071 ;
  assign n37196 = n37193 & n37195 ;
  assign n37198 = n37197 ^ n37196 ;
  assign n37796 = n37199 ^ n37198 ;
  assign n37949 = n37796 ^ n35149 ;
  assign n37950 = n37949 ^ n37255 ;
  assign n37951 = n37950 ^ n37796 ;
  assign n37952 = n37948 & ~n37951 ;
  assign n37953 = n37952 ^ n37949 ;
  assign n37891 = n36676 ^ n35952 ;
  assign n37329 = n36457 ^ n36300 ;
  assign n37892 = n37329 ^ n36676 ;
  assign n37893 = n37891 & ~n37892 ;
  assign n37894 = n37893 ^ n35952 ;
  assign n37813 = n37194 ^ n37193 ;
  assign n37895 = n37894 ^ n37813 ;
  assign n37896 = n36650 ^ n35924 ;
  assign n37316 = n36453 ^ n36306 ;
  assign n37897 = n37316 ^ n36650 ;
  assign n37898 = n37896 & n37897 ;
  assign n37899 = n37898 ^ n35924 ;
  assign n37820 = n37190 ^ n37068 ;
  assign n37900 = n37899 ^ n37820 ;
  assign n37775 = n37176 ^ n37091 ;
  assign n36977 = n36437 ^ n36314 ;
  assign n37771 = n36977 ^ n36096 ;
  assign n37772 = n36096 ^ n34712 ;
  assign n37773 = ~n37771 & ~n37772 ;
  assign n37774 = n37773 ^ n34712 ;
  assign n37776 = n37775 ^ n37774 ;
  assign n36964 = n36434 ^ n36324 ;
  assign n37261 = n36964 ^ n35838 ;
  assign n37262 = n37173 ^ n37101 ;
  assign n37263 = n37262 ^ n35308 ;
  assign n37264 = n37263 ^ n36964 ;
  assign n37265 = n37264 ^ n37262 ;
  assign n37266 = n37261 & ~n37265 ;
  assign n37267 = n37266 ^ n37263 ;
  assign n37508 = n37171 ^ n37102 ;
  assign n37499 = n37168 ^ n37112 ;
  assign n37272 = n37166 ^ n37116 ;
  assign n37268 = n36794 ^ n35846 ;
  assign n37269 = n35846 ^ n34752 ;
  assign n37270 = n37268 & ~n37269 ;
  assign n37271 = n37270 ^ n34752 ;
  assign n37273 = n37272 ^ n37271 ;
  assign n37278 = n37162 ^ n37119 ;
  assign n37274 = n35856 ^ n34760 ;
  assign n37275 = n36590 ^ n34760 ;
  assign n37276 = n37274 & ~n37275 ;
  assign n37277 = n37276 ^ n35856 ;
  assign n37279 = n37278 ^ n37277 ;
  assign n37281 = n36061 ^ n34781 ;
  assign n37282 = n36782 ^ n36061 ;
  assign n37283 = n37281 & ~n37282 ;
  assign n37284 = n37283 ^ n34781 ;
  assign n37280 = n37160 ^ n37123 ;
  assign n37285 = n37284 ^ n37280 ;
  assign n37286 = n36597 ^ n36057 ;
  assign n37287 = n37155 ^ n2124 ;
  assign n37288 = n37287 ^ n37153 ;
  assign n37289 = n37288 ^ n35276 ;
  assign n37290 = n37289 ^ n36597 ;
  assign n37291 = n37290 ^ n37288 ;
  assign n37292 = ~n37286 & n37291 ;
  assign n37293 = n37292 ^ n37289 ;
  assign n37469 = n37148 ^ n37133 ;
  assign n37298 = n36611 ^ n35868 ;
  assign n37299 = n35868 ^ n35259 ;
  assign n37300 = n37298 & n37299 ;
  assign n37301 = n37300 ^ n35259 ;
  assign n37297 = n37145 ^ n37138 ;
  assign n37302 = n37301 ^ n37297 ;
  assign n36577 = n36576 ^ n36535 ;
  assign n36578 = n36577 ^ n36532 ;
  assign n37465 = n37301 ^ n36578 ;
  assign n37307 = n36529 ^ n36492 ;
  assign n37303 = n35876 ^ n34808 ;
  assign n37304 = n36624 ^ n35876 ;
  assign n37305 = ~n37303 & n37304 ;
  assign n37306 = n37305 ^ n34808 ;
  assign n37308 = n37307 ^ n37306 ;
  assign n36941 = n36896 & n36940 ;
  assign n36953 = n36894 ^ n36888 ;
  assign n36954 = n36893 & ~n36953 ;
  assign n36951 = n36431 ^ n36329 ;
  assign n36952 = n36951 ^ n36888 ;
  assign n36955 = n36954 ^ n36952 ;
  assign n36947 = n36220 ^ n34864 ;
  assign n36948 = n36220 ^ n35757 ;
  assign n36949 = ~n36947 & n36948 ;
  assign n36950 = n36949 ^ n34864 ;
  assign n36956 = n36955 ^ n36950 ;
  assign n36942 = n36895 ^ n34027 ;
  assign n36943 = n36895 ^ n36883 ;
  assign n36944 = ~n36942 & n36943 ;
  assign n36945 = n36944 ^ n34027 ;
  assign n36946 = n36945 ^ n34147 ;
  assign n36957 = n36956 ^ n36946 ;
  assign n36958 = ~n36941 & ~n36957 ;
  assign n36970 = n36951 ^ n36950 ;
  assign n36971 = n36955 & ~n36970 ;
  assign n36972 = n36971 ^ n36951 ;
  assign n36963 = n36479 ^ n35807 ;
  assign n36965 = n36964 ^ n34719 ;
  assign n36966 = n36965 ^ n36479 ;
  assign n36967 = n36966 ^ n36964 ;
  assign n36968 = n36963 & ~n36967 ;
  assign n36969 = n36968 ^ n36965 ;
  assign n36973 = n36972 ^ n36969 ;
  assign n36959 = n36956 ^ n36945 ;
  assign n36960 = n36946 & n36959 ;
  assign n36961 = n36960 ^ n34147 ;
  assign n36962 = n36961 ^ n34156 ;
  assign n36974 = n36973 ^ n36962 ;
  assign n36975 = n36958 & n36974 ;
  assign n36988 = n36973 ^ n34156 ;
  assign n36989 = n36973 ^ n36961 ;
  assign n36990 = n36988 & n36989 ;
  assign n36991 = n36990 ^ n34156 ;
  assign n36983 = n36972 ^ n36964 ;
  assign n36984 = ~n36969 & n36983 ;
  assign n36985 = n36984 ^ n36964 ;
  assign n36976 = n36513 ^ n35924 ;
  assign n36978 = n36977 ^ n34062 ;
  assign n36979 = n36978 ^ n36513 ;
  assign n36980 = n36979 ^ n36977 ;
  assign n36981 = n36976 & n36980 ;
  assign n36982 = n36981 ^ n36978 ;
  assign n36986 = n36985 ^ n36982 ;
  assign n36987 = n36986 ^ n34174 ;
  assign n36992 = n36991 ^ n36987 ;
  assign n36993 = n36975 & ~n36992 ;
  assign n37006 = n36441 ^ n36440 ;
  assign n37003 = n36985 ^ n36977 ;
  assign n37004 = n36982 & ~n37003 ;
  assign n36998 = n35952 ^ n35192 ;
  assign n36999 = n36561 ^ n35952 ;
  assign n37000 = n36998 & n36999 ;
  assign n37001 = n37000 ^ n35192 ;
  assign n37002 = n37001 ^ n36977 ;
  assign n37005 = n37004 ^ n37002 ;
  assign n37007 = n37006 ^ n37005 ;
  assign n37008 = n37007 ^ n34227 ;
  assign n36994 = n36991 ^ n36986 ;
  assign n36995 = n36991 ^ n34174 ;
  assign n36996 = ~n36994 & n36995 ;
  assign n36997 = n36996 ^ n36986 ;
  assign n37009 = n37008 ^ n36997 ;
  assign n37010 = ~n36993 & n37009 ;
  assign n37021 = n37006 ^ n37001 ;
  assign n37022 = ~n37005 & n37021 ;
  assign n37023 = n37022 ^ n37001 ;
  assign n37014 = n36650 ^ n35149 ;
  assign n37015 = n36445 ^ n36311 ;
  assign n37016 = n37015 ^ n34045 ;
  assign n37017 = n37016 ^ n36650 ;
  assign n37018 = n37017 ^ n37015 ;
  assign n37019 = n37014 & ~n37018 ;
  assign n37020 = n37019 ^ n37016 ;
  assign n37024 = n37023 ^ n37020 ;
  assign n37025 = n37024 ^ n33211 ;
  assign n37011 = n37007 ^ n36997 ;
  assign n37012 = ~n37008 & n37011 ;
  assign n37013 = n37012 ^ n34227 ;
  assign n37026 = n37025 ^ n37013 ;
  assign n37027 = n37010 & n37026 ;
  assign n37036 = n35155 ^ n34257 ;
  assign n37037 = n36676 ^ n35155 ;
  assign n37038 = ~n37036 & ~n37037 ;
  assign n37039 = n37038 ^ n34257 ;
  assign n37035 = n36447 ^ n36310 ;
  assign n37040 = n37039 ^ n37035 ;
  assign n37032 = n37023 ^ n37015 ;
  assign n37033 = ~n37020 & n37032 ;
  assign n37034 = n37033 ^ n37015 ;
  assign n37041 = n37040 ^ n37034 ;
  assign n37028 = n37024 ^ n37013 ;
  assign n37029 = ~n37025 & n37028 ;
  assign n37030 = n37029 ^ n33211 ;
  assign n37031 = n37030 ^ n33273 ;
  assign n37042 = n37041 ^ n37031 ;
  assign n37224 = n37027 & ~n37042 ;
  assign n37233 = n35143 ^ n34255 ;
  assign n37234 = n35732 ^ n35143 ;
  assign n37235 = ~n37233 & n37234 ;
  assign n37236 = n37235 ^ n34255 ;
  assign n37232 = n36450 ^ n36308 ;
  assign n37237 = n37236 ^ n37232 ;
  assign n37229 = n37035 ^ n37034 ;
  assign n37230 = ~n37040 & ~n37229 ;
  assign n37231 = n37230 ^ n37039 ;
  assign n37238 = n37237 ^ n37231 ;
  assign n37239 = n37238 ^ n33312 ;
  assign n37225 = n37041 ^ n33273 ;
  assign n37226 = n37041 ^ n37030 ;
  assign n37227 = n37225 & n37226 ;
  assign n37228 = n37227 ^ n33273 ;
  assign n37240 = n37239 ^ n37228 ;
  assign n37341 = n37224 & ~n37240 ;
  assign n37318 = n37232 ^ n37231 ;
  assign n37319 = ~n37237 & n37318 ;
  assign n37320 = n37319 ^ n37236 ;
  assign n37312 = n35141 ^ n34248 ;
  assign n37313 = n35775 ^ n35141 ;
  assign n37314 = n37312 & ~n37313 ;
  assign n37315 = n37314 ^ n34248 ;
  assign n37317 = n37316 ^ n37315 ;
  assign n37335 = n37320 ^ n37317 ;
  assign n37331 = n37238 ^ n37228 ;
  assign n37332 = ~n37239 & n37331 ;
  assign n37333 = n37332 ^ n33312 ;
  assign n37334 = n37333 ^ n33478 ;
  assign n37342 = n37335 ^ n37334 ;
  assign n37343 = ~n37341 & n37342 ;
  assign n37336 = n37335 ^ n37333 ;
  assign n37337 = n37334 & n37336 ;
  assign n37338 = n37337 ^ n33478 ;
  assign n37339 = n37338 ^ n33472 ;
  assign n37311 = n35812 ^ n35204 ;
  assign n37321 = n37320 ^ n37315 ;
  assign n37322 = ~n37317 & n37321 ;
  assign n37323 = n37322 ^ n37316 ;
  assign n37324 = n37323 ^ n34242 ;
  assign n37325 = n37324 ^ n35812 ;
  assign n37326 = n37325 ^ n37323 ;
  assign n37327 = n37311 & n37326 ;
  assign n37328 = n37327 ^ n37324 ;
  assign n37330 = n37329 ^ n37328 ;
  assign n37340 = n37339 ^ n37330 ;
  assign n37384 = n37343 ^ n37340 ;
  assign n37388 = n37387 ^ n37384 ;
  assign n37390 = n35047 ^ n26581 ;
  assign n37391 = n37390 ^ n2651 ;
  assign n37392 = n37391 ^ n3215 ;
  assign n37389 = n37342 ^ n37341 ;
  assign n37393 = n37392 ^ n37389 ;
  assign n37043 = n37042 ^ n37027 ;
  assign n37047 = n37046 ^ n37043 ;
  assign n37056 = n37026 ^ n37010 ;
  assign n37053 = n26450 ^ n1399 ;
  assign n37054 = n37053 ^ n30643 ;
  assign n37055 = n37054 ^ n2822 ;
  assign n37057 = n37056 ^ n37055 ;
  assign n37058 = n37009 ^ n36993 ;
  assign n37059 = n37058 ^ n2798 ;
  assign n1317 = n1277 ^ n1220 ;
  assign n1318 = n1317 ^ n1314 ;
  assign n1322 = n1321 ^ n1318 ;
  assign n37214 = n2798 ^ n1322 ;
  assign n37060 = n36992 ^ n36975 ;
  assign n37061 = n37060 ^ n1322 ;
  assign n37062 = n36974 ^ n36958 ;
  assign n1290 = n1205 ^ n1134 ;
  assign n1300 = n1299 ^ n1290 ;
  assign n1307 = n1306 ^ n1300 ;
  assign n37063 = n37062 ^ n1307 ;
  assign n1697 = n1678 ^ n1103 ;
  assign n1698 = n1697 ^ n1694 ;
  assign n1699 = n1698 ^ n1297 ;
  assign n37208 = n1699 ^ n1307 ;
  assign n37201 = n1699 ^ n1690 ;
  assign n37200 = n37199 ^ n1699 ;
  assign n37202 = n37201 ^ n37200 ;
  assign n37203 = n37198 & ~n37202 ;
  assign n37204 = n37203 ^ n37201 ;
  assign n37205 = n36957 ^ n36941 ;
  assign n37206 = n37205 ^ n1699 ;
  assign n37207 = n37204 & n37206 ;
  assign n37209 = n37208 ^ n37207 ;
  assign n37210 = n37063 & ~n37209 ;
  assign n37211 = n37210 ^ n37062 ;
  assign n37212 = n37211 ^ n1322 ;
  assign n37213 = ~n37061 & n37212 ;
  assign n37215 = n37214 ^ n37213 ;
  assign n37216 = n37059 & ~n37215 ;
  assign n37217 = n37216 ^ n37058 ;
  assign n37218 = n37217 ^ n37055 ;
  assign n37219 = ~n37057 & ~n37218 ;
  assign n37220 = n37219 ^ n37056 ;
  assign n37048 = n35051 ^ n26443 ;
  assign n37049 = n37048 ^ n30639 ;
  assign n37050 = n37049 ^ n2570 ;
  assign n37051 = n37050 ^ n37046 ;
  assign n37052 = n37051 ^ n37050 ;
  assign n37221 = n37220 ^ n37052 ;
  assign n37222 = n37047 & ~n37221 ;
  assign n37223 = n37222 ^ n37051 ;
  assign n37241 = n37240 ^ n37224 ;
  assign n37396 = n37241 ^ n37050 ;
  assign n37397 = ~n37223 & n37396 ;
  assign n37398 = n37397 ^ n37241 ;
  assign n37399 = n37398 ^ n37392 ;
  assign n37400 = ~n37393 & n37399 ;
  assign n37394 = n37392 ^ n37387 ;
  assign n37401 = n37400 ^ n37394 ;
  assign n37402 = n37388 & n37401 ;
  assign n37403 = n37402 ^ n37387 ;
  assign n37354 = n34130 ^ n34055 ;
  assign n37355 = n35977 ^ n34055 ;
  assign n37356 = ~n37354 & ~n37355 ;
  assign n37357 = n37356 ^ n34130 ;
  assign n37350 = n37329 ^ n37255 ;
  assign n37349 = n37323 ^ n37255 ;
  assign n37351 = n37350 ^ n37349 ;
  assign n37352 = n37328 & ~n37351 ;
  assign n37353 = n37352 ^ n37350 ;
  assign n37358 = n37357 ^ n37353 ;
  assign n37345 = n37338 ^ n37330 ;
  assign n37346 = ~n37339 & ~n37345 ;
  assign n37347 = n37346 ^ n33472 ;
  assign n37348 = n37347 ^ n33424 ;
  assign n37359 = n37358 ^ n37348 ;
  assign n37344 = n37340 & n37343 ;
  assign n37382 = n37359 ^ n37344 ;
  assign n37371 = n35042 ^ n26755 ;
  assign n37372 = n37371 ^ n30900 ;
  assign n37373 = n37372 ^ n3168 ;
  assign n37383 = n37382 ^ n37373 ;
  assign n37411 = n37403 ^ n37383 ;
  assign n37407 = n35896 ^ n34827 ;
  assign n37408 = n36633 ^ n35896 ;
  assign n37409 = n37407 & ~n37408 ;
  assign n37410 = n37409 ^ n34827 ;
  assign n37412 = n37411 ^ n37410 ;
  assign n37418 = n37398 ^ n37393 ;
  assign n36581 = n36580 ^ n36012 ;
  assign n36582 = n36012 ^ n34839 ;
  assign n36583 = ~n36581 & ~n36582 ;
  assign n36584 = n36583 ^ n34839 ;
  assign n37242 = n37241 ^ n37223 ;
  assign n37417 = ~n36584 & n37242 ;
  assign n37419 = n37418 ^ n37417 ;
  assign n37420 = n36723 ^ n35908 ;
  assign n37421 = n37417 ^ n35218 ;
  assign n37422 = n37421 ^ n36723 ;
  assign n37423 = n37422 ^ n37417 ;
  assign n37424 = ~n37420 & n37423 ;
  assign n37425 = n37424 ^ n37421 ;
  assign n37426 = ~n37419 & n37425 ;
  assign n37427 = n37426 ^ n37418 ;
  assign n37413 = n35902 ^ n34833 ;
  assign n37414 = n35902 ^ n35825 ;
  assign n37415 = ~n37413 & ~n37414 ;
  assign n37416 = n37415 ^ n34833 ;
  assign n37428 = n37427 ^ n37416 ;
  assign n37429 = n37401 ^ n37384 ;
  assign n37538 = n37429 ^ n37416 ;
  assign n37433 = n37428 & n37538 ;
  assign n37430 = n37429 ^ n37410 ;
  assign n37434 = n37433 ^ n37430 ;
  assign n37435 = ~n37412 & ~n37434 ;
  assign n37436 = n37435 ^ n37411 ;
  assign n37404 = n37403 ^ n37373 ;
  assign n37405 = ~n37383 & n37404 ;
  assign n37378 = n37357 ^ n37255 ;
  assign n37379 = ~n37353 & ~n37378 ;
  assign n3162 = n3161 ^ n3158 ;
  assign n3172 = n3171 ^ n3162 ;
  assign n3173 = n3172 ^ n2772 ;
  assign n37374 = n37373 ^ n3173 ;
  assign n37368 = n37357 ^ n34280 ;
  assign n37253 = n36462 ^ n36289 ;
  assign n37369 = n37368 ^ n37253 ;
  assign n37367 = n33424 ^ n33418 ;
  assign n37370 = n37369 ^ n37367 ;
  assign n37375 = n37374 ^ n37370 ;
  assign n37364 = n35965 ^ n34845 ;
  assign n37365 = n34845 ^ n34280 ;
  assign n37366 = ~n37364 & ~n37365 ;
  assign n37376 = n37375 ^ n37366 ;
  assign n37361 = n37358 ^ n37347 ;
  assign n37362 = n37358 ^ n33424 ;
  assign n37363 = n37361 & ~n37362 ;
  assign n37377 = n37376 ^ n37363 ;
  assign n37380 = n37379 ^ n37377 ;
  assign n37360 = n37344 & ~n37359 ;
  assign n37381 = n37380 ^ n37360 ;
  assign n37406 = n37405 ^ n37381 ;
  assign n37437 = n37436 ^ n37406 ;
  assign n37438 = n36626 ^ n35893 ;
  assign n37439 = n37406 ^ n34821 ;
  assign n37440 = n37439 ^ n36626 ;
  assign n37441 = n37440 ^ n37406 ;
  assign n37442 = n37438 & ~n37441 ;
  assign n37443 = n37442 ^ n37439 ;
  assign n37444 = ~n37437 & ~n37443 ;
  assign n37445 = n37444 ^ n37436 ;
  assign n37446 = n37445 ^ n37309 ;
  assign n37447 = n36741 ^ n35883 ;
  assign n37448 = n37309 ^ n34811 ;
  assign n37449 = n37448 ^ n36741 ;
  assign n37450 = n37449 ^ n37309 ;
  assign n37451 = ~n37447 & n37450 ;
  assign n37452 = n37451 ^ n37448 ;
  assign n37453 = ~n37446 & n37452 ;
  assign n37310 = n37309 ^ n37306 ;
  assign n37454 = n37453 ^ n37310 ;
  assign n37455 = n37308 & n37454 ;
  assign n37456 = n37455 ^ n37307 ;
  assign n37457 = n37456 ^ n36578 ;
  assign n37458 = n36614 ^ n34802 ;
  assign n37459 = n36578 ^ n35874 ;
  assign n37460 = n37459 ^ n36578 ;
  assign n37461 = n37460 ^ n34802 ;
  assign n37462 = ~n37458 & n37461 ;
  assign n37463 = n37462 ^ n37459 ;
  assign n37464 = n37457 & n37463 ;
  assign n37466 = n37465 ^ n37464 ;
  assign n37467 = ~n37302 & n37466 ;
  assign n37468 = n37467 ^ n37301 ;
  assign n37470 = n37469 ^ n37468 ;
  assign n37471 = n36600 ^ n35269 ;
  assign n37472 = n37469 ^ n35858 ;
  assign n37473 = n37472 ^ n37469 ;
  assign n37474 = n37473 ^ n35269 ;
  assign n37475 = ~n37471 & n37474 ;
  assign n37476 = n37475 ^ n37472 ;
  assign n37477 = n37470 & n37476 ;
  assign n37478 = n37477 ^ n37469 ;
  assign n37296 = n37151 ^ n37125 ;
  assign n37479 = n37478 ^ n37296 ;
  assign n37480 = n36606 ^ n34789 ;
  assign n37481 = n37296 ^ n36043 ;
  assign n37482 = n37481 ^ n36606 ;
  assign n37483 = n37482 ^ n37296 ;
  assign n37484 = ~n37480 & ~n37483 ;
  assign n37485 = n37484 ^ n37481 ;
  assign n37486 = n37479 & n37485 ;
  assign n37487 = n37486 ^ n37478 ;
  assign n37488 = n37487 ^ n37288 ;
  assign n37489 = ~n37293 & ~n37488 ;
  assign n37294 = n37288 ^ n37284 ;
  assign n37490 = n37489 ^ n37294 ;
  assign n37491 = n37285 & n37490 ;
  assign n37492 = n37491 ^ n37284 ;
  assign n37493 = n37492 ^ n37278 ;
  assign n37494 = n37279 & n37493 ;
  assign n37495 = n37494 ^ n37492 ;
  assign n37496 = n37495 ^ n37271 ;
  assign n37497 = ~n37273 & ~n37496 ;
  assign n37498 = n37497 ^ n37272 ;
  assign n37500 = n37499 ^ n37498 ;
  assign n37501 = n36894 ^ n35844 ;
  assign n37502 = n36894 ^ n34744 ;
  assign n37503 = ~n37501 & ~n37502 ;
  assign n37504 = n37503 ^ n35844 ;
  assign n37505 = n37504 ^ n37498 ;
  assign n37506 = ~n37500 & n37505 ;
  assign n37507 = n37506 ^ n37499 ;
  assign n37509 = n37508 ^ n37507 ;
  assign n37510 = n36951 ^ n36080 ;
  assign n37511 = n37508 ^ n34735 ;
  assign n37512 = n37511 ^ n36951 ;
  assign n37513 = n37512 ^ n37508 ;
  assign n37514 = n37510 & n37513 ;
  assign n37515 = n37514 ^ n37511 ;
  assign n37516 = n37509 & n37515 ;
  assign n37517 = n37516 ^ n37508 ;
  assign n37768 = n37517 ^ n37262 ;
  assign n37769 = ~n37267 & n37768 ;
  assign n37770 = n37769 ^ n37262 ;
  assign n37901 = n37774 ^ n37770 ;
  assign n37902 = n37776 & ~n37901 ;
  assign n37903 = n37902 ^ n37775 ;
  assign n37849 = n37178 ^ n37090 ;
  assign n37904 = n37903 ^ n37849 ;
  assign n37905 = n37006 ^ n36220 ;
  assign n37906 = n37903 ^ n35458 ;
  assign n37907 = n37906 ^ n37006 ;
  assign n37908 = n37907 ^ n37903 ;
  assign n37909 = ~n37905 & ~n37908 ;
  assign n37910 = n37909 ^ n37906 ;
  assign n37911 = n37904 & n37910 ;
  assign n37912 = n37911 ^ n37849 ;
  assign n37842 = n37182 ^ n37084 ;
  assign n37913 = n37912 ^ n37842 ;
  assign n37914 = n37015 ^ n36479 ;
  assign n37915 = n37842 ^ n35717 ;
  assign n37916 = n37915 ^ n37015 ;
  assign n37917 = n37916 ^ n37842 ;
  assign n37918 = ~n37914 & n37917 ;
  assign n37919 = n37918 ^ n37915 ;
  assign n37920 = n37913 & n37919 ;
  assign n37921 = n37920 ^ n37842 ;
  assign n37835 = n37185 ^ n37078 ;
  assign n37922 = n37921 ^ n37835 ;
  assign n37923 = n37035 ^ n35757 ;
  assign n37924 = n37835 ^ n36513 ;
  assign n37925 = n37924 ^ n37835 ;
  assign n37926 = n37925 ^ n35757 ;
  assign n37927 = n37923 & n37926 ;
  assign n37928 = n37927 ^ n37924 ;
  assign n37929 = n37922 & ~n37928 ;
  assign n37930 = n37929 ^ n37835 ;
  assign n37825 = n37187 ^ n37075 ;
  assign n37931 = n37930 ^ n37825 ;
  assign n37932 = n37232 ^ n36561 ;
  assign n37933 = n37825 ^ n35807 ;
  assign n37934 = n37933 ^ n37232 ;
  assign n37935 = n37934 ^ n37825 ;
  assign n37936 = n37932 & ~n37935 ;
  assign n37937 = n37936 ^ n37933 ;
  assign n37938 = ~n37931 & n37937 ;
  assign n37939 = n37938 ^ n37825 ;
  assign n37940 = n37939 ^ n37894 ;
  assign n37941 = n37940 ^ n37820 ;
  assign n37942 = n37941 ^ n37894 ;
  assign n37943 = n37900 & n37942 ;
  assign n37944 = n37943 ^ n37940 ;
  assign n37945 = n37895 & ~n37944 ;
  assign n37946 = n37945 ^ n37894 ;
  assign n37972 = n37953 ^ n37946 ;
  assign n37973 = n37972 ^ n34045 ;
  assign n37975 = n37939 ^ n37900 ;
  assign n37976 = n37975 ^ n34062 ;
  assign n37996 = n37937 ^ n37930 ;
  assign n37981 = n37910 ^ n37849 ;
  assign n37777 = n37776 ^ n37770 ;
  assign n37977 = n37777 ^ n34761 ;
  assign n37518 = n37517 ^ n37267 ;
  assign n37519 = n37518 ^ n34777 ;
  assign n37520 = n37515 ^ n37507 ;
  assign n37521 = n37520 ^ n34913 ;
  assign n37524 = n37495 ^ n37273 ;
  assign n37525 = n37524 ^ n34882 ;
  assign n37526 = n37492 ^ n37279 ;
  assign n37527 = n37526 ^ n34680 ;
  assign n37585 = n37490 ^ n37280 ;
  assign n37528 = n37487 ^ n37293 ;
  assign n37529 = n37528 ^ n34489 ;
  assign n37577 = n37485 ^ n37478 ;
  assign n37530 = n37476 ^ n37468 ;
  assign n37531 = n37530 ^ n34064 ;
  assign n37569 = n37466 ^ n37297 ;
  assign n37532 = n37463 ^ n37456 ;
  assign n37533 = n37532 ^ n34081 ;
  assign n37534 = n37452 ^ n37445 ;
  assign n37535 = n37534 ^ n34094 ;
  assign n37536 = n37434 ^ n37411 ;
  assign n37537 = n37536 ^ n34095 ;
  assign n37243 = n37242 ^ n36584 ;
  assign n37540 = ~n33325 & ~n37243 ;
  assign n37541 = n37540 ^ n34109 ;
  assign n37542 = n37425 ^ n37418 ;
  assign n37543 = n37542 ^ n37540 ;
  assign n37544 = ~n37541 & ~n37543 ;
  assign n37545 = n37544 ^ n34109 ;
  assign n37539 = n37538 ^ n37427 ;
  assign n37546 = n37545 ^ n37539 ;
  assign n37547 = n37545 ^ n34113 ;
  assign n37548 = ~n37546 & n37547 ;
  assign n37549 = n37548 ^ n34113 ;
  assign n37550 = n37549 ^ n37536 ;
  assign n37551 = ~n37537 & ~n37550 ;
  assign n37552 = n37551 ^ n34095 ;
  assign n37553 = n37552 ^ n34118 ;
  assign n37554 = n37443 ^ n37436 ;
  assign n37555 = n37554 ^ n37552 ;
  assign n37556 = ~n37553 & n37555 ;
  assign n37557 = n37556 ^ n34118 ;
  assign n37558 = n37557 ^ n37534 ;
  assign n37559 = ~n37535 & ~n37558 ;
  assign n37560 = n37559 ^ n34094 ;
  assign n37561 = n37560 ^ n34088 ;
  assign n37562 = n37454 ^ n37307 ;
  assign n37563 = n37562 ^ n37560 ;
  assign n37564 = ~n37561 & ~n37563 ;
  assign n37565 = n37564 ^ n34088 ;
  assign n37566 = n37565 ^ n37532 ;
  assign n37567 = n37533 & ~n37566 ;
  assign n37568 = n37567 ^ n34081 ;
  assign n37570 = n37569 ^ n37568 ;
  assign n37571 = n37569 ^ n34075 ;
  assign n37572 = n37570 & ~n37571 ;
  assign n37573 = n37572 ^ n34075 ;
  assign n37574 = n37573 ^ n37530 ;
  assign n37575 = n37531 & ~n37574 ;
  assign n37576 = n37575 ^ n34064 ;
  assign n37578 = n37577 ^ n37576 ;
  assign n37579 = n37577 ^ n34329 ;
  assign n37580 = n37578 & ~n37579 ;
  assign n37581 = n37580 ^ n34329 ;
  assign n37582 = n37581 ^ n37528 ;
  assign n37583 = ~n37529 & n37582 ;
  assign n37584 = n37583 ^ n34489 ;
  assign n37586 = n37585 ^ n37584 ;
  assign n37587 = n37585 ^ n34503 ;
  assign n37588 = n37586 & n37587 ;
  assign n37589 = n37588 ^ n34503 ;
  assign n37590 = n37589 ^ n37526 ;
  assign n37591 = n37527 & n37590 ;
  assign n37592 = n37591 ^ n34680 ;
  assign n37593 = n37592 ^ n37524 ;
  assign n37594 = ~n37525 & ~n37593 ;
  assign n37595 = n37594 ^ n34882 ;
  assign n37522 = n37504 ^ n37499 ;
  assign n37523 = n37522 ^ n37498 ;
  assign n37596 = n37595 ^ n37523 ;
  assign n37597 = n37595 ^ n34784 ;
  assign n37598 = n37596 & ~n37597 ;
  assign n37599 = n37598 ^ n34784 ;
  assign n37600 = n37599 ^ n37520 ;
  assign n37601 = n37521 & n37600 ;
  assign n37602 = n37601 ^ n34913 ;
  assign n37778 = n37602 ^ n37518 ;
  assign n37779 = ~n37519 & ~n37778 ;
  assign n37780 = n37779 ^ n37602 ;
  assign n37978 = n37780 ^ n37777 ;
  assign n37979 = ~n37977 & ~n37978 ;
  assign n37980 = n37979 ^ n34761 ;
  assign n37982 = n37981 ^ n37980 ;
  assign n37983 = n37980 ^ n34750 ;
  assign n37984 = n37982 & ~n37983 ;
  assign n37985 = n37984 ^ n37981 ;
  assign n37986 = n37985 ^ n34727 ;
  assign n37987 = n37919 ^ n37912 ;
  assign n37988 = n37987 ^ n37985 ;
  assign n37989 = ~n37986 & n37988 ;
  assign n37990 = n37989 ^ n34727 ;
  assign n37991 = n37990 ^ n34864 ;
  assign n37992 = n37928 ^ n37921 ;
  assign n37993 = n37992 ^ n37990 ;
  assign n37994 = ~n37991 & n37993 ;
  assign n37995 = n37994 ^ n34864 ;
  assign n37997 = n37996 ^ n37995 ;
  assign n37998 = n37996 ^ n34719 ;
  assign n37999 = n37997 & ~n37998 ;
  assign n38000 = n37999 ^ n34719 ;
  assign n38001 = n38000 ^ n37975 ;
  assign n38002 = ~n37976 & n38001 ;
  assign n38003 = n38002 ^ n34062 ;
  assign n37974 = n37944 ^ n37813 ;
  assign n38004 = n38003 ^ n37974 ;
  assign n38005 = n38003 ^ n35192 ;
  assign n38006 = ~n38004 & ~n38005 ;
  assign n38007 = n38006 ^ n35192 ;
  assign n38008 = n38007 ^ n37972 ;
  assign n38009 = ~n37973 & ~n38008 ;
  assign n38010 = n38009 ^ n34045 ;
  assign n38056 = n38010 ^ n34257 ;
  assign n37947 = n37946 ^ n37796 ;
  assign n37954 = ~n37947 & ~n37953 ;
  assign n37955 = n37954 ^ n37946 ;
  assign n37879 = n37253 ^ n35775 ;
  assign n37805 = n37205 ^ n37204 ;
  assign n37880 = n37805 ^ n35155 ;
  assign n37881 = n37880 ^ n37253 ;
  assign n37882 = n37881 ^ n37805 ;
  assign n37883 = n37879 & ~n37882 ;
  assign n37884 = n37883 ^ n37880 ;
  assign n38011 = n37955 ^ n37884 ;
  assign n38057 = n38056 ^ n38011 ;
  assign n37781 = n37780 ^ n34761 ;
  assign n37782 = n37781 ^ n37777 ;
  assign n37603 = n37602 ^ n37519 ;
  assign n37604 = n37584 ^ n34503 ;
  assign n37605 = n37604 ^ n37585 ;
  assign n37606 = n37562 ^ n37561 ;
  assign n37607 = n37557 ^ n37535 ;
  assign n37608 = n37547 ^ n37539 ;
  assign n37609 = n37549 ^ n37537 ;
  assign n37610 = n37608 & ~n37609 ;
  assign n37611 = n37554 ^ n37553 ;
  assign n37612 = n37610 & ~n37611 ;
  assign n37613 = n37607 & ~n37612 ;
  assign n37614 = n37606 & ~n37613 ;
  assign n37615 = n37565 ^ n37533 ;
  assign n37616 = n37614 & n37615 ;
  assign n37617 = n37568 ^ n34075 ;
  assign n37618 = n37617 ^ n37569 ;
  assign n37619 = ~n37616 & n37618 ;
  assign n37620 = n37573 ^ n37531 ;
  assign n37621 = n37619 & ~n37620 ;
  assign n37622 = n37576 ^ n34329 ;
  assign n37623 = n37622 ^ n37577 ;
  assign n37624 = ~n37621 & ~n37623 ;
  assign n37625 = n37581 ^ n37529 ;
  assign n37626 = n37624 & ~n37625 ;
  assign n37627 = n37605 & n37626 ;
  assign n37628 = n37589 ^ n37527 ;
  assign n37629 = n37627 & ~n37628 ;
  assign n37630 = n37592 ^ n34882 ;
  assign n37631 = n37630 ^ n37524 ;
  assign n37632 = ~n37629 & n37631 ;
  assign n37633 = n37523 ^ n34784 ;
  assign n37634 = n37633 ^ n37595 ;
  assign n37635 = ~n37632 & ~n37634 ;
  assign n37636 = n37599 ^ n37521 ;
  assign n37637 = n37635 & n37636 ;
  assign n37783 = ~n37603 & n37637 ;
  assign n38037 = ~n37782 & ~n37783 ;
  assign n38038 = n37981 ^ n34750 ;
  assign n38039 = n38038 ^ n37980 ;
  assign n38040 = ~n38037 & n38039 ;
  assign n38041 = n37987 ^ n37986 ;
  assign n38042 = n38040 & n38041 ;
  assign n38043 = n37992 ^ n34864 ;
  assign n38044 = n38043 ^ n37990 ;
  assign n38045 = ~n38042 & n38044 ;
  assign n38046 = n37995 ^ n34719 ;
  assign n38047 = n38046 ^ n37996 ;
  assign n38048 = n38045 & n38047 ;
  assign n38049 = n38000 ^ n37976 ;
  assign n38050 = n38048 & n38049 ;
  assign n38051 = n37974 ^ n35192 ;
  assign n38052 = n38051 ^ n38003 ;
  assign n38053 = ~n38050 & ~n38052 ;
  assign n38054 = n38007 ^ n37973 ;
  assign n38055 = n38053 & n38054 ;
  assign n38078 = n38057 ^ n38055 ;
  assign n2875 = n2867 ^ n2850 ;
  assign n2888 = n2887 ^ n2875 ;
  assign n2895 = n2894 ^ n2888 ;
  assign n38079 = n38078 ^ n2895 ;
  assign n38081 = n35529 ^ n2811 ;
  assign n38082 = n38081 ^ n2882 ;
  assign n38083 = n38082 ^ n31522 ;
  assign n38080 = n38054 ^ n38053 ;
  assign n38084 = n38083 ^ n38080 ;
  assign n38086 = n35534 ^ n1435 ;
  assign n38087 = n38086 ^ n1385 ;
  assign n38088 = n38087 ^ n1773 ;
  assign n38085 = n38052 ^ n38050 ;
  assign n38089 = n38088 ^ n38085 ;
  assign n38090 = n38049 ^ n38048 ;
  assign n1761 = n1739 ^ n1410 ;
  assign n1762 = n1761 ^ n1160 ;
  assign n1766 = n1765 ^ n1762 ;
  assign n38091 = n38090 ^ n1766 ;
  assign n38092 = n38047 ^ n38045 ;
  assign n1752 = n1730 ^ n1418 ;
  assign n1756 = n1755 ^ n1752 ;
  assign n1757 = n1756 ^ n1151 ;
  assign n38093 = n38092 ^ n1757 ;
  assign n38094 = n38044 ^ n38042 ;
  assign n984 = n983 ^ n929 ;
  assign n997 = n996 ^ n984 ;
  assign n1004 = n1003 ^ n997 ;
  assign n38095 = n38094 ^ n1004 ;
  assign n38099 = n38041 ^ n38040 ;
  assign n38096 = n35545 ^ n1707 ;
  assign n38097 = n38096 ^ n892 ;
  assign n38098 = n38097 ^ n991 ;
  assign n38100 = n38099 ^ n38098 ;
  assign n38101 = n38039 ^ n38037 ;
  assign n38102 = n38101 ^ n885 ;
  assign n37784 = n37783 ^ n37782 ;
  assign n37785 = n37784 ^ n37767 ;
  assign n37638 = n37637 ^ n37603 ;
  assign n37639 = n37638 ^ n1595 ;
  assign n37640 = n37636 ^ n37635 ;
  assign n37644 = n37643 ^ n37640 ;
  assign n37645 = n35558 ^ n1548 ;
  assign n37646 = n37645 ^ n31390 ;
  assign n37647 = n37646 ^ n2960 ;
  assign n37758 = n37647 ^ n37640 ;
  assign n37648 = n37634 ^ n37632 ;
  assign n37649 = n37648 ^ n37647 ;
  assign n37653 = n37631 ^ n37629 ;
  assign n37650 = n35568 ^ n27195 ;
  assign n37651 = n37650 ^ n2948 ;
  assign n37652 = n37651 ^ n25814 ;
  assign n37654 = n37653 ^ n37652 ;
  assign n37655 = n37628 ^ n37627 ;
  assign n37659 = n37658 ^ n37655 ;
  assign n37663 = n35573 ^ n2930 ;
  assign n37664 = n37663 ^ n25823 ;
  assign n37665 = n37664 ^ n31403 ;
  assign n37662 = n37626 ^ n37605 ;
  assign n37666 = n37665 ^ n37662 ;
  assign n37671 = n37625 ^ n37624 ;
  assign n37667 = n35578 ^ n27208 ;
  assign n37668 = n37667 ^ n31461 ;
  assign n37669 = n37668 ^ n25827 ;
  assign n37672 = n37671 ^ n37669 ;
  assign n37676 = n37623 ^ n37621 ;
  assign n37673 = n27212 ^ n2391 ;
  assign n37674 = n37673 ^ n31407 ;
  assign n37675 = n37674 ^ n25832 ;
  assign n37677 = n37676 ^ n37675 ;
  assign n37678 = n37620 ^ n37619 ;
  assign n2358 = n2314 ^ n2278 ;
  assign n2357 = n2356 ^ n2348 ;
  assign n2359 = n2358 ^ n2357 ;
  assign n37679 = n37678 ^ n2359 ;
  assign n37680 = n37618 ^ n37616 ;
  assign n2318 = n2305 ^ n2260 ;
  assign n2334 = n2333 ^ n2318 ;
  assign n2341 = n2340 ^ n2334 ;
  assign n37681 = n37680 ^ n2341 ;
  assign n37684 = n35594 ^ n31423 ;
  assign n37685 = n37684 ^ n2180 ;
  assign n37686 = n37685 ^ n25842 ;
  assign n37683 = n37613 ^ n37606 ;
  assign n37687 = n37686 ^ n37683 ;
  assign n37689 = n35624 ^ n27222 ;
  assign n37690 = n37689 ^ n31428 ;
  assign n37691 = n37690 ^ n25868 ;
  assign n37688 = n37612 ^ n37607 ;
  assign n37692 = n37691 ^ n37688 ;
  assign n37716 = n37611 ^ n37610 ;
  assign n37693 = n35612 ^ n27240 ;
  assign n37694 = n37693 ^ n25850 ;
  assign n37695 = n37694 ^ n1895 ;
  assign n37696 = n37695 ^ n37609 ;
  assign n37697 = n37696 ^ n37608 ;
  assign n37698 = n35599 ^ n1890 ;
  assign n37699 = n37698 ^ n27230 ;
  assign n37700 = n37699 ^ n30821 ;
  assign n37701 = n37700 ^ n37608 ;
  assign n37244 = n37243 ^ n33325 ;
  assign n37245 = n35958 ^ n3183 ;
  assign n37246 = n37245 ^ n3200 ;
  assign n37247 = n37246 ^ n2705 ;
  assign n37705 = n37244 & n37247 ;
  assign n37706 = n37705 ^ n37704 ;
  assign n37707 = n37542 ^ n37541 ;
  assign n37708 = n37707 ^ n37704 ;
  assign n37709 = n37706 & n37708 ;
  assign n37710 = n37709 ^ n37705 ;
  assign n37711 = n37710 ^ n37700 ;
  assign n37712 = n37701 & ~n37711 ;
  assign n37713 = n37712 ^ n37609 ;
  assign n37714 = n37697 & ~n37713 ;
  assign n37715 = n37714 ^ n37695 ;
  assign n37717 = n37716 ^ n37715 ;
  assign n37718 = n35616 ^ n27226 ;
  assign n37719 = n37718 ^ n31435 ;
  assign n37720 = n37719 ^ n1943 ;
  assign n37721 = n37720 ^ n37715 ;
  assign n37722 = n37717 & ~n37721 ;
  assign n37723 = n37722 ^ n37716 ;
  assign n37724 = n37723 ^ n37688 ;
  assign n37725 = ~n37692 & n37724 ;
  assign n37726 = n37725 ^ n37691 ;
  assign n37727 = n37726 ^ n37686 ;
  assign n37728 = n37687 & n37727 ;
  assign n37729 = n37728 ^ n37686 ;
  assign n37736 = n37729 ^ n37680 ;
  assign n37682 = n37615 ^ n37614 ;
  assign n37730 = n37729 ^ n37682 ;
  assign n37731 = n35590 ^ n2192 ;
  assign n37732 = n37731 ^ n31418 ;
  assign n37733 = n37732 ^ n2330 ;
  assign n37734 = n37733 ^ n37682 ;
  assign n37735 = ~n37730 & n37734 ;
  assign n37737 = n37736 ^ n37735 ;
  assign n37738 = ~n37681 & n37737 ;
  assign n37739 = n37738 ^ n2341 ;
  assign n37740 = n37739 ^ n2359 ;
  assign n37741 = ~n37679 & ~n37740 ;
  assign n37742 = n37741 ^ n37678 ;
  assign n37743 = n37742 ^ n37675 ;
  assign n37744 = ~n37677 & ~n37743 ;
  assign n37745 = n37744 ^ n37675 ;
  assign n37746 = n37745 ^ n37669 ;
  assign n37747 = n37672 & n37746 ;
  assign n37670 = n37669 ^ n37662 ;
  assign n37748 = n37747 ^ n37670 ;
  assign n37749 = ~n37666 & n37748 ;
  assign n37750 = n37749 ^ n37665 ;
  assign n37751 = n37750 ^ n37658 ;
  assign n37752 = n37659 & n37751 ;
  assign n37660 = n37658 ^ n37653 ;
  assign n37753 = n37752 ^ n37660 ;
  assign n37754 = ~n37654 & ~n37753 ;
  assign n37755 = n37754 ^ n37653 ;
  assign n37756 = n37755 ^ n37647 ;
  assign n37757 = ~n37649 & ~n37756 ;
  assign n37759 = n37758 ^ n37757 ;
  assign n37760 = ~n37644 & n37759 ;
  assign n37761 = n37760 ^ n37643 ;
  assign n37762 = n37761 ^ n1595 ;
  assign n37763 = n37639 & ~n37762 ;
  assign n37764 = n37763 ^ n37638 ;
  assign n38103 = n37767 ^ n37764 ;
  assign n38104 = n37785 & ~n38103 ;
  assign n38105 = n38104 ^ n37784 ;
  assign n38106 = n38105 ^ n885 ;
  assign n38107 = n38102 & ~n38106 ;
  assign n38108 = n38107 ^ n38101 ;
  assign n38109 = n38108 ^ n38098 ;
  assign n38110 = ~n38100 & ~n38109 ;
  assign n38111 = n38110 ^ n38099 ;
  assign n38112 = n38111 ^ n1004 ;
  assign n38113 = ~n38095 & n38112 ;
  assign n38114 = n38113 ^ n38094 ;
  assign n38115 = n38114 ^ n1757 ;
  assign n38116 = n38093 & n38115 ;
  assign n38117 = n38116 ^ n38092 ;
  assign n38118 = n38117 ^ n38090 ;
  assign n38119 = n38091 & ~n38118 ;
  assign n38120 = n38119 ^ n1766 ;
  assign n38121 = n38120 ^ n38085 ;
  assign n38122 = ~n38089 & n38121 ;
  assign n38123 = n38122 ^ n38088 ;
  assign n38124 = n38123 ^ n38080 ;
  assign n38125 = ~n38084 & n38124 ;
  assign n38126 = n38125 ^ n38083 ;
  assign n38127 = n38126 ^ n2895 ;
  assign n38128 = n38079 & ~n38127 ;
  assign n38129 = n38128 ^ n38078 ;
  assign n38058 = n38055 & ~n38057 ;
  assign n38012 = n38011 ^ n38010 ;
  assign n38013 = n38011 ^ n34257 ;
  assign n38014 = n38012 & ~n38013 ;
  assign n38015 = n38014 ^ n34257 ;
  assign n37885 = n35812 ^ n35143 ;
  assign n37886 = n36485 ^ n35812 ;
  assign n37887 = n37885 & ~n37886 ;
  assign n37888 = n37887 ^ n35143 ;
  assign n37889 = n37888 ^ n37805 ;
  assign n37890 = n37889 ^ n37888 ;
  assign n37956 = n37955 ^ n37890 ;
  assign n37957 = n37884 & n37956 ;
  assign n37958 = n37957 ^ n37889 ;
  assign n37791 = n37209 ^ n37062 ;
  assign n37970 = n37958 ^ n37791 ;
  assign n37971 = n37970 ^ n34255 ;
  assign n38036 = n38015 ^ n37971 ;
  assign n38074 = n38058 ^ n38036 ;
  assign n38071 = n34061 ^ n27168 ;
  assign n38072 = n38071 ^ n2902 ;
  assign n38073 = n38072 ^ n3116 ;
  assign n38075 = n38074 ^ n38073 ;
  assign n38167 = n38129 ^ n38075 ;
  assign n38365 = n38171 ^ n38167 ;
  assign n38640 = n38365 ^ n34839 ;
  assign n2758 = n2750 ^ n2724 ;
  assign n2768 = n2767 ^ n2758 ;
  assign n2775 = n2774 ^ n2768 ;
  assign n38935 = n38640 ^ n2775 ;
  assign n38247 = n37710 ^ n37701 ;
  assign n39679 = n38935 ^ n38247 ;
  assign n39680 = n38935 ^ n36578 ;
  assign n39681 = n39679 & n39680 ;
  assign n39682 = n39681 ^ n36578 ;
  assign n38951 = n38123 ^ n38084 ;
  assign n39513 = n38951 ^ n37242 ;
  assign n37819 = n37015 ^ n36096 ;
  assign n37821 = n37820 ^ n37015 ;
  assign n37822 = ~n37819 & n37821 ;
  assign n37823 = n37822 ^ n36096 ;
  assign n37818 = n37750 ^ n37659 ;
  assign n37824 = n37823 ^ n37818 ;
  assign n37826 = n37825 ^ n37006 ;
  assign n37827 = n37748 ^ n37665 ;
  assign n37828 = n37827 ^ n35838 ;
  assign n37829 = n37828 ^ n37825 ;
  assign n37830 = n37829 ^ n37827 ;
  assign n37831 = n37826 & n37830 ;
  assign n37832 = n37831 ^ n37828 ;
  assign n37834 = n36977 ^ n36080 ;
  assign n37836 = n37835 ^ n36977 ;
  assign n37837 = n37834 & n37836 ;
  assign n37838 = n37837 ^ n36080 ;
  assign n37833 = n37745 ^ n37672 ;
  assign n37839 = n37838 ^ n37833 ;
  assign n37841 = n36964 ^ n35844 ;
  assign n37843 = n37842 ^ n36964 ;
  assign n37844 = n37841 & ~n37843 ;
  assign n37845 = n37844 ^ n35844 ;
  assign n37840 = n37742 ^ n37677 ;
  assign n37846 = n37845 ^ n37840 ;
  assign n37848 = n36951 ^ n35846 ;
  assign n37850 = n37849 ^ n36951 ;
  assign n37851 = ~n37848 & ~n37850 ;
  assign n37852 = n37851 ^ n35846 ;
  assign n37847 = n37739 ^ n37679 ;
  assign n37853 = n37852 ^ n37847 ;
  assign n38280 = n37737 ^ n2341 ;
  assign n37855 = n36794 ^ n36061 ;
  assign n37856 = n37262 ^ n36794 ;
  assign n37857 = n37855 & ~n37856 ;
  assign n37858 = n37857 ^ n36061 ;
  assign n37854 = n37734 ^ n37729 ;
  assign n37859 = n37858 ^ n37854 ;
  assign n37860 = n37508 ^ n36590 ;
  assign n37861 = n37726 ^ n37687 ;
  assign n37862 = n37861 ^ n36057 ;
  assign n37863 = n37862 ^ n37508 ;
  assign n37864 = n37863 ^ n37861 ;
  assign n37865 = n37860 & ~n37864 ;
  assign n37866 = n37865 ^ n37862 ;
  assign n37873 = n37723 ^ n37692 ;
  assign n37869 = n36782 ^ n36043 ;
  assign n37870 = n37499 ^ n36782 ;
  assign n37871 = n37869 & ~n37870 ;
  assign n37872 = n37871 ^ n36043 ;
  assign n37874 = n37873 ^ n37872 ;
  assign n38267 = n37720 ^ n37716 ;
  assign n38268 = n38267 ^ n37715 ;
  assign n38271 = n38268 ^ n37872 ;
  assign n38222 = n37296 ^ n36614 ;
  assign n38223 = n36614 ^ n35883 ;
  assign n38224 = ~n38222 & ~n38223 ;
  assign n38225 = n38224 ^ n35883 ;
  assign n37959 = n35977 ^ n35141 ;
  assign n37960 = n36525 ^ n35977 ;
  assign n37961 = n37959 & n37960 ;
  assign n37962 = n37961 ^ n35141 ;
  assign n37964 = n37962 ^ n37888 ;
  assign n37963 = n37962 ^ n37791 ;
  assign n37965 = n37964 ^ n37963 ;
  assign n37966 = n37958 & n37965 ;
  assign n37967 = n37966 ^ n37964 ;
  assign n38023 = n36566 ^ n35965 ;
  assign n38024 = n35965 ^ n35204 ;
  assign n38025 = ~n38023 & n38024 ;
  assign n38026 = n38025 ^ n35204 ;
  assign n38028 = n38026 ^ n37962 ;
  assign n37257 = n37211 ^ n37061 ;
  assign n38027 = n38026 ^ n37257 ;
  assign n38029 = n38028 ^ n38027 ;
  assign n38030 = n37967 & ~n38029 ;
  assign n38031 = n38030 ^ n38028 ;
  assign n38147 = n37217 ^ n37057 ;
  assign n38149 = n38147 ^ n38026 ;
  assign n37252 = n37215 ^ n37058 ;
  assign n38148 = n38147 ^ n37252 ;
  assign n38150 = n38149 ^ n38148 ;
  assign n38151 = n38031 & ~n38150 ;
  assign n38152 = n38151 ^ n38148 ;
  assign n38143 = n35830 ^ n34055 ;
  assign n38144 = n36699 ^ n34055 ;
  assign n38145 = n38143 & n38144 ;
  assign n38146 = n38145 ^ n35830 ;
  assign n38153 = n38152 ^ n38146 ;
  assign n37968 = n37967 ^ n37257 ;
  assign n37969 = n37968 ^ n34248 ;
  assign n38016 = n38015 ^ n37970 ;
  assign n38017 = ~n37971 & n38016 ;
  assign n38018 = n38017 ^ n34255 ;
  assign n38019 = n38018 ^ n37968 ;
  assign n38020 = ~n37969 & ~n38019 ;
  assign n38021 = n38020 ^ n34248 ;
  assign n38022 = n38021 ^ n34242 ;
  assign n38032 = n38031 ^ n37252 ;
  assign n38139 = n38032 ^ n38021 ;
  assign n38140 = n38022 & n38139 ;
  assign n38141 = n38140 ^ n34242 ;
  assign n38142 = n38141 ^ n34130 ;
  assign n38154 = n38153 ^ n38142 ;
  assign n38033 = n38032 ^ n38022 ;
  assign n38034 = n38018 ^ n34248 ;
  assign n38035 = n38034 ^ n37968 ;
  assign n38059 = ~n38036 & n38058 ;
  assign n38060 = n38035 & ~n38059 ;
  assign n38138 = ~n38033 & n38060 ;
  assign n38155 = n38154 ^ n38138 ;
  assign n2658 = n2657 ^ n2522 ;
  assign n2659 = n2658 ^ n2636 ;
  assign n2660 = n2659 ^ n2612 ;
  assign n38156 = n38155 ^ n2660 ;
  assign n38062 = n35773 ^ n3218 ;
  assign n38063 = n38062 ^ n31774 ;
  assign n38064 = n38063 ^ n2607 ;
  assign n38061 = n38060 ^ n38033 ;
  assign n38065 = n38064 ^ n38061 ;
  assign n38067 = n35731 ^ n2582 ;
  assign n38068 = n38067 ^ n25949 ;
  assign n38069 = n38068 ^ n31577 ;
  assign n38066 = n38059 ^ n38035 ;
  assign n38070 = n38069 ^ n38066 ;
  assign n38130 = n38129 ^ n38073 ;
  assign n38131 = n38075 & n38130 ;
  assign n38076 = n38073 ^ n38066 ;
  assign n38132 = n38131 ^ n38076 ;
  assign n38133 = ~n38070 & n38132 ;
  assign n38134 = n38133 ^ n38069 ;
  assign n38135 = n38134 ^ n38064 ;
  assign n38136 = ~n38065 & n38135 ;
  assign n38137 = n38136 ^ n38064 ;
  assign n38211 = n38137 ^ n2660 ;
  assign n38212 = n38156 & n38211 ;
  assign n38206 = n36001 ^ n34845 ;
  assign n38207 = n36697 ^ n36001 ;
  assign n38208 = ~n38206 & n38207 ;
  assign n38202 = n38201 ^ n2660 ;
  assign n38197 = n34280 ^ n34130 ;
  assign n38195 = n37220 ^ n37047 ;
  assign n38194 = n38147 ^ n34845 ;
  assign n38196 = n38195 ^ n38194 ;
  assign n38198 = n38197 ^ n38196 ;
  assign n38203 = n38202 ^ n38198 ;
  assign n38192 = n38147 ^ n38146 ;
  assign n38193 = ~n38152 & ~n38192 ;
  assign n38204 = n38203 ^ n38193 ;
  assign n38189 = n38153 ^ n38141 ;
  assign n38190 = n38153 ^ n34130 ;
  assign n38191 = n38189 & n38190 ;
  assign n38205 = n38204 ^ n38191 ;
  assign n38209 = n38208 ^ n38205 ;
  assign n38188 = n38138 & n38154 ;
  assign n38210 = n38209 ^ n38188 ;
  assign n38213 = n38212 ^ n38210 ;
  assign n38226 = n38225 ^ n38213 ;
  assign n38157 = n38156 ^ n38137 ;
  assign n37875 = n37297 ^ n36741 ;
  assign n37876 = n37297 ^ n35896 ;
  assign n37877 = ~n37875 & n37876 ;
  assign n37878 = n37877 ^ n35896 ;
  assign n38158 = n38157 ^ n37878 ;
  assign n38160 = n38134 ^ n38065 ;
  assign n38184 = n38160 ^ n37878 ;
  assign n38159 = n36626 ^ n36578 ;
  assign n38161 = n38160 ^ n35902 ;
  assign n38162 = n38161 ^ n36626 ;
  assign n38163 = n38162 ^ n38160 ;
  assign n38164 = ~n38159 & n38163 ;
  assign n38165 = n38164 ^ n38161 ;
  assign n38172 = n38167 & n38171 ;
  assign n38166 = n38132 ^ n38069 ;
  assign n38173 = n38172 ^ n38166 ;
  assign n38174 = n37307 ^ n36633 ;
  assign n38175 = n38172 ^ n35908 ;
  assign n38176 = n38175 ^ n36633 ;
  assign n38177 = n38176 ^ n38172 ;
  assign n38178 = n38174 & ~n38177 ;
  assign n38179 = n38178 ^ n38175 ;
  assign n38180 = ~n38173 & ~n38179 ;
  assign n38181 = n38180 ^ n38172 ;
  assign n38182 = n38181 ^ n38160 ;
  assign n38183 = n38165 & ~n38182 ;
  assign n38185 = n38184 ^ n38183 ;
  assign n38186 = n38158 & n38185 ;
  assign n38187 = n38186 ^ n38157 ;
  assign n38214 = n38213 ^ n38187 ;
  assign n38215 = n37469 ^ n36624 ;
  assign n38216 = n38213 ^ n35893 ;
  assign n38217 = n38216 ^ n36624 ;
  assign n38218 = n38217 ^ n38213 ;
  assign n38219 = ~n38215 & ~n38218 ;
  assign n38220 = n38219 ^ n38216 ;
  assign n38221 = ~n38214 & ~n38220 ;
  assign n38227 = n38226 ^ n38221 ;
  assign n38228 = n37288 ^ n36611 ;
  assign n38229 = n37288 ^ n35876 ;
  assign n38230 = ~n38228 & n38229 ;
  assign n38231 = n38230 ^ n35876 ;
  assign n38232 = n38231 ^ n38225 ;
  assign n38233 = n38232 ^ n38231 ;
  assign n37248 = n37247 ^ n37244 ;
  assign n38234 = n38233 ^ n37248 ;
  assign n38235 = ~n38227 & n38234 ;
  assign n38236 = n38235 ^ n38232 ;
  assign n38238 = n36600 ^ n35874 ;
  assign n38239 = n37280 ^ n36600 ;
  assign n38240 = n38238 & n38239 ;
  assign n38241 = n38240 ^ n35874 ;
  assign n38243 = n38241 ^ n38231 ;
  assign n38237 = n37707 ^ n37706 ;
  assign n38242 = n38241 ^ n38237 ;
  assign n38244 = n38243 ^ n38242 ;
  assign n38245 = n38236 & ~n38244 ;
  assign n38246 = n38245 ^ n38243 ;
  assign n38248 = n36606 ^ n35868 ;
  assign n38249 = n37278 ^ n36606 ;
  assign n38250 = n38248 & n38249 ;
  assign n38251 = n38250 ^ n35868 ;
  assign n38253 = n38251 ^ n38241 ;
  assign n38252 = n38251 ^ n38247 ;
  assign n38254 = n38253 ^ n38252 ;
  assign n38255 = ~n38246 & ~n38254 ;
  assign n38256 = n38255 ^ n38253 ;
  assign n38262 = n37713 ^ n37695 ;
  assign n38257 = n36597 ^ n35858 ;
  assign n38258 = n37272 ^ n36597 ;
  assign n38259 = n38257 & ~n38258 ;
  assign n38260 = n38259 ^ n35858 ;
  assign n38261 = n38260 ^ n38251 ;
  assign n38263 = n38262 ^ n38261 ;
  assign n38264 = n38263 ^ n38260 ;
  assign n38265 = n38256 & ~n38264 ;
  assign n38266 = n38265 ^ n38261 ;
  assign n38269 = n38268 ^ n38260 ;
  assign n38270 = ~n38266 & ~n38269 ;
  assign n38272 = n38271 ^ n38270 ;
  assign n38273 = ~n37874 & ~n38272 ;
  assign n38274 = n38273 ^ n37873 ;
  assign n38275 = n38274 ^ n37861 ;
  assign n38276 = ~n37866 & ~n38275 ;
  assign n37867 = n37861 ^ n37858 ;
  assign n38277 = n38276 ^ n37867 ;
  assign n38278 = ~n37859 & n38277 ;
  assign n38279 = n38278 ^ n37858 ;
  assign n38281 = n38280 ^ n38279 ;
  assign n38282 = n37775 ^ n36894 ;
  assign n38283 = n38280 ^ n35856 ;
  assign n38284 = n38283 ^ n37775 ;
  assign n38285 = n38284 ^ n38280 ;
  assign n38286 = n38282 & ~n38285 ;
  assign n38287 = n38286 ^ n38283 ;
  assign n38288 = ~n38281 & n38287 ;
  assign n38289 = n38288 ^ n38280 ;
  assign n38290 = n38289 ^ n37847 ;
  assign n38291 = n37853 & ~n38290 ;
  assign n38292 = n38291 ^ n37852 ;
  assign n38293 = n38292 ^ n37840 ;
  assign n38294 = n37846 & n38293 ;
  assign n38295 = n38294 ^ n37845 ;
  assign n38296 = n38295 ^ n37833 ;
  assign n38297 = ~n37839 & ~n38296 ;
  assign n38298 = n38297 ^ n37838 ;
  assign n38299 = n38298 ^ n37827 ;
  assign n38300 = n37832 & n38299 ;
  assign n38301 = n38300 ^ n37827 ;
  assign n38302 = n38301 ^ n37818 ;
  assign n38303 = ~n37824 & n38302 ;
  assign n38304 = n38303 ^ n37823 ;
  assign n37812 = n37035 ^ n36220 ;
  assign n37814 = n37813 ^ n37035 ;
  assign n37815 = n37812 & ~n37814 ;
  assign n37816 = n37815 ^ n36220 ;
  assign n37811 = n37753 ^ n37652 ;
  assign n37817 = n37816 ^ n37811 ;
  assign n38442 = n38304 ^ n37817 ;
  assign n38444 = n38442 ^ n35458 ;
  assign n38348 = n38301 ^ n37824 ;
  assign n38349 = n38348 ^ n34712 ;
  assign n38434 = n38298 ^ n37832 ;
  assign n38350 = n38295 ^ n37839 ;
  assign n38351 = n38350 ^ n34735 ;
  assign n38426 = n38292 ^ n37846 ;
  assign n38352 = n38289 ^ n37853 ;
  assign n38353 = n38352 ^ n34752 ;
  assign n38355 = n38277 ^ n37854 ;
  assign n38356 = n38355 ^ n34781 ;
  assign n38357 = n38274 ^ n37866 ;
  assign n38358 = n38357 ^ n35276 ;
  assign n38407 = n38272 ^ n37873 ;
  assign n38359 = n38268 ^ n38266 ;
  assign n38360 = n38359 ^ n35269 ;
  assign n38398 = n38262 ^ n38256 ;
  assign n38393 = n38247 ^ n38246 ;
  assign n38361 = n38237 ^ n38236 ;
  assign n38362 = n38361 ^ n34808 ;
  assign n38385 = n38227 ^ n37248 ;
  assign n38363 = n38220 ^ n38187 ;
  assign n38364 = n38363 ^ n34821 ;
  assign n38377 = n38185 ^ n38157 ;
  assign n38372 = n38181 ^ n38165 ;
  assign n38367 = n38179 ^ n38166 ;
  assign n38366 = ~n34839 & n38365 ;
  assign n38368 = n38367 ^ n38366 ;
  assign n38369 = n38367 ^ n35218 ;
  assign n38370 = ~n38368 & ~n38369 ;
  assign n38371 = n38370 ^ n35218 ;
  assign n38373 = n38372 ^ n38371 ;
  assign n38374 = n38372 ^ n34833 ;
  assign n38375 = n38373 & n38374 ;
  assign n38376 = n38375 ^ n34833 ;
  assign n38378 = n38377 ^ n38376 ;
  assign n38379 = n38377 ^ n34827 ;
  assign n38380 = n38378 & ~n38379 ;
  assign n38381 = n38380 ^ n34827 ;
  assign n38382 = n38381 ^ n38363 ;
  assign n38383 = ~n38364 & n38382 ;
  assign n38384 = n38383 ^ n34821 ;
  assign n38386 = n38385 ^ n38384 ;
  assign n38387 = n38385 ^ n34811 ;
  assign n38388 = n38386 & ~n38387 ;
  assign n38389 = n38388 ^ n34811 ;
  assign n38390 = n38389 ^ n38361 ;
  assign n38391 = n38362 & n38390 ;
  assign n38392 = n38391 ^ n34808 ;
  assign n38394 = n38393 ^ n38392 ;
  assign n38395 = n38392 ^ n34802 ;
  assign n38396 = n38394 & ~n38395 ;
  assign n38397 = n38396 ^ n38393 ;
  assign n38399 = n38398 ^ n38397 ;
  assign n38400 = n35269 ^ n35259 ;
  assign n38401 = n38400 ^ n35269 ;
  assign n38402 = n38401 ^ n38397 ;
  assign n38403 = n38399 & n38402 ;
  assign n38404 = n38403 ^ n38400 ;
  assign n38405 = ~n38360 & ~n38404 ;
  assign n38406 = n38405 ^ n38359 ;
  assign n38408 = n38407 ^ n38406 ;
  assign n38409 = n38407 ^ n34789 ;
  assign n38410 = n38408 & n38409 ;
  assign n38411 = n38410 ^ n34789 ;
  assign n38412 = n38411 ^ n38357 ;
  assign n38413 = ~n38358 & n38412 ;
  assign n38414 = n38413 ^ n35276 ;
  assign n38415 = n38414 ^ n38355 ;
  assign n38416 = ~n38356 & ~n38415 ;
  assign n38417 = n38416 ^ n34781 ;
  assign n38354 = n38287 ^ n38279 ;
  assign n38418 = n38417 ^ n38354 ;
  assign n38419 = n38352 ^ n34760 ;
  assign n38420 = n38419 ^ n38352 ;
  assign n38421 = n38420 ^ n38354 ;
  assign n38422 = ~n38418 & ~n38421 ;
  assign n38423 = n38422 ^ n38419 ;
  assign n38424 = ~n38353 & ~n38423 ;
  assign n38425 = n38424 ^ n34752 ;
  assign n38427 = n38426 ^ n38425 ;
  assign n38428 = n38425 ^ n34744 ;
  assign n38429 = ~n38427 & n38428 ;
  assign n38430 = n38429 ^ n38426 ;
  assign n38431 = n38430 ^ n38350 ;
  assign n38432 = ~n38351 & ~n38431 ;
  assign n38433 = n38432 ^ n34735 ;
  assign n38435 = n38434 ^ n38433 ;
  assign n38436 = n38434 ^ n35308 ;
  assign n38437 = n38435 & n38436 ;
  assign n38438 = n38437 ^ n35308 ;
  assign n38439 = n38438 ^ n38348 ;
  assign n38440 = n38349 & n38439 ;
  assign n38441 = n38440 ^ n34712 ;
  assign n38520 = n38444 ^ n38441 ;
  assign n38480 = n38436 ^ n38433 ;
  assign n38481 = n38430 ^ n38351 ;
  assign n38482 = n38423 ^ n34752 ;
  assign n38483 = n38371 ^ n34833 ;
  assign n38484 = n38483 ^ n38372 ;
  assign n38485 = n38379 ^ n38376 ;
  assign n38486 = n38484 & n38485 ;
  assign n38487 = n38381 ^ n34821 ;
  assign n38488 = n38487 ^ n38363 ;
  assign n38489 = n38486 & n38488 ;
  assign n38490 = n38387 ^ n38384 ;
  assign n38491 = ~n38489 & ~n38490 ;
  assign n38492 = n38389 ^ n34808 ;
  assign n38493 = n38492 ^ n38361 ;
  assign n38494 = ~n38491 & ~n38493 ;
  assign n38495 = n38395 ^ n38393 ;
  assign n38496 = n38494 & n38495 ;
  assign n38497 = n38397 ^ n35259 ;
  assign n38498 = n38497 ^ n38398 ;
  assign n38499 = ~n38496 & n38498 ;
  assign n38500 = n38404 ^ n38359 ;
  assign n38501 = n38499 & n38500 ;
  assign n38502 = n38406 ^ n34789 ;
  assign n38503 = n38502 ^ n38407 ;
  assign n38504 = ~n38501 & ~n38503 ;
  assign n38505 = n38411 ^ n38358 ;
  assign n38506 = n38504 & ~n38505 ;
  assign n38507 = n38414 ^ n38356 ;
  assign n38508 = n38506 & ~n38507 ;
  assign n38509 = n38354 ^ n34760 ;
  assign n38510 = n38509 ^ n38417 ;
  assign n38511 = n38508 & n38510 ;
  assign n38512 = n38482 & ~n38511 ;
  assign n38513 = n38426 ^ n34744 ;
  assign n38514 = n38513 ^ n38425 ;
  assign n38515 = ~n38512 & ~n38514 ;
  assign n38516 = ~n38481 & n38515 ;
  assign n38517 = ~n38480 & n38516 ;
  assign n38518 = n38438 ^ n38349 ;
  assign n38519 = ~n38517 & ~n38518 ;
  assign n38562 = n38520 ^ n38519 ;
  assign n38563 = n38562 ^ n1653 ;
  assign n38567 = n38518 ^ n38517 ;
  assign n38568 = n38567 ^ n38566 ;
  assign n38572 = n38516 ^ n38480 ;
  assign n38573 = n38572 ^ n38571 ;
  assign n38574 = n38515 ^ n38481 ;
  assign n2970 = n2969 ^ n2966 ;
  assign n2971 = n2970 ^ n638 ;
  assign n2975 = n2974 ^ n2971 ;
  assign n38575 = n38574 ^ n2975 ;
  assign n38579 = n38514 ^ n38512 ;
  assign n38580 = n38579 ^ n38578 ;
  assign n38584 = n38511 ^ n38482 ;
  assign n38581 = n36342 ^ n608 ;
  assign n38582 = n38581 ^ n32003 ;
  assign n38583 = n38582 ^ n26525 ;
  assign n38585 = n38584 ^ n38583 ;
  assign n38587 = n36347 ^ n27794 ;
  assign n38588 = n38587 ^ n32008 ;
  assign n38589 = n38588 ^ n1499 ;
  assign n38685 = n38589 ^ n38584 ;
  assign n38586 = n38510 ^ n38508 ;
  assign n38590 = n38589 ^ n38586 ;
  assign n38594 = n38507 ^ n38506 ;
  assign n38591 = n36351 ^ n27799 ;
  assign n38592 = n38591 ^ n32014 ;
  assign n38593 = n38592 ^ n26517 ;
  assign n38595 = n38594 ^ n38593 ;
  assign n38597 = n36357 ^ n27803 ;
  assign n38598 = n38597 ^ n32019 ;
  assign n38599 = n38598 ^ n26472 ;
  assign n38679 = n38599 ^ n38594 ;
  assign n38596 = n38505 ^ n38504 ;
  assign n38600 = n38599 ^ n38596 ;
  assign n38602 = n36362 ^ n2439 ;
  assign n38603 = n38602 ^ n32024 ;
  assign n38604 = n38603 ^ n26481 ;
  assign n38601 = n38503 ^ n38501 ;
  assign n38605 = n38604 ^ n38601 ;
  assign n38610 = n38500 ^ n38499 ;
  assign n38606 = n32029 ^ n2421 ;
  assign n38607 = n38606 ^ n36367 ;
  assign n38608 = n38607 ^ n26486 ;
  assign n38611 = n38610 ^ n38608 ;
  assign n38615 = n38498 ^ n38496 ;
  assign n38612 = n36372 ^ n2411 ;
  assign n38613 = n38612 ^ n32033 ;
  assign n38614 = n38613 ^ n2216 ;
  assign n38616 = n38615 ^ n38614 ;
  assign n38618 = n36402 ^ n27436 ;
  assign n38619 = n38618 ^ n2096 ;
  assign n38620 = n38619 ^ n26497 ;
  assign n38668 = n38620 ^ n38615 ;
  assign n38617 = n38495 ^ n38494 ;
  assign n38621 = n38620 ^ n38617 ;
  assign n38625 = n38493 ^ n38491 ;
  assign n38622 = n36377 ^ n27469 ;
  assign n38623 = n38622 ^ n32040 ;
  assign n38624 = n38623 ^ n2091 ;
  assign n38626 = n38625 ^ n38624 ;
  assign n38627 = n38490 ^ n38489 ;
  assign n1989 = n1988 ^ n1970 ;
  assign n2008 = n2007 ^ n1989 ;
  assign n2015 = n2014 ^ n2008 ;
  assign n38628 = n38627 ^ n2015 ;
  assign n38630 = n36384 ^ n27448 ;
  assign n38631 = n38630 ^ n32048 ;
  assign n38632 = n38631 ^ n2002 ;
  assign n38629 = n38488 ^ n38486 ;
  assign n38633 = n38632 ^ n38629 ;
  assign n38637 = n38485 ^ n38484 ;
  assign n38634 = n35785 ^ n1923 ;
  assign n38635 = n38634 ^ n32052 ;
  assign n38636 = n38635 ^ n26112 ;
  assign n38638 = n38637 ^ n38636 ;
  assign n3033 = n3032 ^ n3023 ;
  assign n3046 = n3045 ^ n3033 ;
  assign n3053 = n3052 ^ n3046 ;
  assign n38639 = n38484 ^ n3053 ;
  assign n38642 = n3240 ^ n3230 ;
  assign n38643 = n38642 ^ n3040 ;
  assign n38644 = n38643 ^ n2782 ;
  assign n38641 = n2775 & ~n38640 ;
  assign n38645 = n38644 ^ n38641 ;
  assign n38646 = n38366 ^ n35218 ;
  assign n38647 = n38646 ^ n38367 ;
  assign n38648 = n38647 ^ n38644 ;
  assign n38649 = ~n38645 & ~n38648 ;
  assign n38650 = n38649 ^ n38647 ;
  assign n38651 = n38650 ^ n3053 ;
  assign n38652 = n38639 & n38651 ;
  assign n38653 = n38652 ^ n38484 ;
  assign n38654 = n38653 ^ n38636 ;
  assign n38655 = ~n38638 & ~n38654 ;
  assign n38656 = n38655 ^ n38637 ;
  assign n38657 = n38656 ^ n38629 ;
  assign n38658 = ~n38633 & ~n38657 ;
  assign n38659 = n38658 ^ n38632 ;
  assign n38660 = n38659 ^ n2015 ;
  assign n38661 = n38628 & ~n38660 ;
  assign n38662 = n38661 ^ n38627 ;
  assign n38663 = n38662 ^ n38624 ;
  assign n38664 = ~n38626 & ~n38663 ;
  assign n38665 = n38664 ^ n38625 ;
  assign n38666 = n38665 ^ n38620 ;
  assign n38667 = ~n38621 & ~n38666 ;
  assign n38669 = n38668 ^ n38667 ;
  assign n38670 = ~n38616 & ~n38669 ;
  assign n38671 = n38670 ^ n38615 ;
  assign n38672 = n38671 ^ n38608 ;
  assign n38673 = n38611 & ~n38672 ;
  assign n38609 = n38608 ^ n38601 ;
  assign n38674 = n38673 ^ n38609 ;
  assign n38675 = ~n38605 & n38674 ;
  assign n38676 = n38675 ^ n38604 ;
  assign n38677 = n38676 ^ n38599 ;
  assign n38678 = n38600 & n38677 ;
  assign n38680 = n38679 ^ n38678 ;
  assign n38681 = n38595 & n38680 ;
  assign n38682 = n38681 ^ n38594 ;
  assign n38683 = n38682 ^ n38589 ;
  assign n38684 = ~n38590 & n38683 ;
  assign n38686 = n38685 ^ n38684 ;
  assign n38687 = ~n38585 & ~n38686 ;
  assign n38688 = n38687 ^ n38584 ;
  assign n38689 = n38688 ^ n38578 ;
  assign n38690 = ~n38580 & n38689 ;
  assign n38691 = n38690 ^ n38579 ;
  assign n38692 = n38691 ^ n2975 ;
  assign n38693 = n38575 & n38692 ;
  assign n38694 = n38693 ^ n38574 ;
  assign n38695 = n38694 ^ n38571 ;
  assign n38696 = n38573 & ~n38695 ;
  assign n38697 = n38696 ^ n38572 ;
  assign n38698 = n38697 ^ n38566 ;
  assign n38699 = n38568 & ~n38698 ;
  assign n38700 = n38699 ^ n38567 ;
  assign n38701 = n38700 ^ n1653 ;
  assign n38702 = n38563 & ~n38701 ;
  assign n38703 = n38702 ^ n38562 ;
  assign n38521 = ~n38519 & n38520 ;
  assign n38443 = n38442 ^ n38441 ;
  assign n38445 = ~n38443 & ~n38444 ;
  assign n38446 = n38445 ^ n35458 ;
  assign n38305 = n38304 ^ n37811 ;
  assign n38306 = ~n37817 & ~n38305 ;
  assign n38307 = n38306 ^ n37816 ;
  assign n37797 = n37796 ^ n37232 ;
  assign n37798 = n37755 ^ n37649 ;
  assign n37799 = n37798 ^ n36479 ;
  assign n37800 = n37799 ^ n37796 ;
  assign n37801 = n37800 ^ n37798 ;
  assign n37802 = n37797 & ~n37801 ;
  assign n37803 = n37802 ^ n37799 ;
  assign n38346 = n38307 ^ n37803 ;
  assign n38347 = n38346 ^ n35717 ;
  assign n38479 = n38446 ^ n38347 ;
  assign n38560 = n38521 ^ n38479 ;
  assign n38561 = n38560 ^ n38559 ;
  assign n39416 = n38703 ^ n38561 ;
  assign n39514 = n39416 ^ n36485 ;
  assign n39515 = n39514 ^ n38951 ;
  assign n39516 = n39515 ^ n39416 ;
  assign n39517 = n39513 & ~n39516 ;
  assign n39518 = n39517 ^ n39514 ;
  assign n39492 = n38195 ^ n37253 ;
  assign n38817 = n38120 ^ n38089 ;
  assign n39493 = n38817 ^ n38195 ;
  assign n39494 = n39492 & ~n39493 ;
  assign n39495 = n39494 ^ n37253 ;
  assign n39424 = n38700 ^ n38563 ;
  assign n39496 = n39495 ^ n39424 ;
  assign n39431 = n38697 ^ n38568 ;
  assign n39508 = n39495 ^ n39431 ;
  assign n38777 = n38117 ^ n38091 ;
  assign n39497 = n38777 ^ n38147 ;
  assign n39498 = n39431 ^ n37255 ;
  assign n39499 = n39498 ^ n38777 ;
  assign n39500 = n39499 ^ n39431 ;
  assign n39501 = n39497 & n39500 ;
  assign n39502 = n39501 ^ n39498 ;
  assign n39357 = n37329 ^ n37252 ;
  assign n38735 = n38114 ^ n38093 ;
  assign n39358 = n38735 ^ n37252 ;
  assign n39359 = n39357 & n39358 ;
  assign n39360 = n39359 ^ n37329 ;
  assign n39356 = n38694 ^ n38573 ;
  assign n39361 = n39360 ^ n39356 ;
  assign n39068 = n37316 ^ n37257 ;
  assign n38476 = n38111 ^ n38095 ;
  assign n39069 = n38476 ^ n37257 ;
  assign n39070 = n39068 & n39069 ;
  assign n39071 = n39070 ^ n37316 ;
  assign n39067 = n38691 ^ n38575 ;
  assign n39072 = n39071 ^ n39067 ;
  assign n38851 = n38688 ^ n38580 ;
  assign n38847 = n37791 ^ n37232 ;
  assign n38336 = n38108 ^ n38100 ;
  assign n38848 = n38336 ^ n37791 ;
  assign n38849 = n38847 & n38848 ;
  assign n38850 = n38849 ^ n37232 ;
  assign n38852 = n38851 ^ n38850 ;
  assign n38857 = n38686 ^ n38583 ;
  assign n38853 = n37805 ^ n37035 ;
  assign n38331 = n38105 ^ n38102 ;
  assign n38854 = n38331 ^ n37805 ;
  assign n38855 = n38853 & ~n38854 ;
  assign n38856 = n38855 ^ n37035 ;
  assign n38858 = n38857 ^ n38856 ;
  assign n37786 = n37785 ^ n37764 ;
  assign n38859 = n37796 ^ n37786 ;
  assign n38860 = n38682 ^ n38590 ;
  assign n38861 = n38860 ^ n37015 ;
  assign n38862 = n38861 ^ n37786 ;
  assign n38863 = n38862 ^ n38860 ;
  assign n38864 = n38859 & n38863 ;
  assign n38865 = n38864 ^ n38861 ;
  assign n38870 = n38680 ^ n38593 ;
  assign n38866 = n37813 ^ n37006 ;
  assign n37788 = n37761 ^ n37639 ;
  assign n38867 = n37813 ^ n37788 ;
  assign n38868 = n38866 & ~n38867 ;
  assign n38869 = n38868 ^ n37006 ;
  assign n38871 = n38870 ^ n38869 ;
  assign n38876 = n38676 ^ n38600 ;
  assign n38312 = n37759 ^ n37643 ;
  assign n38872 = n38312 ^ n37820 ;
  assign n38873 = n37820 ^ n36977 ;
  assign n38874 = ~n38872 & n38873 ;
  assign n38875 = n38874 ^ n36977 ;
  assign n38877 = n38876 ^ n38875 ;
  assign n38884 = n38671 ^ n38611 ;
  assign n38880 = n37835 ^ n36951 ;
  assign n38881 = n37835 ^ n37811 ;
  assign n38882 = n38880 & n38881 ;
  assign n38883 = n38882 ^ n36951 ;
  assign n38885 = n38884 ^ n38883 ;
  assign n38890 = n38669 ^ n38614 ;
  assign n38886 = n37842 ^ n36894 ;
  assign n38887 = n37842 ^ n37818 ;
  assign n38888 = ~n38886 & ~n38887 ;
  assign n38889 = n38888 ^ n36894 ;
  assign n38891 = n38890 ^ n38889 ;
  assign n38896 = n38665 ^ n38621 ;
  assign n38892 = n37849 ^ n37827 ;
  assign n38893 = n37849 ^ n36794 ;
  assign n38894 = n38892 & n38893 ;
  assign n38895 = n38894 ^ n36794 ;
  assign n38897 = n38896 ^ n38895 ;
  assign n38902 = n38662 ^ n38626 ;
  assign n38898 = n37833 ^ n37775 ;
  assign n38899 = n37775 ^ n36590 ;
  assign n38900 = ~n38898 & ~n38899 ;
  assign n38901 = n38900 ^ n36590 ;
  assign n38903 = n38902 ^ n38901 ;
  assign n38908 = n38659 ^ n38628 ;
  assign n38904 = n37840 ^ n37262 ;
  assign n38905 = n37262 ^ n36782 ;
  assign n38906 = ~n38904 & n38905 ;
  assign n38907 = n38906 ^ n36782 ;
  assign n38909 = n38908 ^ n38907 ;
  assign n38910 = n37508 ^ n36597 ;
  assign n38911 = n37847 ^ n37508 ;
  assign n38912 = ~n38910 & n38911 ;
  assign n38913 = n38912 ^ n36597 ;
  assign n38841 = n38656 ^ n38633 ;
  assign n38914 = n38913 ^ n38841 ;
  assign n38916 = n38280 ^ n37499 ;
  assign n38917 = n37499 ^ n36606 ;
  assign n38918 = n38916 & ~n38917 ;
  assign n38919 = n38918 ^ n36606 ;
  assign n38915 = n38653 ^ n38638 ;
  assign n38920 = n38919 ^ n38915 ;
  assign n38921 = n37854 ^ n37272 ;
  assign n38922 = n38650 ^ n38639 ;
  assign n38923 = n38922 ^ n36600 ;
  assign n38924 = n38923 ^ n37854 ;
  assign n38925 = n38924 ^ n38922 ;
  assign n38926 = ~n38921 & n38925 ;
  assign n38927 = n38926 ^ n38923 ;
  assign n39020 = n38922 ^ n38919 ;
  assign n38932 = n38647 ^ n38645 ;
  assign n38928 = n37861 ^ n37278 ;
  assign n38929 = n37278 ^ n36611 ;
  assign n38930 = ~n38928 & n38929 ;
  assign n38931 = n38930 ^ n36611 ;
  assign n38933 = n38932 ^ n38931 ;
  assign n39015 = n38935 ^ n38931 ;
  assign n38934 = n37873 ^ n37280 ;
  assign n38936 = n38935 ^ n36614 ;
  assign n38937 = n38936 ^ n37873 ;
  assign n38938 = n38937 ^ n38935 ;
  assign n38939 = n38934 & n38938 ;
  assign n38940 = n38939 ^ n38936 ;
  assign n38823 = n37429 ^ n36697 ;
  assign n38824 = n36697 ^ n35965 ;
  assign n38825 = n38823 & n38824 ;
  assign n38826 = n38825 ^ n35965 ;
  assign n37254 = n37253 ^ n37252 ;
  assign n37256 = n37255 ^ n36650 ;
  assign n37258 = n37257 ^ n37255 ;
  assign n37259 = n37256 & n37258 ;
  assign n37260 = n37259 ^ n36650 ;
  assign n37787 = n37786 ^ n37260 ;
  assign n37790 = n37329 ^ n36561 ;
  assign n37792 = n37791 ^ n37329 ;
  assign n37793 = ~n37790 & ~n37792 ;
  assign n37794 = n37793 ^ n36561 ;
  assign n37795 = n37794 ^ n37788 ;
  assign n37804 = n37316 ^ n36513 ;
  assign n37806 = n37805 ^ n37316 ;
  assign n37807 = n37804 & n37806 ;
  assign n37808 = n37807 ^ n36513 ;
  assign n37809 = n37808 ^ n37798 ;
  assign n37810 = n37809 ^ n37808 ;
  assign n38308 = n38307 ^ n37810 ;
  assign n38309 = n37803 & n38308 ;
  assign n38310 = n38309 ^ n37809 ;
  assign n38313 = n38312 ^ n37788 ;
  assign n38311 = n37808 ^ n37788 ;
  assign n38314 = n38313 ^ n38311 ;
  assign n38315 = ~n38310 & n38314 ;
  assign n38316 = n38315 ^ n38311 ;
  assign n38317 = ~n37795 & ~n38316 ;
  assign n37789 = n37788 ^ n37260 ;
  assign n38318 = n38317 ^ n37789 ;
  assign n38319 = n37787 & ~n38318 ;
  assign n38320 = n38319 ^ n37786 ;
  assign n38321 = n38320 ^ n36676 ;
  assign n38322 = n38321 ^ n37252 ;
  assign n38323 = n38322 ^ n38320 ;
  assign n38324 = n37254 & n38323 ;
  assign n38325 = n38324 ^ n38321 ;
  assign n38326 = n36485 ^ n35732 ;
  assign n38327 = n38147 ^ n36485 ;
  assign n38328 = ~n38326 & n38327 ;
  assign n38329 = n38328 ^ n35732 ;
  assign n38332 = n38331 ^ n38329 ;
  assign n38330 = n38329 ^ n38320 ;
  assign n38333 = n38332 ^ n38330 ;
  assign n38334 = ~n38325 & n38333 ;
  assign n38335 = n38334 ^ n38332 ;
  assign n38467 = n36525 ^ n35775 ;
  assign n38468 = n38195 ^ n36525 ;
  assign n38469 = ~n38467 & ~n38468 ;
  assign n38470 = n38469 ^ n35775 ;
  assign n38472 = n38470 ^ n38329 ;
  assign n38471 = n38470 ^ n38336 ;
  assign n38473 = n38472 ^ n38471 ;
  assign n38474 = ~n38335 & n38473 ;
  assign n38475 = n38474 ^ n38472 ;
  assign n38726 = n36566 ^ n35812 ;
  assign n38727 = n37242 ^ n36566 ;
  assign n38728 = ~n38726 & n38727 ;
  assign n38729 = n38728 ^ n35812 ;
  assign n38731 = n38729 ^ n38470 ;
  assign n38730 = n38729 ^ n38476 ;
  assign n38732 = n38731 ^ n38730 ;
  assign n38733 = ~n38475 & n38732 ;
  assign n38734 = n38733 ^ n38731 ;
  assign n38768 = n36699 ^ n35977 ;
  assign n38769 = n37418 ^ n36699 ;
  assign n38770 = ~n38768 & ~n38769 ;
  assign n38771 = n38770 ^ n35977 ;
  assign n38773 = n38771 ^ n38729 ;
  assign n38772 = n38771 ^ n38735 ;
  assign n38774 = n38773 ^ n38772 ;
  assign n38775 = n38734 & ~n38774 ;
  assign n38776 = n38775 ^ n38773 ;
  assign n38819 = n38817 ^ n38771 ;
  assign n38818 = n38817 ^ n38777 ;
  assign n38820 = n38819 ^ n38818 ;
  assign n38821 = n38776 & n38820 ;
  assign n38822 = n38821 ^ n38819 ;
  assign n38827 = n38826 ^ n38822 ;
  assign n38477 = n38476 ^ n38475 ;
  assign n38737 = n38477 ^ n35155 ;
  assign n38337 = n38336 ^ n38335 ;
  assign n38338 = n38337 ^ n35149 ;
  assign n38339 = n38331 ^ n38325 ;
  assign n38340 = n38339 ^ n35952 ;
  assign n38341 = n38318 ^ n37786 ;
  assign n38342 = n38341 ^ n35924 ;
  assign n38343 = n38316 ^ n37794 ;
  assign n38344 = n38343 ^ n35807 ;
  assign n38447 = n38446 ^ n38346 ;
  assign n38448 = n38347 & n38447 ;
  assign n38449 = n38448 ^ n35717 ;
  assign n38345 = n38312 ^ n38310 ;
  assign n38450 = n38449 ^ n38345 ;
  assign n38451 = n38345 ^ n35757 ;
  assign n38452 = n38450 & n38451 ;
  assign n38453 = n38452 ^ n38449 ;
  assign n38454 = n38453 ^ n38343 ;
  assign n38455 = ~n38344 & ~n38454 ;
  assign n38456 = n38455 ^ n35807 ;
  assign n38457 = n38456 ^ n38341 ;
  assign n38458 = n38342 & n38457 ;
  assign n38459 = n38458 ^ n35924 ;
  assign n38460 = n38459 ^ n38339 ;
  assign n38461 = n38340 & ~n38460 ;
  assign n38462 = n38461 ^ n35952 ;
  assign n38463 = n38462 ^ n38337 ;
  assign n38464 = ~n38338 & ~n38463 ;
  assign n38465 = n38464 ^ n35149 ;
  assign n38738 = n38477 ^ n38465 ;
  assign n38739 = ~n38737 & ~n38738 ;
  assign n38740 = n38739 ^ n35155 ;
  assign n38741 = n38740 ^ n35143 ;
  assign n38736 = n38735 ^ n38734 ;
  assign n38764 = n38740 ^ n38736 ;
  assign n38765 = n38741 & n38764 ;
  assign n38766 = n38765 ^ n35143 ;
  assign n38767 = n38766 ^ n35141 ;
  assign n38778 = n38777 ^ n38776 ;
  assign n38813 = n38778 ^ n38766 ;
  assign n38814 = n38767 & ~n38813 ;
  assign n38815 = n38814 ^ n35141 ;
  assign n38816 = n38815 ^ n35204 ;
  assign n38828 = n38827 ^ n38816 ;
  assign n38779 = n38778 ^ n38767 ;
  assign n38466 = n38465 ^ n35155 ;
  assign n38478 = n38477 ^ n38466 ;
  assign n38522 = n38479 & n38521 ;
  assign n38523 = n38451 ^ n38449 ;
  assign n38524 = ~n38522 & ~n38523 ;
  assign n38525 = n38453 ^ n35807 ;
  assign n38526 = n38525 ^ n38343 ;
  assign n38527 = n38524 & ~n38526 ;
  assign n38528 = n38456 ^ n35924 ;
  assign n38529 = n38528 ^ n38341 ;
  assign n38530 = n38527 & ~n38529 ;
  assign n38531 = n38459 ^ n38340 ;
  assign n38532 = ~n38530 & ~n38531 ;
  assign n38533 = n38462 ^ n35149 ;
  assign n38534 = n38533 ^ n38337 ;
  assign n38535 = n38532 & n38534 ;
  assign n38725 = ~n38478 & n38535 ;
  assign n38742 = n38741 ^ n38736 ;
  assign n38780 = n38725 & n38742 ;
  assign n38829 = n38779 & ~n38780 ;
  assign n38950 = ~n38828 & n38829 ;
  assign n38962 = n38827 ^ n38815 ;
  assign n38963 = ~n38816 & ~n38962 ;
  assign n38964 = n38963 ^ n35204 ;
  assign n38965 = n38964 ^ n34055 ;
  assign n38957 = n36580 ^ n35830 ;
  assign n38958 = n37411 ^ n36580 ;
  assign n38959 = n38957 & n38958 ;
  assign n38960 = n38959 ^ n35830 ;
  assign n38953 = n38951 ^ n38817 ;
  assign n38952 = n38951 ^ n38826 ;
  assign n38954 = n38953 ^ n38952 ;
  assign n38955 = ~n38822 & n38954 ;
  assign n38956 = n38955 ^ n38953 ;
  assign n38961 = n38960 ^ n38956 ;
  assign n38966 = n38965 ^ n38961 ;
  assign n39001 = n38950 & ~n38966 ;
  assign n38996 = n38960 ^ n38951 ;
  assign n38997 = n38956 & ~n38996 ;
  assign n38991 = n36683 ^ n2683 ;
  assign n38992 = n38991 ^ n2772 ;
  assign n38993 = n38992 ^ n32501 ;
  assign n38947 = n36545 ^ n2671 ;
  assign n38948 = n38947 ^ n26755 ;
  assign n38949 = n38948 ^ n3143 ;
  assign n38994 = n38993 ^ n38949 ;
  assign n38989 = n34845 ^ n34055 ;
  assign n38987 = n38951 ^ n36001 ;
  assign n38986 = n38126 ^ n38079 ;
  assign n38988 = n38987 ^ n38986 ;
  assign n38990 = n38989 ^ n38988 ;
  assign n38995 = n38994 ^ n38990 ;
  assign n38998 = n38997 ^ n38995 ;
  assign n38984 = n38964 ^ n38961 ;
  assign n38985 = ~n38965 & n38984 ;
  assign n38999 = n38998 ^ n38985 ;
  assign n38981 = n36723 ^ n36001 ;
  assign n38982 = n37406 ^ n36723 ;
  assign n38983 = ~n38981 & n38982 ;
  assign n39000 = n38999 ^ n38983 ;
  assign n39002 = n39001 ^ n39000 ;
  assign n38967 = n38966 ^ n38950 ;
  assign n38968 = n38967 ^ n38949 ;
  assign n38830 = n38829 ^ n38828 ;
  assign n38810 = n36502 ^ n27927 ;
  assign n38811 = n38810 ^ n32512 ;
  assign n38812 = n38811 ^ n3138 ;
  assign n38831 = n38830 ^ n38812 ;
  assign n38781 = n38780 ^ n38779 ;
  assign n38761 = n36292 ^ n3122 ;
  assign n38762 = n38761 ^ n26581 ;
  assign n38763 = n38762 ^ n32518 ;
  assign n38782 = n38781 ^ n38763 ;
  assign n38744 = n36288 ^ n27522 ;
  assign n38745 = n38744 ^ n32523 ;
  assign n38746 = n38745 ^ n26443 ;
  assign n38743 = n38742 ^ n38725 ;
  assign n38747 = n38746 ^ n38743 ;
  assign n38537 = n36298 ^ n27867 ;
  assign n38538 = n38537 ^ n32527 ;
  assign n38539 = n38538 ^ n2645 ;
  assign n38536 = n38535 ^ n38478 ;
  assign n38540 = n38539 ^ n38536 ;
  assign n38542 = n27861 ^ n1388 ;
  assign n38543 = n38542 ^ n32533 ;
  assign n38544 = n38543 ^ n26450 ;
  assign n38541 = n38534 ^ n38532 ;
  assign n38545 = n38544 ^ n38541 ;
  assign n38546 = n36304 ^ n27856 ;
  assign n38547 = n38546 ^ n1285 ;
  assign n38548 = n38547 ^ n2789 ;
  assign n38718 = n38548 ^ n38541 ;
  assign n38549 = n38531 ^ n38530 ;
  assign n38550 = n38549 ^ n38548 ;
  assign n38551 = n38529 ^ n38527 ;
  assign n38552 = n38551 ^ n1278 ;
  assign n38553 = n38526 ^ n38524 ;
  assign n1127 = n1090 ^ n1048 ;
  assign n1128 = n1127 ^ n1124 ;
  assign n1135 = n1134 ^ n1128 ;
  assign n38554 = n38553 ^ n1135 ;
  assign n38555 = n38523 ^ n38522 ;
  assign n1094 = n1078 ^ n1030 ;
  assign n1104 = n1103 ^ n1094 ;
  assign n1117 = n1116 ^ n1104 ;
  assign n38556 = n38555 ^ n1117 ;
  assign n38704 = n38703 ^ n38559 ;
  assign n38705 = ~n38561 & ~n38704 ;
  assign n38706 = n38705 ^ n38560 ;
  assign n38707 = n38706 ^ n1117 ;
  assign n38708 = n38556 & n38707 ;
  assign n38709 = n38708 ^ n38555 ;
  assign n38710 = n38709 ^ n1135 ;
  assign n38711 = ~n38554 & ~n38710 ;
  assign n38712 = n38711 ^ n38553 ;
  assign n38713 = n38712 ^ n1278 ;
  assign n38714 = ~n38552 & n38713 ;
  assign n38715 = n38714 ^ n38551 ;
  assign n38716 = n38715 ^ n38548 ;
  assign n38717 = ~n38550 & ~n38716 ;
  assign n38719 = n38718 ^ n38717 ;
  assign n38720 = ~n38545 & n38719 ;
  assign n38721 = n38720 ^ n38544 ;
  assign n38722 = n38721 ^ n38536 ;
  assign n38723 = n38540 & ~n38722 ;
  assign n38724 = n38723 ^ n38539 ;
  assign n38758 = n38743 ^ n38724 ;
  assign n38759 = ~n38747 & n38758 ;
  assign n38760 = n38759 ^ n38746 ;
  assign n38807 = n38763 ^ n38760 ;
  assign n38808 = ~n38782 & ~n38807 ;
  assign n38809 = n38808 ^ n38781 ;
  assign n38944 = n38812 ^ n38809 ;
  assign n38945 = ~n38831 & n38944 ;
  assign n38946 = n38945 ^ n38830 ;
  assign n38979 = n38949 ^ n38946 ;
  assign n38980 = ~n38968 & ~n38979 ;
  assign n39003 = n39002 ^ n38980 ;
  assign n38969 = n38968 ^ n38946 ;
  assign n36579 = n36578 ^ n35825 ;
  assign n37249 = n37248 ^ n35825 ;
  assign n37250 = n36579 & n37249 ;
  assign n37251 = n37250 ^ n36578 ;
  assign n38748 = n38747 ^ n38724 ;
  assign n38788 = ~n37251 & ~n38748 ;
  assign n38784 = n37297 ^ n36633 ;
  assign n38785 = n38237 ^ n37297 ;
  assign n38786 = n38784 & n38785 ;
  assign n38787 = n38786 ^ n36633 ;
  assign n38789 = n38788 ^ n38787 ;
  assign n38798 = n37469 ^ n36626 ;
  assign n38799 = n38247 ^ n36626 ;
  assign n38800 = n38798 & n38799 ;
  assign n38801 = n38800 ^ n37469 ;
  assign n38783 = n38782 ^ n38760 ;
  assign n38802 = n38801 ^ n38783 ;
  assign n38803 = n38802 ^ n38801 ;
  assign n38804 = n38803 ^ n38787 ;
  assign n38805 = ~n38789 & ~n38804 ;
  assign n38806 = n38805 ^ n38802 ;
  assign n38832 = n38831 ^ n38809 ;
  assign n38941 = n38832 ^ n38801 ;
  assign n38942 = ~n38806 & ~n38941 ;
  assign n38943 = n38942 ^ n38832 ;
  assign n38970 = n38969 ^ n38943 ;
  assign n38971 = n38262 ^ n37296 ;
  assign n38972 = n38943 ^ n36741 ;
  assign n38973 = n38972 ^ n38262 ;
  assign n38974 = n38973 ^ n38943 ;
  assign n38975 = n38971 & n38974 ;
  assign n38976 = n38975 ^ n38972 ;
  assign n38977 = n38970 & ~n38976 ;
  assign n38978 = n38977 ^ n38969 ;
  assign n39004 = n39003 ^ n38978 ;
  assign n39005 = n38268 ^ n36624 ;
  assign n39006 = n39003 ^ n37288 ;
  assign n39007 = n39006 ^ n38268 ;
  assign n39008 = n39007 ^ n39003 ;
  assign n39009 = n39005 & n39008 ;
  assign n39010 = n39009 ^ n39006 ;
  assign n39011 = ~n39004 & ~n39010 ;
  assign n39012 = n39011 ^ n39003 ;
  assign n39013 = n39012 ^ n38935 ;
  assign n39014 = n38940 & n39013 ;
  assign n39016 = n39015 ^ n39014 ;
  assign n39017 = ~n38933 & n39016 ;
  assign n39018 = n39017 ^ n38932 ;
  assign n39019 = n39018 ^ n38919 ;
  assign n39021 = n39020 ^ n39019 ;
  assign n39022 = n38927 & n39021 ;
  assign n39023 = n39022 ^ n39020 ;
  assign n39024 = n38920 & n39023 ;
  assign n39025 = n39024 ^ n38919 ;
  assign n39026 = n39025 ^ n38841 ;
  assign n39027 = ~n38914 & ~n39026 ;
  assign n39028 = n39027 ^ n38841 ;
  assign n39029 = n39028 ^ n38907 ;
  assign n39030 = n38909 & ~n39029 ;
  assign n39031 = n39030 ^ n38908 ;
  assign n39032 = n39031 ^ n38901 ;
  assign n39033 = n38903 & n39032 ;
  assign n39034 = n39033 ^ n38902 ;
  assign n39035 = n39034 ^ n38895 ;
  assign n39036 = n38897 & n39035 ;
  assign n39037 = n39036 ^ n38896 ;
  assign n39038 = n39037 ^ n38889 ;
  assign n39039 = n38891 & n39038 ;
  assign n39040 = n39039 ^ n38890 ;
  assign n39041 = n39040 ^ n38883 ;
  assign n39042 = ~n38885 & n39041 ;
  assign n39043 = n39042 ^ n38884 ;
  assign n38878 = n38674 ^ n38604 ;
  assign n39044 = n39043 ^ n38878 ;
  assign n39045 = n37825 ^ n37798 ;
  assign n39046 = n38878 ^ n36964 ;
  assign n39047 = n39046 ^ n37798 ;
  assign n39048 = n39047 ^ n38878 ;
  assign n39049 = n39045 & n39048 ;
  assign n39050 = n39049 ^ n39046 ;
  assign n39051 = n39044 & ~n39050 ;
  assign n38879 = n38878 ^ n38875 ;
  assign n39052 = n39051 ^ n38879 ;
  assign n39053 = ~n38877 & ~n39052 ;
  assign n39054 = n39053 ^ n38876 ;
  assign n39055 = n39054 ^ n38869 ;
  assign n39056 = n38871 & ~n39055 ;
  assign n39057 = n39056 ^ n38870 ;
  assign n39058 = n39057 ^ n38860 ;
  assign n39059 = ~n38865 & ~n39058 ;
  assign n39060 = n39059 ^ n38860 ;
  assign n39061 = n39060 ^ n38856 ;
  assign n39062 = ~n38858 & n39061 ;
  assign n39063 = n39062 ^ n38857 ;
  assign n39064 = n39063 ^ n38850 ;
  assign n39065 = n38852 & n39064 ;
  assign n39066 = n39065 ^ n38851 ;
  assign n39353 = n39067 ^ n39066 ;
  assign n39354 = n39072 & n39353 ;
  assign n39355 = n39354 ^ n39071 ;
  assign n39503 = n39356 ^ n39355 ;
  assign n39504 = n39361 & n39503 ;
  assign n39505 = n39504 ^ n39360 ;
  assign n39506 = n39505 ^ n39431 ;
  assign n39507 = n39502 & n39506 ;
  assign n39509 = n39508 ^ n39507 ;
  assign n39510 = ~n39496 & n39509 ;
  assign n39511 = n39510 ^ n39424 ;
  assign n39559 = n39518 ^ n39511 ;
  assign n39546 = n39509 ^ n39424 ;
  assign n39547 = n39546 ^ n36676 ;
  assign n39551 = n39505 ^ n39502 ;
  assign n39362 = n39361 ^ n39355 ;
  assign n39363 = n39362 ^ n36561 ;
  assign n39073 = n39072 ^ n39066 ;
  assign n39074 = n39073 ^ n36513 ;
  assign n39075 = n39063 ^ n38852 ;
  assign n39076 = n39075 ^ n36479 ;
  assign n39077 = n39060 ^ n38858 ;
  assign n39078 = n39077 ^ n36220 ;
  assign n39158 = n39057 ^ n38865 ;
  assign n39079 = n39054 ^ n38871 ;
  assign n39080 = n39079 ^ n35838 ;
  assign n39081 = n39052 ^ n38876 ;
  assign n39082 = n39081 ^ n36080 ;
  assign n39084 = n39040 ^ n38885 ;
  assign n39085 = n39084 ^ n35846 ;
  assign n39140 = n39037 ^ n38891 ;
  assign n39086 = n39034 ^ n38897 ;
  assign n39087 = n39086 ^ n36061 ;
  assign n39088 = n39031 ^ n38903 ;
  assign n39089 = n39088 ^ n36057 ;
  assign n39090 = n39028 ^ n38909 ;
  assign n39091 = n39090 ^ n36043 ;
  assign n39092 = n39025 ^ n38914 ;
  assign n39093 = n39092 ^ n35858 ;
  assign n39095 = n39018 ^ n38927 ;
  assign n39096 = n39095 ^ n35874 ;
  assign n39116 = n39016 ^ n38932 ;
  assign n39097 = n39012 ^ n38940 ;
  assign n39098 = n39097 ^ n35883 ;
  assign n39108 = n39010 ^ n38978 ;
  assign n39099 = n38976 ^ n38969 ;
  assign n39100 = n39099 ^ n35896 ;
  assign n38749 = n38748 ^ n37251 ;
  assign n38756 = n36012 & n38749 ;
  assign n38757 = n38756 ^ n35908 ;
  assign n38790 = n38789 ^ n38783 ;
  assign n38835 = n38790 ^ n38756 ;
  assign n38836 = ~n38757 & n38835 ;
  assign n38837 = n38836 ^ n35908 ;
  assign n38833 = n38832 ^ n38806 ;
  assign n39101 = n38837 ^ n38833 ;
  assign n39102 = n38837 ^ n35902 ;
  assign n39103 = n39101 & n39102 ;
  assign n39104 = n39103 ^ n35902 ;
  assign n39105 = n39104 ^ n39099 ;
  assign n39106 = n39100 & n39105 ;
  assign n39107 = n39106 ^ n35896 ;
  assign n39109 = n39108 ^ n39107 ;
  assign n39110 = n39108 ^ n35893 ;
  assign n39111 = n39109 & ~n39110 ;
  assign n39112 = n39111 ^ n35893 ;
  assign n39113 = n39112 ^ n39097 ;
  assign n39114 = ~n39098 & n39113 ;
  assign n39115 = n39114 ^ n35883 ;
  assign n39117 = n39116 ^ n39115 ;
  assign n39118 = n39116 ^ n35876 ;
  assign n39119 = ~n39117 & n39118 ;
  assign n39120 = n39119 ^ n35876 ;
  assign n39121 = n39120 ^ n39095 ;
  assign n39122 = n39096 & n39121 ;
  assign n39123 = n39122 ^ n35874 ;
  assign n39094 = n39023 ^ n38915 ;
  assign n39124 = n39123 ^ n39094 ;
  assign n39125 = n39123 ^ n35868 ;
  assign n39126 = ~n39124 & n39125 ;
  assign n39127 = n39126 ^ n35868 ;
  assign n39128 = n39127 ^ n39092 ;
  assign n39129 = ~n39093 & n39128 ;
  assign n39130 = n39129 ^ n35858 ;
  assign n39131 = n39130 ^ n39090 ;
  assign n39132 = n39091 & n39131 ;
  assign n39133 = n39132 ^ n36043 ;
  assign n39134 = n39133 ^ n39088 ;
  assign n39135 = ~n39089 & ~n39134 ;
  assign n39136 = n39135 ^ n36057 ;
  assign n39137 = n39136 ^ n39086 ;
  assign n39138 = ~n39087 & ~n39137 ;
  assign n39139 = n39138 ^ n36061 ;
  assign n39141 = n39140 ^ n39139 ;
  assign n39142 = n39140 ^ n35856 ;
  assign n39143 = ~n39141 & ~n39142 ;
  assign n39144 = n39143 ^ n35856 ;
  assign n39145 = n39144 ^ n39084 ;
  assign n39146 = ~n39085 & n39145 ;
  assign n39147 = n39146 ^ n35846 ;
  assign n39083 = n39050 ^ n39043 ;
  assign n39148 = n39147 ^ n39083 ;
  assign n39149 = n39147 ^ n35844 ;
  assign n39150 = n39148 & ~n39149 ;
  assign n39151 = n39150 ^ n35844 ;
  assign n39152 = n39151 ^ n39081 ;
  assign n39153 = ~n39082 & ~n39152 ;
  assign n39154 = n39153 ^ n36080 ;
  assign n39155 = n39154 ^ n39079 ;
  assign n39156 = ~n39080 & n39155 ;
  assign n39157 = n39156 ^ n35838 ;
  assign n39159 = n39158 ^ n39157 ;
  assign n39160 = n39158 ^ n36096 ;
  assign n39161 = ~n39159 & n39160 ;
  assign n39162 = n39161 ^ n36096 ;
  assign n39163 = n39162 ^ n39077 ;
  assign n39164 = n39078 & n39163 ;
  assign n39165 = n39164 ^ n36220 ;
  assign n39166 = n39165 ^ n39075 ;
  assign n39167 = ~n39076 & n39166 ;
  assign n39168 = n39167 ^ n36479 ;
  assign n39350 = n39168 ^ n39073 ;
  assign n39351 = ~n39074 & ~n39350 ;
  assign n39352 = n39351 ^ n36513 ;
  assign n39548 = n39362 ^ n39352 ;
  assign n39549 = n39363 & ~n39548 ;
  assign n39550 = n39549 ^ n36561 ;
  assign n39552 = n39551 ^ n39550 ;
  assign n39553 = n39551 ^ n36650 ;
  assign n39554 = n39552 & n39553 ;
  assign n39555 = n39554 ^ n36650 ;
  assign n39556 = n39555 ^ n39546 ;
  assign n39557 = ~n39547 & n39556 ;
  assign n39558 = n39557 ^ n36676 ;
  assign n39560 = n39559 ^ n39558 ;
  assign n39561 = n39559 ^ n35732 ;
  assign n39562 = n39560 & n39561 ;
  assign n39563 = n39562 ^ n35732 ;
  assign n39522 = n38986 ^ n37418 ;
  assign n39410 = n38706 ^ n38556 ;
  assign n39523 = n39410 ^ n36525 ;
  assign n39524 = n39523 ^ n38986 ;
  assign n39525 = n39524 ^ n39410 ;
  assign n39526 = n39522 & ~n39525 ;
  assign n39527 = n39526 ^ n39523 ;
  assign n39512 = n39511 ^ n39416 ;
  assign n39519 = ~n39512 & ~n39518 ;
  assign n39520 = n39519 ^ n39416 ;
  assign n39544 = n39527 ^ n39520 ;
  assign n39545 = n39544 ^ n35775 ;
  assign n39585 = n39563 ^ n39545 ;
  assign n39364 = n39363 ^ n39352 ;
  assign n39169 = n39168 ^ n39074 ;
  assign n39170 = n39162 ^ n39078 ;
  assign n39171 = n39160 ^ n39157 ;
  assign n39172 = n39151 ^ n39082 ;
  assign n39173 = n39083 ^ n35844 ;
  assign n39174 = n39173 ^ n39147 ;
  assign n39175 = n39144 ^ n39085 ;
  assign n39176 = n39142 ^ n39139 ;
  assign n39177 = n39130 ^ n39091 ;
  assign n39178 = n39094 ^ n35868 ;
  assign n39179 = n39178 ^ n39123 ;
  assign n38834 = n38833 ^ n35902 ;
  assign n38838 = n38837 ^ n38834 ;
  assign n39180 = n39104 ^ n39100 ;
  assign n39181 = ~n38838 & n39180 ;
  assign n39182 = n39110 ^ n39107 ;
  assign n39183 = n39181 & n39182 ;
  assign n39184 = n39112 ^ n39098 ;
  assign n39185 = ~n39183 & ~n39184 ;
  assign n39186 = n39118 ^ n39115 ;
  assign n39187 = ~n39185 & ~n39186 ;
  assign n39188 = n39120 ^ n39096 ;
  assign n39189 = n39187 & ~n39188 ;
  assign n39190 = ~n39179 & ~n39189 ;
  assign n39191 = n39127 ^ n39093 ;
  assign n39192 = n39190 & n39191 ;
  assign n39193 = n39177 & ~n39192 ;
  assign n39194 = n39133 ^ n39089 ;
  assign n39195 = n39193 & n39194 ;
  assign n39196 = n39136 ^ n39087 ;
  assign n39197 = n39195 & ~n39196 ;
  assign n39198 = n39176 & n39197 ;
  assign n39199 = n39175 & ~n39198 ;
  assign n39200 = n39174 & ~n39199 ;
  assign n39201 = n39172 & n39200 ;
  assign n39202 = n39154 ^ n39080 ;
  assign n39203 = n39201 & ~n39202 ;
  assign n39204 = ~n39171 & ~n39203 ;
  assign n39205 = n39170 & ~n39204 ;
  assign n39206 = n39165 ^ n39076 ;
  assign n39207 = n39205 & n39206 ;
  assign n39365 = ~n39169 & ~n39207 ;
  assign n39578 = ~n39364 & n39365 ;
  assign n39579 = n39553 ^ n39550 ;
  assign n39580 = n39578 & ~n39579 ;
  assign n39581 = n39555 ^ n39547 ;
  assign n39582 = ~n39580 & n39581 ;
  assign n39583 = n39561 ^ n39558 ;
  assign n39584 = n39582 & ~n39583 ;
  assign n39610 = n39585 ^ n39584 ;
  assign n39607 = n37055 ^ n28598 ;
  assign n39608 = n39607 ^ n32973 ;
  assign n39609 = n39608 ^ n2867 ;
  assign n39611 = n39610 ^ n39609 ;
  assign n39612 = n39583 ^ n39582 ;
  assign n39613 = n39612 ^ n2813 ;
  assign n39615 = n39581 ^ n39580 ;
  assign n1431 = n1369 ^ n1322 ;
  assign n1432 = n1431 ^ n1428 ;
  assign n1436 = n1435 ^ n1432 ;
  assign n39616 = n39615 ^ n1436 ;
  assign n39617 = n39579 ^ n39578 ;
  assign n1404 = n1307 ^ n1230 ;
  assign n1411 = n1410 ^ n1404 ;
  assign n1421 = n1420 ^ n1411 ;
  assign n39618 = n39617 ^ n1421 ;
  assign n39366 = n39365 ^ n39364 ;
  assign n1718 = n1699 ^ n1212 ;
  assign n1719 = n1718 ^ n1715 ;
  assign n1720 = n1719 ^ n1418 ;
  assign n39367 = n39366 ^ n1720 ;
  assign n39208 = n39207 ^ n39169 ;
  assign n1703 = n1690 ^ n1197 ;
  assign n1710 = n1709 ^ n1703 ;
  assign n1711 = n1710 ^ n983 ;
  assign n39209 = n39208 ^ n1711 ;
  assign n39213 = n39206 ^ n39205 ;
  assign n39210 = n37071 ^ n1673 ;
  assign n39211 = n39210 ^ n857 ;
  assign n39212 = n39211 ^ n1707 ;
  assign n39214 = n39213 ^ n39212 ;
  assign n39218 = n39204 ^ n39170 ;
  assign n39215 = n37067 ^ n1666 ;
  assign n39216 = n39215 ^ n33051 ;
  assign n39217 = n39216 ^ n852 ;
  assign n39219 = n39218 ^ n39217 ;
  assign n39220 = n39203 ^ n39171 ;
  assign n744 = n743 ^ n722 ;
  assign n763 = n762 ^ n744 ;
  assign n770 = n769 ^ n763 ;
  assign n39221 = n39220 ^ n770 ;
  assign n39222 = n37078 ^ n2983 ;
  assign n39223 = n39222 ^ n33055 ;
  assign n39224 = n39223 ^ n757 ;
  assign n39337 = n39224 ^ n39220 ;
  assign n39225 = n39202 ^ n39201 ;
  assign n39226 = n39225 ^ n39224 ;
  assign n39230 = n39200 ^ n39172 ;
  assign n39231 = n39230 ^ n39229 ;
  assign n39236 = n39199 ^ n39174 ;
  assign n39237 = n39236 ^ n39234 ;
  assign n39239 = n37094 ^ n1517 ;
  assign n39240 = n39239 ^ n33092 ;
  assign n39241 = n39240 ^ n27195 ;
  assign n39238 = n39198 ^ n39175 ;
  assign n39242 = n39241 ^ n39238 ;
  assign n39244 = n37098 ^ n28629 ;
  assign n39245 = n39244 ^ n27201 ;
  assign n39246 = n39245 ^ n33097 ;
  assign n39326 = n39246 ^ n39238 ;
  assign n39243 = n39197 ^ n39176 ;
  assign n39247 = n39246 ^ n39243 ;
  assign n39249 = n37105 ^ n28679 ;
  assign n39250 = n39249 ^ n33103 ;
  assign n39251 = n39250 ^ n2930 ;
  assign n39248 = n39196 ^ n39195 ;
  assign n39252 = n39251 ^ n39248 ;
  assign n39257 = n39194 ^ n39193 ;
  assign n39253 = n37109 ^ n28636 ;
  assign n39254 = n39253 ^ n33107 ;
  assign n39255 = n39254 ^ n27208 ;
  assign n39258 = n39257 ^ n39255 ;
  assign n39262 = n39192 ^ n39177 ;
  assign n39259 = n37115 ^ n28665 ;
  assign n39260 = n39259 ^ n33112 ;
  assign n39261 = n39260 ^ n27212 ;
  assign n39263 = n39262 ^ n39261 ;
  assign n39264 = n39191 ^ n39190 ;
  assign n2298 = n2297 ^ n2234 ;
  assign n2311 = n2310 ^ n2298 ;
  assign n2315 = n2314 ^ n2311 ;
  assign n39265 = n39264 ^ n2315 ;
  assign n39269 = n39189 ^ n39179 ;
  assign n39266 = n37122 ^ n28641 ;
  assign n39267 = n39266 ^ n2200 ;
  assign n39268 = n39267 ^ n2305 ;
  assign n39270 = n39269 ^ n39268 ;
  assign n39275 = n39186 ^ n39185 ;
  assign n39272 = n37128 ^ n2071 ;
  assign n39273 = n39272 ^ n33124 ;
  assign n39274 = n39273 ^ n2180 ;
  assign n39276 = n39275 ^ n39274 ;
  assign n39280 = n39184 ^ n39183 ;
  assign n39277 = n37132 ^ n2056 ;
  assign n39278 = n39277 ^ n33128 ;
  assign n39279 = n39278 ^ n27222 ;
  assign n39281 = n39280 ^ n39279 ;
  assign n39292 = n39182 ^ n39181 ;
  assign n39282 = n36535 ^ n3088 ;
  assign n39283 = n39282 ^ n27240 ;
  assign n39284 = n39283 ^ n33138 ;
  assign n39285 = n39284 ^ n39180 ;
  assign n39286 = n39285 ^ n38838 ;
  assign n38795 = n36491 ^ n27230 ;
  assign n38796 = n38795 ^ n3076 ;
  assign n38797 = n38796 ^ n33147 ;
  assign n38839 = n38838 ^ n38797 ;
  assign n38752 = n35828 ^ n28017 ;
  assign n38753 = n38752 ^ n1850 ;
  assign n38754 = n38753 ^ n33142 ;
  assign n3180 = n3179 ^ n3173 ;
  assign n3184 = n3183 ^ n3180 ;
  assign n3194 = n3193 ^ n3184 ;
  assign n38750 = n38749 ^ n36012 ;
  assign n38751 = n3194 & n38750 ;
  assign n38755 = n38754 ^ n38751 ;
  assign n38791 = n38790 ^ n38757 ;
  assign n38792 = n38791 ^ n38754 ;
  assign n38793 = n38755 & n38792 ;
  assign n38794 = n38793 ^ n38754 ;
  assign n39287 = n38797 ^ n38794 ;
  assign n39288 = ~n38839 & ~n39287 ;
  assign n39289 = n39288 ^ n39180 ;
  assign n39290 = n39286 & n39289 ;
  assign n39291 = n39290 ^ n39284 ;
  assign n39293 = n39292 ^ n39291 ;
  assign n39294 = n37137 ^ n28012 ;
  assign n39295 = n39294 ^ n33134 ;
  assign n39296 = n39295 ^ n27226 ;
  assign n39297 = n39296 ^ n39291 ;
  assign n39298 = ~n39293 & ~n39297 ;
  assign n39299 = n39298 ^ n39292 ;
  assign n39300 = n39299 ^ n39279 ;
  assign n39301 = n39281 & n39300 ;
  assign n39302 = n39301 ^ n39280 ;
  assign n39303 = n39302 ^ n39274 ;
  assign n39304 = ~n39276 & n39303 ;
  assign n39305 = n39304 ^ n39274 ;
  assign n39309 = n39305 ^ n39269 ;
  assign n39271 = n39188 ^ n39187 ;
  assign n39306 = n39305 ^ n39271 ;
  assign n2167 = n2160 ^ n2124 ;
  assign n2186 = n2185 ^ n2167 ;
  assign n2193 = n2192 ^ n2186 ;
  assign n39307 = n39271 ^ n2193 ;
  assign n39308 = n39306 & ~n39307 ;
  assign n39310 = n39309 ^ n39308 ;
  assign n39311 = n39270 & n39310 ;
  assign n39312 = n39311 ^ n39269 ;
  assign n39313 = n39312 ^ n2315 ;
  assign n39314 = n39265 & ~n39313 ;
  assign n39315 = n39314 ^ n39264 ;
  assign n39316 = n39315 ^ n39261 ;
  assign n39317 = n39263 & ~n39316 ;
  assign n39318 = n39317 ^ n39262 ;
  assign n39319 = n39318 ^ n39255 ;
  assign n39320 = ~n39258 & n39319 ;
  assign n39256 = n39255 ^ n39248 ;
  assign n39321 = n39320 ^ n39256 ;
  assign n39322 = n39252 & ~n39321 ;
  assign n39323 = n39322 ^ n39251 ;
  assign n39324 = n39323 ^ n39246 ;
  assign n39325 = ~n39247 & n39324 ;
  assign n39327 = n39326 ^ n39325 ;
  assign n39328 = ~n39242 & n39327 ;
  assign n39329 = n39328 ^ n39241 ;
  assign n39330 = n39329 ^ n39234 ;
  assign n39331 = n39237 & n39330 ;
  assign n39235 = n39234 ^ n39230 ;
  assign n39332 = n39331 ^ n39235 ;
  assign n39333 = ~n39231 & ~n39332 ;
  assign n39334 = n39333 ^ n39230 ;
  assign n39335 = n39334 ^ n39224 ;
  assign n39336 = n39226 & ~n39335 ;
  assign n39338 = n39337 ^ n39336 ;
  assign n39339 = n39221 & n39338 ;
  assign n39340 = n39339 ^ n39220 ;
  assign n39341 = n39340 ^ n39217 ;
  assign n39342 = n39219 & ~n39341 ;
  assign n39343 = n39342 ^ n39218 ;
  assign n39344 = n39343 ^ n39212 ;
  assign n39345 = ~n39214 & ~n39344 ;
  assign n39346 = n39345 ^ n39213 ;
  assign n39347 = n39346 ^ n39208 ;
  assign n39348 = n39209 & n39347 ;
  assign n39349 = n39348 ^ n1711 ;
  assign n39619 = n39349 ^ n1720 ;
  assign n39620 = ~n39367 & ~n39619 ;
  assign n39621 = n39620 ^ n39366 ;
  assign n39622 = n39621 ^ n1421 ;
  assign n39623 = ~n39618 & n39622 ;
  assign n39624 = n39623 ^ n39617 ;
  assign n39625 = n39624 ^ n1436 ;
  assign n39626 = n39616 & ~n39625 ;
  assign n39614 = n39612 ^ n1436 ;
  assign n39627 = n39626 ^ n39614 ;
  assign n39628 = n39613 & n39627 ;
  assign n39629 = n39628 ^ n39612 ;
  assign n39630 = n39629 ^ n39609 ;
  assign n39631 = n39611 & ~n39630 ;
  assign n39632 = n39631 ^ n39610 ;
  assign n39601 = n37046 ^ n2648 ;
  assign n39602 = n39601 ^ n27168 ;
  assign n39603 = n39602 ^ n2873 ;
  assign n39564 = n39563 ^ n39544 ;
  assign n39565 = ~n39545 & ~n39564 ;
  assign n39566 = n39565 ^ n35775 ;
  assign n39521 = n39520 ^ n39410 ;
  assign n39528 = n39521 & n39527 ;
  assign n39529 = n39528 ^ n39410 ;
  assign n39487 = n37429 ^ n36566 ;
  assign n39488 = n38167 ^ n37429 ;
  assign n39489 = ~n39487 & ~n39488 ;
  assign n39490 = n39489 ^ n36566 ;
  assign n39403 = n38709 ^ n38554 ;
  assign n39491 = n39490 ^ n39403 ;
  assign n39542 = n39529 ^ n39491 ;
  assign n39543 = n39542 ^ n35812 ;
  assign n39587 = n39566 ^ n39543 ;
  assign n39586 = n39584 & ~n39585 ;
  assign n39600 = n39587 ^ n39586 ;
  assign n39604 = n39603 ^ n39600 ;
  assign n39678 = n39632 ^ n39604 ;
  assign n39891 = n39682 ^ n39678 ;
  assign n39892 = ~n35825 & n39891 ;
  assign n39893 = n39892 ^ n36633 ;
  assign n39685 = n38932 ^ n38262 ;
  assign n39683 = ~n39678 & ~n39682 ;
  assign n39686 = n39683 ^ n37297 ;
  assign n39687 = n39686 ^ n38262 ;
  assign n39688 = n39687 ^ n39683 ;
  assign n39689 = n39685 & n39688 ;
  assign n39690 = n39689 ^ n39686 ;
  assign n39588 = n39586 & n39587 ;
  assign n39530 = n39529 ^ n39403 ;
  assign n39531 = n39491 & ~n39530 ;
  assign n39532 = n39531 ^ n39490 ;
  assign n39478 = n38166 ^ n37411 ;
  assign n39394 = n38712 ^ n38552 ;
  assign n39479 = n39394 ^ n36699 ;
  assign n39480 = n39479 ^ n38166 ;
  assign n39481 = n39480 ^ n39394 ;
  assign n39482 = ~n39478 & n39481 ;
  assign n39483 = n39482 ^ n39479 ;
  assign n39541 = n39532 ^ n39483 ;
  assign n39576 = n39541 ^ n35977 ;
  assign n39567 = n39566 ^ n39542 ;
  assign n39568 = ~n39543 & n39567 ;
  assign n39569 = n39568 ^ n35812 ;
  assign n39577 = n39576 ^ n39569 ;
  assign n39598 = n39588 ^ n39577 ;
  assign n39605 = n39603 ^ n39598 ;
  assign n39606 = n39605 ^ n39598 ;
  assign n39633 = n39632 ^ n39606 ;
  assign n39634 = ~n39604 & n39633 ;
  assign n39635 = n39634 ^ n39605 ;
  assign n39595 = n37050 ^ n2582 ;
  assign n39596 = n39595 ^ n28589 ;
  assign n39597 = n39596 ^ n33006 ;
  assign n39677 = n39635 ^ n39597 ;
  assign n39894 = n39690 ^ n39677 ;
  assign n39895 = n39894 ^ n39892 ;
  assign n39896 = n39893 & n39895 ;
  assign n39897 = n39896 ^ n36633 ;
  assign n39684 = n39683 ^ n39677 ;
  assign n39691 = ~n39684 & n39690 ;
  assign n39692 = n39691 ^ n39683 ;
  assign n39668 = n38922 ^ n38268 ;
  assign n39599 = n39598 ^ n39597 ;
  assign n39636 = ~n39599 & ~n39635 ;
  assign n39637 = n39636 ^ n39598 ;
  assign n39591 = n37392 ^ n28582 ;
  assign n39592 = n39591 ^ n2654 ;
  assign n39593 = n39592 ^ n3218 ;
  assign n39589 = n39577 & ~n39588 ;
  assign n39573 = n35977 ^ n35965 ;
  assign n39570 = n39569 ^ n39541 ;
  assign n39571 = n39569 ^ n35977 ;
  assign n39572 = ~n39570 & n39571 ;
  assign n39574 = n39573 ^ n39572 ;
  assign n39536 = n38160 ^ n37406 ;
  assign n39537 = n37406 ^ n36697 ;
  assign n39538 = n39536 & ~n39537 ;
  assign n39539 = n39538 ^ n36697 ;
  assign n39484 = n38715 ^ n38550 ;
  assign n39485 = n39484 ^ n39394 ;
  assign n39486 = n39485 ^ n39484 ;
  assign n39533 = n39532 ^ n39486 ;
  assign n39534 = ~n39483 & ~n39533 ;
  assign n39535 = n39534 ^ n39485 ;
  assign n39540 = n39539 ^ n39535 ;
  assign n39575 = n39574 ^ n39540 ;
  assign n39590 = n39589 ^ n39575 ;
  assign n39594 = n39593 ^ n39590 ;
  assign n39669 = n39637 ^ n39594 ;
  assign n39670 = n39669 ^ n37469 ;
  assign n39671 = n39670 ^ n38922 ;
  assign n39672 = n39671 ^ n39669 ;
  assign n39673 = n39668 & n39672 ;
  assign n39674 = n39673 ^ n39670 ;
  assign n39889 = n39692 ^ n39674 ;
  assign n39890 = n39889 ^ n36626 ;
  assign n40007 = n39897 ^ n39890 ;
  assign n40166 = n40165 ^ n40007 ;
  assign n40173 = n39891 ^ n35825 ;
  assign n40174 = n40172 & ~n40173 ;
  assign n40167 = n37247 ^ n3240 ;
  assign n40168 = n40167 ^ n2756 ;
  assign n40169 = n40168 ^ n28904 ;
  assign n40175 = n40174 ^ n40169 ;
  assign n40176 = n39894 ^ n39893 ;
  assign n40177 = n40176 ^ n40169 ;
  assign n40178 = n40175 & n40177 ;
  assign n40179 = n40178 ^ n40174 ;
  assign n40180 = n40179 ^ n40165 ;
  assign n40181 = n40166 & ~n40180 ;
  assign n39693 = n39692 ^ n39669 ;
  assign n39694 = n39674 & ~n39693 ;
  assign n39663 = n37873 ^ n37296 ;
  assign n39664 = n38915 ^ n37873 ;
  assign n39665 = n39663 & ~n39664 ;
  assign n39666 = n39665 ^ n37296 ;
  assign n39675 = n39669 ^ n39666 ;
  assign n39695 = n39694 ^ n39675 ;
  assign n39650 = n37309 ^ n36580 ;
  assign n39651 = n38157 ^ n37309 ;
  assign n39652 = n39650 & ~n39651 ;
  assign n39653 = n39652 ^ n36580 ;
  assign n39389 = n38719 ^ n38544 ;
  assign n39646 = n39484 ^ n39389 ;
  assign n39645 = n39539 ^ n39389 ;
  assign n39647 = n39646 ^ n39645 ;
  assign n39648 = n39535 & ~n39647 ;
  assign n39649 = n39648 ^ n39646 ;
  assign n39654 = n39653 ^ n39649 ;
  assign n39655 = n39654 ^ n35830 ;
  assign n39642 = n39540 ^ n35965 ;
  assign n39643 = ~n39574 & n39642 ;
  assign n39644 = n39643 ^ n35965 ;
  assign n39656 = n39655 ^ n39644 ;
  assign n39641 = n39575 & n39589 ;
  assign n39657 = n39656 ^ n39641 ;
  assign n39661 = n39660 ^ n39657 ;
  assign n39638 = n39637 ^ n39593 ;
  assign n39639 = n39594 & ~n39638 ;
  assign n39640 = n39639 ^ n39593 ;
  assign n39662 = n39661 ^ n39640 ;
  assign n39901 = n39695 ^ n39662 ;
  assign n39903 = n39901 ^ n36741 ;
  assign n39898 = n39897 ^ n39889 ;
  assign n39899 = ~n39890 & ~n39898 ;
  assign n39900 = n39899 ^ n36626 ;
  assign n40008 = n39903 ^ n39900 ;
  assign n40182 = n40181 ^ n40008 ;
  assign n40186 = n40008 ^ n40007 ;
  assign n40183 = n33281 ^ n28915 ;
  assign n40184 = n40183 ^ n37700 ;
  assign n40185 = n40184 ^ n1923 ;
  assign n40187 = n40186 ^ n40185 ;
  assign n40188 = n40182 & ~n40187 ;
  assign n40189 = n40188 ^ n40185 ;
  assign n40159 = n37695 ^ n28899 ;
  assign n40160 = n40159 ^ n1928 ;
  assign n40161 = n40160 ^ n27448 ;
  assign n40009 = n40007 & n40008 ;
  assign n39723 = n38841 ^ n37861 ;
  assign n39712 = n37373 ^ n28571 ;
  assign n39713 = n39712 ^ n33445 ;
  assign n39714 = n39713 ^ n3190 ;
  assign n39715 = n39714 ^ n39660 ;
  assign n39710 = n36001 ^ n35830 ;
  assign n39708 = n39389 ^ n36723 ;
  assign n39381 = n38721 ^ n38540 ;
  assign n39709 = n39708 ^ n39381 ;
  assign n39711 = n39710 ^ n39709 ;
  assign n39716 = n39715 ^ n39711 ;
  assign n39706 = n39653 ^ n39389 ;
  assign n39707 = ~n39649 & ~n39706 ;
  assign n39717 = n39716 ^ n39707 ;
  assign n39704 = n39654 ^ n39644 ;
  assign n39705 = ~n39655 & ~n39704 ;
  assign n39718 = n39717 ^ n39705 ;
  assign n39701 = n37307 ^ n36723 ;
  assign n39702 = n38213 ^ n36723 ;
  assign n39703 = n39701 & n39702 ;
  assign n39719 = n39718 ^ n39703 ;
  assign n39700 = n39641 & n39656 ;
  assign n39720 = n39719 ^ n39700 ;
  assign n39698 = n39660 ^ n39640 ;
  assign n39699 = n39661 & n39698 ;
  assign n39721 = n39720 ^ n39699 ;
  assign n39724 = n39721 ^ n37288 ;
  assign n39725 = n39724 ^ n38841 ;
  assign n39726 = n39725 ^ n39721 ;
  assign n39727 = ~n39723 & n39726 ;
  assign n39728 = n39727 ^ n39724 ;
  assign n39667 = n39666 ^ n39662 ;
  assign n39696 = ~n39667 & n39695 ;
  assign n39697 = n39696 ^ n39666 ;
  assign n39888 = n39728 ^ n39697 ;
  assign n40005 = n39888 ^ n36624 ;
  assign n39902 = n39901 ^ n39900 ;
  assign n39904 = n39902 & n39903 ;
  assign n39905 = n39904 ^ n36741 ;
  assign n40006 = n40005 ^ n39905 ;
  assign n40158 = n40009 ^ n40006 ;
  assign n40162 = n40161 ^ n40158 ;
  assign n40522 = n40189 ^ n40162 ;
  assign n40494 = n40185 ^ n40182 ;
  assign n40490 = n38878 ^ n37840 ;
  assign n39784 = n39310 ^ n39268 ;
  assign n40491 = n39784 ^ n38878 ;
  assign n40492 = ~n40490 & n40491 ;
  assign n40493 = n40492 ^ n37840 ;
  assign n40495 = n40494 ^ n40493 ;
  assign n39451 = n39299 ^ n39281 ;
  assign n40431 = n39451 ^ n38896 ;
  assign n40432 = n40173 ^ n40172 ;
  assign n40433 = n40432 ^ n37854 ;
  assign n40434 = n40433 ^ n39451 ;
  assign n40435 = n40434 ^ n40432 ;
  assign n40436 = n40431 & n40435 ;
  assign n40437 = n40436 ^ n40433 ;
  assign n40500 = n38890 ^ n38280 ;
  assign n39448 = n39302 ^ n39276 ;
  assign n40501 = n39448 ^ n38890 ;
  assign n40502 = n40500 & ~n40501 ;
  assign n40503 = n40502 ^ n38280 ;
  assign n40504 = n40503 ^ n40432 ;
  assign n40505 = n40504 ^ n40503 ;
  assign n40329 = n37309 ^ n37248 ;
  assign n40330 = n38969 ^ n37248 ;
  assign n40331 = n40329 & ~n40330 ;
  assign n40332 = n40331 ^ n37309 ;
  assign n38846 = n38748 ^ n38160 ;
  assign n39368 = n39367 ^ n39349 ;
  assign n39369 = n39368 ^ n37429 ;
  assign n39370 = n39369 ^ n38748 ;
  assign n39371 = n39370 ^ n39368 ;
  assign n39372 = ~n38846 & ~n39371 ;
  assign n39373 = n39372 ^ n39369 ;
  assign n39385 = n39346 ^ n39209 ;
  assign n39380 = n38166 ^ n37418 ;
  assign n39382 = n39381 ^ n38166 ;
  assign n39383 = n39380 & n39382 ;
  assign n39384 = n39383 ^ n37418 ;
  assign n39386 = n39385 ^ n39384 ;
  assign n39388 = n38167 ^ n37242 ;
  assign n39390 = n39389 ^ n38167 ;
  assign n39391 = n39388 & n39390 ;
  assign n39392 = n39391 ^ n37242 ;
  assign n39387 = n39343 ^ n39214 ;
  assign n39393 = n39392 ^ n39387 ;
  assign n39831 = n38986 ^ n38195 ;
  assign n39832 = n39484 ^ n38986 ;
  assign n39833 = ~n39831 & ~n39832 ;
  assign n39834 = n39833 ^ n38195 ;
  assign n39843 = n39834 ^ n39387 ;
  assign n39395 = n39394 ^ n38951 ;
  assign n39396 = n39338 ^ n770 ;
  assign n39397 = n39396 ^ n38147 ;
  assign n39398 = n39397 ^ n39394 ;
  assign n39399 = n39398 ^ n39396 ;
  assign n39400 = n39395 & ~n39399 ;
  assign n39401 = n39400 ^ n39397 ;
  assign n39836 = n39834 ^ n39396 ;
  assign n39407 = n39334 ^ n39226 ;
  assign n39402 = n38817 ^ n37252 ;
  assign n39404 = n39403 ^ n38817 ;
  assign n39405 = ~n39402 & ~n39404 ;
  assign n39406 = n39405 ^ n37252 ;
  assign n39408 = n39407 ^ n39406 ;
  assign n39414 = n39332 ^ n39229 ;
  assign n39409 = n38777 ^ n37257 ;
  assign n39411 = n39410 ^ n38777 ;
  assign n39412 = ~n39409 & n39411 ;
  assign n39413 = n39412 ^ n37257 ;
  assign n39415 = n39414 ^ n39413 ;
  assign n39421 = n39329 ^ n39237 ;
  assign n39417 = n39416 ^ n38735 ;
  assign n39418 = n38735 ^ n37791 ;
  assign n39419 = ~n39417 & ~n39418 ;
  assign n39420 = n39419 ^ n37791 ;
  assign n39422 = n39421 ^ n39420 ;
  assign n39425 = n39424 ^ n38476 ;
  assign n39426 = n38476 ^ n37805 ;
  assign n39427 = ~n39425 & n39426 ;
  assign n39428 = n39427 ^ n37805 ;
  assign n39423 = n39327 ^ n39241 ;
  assign n39429 = n39428 ^ n39423 ;
  assign n39432 = n39431 ^ n38336 ;
  assign n39433 = n38336 ^ n37796 ;
  assign n39434 = n39432 & n39433 ;
  assign n39435 = n39434 ^ n37796 ;
  assign n39430 = n39323 ^ n39247 ;
  assign n39436 = n39435 ^ n39430 ;
  assign n39438 = n39356 ^ n38331 ;
  assign n39439 = n38331 ^ n37813 ;
  assign n39440 = ~n39438 & n39439 ;
  assign n39441 = n39440 ^ n37813 ;
  assign n39437 = n39321 ^ n39251 ;
  assign n39442 = n39441 ^ n39437 ;
  assign n39803 = n39318 ^ n39258 ;
  assign n39793 = n39315 ^ n39263 ;
  assign n39443 = n38870 ^ n37811 ;
  assign n39444 = n38876 ^ n37818 ;
  assign n39445 = n37818 ^ n37775 ;
  assign n39446 = ~n39444 & n39445 ;
  assign n39447 = n39446 ^ n37775 ;
  assign n39449 = n39448 ^ n39447 ;
  assign n39450 = n38878 ^ n37827 ;
  assign n39452 = n39451 ^ n37262 ;
  assign n39453 = n39452 ^ n38878 ;
  assign n39454 = n39453 ^ n39451 ;
  assign n39455 = ~n39450 & ~n39454 ;
  assign n39456 = n39455 ^ n39452 ;
  assign n39758 = n39451 ^ n39447 ;
  assign n39457 = n38884 ^ n37833 ;
  assign n39458 = n39296 ^ n39292 ;
  assign n39459 = n39458 ^ n39291 ;
  assign n39460 = n39459 ^ n37508 ;
  assign n39461 = n39460 ^ n38884 ;
  assign n39462 = n39461 ^ n39459 ;
  assign n39463 = n39457 & ~n39462 ;
  assign n39464 = n39463 ^ n39460 ;
  assign n39466 = n38890 ^ n37840 ;
  assign n39467 = n37840 ^ n37499 ;
  assign n39468 = n39466 & n39467 ;
  assign n39469 = n39468 ^ n37499 ;
  assign n39465 = n39289 ^ n39284 ;
  assign n39470 = n39469 ^ n39465 ;
  assign n38840 = n38839 ^ n38794 ;
  assign n39750 = n39469 ^ n38840 ;
  assign n39739 = n38791 ^ n38755 ;
  assign n39742 = n39739 ^ n38840 ;
  assign n39471 = n38902 ^ n38280 ;
  assign n39473 = n38908 ^ n37854 ;
  assign n39474 = n37854 ^ n37280 ;
  assign n39475 = n39473 & ~n39474 ;
  assign n39476 = n39475 ^ n37280 ;
  assign n39472 = n38750 ^ n3194 ;
  assign n39477 = n39476 ^ n39472 ;
  assign n39722 = n39721 ^ n39697 ;
  assign n39729 = n39722 & ~n39728 ;
  assign n39730 = n39729 ^ n39721 ;
  assign n39731 = n39730 ^ n39472 ;
  assign n39732 = n39477 & n39731 ;
  assign n39733 = n39732 ^ n39476 ;
  assign n39734 = n39733 ^ n37278 ;
  assign n39735 = n39734 ^ n38902 ;
  assign n39736 = n39735 ^ n39733 ;
  assign n39737 = ~n39471 & ~n39736 ;
  assign n39738 = n39737 ^ n39734 ;
  assign n39740 = n39739 ^ n39733 ;
  assign n39741 = ~n39738 & n39740 ;
  assign n39743 = n39742 ^ n39741 ;
  assign n39744 = n38896 ^ n37847 ;
  assign n39745 = n37847 ^ n37272 ;
  assign n39746 = n39744 & n39745 ;
  assign n39747 = n39746 ^ n37272 ;
  assign n39748 = n39747 ^ n38840 ;
  assign n39749 = ~n39743 & n39748 ;
  assign n39751 = n39750 ^ n39749 ;
  assign n39752 = ~n39470 & ~n39751 ;
  assign n39753 = n39752 ^ n39469 ;
  assign n39754 = n39753 ^ n39459 ;
  assign n39755 = ~n39464 & ~n39754 ;
  assign n39756 = n39755 ^ n39459 ;
  assign n39757 = n39756 ^ n39447 ;
  assign n39759 = n39758 ^ n39757 ;
  assign n39760 = ~n39456 & n39759 ;
  assign n39761 = n39760 ^ n39758 ;
  assign n39762 = ~n39449 & n39761 ;
  assign n39763 = n39762 ^ n39448 ;
  assign n39764 = n39763 ^ n37849 ;
  assign n39765 = n39764 ^ n38870 ;
  assign n39766 = n39765 ^ n39763 ;
  assign n39767 = n39443 & n39766 ;
  assign n39768 = n39767 ^ n39764 ;
  assign n39774 = n39307 ^ n39305 ;
  assign n39769 = n37842 ^ n37798 ;
  assign n39770 = n38860 ^ n37798 ;
  assign n39771 = n39769 & n39770 ;
  assign n39772 = n39771 ^ n37842 ;
  assign n39775 = n39774 ^ n39772 ;
  assign n39773 = n39772 ^ n39763 ;
  assign n39776 = n39775 ^ n39773 ;
  assign n39777 = n39768 & ~n39776 ;
  assign n39778 = n39777 ^ n39775 ;
  assign n39779 = n38312 ^ n37835 ;
  assign n39780 = n38857 ^ n38312 ;
  assign n39781 = ~n39779 & ~n39780 ;
  assign n39782 = n39781 ^ n37835 ;
  assign n39785 = n39784 ^ n39782 ;
  assign n39783 = n39782 ^ n39772 ;
  assign n39786 = n39785 ^ n39783 ;
  assign n39787 = ~n39778 & n39786 ;
  assign n39788 = n39787 ^ n39785 ;
  assign n39789 = n39312 ^ n39265 ;
  assign n39790 = n39789 ^ n39782 ;
  assign n39791 = ~n39788 & n39790 ;
  assign n39792 = n39791 ^ n39789 ;
  assign n39794 = n39793 ^ n39792 ;
  assign n39795 = n38851 ^ n37788 ;
  assign n39796 = n39793 ^ n37825 ;
  assign n39797 = n39796 ^ n38851 ;
  assign n39798 = n39797 ^ n39793 ;
  assign n39799 = ~n39795 & ~n39798 ;
  assign n39800 = n39799 ^ n39796 ;
  assign n39801 = n39794 & ~n39800 ;
  assign n39802 = n39801 ^ n39793 ;
  assign n39804 = n39803 ^ n39802 ;
  assign n39805 = n39067 ^ n37786 ;
  assign n39806 = n39803 ^ n37820 ;
  assign n39807 = n39806 ^ n39067 ;
  assign n39808 = n39807 ^ n39803 ;
  assign n39809 = n39805 & n39808 ;
  assign n39810 = n39809 ^ n39806 ;
  assign n39811 = ~n39804 & n39810 ;
  assign n39812 = n39811 ^ n39803 ;
  assign n39813 = n39812 ^ n39437 ;
  assign n39814 = n39442 & n39813 ;
  assign n39815 = n39814 ^ n39441 ;
  assign n39816 = n39815 ^ n39430 ;
  assign n39817 = n39436 & n39816 ;
  assign n39818 = n39817 ^ n39435 ;
  assign n39819 = n39818 ^ n39423 ;
  assign n39820 = ~n39429 & ~n39819 ;
  assign n39821 = n39820 ^ n39428 ;
  assign n39822 = n39821 ^ n39420 ;
  assign n39823 = n39422 & ~n39822 ;
  assign n39824 = n39823 ^ n39421 ;
  assign n39825 = n39824 ^ n39413 ;
  assign n39826 = n39415 & n39825 ;
  assign n39827 = n39826 ^ n39414 ;
  assign n39828 = n39827 ^ n39406 ;
  assign n39829 = ~n39408 & n39828 ;
  assign n39830 = n39829 ^ n39407 ;
  assign n39835 = n39834 ^ n39830 ;
  assign n39837 = n39836 ^ n39835 ;
  assign n39838 = ~n39401 & ~n39837 ;
  assign n39839 = n39838 ^ n39836 ;
  assign n39840 = n39340 ^ n39219 ;
  assign n39841 = n39840 ^ n39834 ;
  assign n39842 = ~n39839 & ~n39841 ;
  assign n39844 = n39843 ^ n39842 ;
  assign n39845 = ~n39393 & ~n39844 ;
  assign n39846 = n39845 ^ n39392 ;
  assign n39847 = n39846 ^ n39384 ;
  assign n39848 = n39386 & n39847 ;
  assign n39849 = n39848 ^ n39385 ;
  assign n39374 = n38157 ^ n37411 ;
  assign n39375 = n38783 ^ n38157 ;
  assign n39376 = ~n39374 & n39375 ;
  assign n39377 = n39376 ^ n37411 ;
  assign n39378 = n39377 ^ n39368 ;
  assign n39379 = n39378 ^ n39377 ;
  assign n39850 = n39849 ^ n39379 ;
  assign n39851 = ~n39373 & n39850 ;
  assign n39852 = n39851 ^ n39378 ;
  assign n40265 = n38213 ^ n37406 ;
  assign n40266 = n38832 ^ n38213 ;
  assign n40267 = ~n40265 & n40266 ;
  assign n40268 = n40267 ^ n37406 ;
  assign n40270 = n40268 ^ n39377 ;
  assign n39853 = n39621 ^ n39618 ;
  assign n40269 = n40268 ^ n39853 ;
  assign n40271 = n40270 ^ n40269 ;
  assign n40272 = n39852 & ~n40271 ;
  assign n40273 = n40272 ^ n40270 ;
  assign n40323 = n39627 ^ n2813 ;
  assign n40325 = n40323 ^ n40268 ;
  assign n40274 = n39624 ^ n39616 ;
  assign n40324 = n40323 ^ n40274 ;
  assign n40326 = n40325 ^ n40324 ;
  assign n40327 = ~n40273 & ~n40326 ;
  assign n40328 = n40327 ^ n40325 ;
  assign n40333 = n40332 ^ n40328 ;
  assign n40334 = n40333 ^ n36580 ;
  assign n39854 = n39853 ^ n39852 ;
  assign n39855 = n39854 ^ n36699 ;
  assign n39856 = n39849 ^ n39373 ;
  assign n39857 = n39856 ^ n36566 ;
  assign n39986 = n39846 ^ n39386 ;
  assign n39858 = n39844 ^ n39392 ;
  assign n39859 = n39858 ^ n36485 ;
  assign n39977 = n39840 ^ n39839 ;
  assign n39861 = n39827 ^ n39408 ;
  assign n39862 = n39861 ^ n37329 ;
  assign n39864 = n39821 ^ n39422 ;
  assign n39865 = n39864 ^ n37232 ;
  assign n39867 = n39815 ^ n39436 ;
  assign n39868 = n39867 ^ n37015 ;
  assign n39951 = n39812 ^ n39442 ;
  assign n39870 = n39800 ^ n39792 ;
  assign n39871 = n39870 ^ n36964 ;
  assign n39872 = n39789 ^ n39788 ;
  assign n39873 = n39872 ^ n36951 ;
  assign n39874 = n39784 ^ n39778 ;
  assign n39875 = n39874 ^ n36894 ;
  assign n39876 = n39774 ^ n39768 ;
  assign n39877 = n39876 ^ n36794 ;
  assign n39879 = n39756 ^ n39456 ;
  assign n39880 = n39879 ^ n36782 ;
  assign n39882 = n39751 ^ n39465 ;
  assign n39883 = n39882 ^ n36606 ;
  assign n39884 = n39747 ^ n39743 ;
  assign n39885 = n39884 ^ n36600 ;
  assign n39886 = n39739 ^ n39738 ;
  assign n39887 = n39886 ^ n36611 ;
  assign n39910 = n39730 ^ n39477 ;
  assign n39906 = n39905 ^ n39888 ;
  assign n39907 = n39905 ^ n36624 ;
  assign n39908 = ~n39906 & ~n39907 ;
  assign n39909 = n39908 ^ n36624 ;
  assign n39911 = n39910 ^ n39909 ;
  assign n39912 = n39910 ^ n36614 ;
  assign n39913 = ~n39911 & n39912 ;
  assign n39914 = n39913 ^ n36614 ;
  assign n39915 = n39914 ^ n39886 ;
  assign n39916 = n39887 & n39915 ;
  assign n39917 = n39916 ^ n36611 ;
  assign n39918 = n39917 ^ n39884 ;
  assign n39919 = ~n39885 & ~n39918 ;
  assign n39920 = n39919 ^ n36600 ;
  assign n39921 = n39920 ^ n39882 ;
  assign n39922 = ~n39883 & n39921 ;
  assign n39923 = n39922 ^ n36606 ;
  assign n39881 = n39753 ^ n39464 ;
  assign n39924 = n39923 ^ n39881 ;
  assign n39925 = n39923 ^ n36597 ;
  assign n39926 = ~n39924 & n39925 ;
  assign n39927 = n39926 ^ n36597 ;
  assign n39928 = n39927 ^ n39879 ;
  assign n39929 = n39880 & n39928 ;
  assign n39930 = n39929 ^ n36782 ;
  assign n39878 = n39761 ^ n39448 ;
  assign n39931 = n39930 ^ n39878 ;
  assign n39932 = n39930 ^ n36590 ;
  assign n39933 = ~n39931 & ~n39932 ;
  assign n39934 = n39933 ^ n36590 ;
  assign n39935 = n39934 ^ n39876 ;
  assign n39936 = ~n39877 & ~n39935 ;
  assign n39937 = n39936 ^ n36794 ;
  assign n39938 = n39937 ^ n39874 ;
  assign n39939 = ~n39875 & ~n39938 ;
  assign n39940 = n39939 ^ n36894 ;
  assign n39941 = n39940 ^ n39872 ;
  assign n39942 = n39873 & n39941 ;
  assign n39943 = n39942 ^ n36951 ;
  assign n39944 = n39943 ^ n39870 ;
  assign n39945 = ~n39871 & n39944 ;
  assign n39946 = n39945 ^ n36964 ;
  assign n39869 = n39810 ^ n39802 ;
  assign n39947 = n39946 ^ n39869 ;
  assign n39948 = n39946 ^ n36977 ;
  assign n39949 = ~n39947 & ~n39948 ;
  assign n39950 = n39949 ^ n36977 ;
  assign n39952 = n39951 ^ n39950 ;
  assign n39953 = n39951 ^ n37006 ;
  assign n39954 = ~n39952 & ~n39953 ;
  assign n39955 = n39954 ^ n37006 ;
  assign n39956 = n39955 ^ n39867 ;
  assign n39957 = n39868 & ~n39956 ;
  assign n39958 = n39957 ^ n37015 ;
  assign n39866 = n39818 ^ n39429 ;
  assign n39959 = n39958 ^ n39866 ;
  assign n39960 = n39958 ^ n37035 ;
  assign n39961 = ~n39959 & n39960 ;
  assign n39962 = n39961 ^ n37035 ;
  assign n39963 = n39962 ^ n39864 ;
  assign n39964 = n39865 & ~n39963 ;
  assign n39965 = n39964 ^ n37232 ;
  assign n39863 = n39824 ^ n39415 ;
  assign n39966 = n39965 ^ n39863 ;
  assign n39967 = n39965 ^ n37316 ;
  assign n39968 = ~n39966 & ~n39967 ;
  assign n39969 = n39968 ^ n37316 ;
  assign n39970 = n39969 ^ n39861 ;
  assign n39971 = n39862 & n39970 ;
  assign n39972 = n39971 ^ n37329 ;
  assign n39860 = n39830 ^ n39401 ;
  assign n39973 = n39972 ^ n39860 ;
  assign n39974 = n39972 ^ n37255 ;
  assign n39975 = ~n39973 & n39974 ;
  assign n39976 = n39975 ^ n37255 ;
  assign n39978 = n39977 ^ n39976 ;
  assign n39979 = n39858 ^ n37253 ;
  assign n39980 = n39979 ^ n39858 ;
  assign n39981 = n39980 ^ n39976 ;
  assign n39982 = n39978 & ~n39981 ;
  assign n39983 = n39982 ^ n39979 ;
  assign n39984 = n39859 & n39983 ;
  assign n39985 = n39984 ^ n36485 ;
  assign n39987 = n39986 ^ n39985 ;
  assign n39988 = n39986 ^ n36525 ;
  assign n39989 = ~n39987 & ~n39988 ;
  assign n39990 = n39989 ^ n36525 ;
  assign n39991 = n39990 ^ n39856 ;
  assign n39992 = ~n39857 & n39991 ;
  assign n39993 = n39992 ^ n36566 ;
  assign n40277 = n39993 ^ n39854 ;
  assign n40278 = ~n39855 & n40277 ;
  assign n40279 = n40278 ^ n36699 ;
  assign n40275 = n40274 ^ n40273 ;
  assign n40319 = n40279 ^ n40275 ;
  assign n40320 = n40279 ^ n36697 ;
  assign n40321 = n40319 & n40320 ;
  assign n40322 = n40321 ^ n36697 ;
  assign n40335 = n40334 ^ n40322 ;
  assign n39994 = n39993 ^ n39855 ;
  assign n39995 = n39990 ^ n39857 ;
  assign n39996 = n39988 ^ n39985 ;
  assign n39997 = n39869 ^ n36977 ;
  assign n39998 = n39997 ^ n39946 ;
  assign n39999 = n39943 ^ n39871 ;
  assign n40000 = n39940 ^ n36951 ;
  assign n40001 = n40000 ^ n39872 ;
  assign n40002 = n39937 ^ n39875 ;
  assign n40003 = n39881 ^ n36597 ;
  assign n40004 = n40003 ^ n39923 ;
  assign n40010 = n40006 & n40009 ;
  assign n40011 = n39912 ^ n39909 ;
  assign n40012 = ~n40010 & ~n40011 ;
  assign n40013 = n39914 ^ n39887 ;
  assign n40014 = ~n40012 & n40013 ;
  assign n40015 = n39917 ^ n39885 ;
  assign n40016 = n40014 & n40015 ;
  assign n40017 = n39920 ^ n39883 ;
  assign n40018 = ~n40016 & n40017 ;
  assign n40019 = ~n40004 & n40018 ;
  assign n40020 = n39927 ^ n39880 ;
  assign n40021 = ~n40019 & n40020 ;
  assign n40022 = n39878 ^ n36590 ;
  assign n40023 = n40022 ^ n39930 ;
  assign n40024 = n40021 & n40023 ;
  assign n40025 = n39934 ^ n39877 ;
  assign n40026 = n40024 & ~n40025 ;
  assign n40027 = n40002 & n40026 ;
  assign n40028 = ~n40001 & ~n40027 ;
  assign n40029 = n39999 & ~n40028 ;
  assign n40030 = n39998 & n40029 ;
  assign n40031 = n39953 ^ n39950 ;
  assign n40032 = n40030 & ~n40031 ;
  assign n40033 = n39955 ^ n39868 ;
  assign n40034 = ~n40032 & n40033 ;
  assign n40035 = n39866 ^ n37035 ;
  assign n40036 = n40035 ^ n39958 ;
  assign n40037 = ~n40034 & ~n40036 ;
  assign n40038 = n39962 ^ n39865 ;
  assign n40039 = n40037 & ~n40038 ;
  assign n40040 = n39863 ^ n37316 ;
  assign n40041 = n40040 ^ n39965 ;
  assign n40042 = ~n40039 & ~n40041 ;
  assign n40043 = n39969 ^ n39862 ;
  assign n40044 = n40042 & ~n40043 ;
  assign n40045 = n39860 ^ n37255 ;
  assign n40046 = n40045 ^ n39972 ;
  assign n40047 = n40044 & n40046 ;
  assign n40048 = n39977 ^ n37253 ;
  assign n40049 = n40048 ^ n39976 ;
  assign n40050 = ~n40047 & ~n40049 ;
  assign n40051 = n39983 ^ n36485 ;
  assign n40052 = n40050 & n40051 ;
  assign n40053 = n39996 & n40052 ;
  assign n40054 = ~n39995 & n40053 ;
  assign n40264 = n39994 & ~n40054 ;
  assign n40276 = n40275 ^ n36697 ;
  assign n40280 = n40279 ^ n40276 ;
  assign n40336 = n40264 & n40280 ;
  assign n40412 = ~n40335 & n40336 ;
  assign n40407 = n40332 ^ n40323 ;
  assign n40408 = n40328 & n40407 ;
  assign n40402 = n40323 ^ n37307 ;
  assign n40401 = n39629 ^ n39611 ;
  assign n40403 = n40402 ^ n40401 ;
  assign n40404 = n40403 ^ n36724 ;
  assign n40338 = n38064 ^ n3221 ;
  assign n40339 = n40338 ^ n34215 ;
  assign n40340 = n40339 ^ n2671 ;
  assign n40405 = n40404 ^ n40340 ;
  assign n2661 = n2660 ^ n2534 ;
  assign n2677 = n2676 ^ n2661 ;
  assign n2684 = n2683 ^ n2677 ;
  assign n40406 = n40405 ^ n2684 ;
  assign n40409 = n40408 ^ n40406 ;
  assign n40399 = n40333 ^ n40322 ;
  assign n40400 = n40334 & n40399 ;
  assign n40410 = n40409 ^ n40400 ;
  assign n40396 = n38237 ^ n37307 ;
  assign n40397 = n39003 ^ n38237 ;
  assign n40398 = n40396 & ~n40397 ;
  assign n40411 = n40410 ^ n40398 ;
  assign n40413 = n40412 ^ n40411 ;
  assign n40337 = n40336 ^ n40335 ;
  assign n40341 = n40340 ^ n40337 ;
  assign n40282 = n38069 ^ n2597 ;
  assign n40283 = n40282 ^ n34204 ;
  assign n40284 = n40283 ^ n27927 ;
  assign n40281 = n40280 ^ n40264 ;
  assign n40285 = n40284 ^ n40281 ;
  assign n40055 = n40054 ^ n39994 ;
  assign n38843 = n38073 ^ n29378 ;
  assign n38844 = n38843 ^ n34021 ;
  assign n38845 = n38844 ^ n3122 ;
  assign n40056 = n40055 ^ n38845 ;
  assign n40058 = n29469 ^ n2895 ;
  assign n40059 = n40058 ^ n33828 ;
  assign n40060 = n40059 ^ n27522 ;
  assign n40057 = n40053 ^ n39995 ;
  assign n40061 = n40060 ^ n40057 ;
  assign n40063 = n38083 ^ n2857 ;
  assign n40064 = n40063 ^ n33833 ;
  assign n40065 = n40064 ^ n27867 ;
  assign n40062 = n40052 ^ n39996 ;
  assign n40066 = n40065 ^ n40062 ;
  assign n40068 = n38088 ^ n2842 ;
  assign n40069 = n40068 ^ n33838 ;
  assign n40070 = n40069 ^ n27861 ;
  assign n40067 = n40051 ^ n40050 ;
  assign n40071 = n40070 ^ n40067 ;
  assign n40073 = n29387 ^ n1766 ;
  assign n40074 = n40073 ^ n1262 ;
  assign n40075 = n40074 ^ n27856 ;
  assign n40251 = n40075 ^ n40067 ;
  assign n40072 = n40049 ^ n40047 ;
  assign n40076 = n40075 ^ n40072 ;
  assign n40080 = n40046 ^ n40044 ;
  assign n40077 = n1757 ^ n1746 ;
  assign n40078 = n40077 ^ n33845 ;
  assign n40079 = n40078 ^ n1253 ;
  assign n40081 = n40080 ^ n40079 ;
  assign n40082 = n40043 ^ n40042 ;
  assign n1071 = n1070 ^ n1004 ;
  assign n1084 = n1083 ^ n1071 ;
  assign n1091 = n1090 ^ n1084 ;
  assign n40083 = n40082 ^ n1091 ;
  assign n40087 = n40041 ^ n40039 ;
  assign n40084 = n38098 ^ n1728 ;
  assign n40085 = n40084 ^ n964 ;
  assign n40086 = n40085 ^ n1078 ;
  assign n40088 = n40087 ^ n40086 ;
  assign n40089 = n40038 ^ n40037 ;
  assign n40090 = n40089 ^ n957 ;
  assign n40236 = n40093 ^ n40089 ;
  assign n40094 = n40036 ^ n40034 ;
  assign n40095 = n40094 ^ n40093 ;
  assign n40096 = n40033 ^ n40032 ;
  assign n40097 = n40096 ^ n1616 ;
  assign n40102 = n40031 ^ n40030 ;
  assign n40103 = n40102 ^ n40100 ;
  assign n40107 = n40029 ^ n39998 ;
  assign n40104 = n37647 ^ n1572 ;
  assign n40105 = n40104 ^ n33909 ;
  assign n40106 = n40105 ^ n2969 ;
  assign n40108 = n40107 ^ n40106 ;
  assign n40112 = n40028 ^ n39999 ;
  assign n40109 = n37652 ^ n29411 ;
  assign n40110 = n40109 ^ n2957 ;
  assign n40111 = n40110 ^ n27786 ;
  assign n40113 = n40112 ^ n40111 ;
  assign n40114 = n40027 ^ n40001 ;
  assign n40118 = n40117 ^ n40114 ;
  assign n40120 = n37665 ^ n2939 ;
  assign n40121 = n40120 ^ n33922 ;
  assign n40122 = n40121 ^ n27794 ;
  assign n40219 = n40122 ^ n40114 ;
  assign n40119 = n40026 ^ n40002 ;
  assign n40123 = n40122 ^ n40119 ;
  assign n40127 = n40025 ^ n40024 ;
  assign n40124 = n37669 ^ n28963 ;
  assign n40125 = n40124 ^ n33926 ;
  assign n40126 = n40125 ^ n27799 ;
  assign n40128 = n40127 ^ n40126 ;
  assign n40132 = n40023 ^ n40021 ;
  assign n40129 = n37675 ^ n28875 ;
  assign n40130 = n40129 ^ n33931 ;
  assign n40131 = n40130 ^ n27803 ;
  assign n40133 = n40132 ^ n40131 ;
  assign n40134 = n40020 ^ n40019 ;
  assign n2432 = n2395 ^ n2359 ;
  assign n2433 = n2432 ^ n2429 ;
  assign n2440 = n2439 ^ n2433 ;
  assign n40135 = n40134 ^ n2440 ;
  assign n40136 = n40018 ^ n40004 ;
  assign n2399 = n2386 ^ n2341 ;
  assign n2415 = n2414 ^ n2399 ;
  assign n2422 = n2421 ^ n2415 ;
  assign n40137 = n40136 ^ n2422 ;
  assign n40139 = n37733 ^ n2267 ;
  assign n40140 = n40139 ^ n33941 ;
  assign n40141 = n40140 ^ n2411 ;
  assign n40138 = n40017 ^ n40016 ;
  assign n40142 = n40141 ^ n40138 ;
  assign n40144 = n37686 ^ n2252 ;
  assign n40145 = n40144 ^ n33946 ;
  assign n40146 = n40145 ^ n27436 ;
  assign n40201 = n40146 ^ n40138 ;
  assign n40143 = n40015 ^ n40014 ;
  assign n40147 = n40146 ^ n40143 ;
  assign n40149 = n37691 ^ n28890 ;
  assign n40150 = n40149 ^ n33951 ;
  assign n40151 = n40150 ^ n27469 ;
  assign n40148 = n40013 ^ n40012 ;
  assign n40152 = n40151 ^ n40148 ;
  assign n40156 = n40011 ^ n40010 ;
  assign n40153 = n37720 ^ n28894 ;
  assign n40154 = n40153 ^ n33955 ;
  assign n40155 = n40154 ^ n1988 ;
  assign n40157 = n40156 ^ n40155 ;
  assign n40190 = n40189 ^ n40158 ;
  assign n40191 = ~n40162 & n40190 ;
  assign n40192 = n40191 ^ n40161 ;
  assign n40193 = n40192 ^ n40155 ;
  assign n40194 = n40157 & ~n40193 ;
  assign n40195 = n40194 ^ n40156 ;
  assign n40196 = n40195 ^ n40151 ;
  assign n40197 = n40152 & n40196 ;
  assign n40198 = n40197 ^ n40151 ;
  assign n40199 = n40198 ^ n40146 ;
  assign n40200 = ~n40147 & n40199 ;
  assign n40202 = n40201 ^ n40200 ;
  assign n40203 = ~n40142 & n40202 ;
  assign n40204 = n40203 ^ n40141 ;
  assign n40205 = n40204 ^ n40136 ;
  assign n40206 = ~n40137 & n40205 ;
  assign n40207 = n40206 ^ n2422 ;
  assign n40208 = n40207 ^ n2440 ;
  assign n40209 = n40135 & ~n40208 ;
  assign n40210 = n40209 ^ n40134 ;
  assign n40211 = n40210 ^ n40131 ;
  assign n40212 = ~n40133 & ~n40211 ;
  assign n40213 = n40212 ^ n40132 ;
  assign n40214 = n40213 ^ n40126 ;
  assign n40215 = n40128 & n40214 ;
  assign n40216 = n40215 ^ n40127 ;
  assign n40217 = n40216 ^ n40122 ;
  assign n40218 = ~n40123 & n40217 ;
  assign n40220 = n40219 ^ n40218 ;
  assign n40221 = n40118 & ~n40220 ;
  assign n40222 = n40221 ^ n40117 ;
  assign n40223 = n40222 ^ n40111 ;
  assign n40224 = n40113 & ~n40223 ;
  assign n40225 = n40224 ^ n40112 ;
  assign n40226 = n40225 ^ n40106 ;
  assign n40227 = ~n40108 & ~n40226 ;
  assign n40228 = n40227 ^ n40107 ;
  assign n40229 = n40228 ^ n40100 ;
  assign n40230 = n40103 & ~n40229 ;
  assign n40101 = n40100 ^ n40096 ;
  assign n40231 = n40230 ^ n40101 ;
  assign n40232 = ~n40097 & ~n40231 ;
  assign n40233 = n40232 ^ n40096 ;
  assign n40234 = n40233 ^ n40093 ;
  assign n40235 = ~n40095 & ~n40234 ;
  assign n40237 = n40236 ^ n40235 ;
  assign n40238 = n40090 & n40237 ;
  assign n40239 = n40238 ^ n40089 ;
  assign n40240 = n40239 ^ n40086 ;
  assign n40241 = n40088 & ~n40240 ;
  assign n40242 = n40241 ^ n40087 ;
  assign n40243 = n40242 ^ n1091 ;
  assign n40244 = ~n40083 & ~n40243 ;
  assign n40245 = n40244 ^ n40082 ;
  assign n40246 = n40245 ^ n40079 ;
  assign n40247 = n40081 & n40246 ;
  assign n40248 = n40247 ^ n40080 ;
  assign n40249 = n40248 ^ n40075 ;
  assign n40250 = ~n40076 & n40249 ;
  assign n40252 = n40251 ^ n40250 ;
  assign n40253 = ~n40071 & n40252 ;
  assign n40254 = n40253 ^ n40070 ;
  assign n40255 = n40254 ^ n40062 ;
  assign n40256 = ~n40066 & n40255 ;
  assign n40257 = n40256 ^ n40065 ;
  assign n40258 = n40257 ^ n40057 ;
  assign n40259 = n40061 & ~n40258 ;
  assign n40260 = n40259 ^ n40060 ;
  assign n40261 = n40260 ^ n38845 ;
  assign n40262 = ~n40056 & ~n40261 ;
  assign n40263 = n40262 ^ n40055 ;
  assign n40316 = n40281 ^ n40263 ;
  assign n40317 = n40285 & n40316 ;
  assign n40318 = n40317 ^ n40284 ;
  assign n40394 = n40340 ^ n40318 ;
  assign n40395 = ~n40341 & n40394 ;
  assign n40414 = n40413 ^ n40395 ;
  assign n40390 = n39459 ^ n38902 ;
  assign n40391 = n38902 ^ n37861 ;
  assign n40392 = ~n40390 & ~n40391 ;
  assign n40393 = n40392 ^ n37861 ;
  assign n40415 = n40414 ^ n40393 ;
  assign n40310 = n38908 ^ n37873 ;
  assign n40311 = n39465 ^ n38908 ;
  assign n40312 = ~n40310 & n40311 ;
  assign n40313 = n40312 ^ n37873 ;
  assign n40286 = n40285 ^ n40263 ;
  assign n40314 = n40313 ^ n40286 ;
  assign n38842 = n38841 ^ n38840 ;
  assign n40287 = n40286 ^ n38268 ;
  assign n40288 = n40287 ^ n38840 ;
  assign n40289 = n40288 ^ n40286 ;
  assign n40290 = n38842 & ~n40289 ;
  assign n40291 = n40290 ^ n40287 ;
  assign n40298 = n40260 ^ n40056 ;
  assign n40292 = n38922 ^ n38247 ;
  assign n40293 = n39472 ^ n38922 ;
  assign n40294 = ~n40292 & n40293 ;
  assign n40295 = n40294 ^ n38247 ;
  assign n40296 = n40257 ^ n40061 ;
  assign n40297 = n40295 & n40296 ;
  assign n40299 = n40298 ^ n40297 ;
  assign n40300 = n39739 ^ n38915 ;
  assign n40301 = n40297 ^ n38262 ;
  assign n40302 = n40301 ^ n39739 ;
  assign n40303 = n40302 ^ n40297 ;
  assign n40304 = n40300 & n40303 ;
  assign n40305 = n40304 ^ n40301 ;
  assign n40306 = ~n40299 & ~n40305 ;
  assign n40307 = n40306 ^ n40298 ;
  assign n40308 = n40307 ^ n40286 ;
  assign n40309 = ~n40291 & n40308 ;
  assign n40315 = n40314 ^ n40309 ;
  assign n40342 = n40341 ^ n40318 ;
  assign n40387 = n40342 ^ n40313 ;
  assign n40388 = ~n40315 & n40387 ;
  assign n40389 = n40388 ^ n40342 ;
  assign n40428 = n40393 ^ n40389 ;
  assign n40429 = ~n40415 & n40428 ;
  assign n40430 = n40429 ^ n40414 ;
  assign n40506 = n40505 ^ n40430 ;
  assign n40507 = n40437 & n40506 ;
  assign n40508 = n40507 ^ n40504 ;
  assign n40509 = n40176 ^ n40175 ;
  assign n40510 = n40509 ^ n40503 ;
  assign n40511 = ~n40508 & n40510 ;
  assign n40512 = n40511 ^ n40509 ;
  assign n40496 = n38884 ^ n37847 ;
  assign n40497 = n39774 ^ n38884 ;
  assign n40498 = n40496 & n40497 ;
  assign n40499 = n40498 ^ n37847 ;
  assign n40513 = n40512 ^ n40499 ;
  assign n40514 = n40179 ^ n40166 ;
  assign n40515 = n40514 ^ n40493 ;
  assign n40516 = n40515 ^ n40499 ;
  assign n40517 = n40516 ^ n40493 ;
  assign n40518 = ~n40513 & ~n40517 ;
  assign n40519 = n40518 ^ n40515 ;
  assign n40520 = ~n40495 & ~n40519 ;
  assign n40521 = n40520 ^ n40494 ;
  assign n40523 = n40522 ^ n40521 ;
  assign n40524 = n39789 ^ n37833 ;
  assign n40525 = n39789 ^ n38876 ;
  assign n40526 = n40524 & ~n40525 ;
  assign n40527 = n40526 ^ n37833 ;
  assign n40528 = n40527 ^ n40521 ;
  assign n40529 = n40523 & n40528 ;
  assign n40530 = n40529 ^ n40522 ;
  assign n40488 = n40192 ^ n40157 ;
  assign n40484 = n39793 ^ n38870 ;
  assign n40485 = n38870 ^ n37827 ;
  assign n40486 = ~n40484 & ~n40485 ;
  assign n40487 = n40486 ^ n37827 ;
  assign n40489 = n40488 ^ n40487 ;
  assign n40585 = n40530 ^ n40489 ;
  assign n40662 = n40585 ^ n37262 ;
  assign n40605 = n40527 ^ n40522 ;
  assign n40606 = n40605 ^ n40521 ;
  assign n40586 = n40519 ^ n40494 ;
  assign n40587 = n40586 ^ n37499 ;
  assign n40596 = n40514 ^ n40499 ;
  assign n40597 = n40596 ^ n40512 ;
  assign n40588 = n40509 ^ n40508 ;
  assign n40589 = n40588 ^ n37278 ;
  assign n40438 = n40437 ^ n40430 ;
  assign n40439 = n40438 ^ n37280 ;
  assign n40416 = n40415 ^ n40389 ;
  assign n40417 = n40416 ^ n37288 ;
  assign n40352 = n40307 ^ n40291 ;
  assign n40345 = n40296 ^ n40295 ;
  assign n40346 = ~n36578 & n40345 ;
  assign n40347 = n40346 ^ n37297 ;
  assign n40348 = n40305 ^ n40298 ;
  assign n40349 = n40348 ^ n40346 ;
  assign n40350 = n40347 & n40349 ;
  assign n40351 = n40350 ^ n37297 ;
  assign n40353 = n40352 ^ n40351 ;
  assign n40354 = n40352 ^ n37469 ;
  assign n40355 = ~n40353 & ~n40354 ;
  assign n40356 = n40355 ^ n37469 ;
  assign n40343 = n40342 ^ n40315 ;
  assign n40383 = n40356 ^ n40343 ;
  assign n40384 = n40356 ^ n37296 ;
  assign n40385 = ~n40383 & n40384 ;
  assign n40386 = n40385 ^ n37296 ;
  assign n40440 = n40416 ^ n40386 ;
  assign n40441 = n40417 & n40440 ;
  assign n40442 = n40441 ^ n37288 ;
  assign n40590 = n40442 ^ n40438 ;
  assign n40591 = ~n40439 & n40590 ;
  assign n40592 = n40591 ^ n37280 ;
  assign n40593 = n40592 ^ n40588 ;
  assign n40594 = ~n40589 & n40593 ;
  assign n40595 = n40594 ^ n37278 ;
  assign n40598 = n40597 ^ n40595 ;
  assign n40599 = n40597 ^ n37272 ;
  assign n40600 = ~n40598 & ~n40599 ;
  assign n40601 = n40600 ^ n37272 ;
  assign n40602 = n40601 ^ n40586 ;
  assign n40603 = ~n40587 & ~n40602 ;
  assign n40604 = n40603 ^ n37499 ;
  assign n40607 = n40606 ^ n40604 ;
  assign n40608 = n40606 ^ n37508 ;
  assign n40609 = ~n40607 & n40608 ;
  assign n40610 = n40609 ^ n37508 ;
  assign n40663 = n40662 ^ n40610 ;
  assign n40443 = n40442 ^ n40439 ;
  assign n40418 = n40417 ^ n40386 ;
  assign n40344 = n40343 ^ n37296 ;
  assign n40357 = n40356 ^ n40344 ;
  assign n40359 = n40354 ^ n40351 ;
  assign n40419 = n40357 & n40359 ;
  assign n40444 = n40418 & n40419 ;
  assign n40664 = ~n40443 & ~n40444 ;
  assign n40665 = n40592 ^ n40589 ;
  assign n40666 = ~n40664 & n40665 ;
  assign n40667 = n40599 ^ n40595 ;
  assign n40668 = n40666 & n40667 ;
  assign n40669 = n40601 ^ n40587 ;
  assign n40670 = ~n40668 & n40669 ;
  assign n40671 = n40608 ^ n40604 ;
  assign n40672 = n40670 & n40671 ;
  assign n40673 = ~n40663 & ~n40672 ;
  assign n40611 = n40610 ^ n40585 ;
  assign n40612 = n40610 ^ n37262 ;
  assign n40613 = ~n40611 & n40612 ;
  assign n40614 = n40613 ^ n37262 ;
  assign n40531 = n40530 ^ n40488 ;
  assign n40532 = n40489 & ~n40531 ;
  assign n40533 = n40532 ^ n40530 ;
  assign n40477 = n39803 ^ n38860 ;
  assign n40478 = n40195 ^ n40152 ;
  assign n40479 = n40478 ^ n37818 ;
  assign n40480 = n40479 ^ n39803 ;
  assign n40481 = n40480 ^ n40478 ;
  assign n40482 = ~n40477 & ~n40481 ;
  assign n40483 = n40482 ^ n40479 ;
  assign n40583 = n40533 ^ n40483 ;
  assign n40584 = n40583 ^ n37775 ;
  assign n40674 = n40614 ^ n40584 ;
  assign n40675 = n40673 & n40674 ;
  assign n40472 = n38857 ^ n37811 ;
  assign n40473 = n39437 ^ n38857 ;
  assign n40474 = n40472 & n40473 ;
  assign n40475 = n40474 ^ n37811 ;
  assign n40535 = n40478 ^ n40475 ;
  assign n40534 = n40533 ^ n40475 ;
  assign n40536 = n40535 ^ n40534 ;
  assign n40537 = n40483 & ~n40536 ;
  assign n40538 = n40537 ^ n40535 ;
  assign n40451 = n40198 ^ n40147 ;
  assign n40582 = n40538 ^ n40451 ;
  assign n40676 = n40582 ^ n37849 ;
  assign n40615 = n40614 ^ n40583 ;
  assign n40616 = ~n40584 & n40615 ;
  assign n40617 = n40616 ^ n37775 ;
  assign n40677 = n40676 ^ n40617 ;
  assign n40678 = n40675 & ~n40677 ;
  assign n40476 = n40475 ^ n40451 ;
  assign n40539 = n40476 & ~n40538 ;
  assign n40540 = n40539 ^ n40475 ;
  assign n40467 = n38851 ^ n37798 ;
  assign n40468 = n39430 ^ n38851 ;
  assign n40469 = n40467 & n40468 ;
  assign n40470 = n40469 ^ n37798 ;
  assign n40466 = n40202 ^ n40141 ;
  assign n40471 = n40470 ^ n40466 ;
  assign n40622 = n40540 ^ n40471 ;
  assign n40624 = n40622 ^ n37842 ;
  assign n40618 = n40617 ^ n40582 ;
  assign n40619 = n40617 ^ n37849 ;
  assign n40620 = ~n40618 & n40619 ;
  assign n40621 = n40620 ^ n37849 ;
  assign n40679 = n40624 ^ n40621 ;
  assign n40680 = n40678 & ~n40679 ;
  assign n40623 = n40622 ^ n40621 ;
  assign n40625 = ~n40623 & n40624 ;
  assign n40626 = n40625 ^ n37842 ;
  assign n40541 = n40540 ^ n40466 ;
  assign n40542 = ~n40471 & ~n40541 ;
  assign n40543 = n40542 ^ n40470 ;
  assign n40461 = n39067 ^ n38312 ;
  assign n40462 = n39423 ^ n39067 ;
  assign n40463 = n40461 & ~n40462 ;
  assign n40464 = n40463 ^ n38312 ;
  assign n40460 = n40204 ^ n40137 ;
  assign n40465 = n40464 ^ n40460 ;
  assign n40580 = n40543 ^ n40465 ;
  assign n40581 = n40580 ^ n37835 ;
  assign n40681 = n40626 ^ n40581 ;
  assign n40682 = ~n40680 & n40681 ;
  assign n40544 = n40543 ^ n40460 ;
  assign n40545 = n40465 & n40544 ;
  assign n40546 = n40545 ^ n40464 ;
  assign n40453 = n39421 ^ n39356 ;
  assign n40454 = n40207 ^ n40135 ;
  assign n40455 = n40454 ^ n37788 ;
  assign n40456 = n40455 ^ n39421 ;
  assign n40457 = n40456 ^ n40454 ;
  assign n40458 = ~n40453 & n40457 ;
  assign n40459 = n40458 ^ n40455 ;
  assign n40579 = n40546 ^ n40459 ;
  assign n40683 = n40579 ^ n37825 ;
  assign n40627 = n40626 ^ n40580 ;
  assign n40628 = n40581 & ~n40627 ;
  assign n40629 = n40628 ^ n37835 ;
  assign n40684 = n40683 ^ n40629 ;
  assign n40685 = ~n40682 & ~n40684 ;
  assign n40552 = n39431 ^ n39414 ;
  assign n40550 = n40210 ^ n40133 ;
  assign n40553 = n40550 ^ n37786 ;
  assign n40554 = n40553 ^ n39414 ;
  assign n40555 = n40554 ^ n40550 ;
  assign n40556 = n40552 & ~n40555 ;
  assign n40557 = n40556 ^ n40553 ;
  assign n40547 = n40546 ^ n40454 ;
  assign n40548 = n40459 & ~n40547 ;
  assign n40549 = n40548 ^ n40454 ;
  assign n40634 = n40557 ^ n40549 ;
  assign n40636 = n40634 ^ n37820 ;
  assign n40630 = n40629 ^ n40579 ;
  assign n40631 = n40629 ^ n37825 ;
  assign n40632 = n40630 & ~n40631 ;
  assign n40633 = n40632 ^ n37825 ;
  assign n40661 = n40636 ^ n40633 ;
  assign n40870 = n40685 ^ n40661 ;
  assign n40871 = n40870 ^ n40869 ;
  assign n40875 = n40684 ^ n40682 ;
  assign n40872 = n38583 ^ n620 ;
  assign n40873 = n40872 ^ n34558 ;
  assign n40874 = n40873 ^ n28622 ;
  assign n40876 = n40875 ^ n40874 ;
  assign n40880 = n40681 ^ n40680 ;
  assign n40877 = n38589 ^ n29771 ;
  assign n40878 = n40877 ^ n34563 ;
  assign n40879 = n40878 ^ n1517 ;
  assign n40881 = n40880 ^ n40879 ;
  assign n40885 = n40679 ^ n40678 ;
  assign n40882 = n38593 ^ n29775 ;
  assign n40883 = n40882 ^ n34569 ;
  assign n40884 = n40883 ^ n28629 ;
  assign n40886 = n40885 ^ n40884 ;
  assign n40890 = n40677 ^ n40675 ;
  assign n40887 = n38599 ^ n29780 ;
  assign n40888 = n40887 ^ n34574 ;
  assign n40889 = n40888 ^ n28679 ;
  assign n40891 = n40890 ^ n40889 ;
  assign n40893 = n38604 ^ n29786 ;
  assign n40894 = n40893 ^ n34580 ;
  assign n40895 = n40894 ^ n28636 ;
  assign n40892 = n40674 ^ n40673 ;
  assign n40896 = n40895 ^ n40892 ;
  assign n40900 = n38608 ^ n29850 ;
  assign n40901 = n40900 ^ n34591 ;
  assign n40902 = n40901 ^ n28665 ;
  assign n40899 = n40672 ^ n40663 ;
  assign n40903 = n40902 ^ n40899 ;
  assign n40907 = n40671 ^ n40670 ;
  assign n40904 = n38614 ^ n29791 ;
  assign n40905 = n40904 ^ n34586 ;
  assign n40906 = n40905 ^ n2297 ;
  assign n40908 = n40907 ^ n40906 ;
  assign n40912 = n40669 ^ n40668 ;
  assign n40909 = n38620 ^ n29795 ;
  assign n40910 = n40909 ^ n2165 ;
  assign n40911 = n40910 ^ n28641 ;
  assign n40913 = n40912 ^ n40911 ;
  assign n40917 = n40667 ^ n40666 ;
  assign n40914 = n38624 ^ n29800 ;
  assign n40915 = n40914 ^ n34613 ;
  assign n40916 = n40915 ^ n2160 ;
  assign n40918 = n40917 ^ n40916 ;
  assign n40919 = n40665 ^ n40664 ;
  assign n2037 = n2036 ^ n2015 ;
  assign n2065 = n2064 ^ n2037 ;
  assign n2072 = n2071 ^ n2065 ;
  assign n40920 = n40919 ^ n2072 ;
  assign n40446 = n38632 ^ n29807 ;
  assign n40447 = n40446 ^ n34621 ;
  assign n40448 = n40447 ^ n2056 ;
  assign n40445 = n40444 ^ n40443 ;
  assign n40449 = n40448 ^ n40445 ;
  assign n40420 = n40419 ^ n40418 ;
  assign n3063 = n3062 ^ n3053 ;
  assign n3082 = n3081 ^ n3063 ;
  assign n3089 = n3088 ^ n3082 ;
  assign n40358 = n40357 ^ n3089 ;
  assign n40360 = n40359 ^ n40358 ;
  assign n40361 = n38644 ^ n29816 ;
  assign n40362 = n40361 ^ n34632 ;
  assign n40363 = n40362 ^ n3076 ;
  assign n40364 = n40363 ^ n40359 ;
  assign n40370 = n34054 ^ n3015 ;
  assign n40371 = n40370 ^ n2775 ;
  assign n40372 = n40371 ^ n28017 ;
  assign n40365 = n38993 ^ n2731 ;
  assign n40366 = n40365 ^ n35198 ;
  assign n40367 = n40366 ^ n3179 ;
  assign n40368 = n40345 ^ n36578 ;
  assign n40369 = n40367 & ~n40368 ;
  assign n40373 = n40372 ^ n40369 ;
  assign n40374 = n40348 ^ n40347 ;
  assign n40375 = n40374 ^ n40369 ;
  assign n40376 = n40373 & n40375 ;
  assign n40377 = n40376 ^ n40372 ;
  assign n40378 = n40377 ^ n40363 ;
  assign n40379 = n40364 & ~n40378 ;
  assign n40380 = n40379 ^ n40357 ;
  assign n40381 = ~n40360 & n40380 ;
  assign n40382 = n40381 ^ n3089 ;
  assign n40421 = n40420 ^ n40382 ;
  assign n40422 = n38636 ^ n1962 ;
  assign n40423 = n40422 ^ n34625 ;
  assign n40424 = n40423 ^ n28012 ;
  assign n40425 = n40424 ^ n40382 ;
  assign n40426 = ~n40421 & ~n40425 ;
  assign n40427 = n40426 ^ n40420 ;
  assign n40921 = n40445 ^ n40427 ;
  assign n40922 = n40449 & n40921 ;
  assign n40923 = n40922 ^ n40448 ;
  assign n40924 = n40923 ^ n2072 ;
  assign n40925 = n40920 & n40924 ;
  assign n40926 = n40925 ^ n2072 ;
  assign n40927 = n40926 ^ n40916 ;
  assign n40928 = ~n40918 & ~n40927 ;
  assign n40929 = n40928 ^ n40917 ;
  assign n40930 = n40929 ^ n40911 ;
  assign n40931 = ~n40913 & ~n40930 ;
  assign n40932 = n40931 ^ n40911 ;
  assign n40933 = n40932 ^ n40906 ;
  assign n40934 = n40908 & ~n40933 ;
  assign n40935 = n40934 ^ n40907 ;
  assign n40936 = n40935 ^ n40899 ;
  assign n40937 = ~n40903 & n40936 ;
  assign n40938 = n40937 ^ n40902 ;
  assign n40939 = n40938 ^ n40895 ;
  assign n40940 = ~n40896 & n40939 ;
  assign n40897 = n40895 ^ n40890 ;
  assign n40941 = n40940 ^ n40897 ;
  assign n40942 = n40891 & n40941 ;
  assign n40943 = n40942 ^ n40890 ;
  assign n40944 = n40943 ^ n40884 ;
  assign n40945 = n40886 & ~n40944 ;
  assign n40946 = n40945 ^ n40885 ;
  assign n40947 = n40946 ^ n40879 ;
  assign n40948 = ~n40881 & ~n40947 ;
  assign n40949 = n40948 ^ n40880 ;
  assign n40950 = n40949 ^ n40874 ;
  assign n40951 = ~n40876 & n40950 ;
  assign n40952 = n40951 ^ n40875 ;
  assign n40953 = n40952 ^ n40869 ;
  assign n40954 = ~n40871 & n40953 ;
  assign n40955 = n40954 ^ n40870 ;
  assign n40686 = n40661 & n40685 ;
  assign n40635 = n40634 ^ n40633 ;
  assign n40637 = ~n40635 & n40636 ;
  assign n40638 = n40637 ^ n37820 ;
  assign n40562 = n39424 ^ n39407 ;
  assign n40560 = n40213 ^ n40128 ;
  assign n40563 = n40560 ^ n38331 ;
  assign n40564 = n40563 ^ n39407 ;
  assign n40565 = n40564 ^ n40560 ;
  assign n40566 = n40562 & ~n40565 ;
  assign n40567 = n40566 ^ n40563 ;
  assign n40551 = n40550 ^ n40549 ;
  assign n40558 = ~n40551 & ~n40557 ;
  assign n40559 = n40558 ^ n40550 ;
  assign n40577 = n40567 ^ n40559 ;
  assign n40578 = n40577 ^ n37813 ;
  assign n40660 = n40638 ^ n40578 ;
  assign n40865 = n40686 ^ n40660 ;
  assign n2979 = n2978 ^ n2975 ;
  assign n2980 = n2979 ^ n680 ;
  assign n2984 = n2983 ^ n2980 ;
  assign n40866 = n40865 ^ n2984 ;
  assign n41047 = n40955 ^ n40866 ;
  assign n40773 = n40233 ^ n40095 ;
  assign n42127 = n41047 ^ n40773 ;
  assign n42128 = n40773 ^ n39840 ;
  assign n42129 = ~n42127 & n42128 ;
  assign n42130 = n42129 ^ n39840 ;
  assign n41687 = n39261 ^ n30685 ;
  assign n41688 = n41687 ^ n35578 ;
  assign n41689 = n41688 ^ n28875 ;
  assign n41114 = n39437 ^ n38870 ;
  assign n41115 = n40454 ^ n39437 ;
  assign n41116 = n41114 & ~n41115 ;
  assign n41117 = n41116 ^ n38870 ;
  assign n40450 = n40449 ^ n40427 ;
  assign n41118 = n41117 ^ n40450 ;
  assign n41119 = n40460 ^ n39803 ;
  assign n41006 = n40424 ^ n40420 ;
  assign n41007 = n41006 ^ n40382 ;
  assign n41120 = n41007 ^ n38876 ;
  assign n41121 = n41120 ^ n40460 ;
  assign n41122 = n41121 ^ n41007 ;
  assign n41123 = ~n41119 & ~n41122 ;
  assign n41124 = n41123 ^ n41120 ;
  assign n41126 = n39793 ^ n38878 ;
  assign n41127 = n40466 ^ n39793 ;
  assign n41128 = ~n41126 & n41127 ;
  assign n41129 = n41128 ^ n38878 ;
  assign n41125 = n40380 ^ n3089 ;
  assign n41130 = n41129 ^ n41125 ;
  assign n41131 = n40451 ^ n38884 ;
  assign n41132 = n40377 ^ n40364 ;
  assign n41133 = n41132 ^ n39789 ;
  assign n41134 = n41133 ^ n40451 ;
  assign n41135 = n41134 ^ n41132 ;
  assign n41136 = ~n41131 & ~n41135 ;
  assign n41137 = n41136 ^ n41133 ;
  assign n41294 = n41132 ^ n41129 ;
  assign n41139 = n40478 ^ n39784 ;
  assign n41140 = n39784 ^ n38890 ;
  assign n41141 = ~n41139 & ~n41140 ;
  assign n41142 = n41141 ^ n38890 ;
  assign n41138 = n40374 ^ n40373 ;
  assign n41143 = n41142 ^ n41138 ;
  assign n41144 = n40488 ^ n39774 ;
  assign n41145 = n40368 ^ n40367 ;
  assign n41146 = n41145 ^ n38896 ;
  assign n41147 = n41146 ^ n40488 ;
  assign n41148 = n41147 ^ n41145 ;
  assign n41149 = ~n41144 & n41148 ;
  assign n41150 = n41149 ^ n41146 ;
  assign n41287 = n41145 ^ n41142 ;
  assign n41248 = n40522 ^ n39448 ;
  assign n41249 = n40522 ^ n38902 ;
  assign n41250 = ~n41248 & n41249 ;
  assign n41251 = n41250 ^ n38902 ;
  assign n41242 = n38949 ^ n2719 ;
  assign n41243 = n41242 ^ n3158 ;
  assign n41244 = n41243 ^ n28571 ;
  assign n41151 = n38812 ^ n30193 ;
  assign n41152 = n41151 ^ n35042 ;
  assign n41153 = n41152 ^ n3153 ;
  assign n41245 = n41244 ^ n41153 ;
  assign n41190 = n38935 ^ n37248 ;
  assign n41191 = n39662 ^ n37248 ;
  assign n41192 = ~n41190 & ~n41191 ;
  assign n41193 = n41192 ^ n38935 ;
  assign n41236 = n41193 ^ n37307 ;
  assign n41237 = n41236 ^ n38237 ;
  assign n41019 = n40254 ^ n40066 ;
  assign n41238 = n41237 ^ n41019 ;
  assign n41233 = n38932 ^ n38237 ;
  assign n41234 = n39721 ^ n38237 ;
  assign n41235 = n41233 & n41234 ;
  assign n41239 = n41238 ^ n41235 ;
  assign n41154 = n39669 ^ n39003 ;
  assign n41155 = n38969 ^ n38157 ;
  assign n41156 = n39677 ^ n38969 ;
  assign n41157 = n41155 & n41156 ;
  assign n41158 = n41157 ^ n38157 ;
  assign n41041 = n40245 ^ n40081 ;
  assign n41159 = n41158 ^ n41041 ;
  assign n40693 = n39403 ^ n39387 ;
  assign n40694 = n40222 ^ n40113 ;
  assign n40695 = n40694 ^ n38735 ;
  assign n40696 = n40695 ^ n39387 ;
  assign n40697 = n40696 ^ n40694 ;
  assign n40698 = ~n40693 & n40697 ;
  assign n40699 = n40698 ^ n40695 ;
  assign n40711 = n40225 ^ n40108 ;
  assign n40712 = n40711 ^ n40694 ;
  assign n40713 = n40712 ^ n40711 ;
  assign n40653 = n40220 ^ n40117 ;
  assign n40649 = n39840 ^ n39410 ;
  assign n40650 = n39410 ^ n38476 ;
  assign n40651 = n40649 & ~n40650 ;
  assign n40652 = n40651 ^ n38476 ;
  assign n40654 = n40653 ^ n40652 ;
  assign n40571 = n39416 ^ n39396 ;
  assign n40572 = n39416 ^ n38336 ;
  assign n40573 = n40571 & n40572 ;
  assign n40574 = n40573 ^ n38336 ;
  assign n40570 = n40216 ^ n40123 ;
  assign n40575 = n40574 ^ n40570 ;
  assign n40561 = n40560 ^ n40559 ;
  assign n40568 = n40561 & ~n40567 ;
  assign n40569 = n40568 ^ n40560 ;
  assign n40646 = n40570 ^ n40569 ;
  assign n40647 = n40575 & ~n40646 ;
  assign n40648 = n40647 ^ n40574 ;
  assign n40690 = n40652 ^ n40648 ;
  assign n40691 = n40654 & n40690 ;
  assign n40692 = n40691 ^ n40653 ;
  assign n40714 = n40713 ^ n40692 ;
  assign n40715 = ~n40699 & n40714 ;
  assign n40716 = n40715 ^ n40712 ;
  assign n40729 = n40228 ^ n40103 ;
  assign n40731 = n40729 ^ n40711 ;
  assign n40717 = n39394 ^ n38777 ;
  assign n40718 = n39394 ^ n39385 ;
  assign n40719 = n40717 & n40718 ;
  assign n40720 = n40719 ^ n38777 ;
  assign n40730 = n40729 ^ n40720 ;
  assign n40732 = n40731 ^ n40730 ;
  assign n40733 = ~n40716 & ~n40732 ;
  assign n40734 = n40733 ^ n40731 ;
  assign n40747 = n39389 ^ n38951 ;
  assign n40748 = n39853 ^ n39389 ;
  assign n40749 = n40747 & n40748 ;
  assign n40750 = n40749 ^ n38951 ;
  assign n40752 = n40750 ^ n40729 ;
  assign n40735 = n39484 ^ n38817 ;
  assign n40736 = n39484 ^ n39368 ;
  assign n40737 = ~n40735 & n40736 ;
  assign n40738 = n40737 ^ n38817 ;
  assign n40751 = n40750 ^ n40738 ;
  assign n40753 = n40752 ^ n40751 ;
  assign n40754 = n40734 & n40753 ;
  assign n40755 = n40754 ^ n40752 ;
  assign n40764 = n39381 ^ n38986 ;
  assign n40765 = n40274 ^ n39381 ;
  assign n40766 = n40764 & n40765 ;
  assign n40767 = n40766 ^ n38986 ;
  assign n40769 = n40767 ^ n40750 ;
  assign n40756 = n40231 ^ n1616 ;
  assign n40768 = n40767 ^ n40756 ;
  assign n40770 = n40769 ^ n40768 ;
  assign n40771 = n40755 & n40770 ;
  assign n40772 = n40771 ^ n40769 ;
  assign n40778 = n38748 ^ n38167 ;
  assign n40779 = n40323 ^ n38748 ;
  assign n40780 = ~n40778 & n40779 ;
  assign n40781 = n40780 ^ n38167 ;
  assign n40783 = n40781 ^ n40767 ;
  assign n40782 = n40781 ^ n40773 ;
  assign n40784 = n40783 ^ n40782 ;
  assign n40785 = ~n40772 & n40784 ;
  assign n40786 = n40785 ^ n40783 ;
  assign n40799 = n38783 ^ n38166 ;
  assign n40800 = n40401 ^ n38783 ;
  assign n40801 = n40799 & n40800 ;
  assign n40802 = n40801 ^ n38166 ;
  assign n40804 = n40802 ^ n40781 ;
  assign n40787 = n40237 ^ n957 ;
  assign n40803 = n40802 ^ n40787 ;
  assign n40805 = n40804 ^ n40803 ;
  assign n40806 = n40786 & n40805 ;
  assign n40807 = n40806 ^ n40804 ;
  assign n40820 = n38832 ^ n38160 ;
  assign n40821 = n39678 ^ n38832 ;
  assign n40822 = ~n40820 & n40821 ;
  assign n40823 = n40822 ^ n38160 ;
  assign n40825 = n40823 ^ n40802 ;
  assign n40808 = n40239 ^ n40088 ;
  assign n40824 = n40823 ^ n40808 ;
  assign n40826 = n40825 ^ n40824 ;
  assign n40827 = ~n40807 & ~n40826 ;
  assign n40828 = n40827 ^ n40825 ;
  assign n40829 = n40242 ^ n40083 ;
  assign n41161 = n40829 ^ n40823 ;
  assign n41162 = n40828 & n41161 ;
  assign n41160 = n41158 ^ n40823 ;
  assign n41163 = n41162 ^ n41160 ;
  assign n41164 = ~n41159 & ~n41163 ;
  assign n41165 = n41164 ^ n41158 ;
  assign n41166 = n41165 ^ n38213 ;
  assign n41167 = n41166 ^ n39669 ;
  assign n41168 = n41167 ^ n41165 ;
  assign n41169 = ~n41154 & n41168 ;
  assign n41170 = n41169 ^ n41166 ;
  assign n41035 = n40248 ^ n40076 ;
  assign n41194 = n41193 ^ n41035 ;
  assign n41195 = n41194 ^ n41165 ;
  assign n41196 = n41195 ^ n41193 ;
  assign n41197 = n41170 & ~n41196 ;
  assign n41198 = n41197 ^ n41194 ;
  assign n41025 = n40252 ^ n40070 ;
  assign n41231 = n41193 ^ n41025 ;
  assign n41232 = n41198 & n41231 ;
  assign n41240 = n41239 ^ n41232 ;
  assign n41199 = n41198 ^ n41025 ;
  assign n41176 = n41163 ^ n41041 ;
  assign n40830 = n40829 ^ n40828 ;
  assign n40831 = n40830 ^ n37429 ;
  assign n40809 = n40808 ^ n40807 ;
  assign n40810 = n40809 ^ n37418 ;
  assign n40774 = n40773 ^ n40772 ;
  assign n40775 = n40774 ^ n38195 ;
  assign n40757 = n40756 ^ n40755 ;
  assign n40739 = n40738 ^ n40734 ;
  assign n40721 = n40720 ^ n40716 ;
  assign n40722 = n40721 ^ n37257 ;
  assign n40655 = n40654 ^ n40648 ;
  assign n40656 = n40655 ^ n37805 ;
  assign n40639 = n40638 ^ n40577 ;
  assign n40640 = n40578 & n40639 ;
  assign n40641 = n40640 ^ n37813 ;
  assign n40576 = n40575 ^ n40569 ;
  assign n40642 = n40641 ^ n40576 ;
  assign n40643 = n40641 ^ n37796 ;
  assign n40644 = n40642 & ~n40643 ;
  assign n40645 = n40644 ^ n37796 ;
  assign n40702 = n40655 ^ n40645 ;
  assign n40703 = ~n40656 & ~n40702 ;
  assign n40704 = n40703 ^ n37805 ;
  assign n40700 = n40699 ^ n40692 ;
  assign n40707 = n40704 ^ n40700 ;
  assign n40708 = n40704 ^ n37791 ;
  assign n40709 = n40707 & n40708 ;
  assign n40710 = n40709 ^ n37791 ;
  assign n40725 = n40721 ^ n40710 ;
  assign n40726 = n40722 & n40725 ;
  assign n40727 = n40726 ^ n37257 ;
  assign n40742 = n40739 ^ n40727 ;
  assign n40743 = n40739 ^ n37252 ;
  assign n40744 = ~n40742 & ~n40743 ;
  assign n40745 = n40744 ^ n37252 ;
  assign n40760 = n40757 ^ n40745 ;
  assign n40761 = n40757 ^ n38147 ;
  assign n40762 = n40760 & n40761 ;
  assign n40763 = n40762 ^ n38147 ;
  assign n40790 = n40774 ^ n40763 ;
  assign n40791 = n40775 & ~n40790 ;
  assign n40792 = n40791 ^ n38195 ;
  assign n40788 = n40787 ^ n40786 ;
  assign n40795 = n40792 ^ n40788 ;
  assign n40796 = n40792 ^ n37242 ;
  assign n40797 = n40795 & ~n40796 ;
  assign n40798 = n40797 ^ n37242 ;
  assign n40817 = n40809 ^ n40798 ;
  assign n40818 = n40810 & n40817 ;
  assign n40819 = n40818 ^ n37418 ;
  assign n41173 = n40830 ^ n40819 ;
  assign n41174 = ~n40831 & ~n41173 ;
  assign n41175 = n41174 ^ n37429 ;
  assign n41177 = n41176 ^ n41175 ;
  assign n41178 = n41176 ^ n37411 ;
  assign n41179 = ~n41177 & ~n41178 ;
  assign n41180 = n41179 ^ n37411 ;
  assign n41171 = n41170 ^ n41035 ;
  assign n41172 = n41171 ^ n37406 ;
  assign n41181 = n41180 ^ n41172 ;
  assign n41182 = n41178 ^ n41175 ;
  assign n40832 = n40831 ^ n40819 ;
  assign n40657 = n40656 ^ n40645 ;
  assign n40658 = n40576 ^ n37796 ;
  assign n40659 = n40658 ^ n40641 ;
  assign n40687 = n40660 & n40686 ;
  assign n40688 = n40659 & ~n40687 ;
  assign n40689 = ~n40657 & ~n40688 ;
  assign n40701 = n40700 ^ n37791 ;
  assign n40705 = n40704 ^ n40701 ;
  assign n40706 = n40689 & n40705 ;
  assign n40723 = n40722 ^ n40710 ;
  assign n40724 = ~n40706 & n40723 ;
  assign n40728 = n40727 ^ n37252 ;
  assign n40740 = n40739 ^ n40728 ;
  assign n40741 = n40724 & n40740 ;
  assign n40746 = n40745 ^ n38147 ;
  assign n40758 = n40757 ^ n40746 ;
  assign n40759 = n40741 & n40758 ;
  assign n40776 = n40775 ^ n40763 ;
  assign n40777 = ~n40759 & n40776 ;
  assign n40789 = n40788 ^ n37242 ;
  assign n40793 = n40792 ^ n40789 ;
  assign n40794 = n40777 & n40793 ;
  assign n40811 = n40810 ^ n40798 ;
  assign n40833 = n40794 & ~n40811 ;
  assign n41183 = ~n40832 & n40833 ;
  assign n41184 = ~n41182 & ~n41183 ;
  assign n41185 = ~n41181 & n41184 ;
  assign n41225 = n41199 ^ n41185 ;
  assign n41186 = n41180 ^ n41171 ;
  assign n41187 = n41180 ^ n37406 ;
  assign n41188 = n41186 & ~n41187 ;
  assign n41189 = n41188 ^ n37406 ;
  assign n41228 = n41189 ^ n41185 ;
  assign n41229 = n41225 & ~n41228 ;
  assign n41226 = n41225 ^ n41189 ;
  assign n41227 = ~n37309 & ~n41226 ;
  assign n41230 = n41229 ^ n41227 ;
  assign n41241 = n41240 ^ n41230 ;
  assign n41246 = n41245 ^ n41241 ;
  assign n41200 = n41199 ^ n37309 ;
  assign n41201 = n41200 ^ n41189 ;
  assign n41202 = n41201 ^ n41185 ;
  assign n41203 = n41202 ^ n41153 ;
  assign n41207 = n41184 ^ n41181 ;
  assign n41204 = n38763 ^ n3128 ;
  assign n41205 = n41204 ^ n35115 ;
  assign n41206 = n41205 ^ n28582 ;
  assign n41208 = n41207 ^ n41206 ;
  assign n41210 = n38746 ^ n30200 ;
  assign n41211 = n41210 ^ n35047 ;
  assign n41212 = n41211 ^ n28589 ;
  assign n41209 = n41183 ^ n41182 ;
  assign n41213 = n41212 ^ n41209 ;
  assign n40813 = n38544 ^ n30211 ;
  assign n40814 = n40813 ^ n35057 ;
  assign n40815 = n40814 ^ n28598 ;
  assign n40812 = n40811 ^ n40794 ;
  assign n40816 = n40815 ^ n40812 ;
  assign n40840 = n40793 ^ n40777 ;
  assign n40837 = n38548 ^ n30215 ;
  assign n40838 = n40837 ^ n1399 ;
  assign n40839 = n40838 ^ n2804 ;
  assign n40841 = n40840 ^ n40839 ;
  assign n40979 = n40840 ^ n1370 ;
  assign n40842 = n40776 ^ n40759 ;
  assign n40843 = n40842 ^ n1370 ;
  assign n40844 = n40758 ^ n40741 ;
  assign n1223 = n1183 ^ n1135 ;
  assign n1224 = n1223 ^ n1220 ;
  assign n1231 = n1230 ^ n1224 ;
  assign n40845 = n40844 ^ n1231 ;
  assign n1187 = n1168 ^ n1117 ;
  assign n1206 = n1205 ^ n1187 ;
  assign n1213 = n1212 ^ n1206 ;
  assign n40973 = n40844 ^ n1213 ;
  assign n40846 = n40740 ^ n40724 ;
  assign n40847 = n40846 ^ n1213 ;
  assign n40849 = n38559 ^ n1037 ;
  assign n40850 = n40849 ^ n1678 ;
  assign n40851 = n40850 ^ n1197 ;
  assign n40848 = n40723 ^ n40706 ;
  assign n40852 = n40851 ^ n40848 ;
  assign n40853 = n40705 ^ n40689 ;
  assign n1660 = n1653 ^ n1022 ;
  assign n1670 = n1669 ^ n1660 ;
  assign n1674 = n1673 ^ n1670 ;
  assign n40854 = n40853 ^ n1674 ;
  assign n40855 = n38566 ^ n1636 ;
  assign n40856 = n40855 ^ n34517 ;
  assign n40857 = n40856 ^ n1666 ;
  assign n40964 = n40857 ^ n40853 ;
  assign n40858 = n40688 ^ n40657 ;
  assign n40859 = n40858 ^ n40857 ;
  assign n40863 = n40687 ^ n40659 ;
  assign n40860 = n38571 ^ n1627 ;
  assign n40861 = n40860 ^ n34522 ;
  assign n40862 = n40861 ^ n743 ;
  assign n40864 = n40863 ^ n40862 ;
  assign n40958 = n40863 ^ n2984 ;
  assign n40956 = n40955 ^ n2984 ;
  assign n40957 = ~n40866 & ~n40956 ;
  assign n40959 = n40958 ^ n40957 ;
  assign n40960 = ~n40864 & ~n40959 ;
  assign n40961 = n40960 ^ n40863 ;
  assign n40962 = n40961 ^ n40857 ;
  assign n40963 = ~n40859 & ~n40962 ;
  assign n40965 = n40964 ^ n40963 ;
  assign n40966 = ~n40854 & ~n40965 ;
  assign n40967 = n40966 ^ n40853 ;
  assign n40968 = n40967 ^ n40848 ;
  assign n40969 = ~n40852 & ~n40968 ;
  assign n40970 = n40969 ^ n40851 ;
  assign n40971 = n40970 ^ n1213 ;
  assign n40972 = n40847 & n40971 ;
  assign n40974 = n40973 ^ n40972 ;
  assign n40975 = n40845 & n40974 ;
  assign n40976 = n40975 ^ n40844 ;
  assign n40977 = n40976 ^ n1370 ;
  assign n40978 = n40843 & n40977 ;
  assign n40980 = n40979 ^ n40978 ;
  assign n40981 = ~n40841 & ~n40980 ;
  assign n40982 = n40981 ^ n40840 ;
  assign n40834 = n40833 ^ n40832 ;
  assign n40835 = n40834 ^ n40815 ;
  assign n40836 = n40835 ^ n40834 ;
  assign n40983 = n40982 ^ n40836 ;
  assign n40984 = n40816 & ~n40983 ;
  assign n40985 = n40984 ^ n40835 ;
  assign n40986 = n38539 ^ n30206 ;
  assign n40987 = n40986 ^ n35051 ;
  assign n40988 = n40987 ^ n2648 ;
  assign n41214 = n40988 ^ n40834 ;
  assign n41215 = ~n40985 & n41214 ;
  assign n41216 = n41215 ^ n40988 ;
  assign n41217 = n41216 ^ n41209 ;
  assign n41218 = n41213 & ~n41217 ;
  assign n41219 = n41218 ^ n41212 ;
  assign n41220 = n41219 ^ n41206 ;
  assign n41221 = ~n41208 & ~n41220 ;
  assign n41222 = n41221 ^ n41207 ;
  assign n41223 = n41222 ^ n41153 ;
  assign n41224 = ~n41203 & ~n41223 ;
  assign n41247 = n41246 ^ n41224 ;
  assign n41252 = n41251 ^ n41247 ;
  assign n41257 = n41222 ^ n41203 ;
  assign n41253 = n40494 ^ n39451 ;
  assign n41254 = n39451 ^ n38908 ;
  assign n41255 = ~n41253 & ~n41254 ;
  assign n41256 = n41255 ^ n38908 ;
  assign n41258 = n41257 ^ n41256 ;
  assign n41270 = n41219 ^ n41208 ;
  assign n41279 = n41270 ^ n41256 ;
  assign n41260 = n41216 ^ n41213 ;
  assign n40989 = n40988 ^ n40985 ;
  assign n40990 = n40432 ^ n38840 ;
  assign n40991 = n40432 ^ n38922 ;
  assign n40992 = ~n40990 & n40991 ;
  assign n40993 = n40992 ^ n38922 ;
  assign n41259 = n40989 & ~n40993 ;
  assign n41261 = n41260 ^ n41259 ;
  assign n41262 = n40509 ^ n39465 ;
  assign n41263 = n41259 ^ n38915 ;
  assign n41264 = n41263 ^ n40509 ;
  assign n41265 = n41264 ^ n41259 ;
  assign n41266 = ~n41262 & n41265 ;
  assign n41267 = n41266 ^ n41263 ;
  assign n41268 = n41261 & n41267 ;
  assign n41269 = n41268 ^ n41260 ;
  assign n41271 = n41270 ^ n41269 ;
  assign n41272 = n40514 ^ n39459 ;
  assign n41273 = n41270 ^ n38841 ;
  assign n41274 = n41273 ^ n39459 ;
  assign n41275 = n41274 ^ n41270 ;
  assign n41276 = n41272 & ~n41275 ;
  assign n41277 = n41276 ^ n41273 ;
  assign n41278 = ~n41271 & ~n41277 ;
  assign n41280 = n41279 ^ n41278 ;
  assign n41281 = n41258 & n41280 ;
  assign n41282 = n41281 ^ n41257 ;
  assign n41283 = n41282 ^ n41247 ;
  assign n41284 = ~n41252 & ~n41283 ;
  assign n41285 = n41284 ^ n41251 ;
  assign n41286 = n41285 ^ n41142 ;
  assign n41288 = n41287 ^ n41286 ;
  assign n41289 = ~n41150 & n41288 ;
  assign n41290 = n41289 ^ n41287 ;
  assign n41291 = n41143 & n41290 ;
  assign n41292 = n41291 ^ n41142 ;
  assign n41293 = n41292 ^ n41129 ;
  assign n41295 = n41294 ^ n41293 ;
  assign n41296 = ~n41137 & ~n41295 ;
  assign n41297 = n41296 ^ n41293 ;
  assign n41298 = n41130 & n41297 ;
  assign n41299 = n41298 ^ n41129 ;
  assign n41300 = n41299 ^ n41007 ;
  assign n41301 = ~n41124 & n41300 ;
  assign n41302 = n41301 ^ n41007 ;
  assign n41303 = n41302 ^ n41117 ;
  assign n41304 = ~n41118 & n41303 ;
  assign n41305 = n41304 ^ n40450 ;
  assign n41112 = n40923 ^ n40920 ;
  assign n41108 = n40550 ^ n39430 ;
  assign n41109 = n39430 ^ n38860 ;
  assign n41110 = ~n41108 & n41109 ;
  assign n41111 = n41110 ^ n38860 ;
  assign n41113 = n41112 ^ n41111 ;
  assign n41409 = n41305 ^ n41113 ;
  assign n41410 = n41409 ^ n37818 ;
  assign n41457 = n41302 ^ n41118 ;
  assign n41411 = n41299 ^ n41124 ;
  assign n41412 = n41411 ^ n37833 ;
  assign n41413 = n41297 ^ n41125 ;
  assign n41414 = n41413 ^ n37840 ;
  assign n41416 = n41290 ^ n41138 ;
  assign n41417 = n41416 ^ n38280 ;
  assign n41418 = n41285 ^ n41150 ;
  assign n41419 = n41418 ^ n37854 ;
  assign n41436 = n41282 ^ n41252 ;
  assign n41420 = n41280 ^ n41257 ;
  assign n41421 = n41420 ^ n37873 ;
  assign n41428 = n41277 ^ n41269 ;
  assign n41423 = n41267 ^ n41260 ;
  assign n40994 = n40993 ^ n40989 ;
  assign n41422 = n38247 & ~n40994 ;
  assign n41424 = n41423 ^ n41422 ;
  assign n41425 = n41423 ^ n38262 ;
  assign n41426 = n41424 & ~n41425 ;
  assign n41427 = n41426 ^ n38262 ;
  assign n41429 = n41428 ^ n41427 ;
  assign n41430 = n41428 ^ n38268 ;
  assign n41431 = n41429 & ~n41430 ;
  assign n41432 = n41431 ^ n38268 ;
  assign n41433 = n41432 ^ n41420 ;
  assign n41434 = n41421 & n41433 ;
  assign n41435 = n41434 ^ n37873 ;
  assign n41437 = n41436 ^ n41435 ;
  assign n41438 = n41436 ^ n37861 ;
  assign n41439 = ~n41437 & ~n41438 ;
  assign n41440 = n41439 ^ n37861 ;
  assign n41441 = n41440 ^ n41418 ;
  assign n41442 = ~n41419 & ~n41441 ;
  assign n41443 = n41442 ^ n37854 ;
  assign n41444 = n41443 ^ n41416 ;
  assign n41445 = n41417 & ~n41444 ;
  assign n41446 = n41445 ^ n38280 ;
  assign n41415 = n41292 ^ n41137 ;
  assign n41447 = n41446 ^ n41415 ;
  assign n41448 = n41446 ^ n37847 ;
  assign n41449 = ~n41447 & n41448 ;
  assign n41450 = n41449 ^ n37847 ;
  assign n41451 = n41450 ^ n41413 ;
  assign n41452 = ~n41414 & ~n41451 ;
  assign n41453 = n41452 ^ n37840 ;
  assign n41454 = n41453 ^ n41411 ;
  assign n41455 = n41412 & ~n41454 ;
  assign n41456 = n41455 ^ n37833 ;
  assign n41458 = n41457 ^ n41456 ;
  assign n41459 = n41457 ^ n37827 ;
  assign n41460 = ~n41458 & ~n41459 ;
  assign n41461 = n41460 ^ n37827 ;
  assign n41462 = n41461 ^ n41409 ;
  assign n41463 = n41410 & n41462 ;
  assign n41464 = n41463 ^ n37818 ;
  assign n41306 = n41305 ^ n41111 ;
  assign n41307 = ~n41113 & ~n41306 ;
  assign n41308 = n41307 ^ n41112 ;
  assign n41106 = n40926 ^ n40918 ;
  assign n41102 = n40560 ^ n39423 ;
  assign n41103 = n39423 ^ n38857 ;
  assign n41104 = ~n41102 & n41103 ;
  assign n41105 = n41104 ^ n38857 ;
  assign n41107 = n41106 ^ n41105 ;
  assign n41407 = n41308 ^ n41107 ;
  assign n41408 = n41407 ^ n37811 ;
  assign n41548 = n41464 ^ n41408 ;
  assign n41528 = n41461 ^ n41410 ;
  assign n41529 = n41459 ^ n41456 ;
  assign n41530 = n41415 ^ n37847 ;
  assign n41531 = n41530 ^ n41446 ;
  assign n41532 = n41443 ^ n41417 ;
  assign n41533 = n41440 ^ n41419 ;
  assign n41534 = n41430 ^ n41427 ;
  assign n41535 = n41432 ^ n41421 ;
  assign n41536 = n41534 & ~n41535 ;
  assign n41537 = n41438 ^ n41435 ;
  assign n41538 = n41536 & ~n41537 ;
  assign n41539 = ~n41533 & ~n41538 ;
  assign n41540 = n41532 & ~n41539 ;
  assign n41541 = n41531 & n41540 ;
  assign n41542 = n41450 ^ n41414 ;
  assign n41543 = ~n41541 & n41542 ;
  assign n41544 = n41453 ^ n41412 ;
  assign n41545 = n41543 & n41544 ;
  assign n41546 = n41529 & ~n41545 ;
  assign n41547 = n41528 & n41546 ;
  assign n41681 = n41548 ^ n41547 ;
  assign n41768 = n41689 ^ n41681 ;
  assign n41686 = n41546 ^ n41528 ;
  assign n41690 = n41689 ^ n41686 ;
  assign n41691 = n41545 ^ n41529 ;
  assign n2379 = n2378 ^ n2315 ;
  assign n2392 = n2391 ^ n2379 ;
  assign n2396 = n2395 ^ n2392 ;
  assign n41692 = n41691 ^ n2396 ;
  assign n41696 = n41544 ^ n41543 ;
  assign n41693 = n39268 ^ n30695 ;
  assign n41694 = n41693 ^ n2278 ;
  assign n41695 = n41694 ^ n2386 ;
  assign n41697 = n41696 ^ n41695 ;
  assign n41698 = n41542 ^ n41541 ;
  assign n2236 = n2229 ^ n2193 ;
  assign n2261 = n2260 ^ n2236 ;
  assign n2268 = n2267 ^ n2261 ;
  assign n41699 = n41698 ^ n2268 ;
  assign n41748 = n41540 ^ n41531 ;
  assign n41703 = n41539 ^ n41532 ;
  assign n41700 = n39279 ^ n2116 ;
  assign n41701 = n41700 ^ n35594 ;
  assign n41702 = n41701 ^ n28890 ;
  assign n41704 = n41703 ^ n41702 ;
  assign n41706 = n39296 ^ n30705 ;
  assign n41707 = n41706 ^ n35624 ;
  assign n41708 = n41707 ^ n28894 ;
  assign n41705 = n41538 ^ n41533 ;
  assign n41709 = n41708 ^ n41705 ;
  assign n41734 = n41537 ^ n41536 ;
  assign n41710 = n38797 ^ n30714 ;
  assign n41711 = n41710 ^ n35612 ;
  assign n41712 = n41711 ^ n28915 ;
  assign n41713 = n41712 ^ n41535 ;
  assign n41714 = n41713 ^ n41534 ;
  assign n41715 = n38754 ^ n35599 ;
  assign n41716 = n41715 ^ n30718 ;
  assign n41717 = n41716 ^ n1868 ;
  assign n41718 = n41717 ^ n41534 ;
  assign n40995 = n40994 ^ n38247 ;
  assign n40996 = n39714 ^ n31059 ;
  assign n40997 = n40996 ^ n35958 ;
  assign n40998 = n40997 ^ n3233 ;
  assign n41722 = ~n40995 & n40998 ;
  assign n41719 = n30721 ^ n3194 ;
  assign n41720 = n41719 ^ n35604 ;
  assign n41721 = n41720 ^ n28904 ;
  assign n41723 = n41722 ^ n41721 ;
  assign n41724 = n41422 ^ n38262 ;
  assign n41725 = n41724 ^ n41423 ;
  assign n41726 = n41725 ^ n41721 ;
  assign n41727 = n41723 & n41726 ;
  assign n41728 = n41727 ^ n41722 ;
  assign n41729 = n41728 ^ n41717 ;
  assign n41730 = n41718 & ~n41729 ;
  assign n41731 = n41730 ^ n41535 ;
  assign n41732 = n41714 & ~n41731 ;
  assign n41733 = n41732 ^ n41712 ;
  assign n41735 = n41734 ^ n41733 ;
  assign n41736 = n39284 ^ n30709 ;
  assign n41737 = n41736 ^ n35616 ;
  assign n41738 = n41737 ^ n28899 ;
  assign n41739 = n41738 ^ n41733 ;
  assign n41740 = n41735 & ~n41739 ;
  assign n41741 = n41740 ^ n41734 ;
  assign n41742 = n41741 ^ n41705 ;
  assign n41743 = n41709 & ~n41742 ;
  assign n41744 = n41743 ^ n41708 ;
  assign n41745 = n41744 ^ n41702 ;
  assign n41746 = n41704 & n41745 ;
  assign n41747 = n41746 ^ n41702 ;
  assign n41749 = n41748 ^ n41747 ;
  assign n41750 = n39274 ^ n2131 ;
  assign n41751 = n41750 ^ n35590 ;
  assign n41752 = n41751 ^ n2252 ;
  assign n41753 = n41752 ^ n41698 ;
  assign n41754 = n41753 ^ n41747 ;
  assign n41755 = n41754 ^ n41698 ;
  assign n41756 = n41749 & n41755 ;
  assign n41757 = n41756 ^ n41753 ;
  assign n41758 = ~n41699 & ~n41757 ;
  assign n41759 = n41758 ^ n41698 ;
  assign n41760 = n41759 ^ n41695 ;
  assign n41761 = n41697 & n41760 ;
  assign n41762 = n41761 ^ n41696 ;
  assign n41763 = n41762 ^ n2396 ;
  assign n41764 = n41692 & ~n41763 ;
  assign n41765 = n41764 ^ n41691 ;
  assign n41766 = n41765 ^ n41689 ;
  assign n41767 = ~n41690 & n41766 ;
  assign n41769 = n41768 ^ n41767 ;
  assign n41682 = n39255 ^ n30679 ;
  assign n41683 = n41682 ^ n35573 ;
  assign n41684 = n41683 ^ n28963 ;
  assign n42038 = n41769 ^ n41684 ;
  assign n42131 = n42130 ^ n42038 ;
  assign n41057 = n40952 ^ n40871 ;
  assign n42133 = n41057 ^ n40756 ;
  assign n42134 = n40756 ^ n39396 ;
  assign n42135 = n42133 & ~n42134 ;
  assign n42136 = n42135 ^ n39396 ;
  assign n42132 = n41765 ^ n41690 ;
  assign n42137 = n42136 ^ n42132 ;
  assign n41063 = n40949 ^ n40876 ;
  assign n42198 = n41063 ^ n40729 ;
  assign n42199 = n40729 ^ n39407 ;
  assign n42200 = n42198 & n42199 ;
  assign n42201 = n42200 ^ n39407 ;
  assign n42139 = n40711 ^ n39414 ;
  assign n41069 = n40946 ^ n40881 ;
  assign n42140 = n41069 ^ n40711 ;
  assign n42141 = n42139 & ~n42140 ;
  assign n42142 = n42141 ^ n39414 ;
  assign n42138 = n41759 ^ n41697 ;
  assign n42143 = n42142 ^ n42138 ;
  assign n41324 = n40941 ^ n40889 ;
  assign n42144 = n41324 ^ n40653 ;
  assign n42043 = n41752 ^ n41748 ;
  assign n42044 = n42043 ^ n41747 ;
  assign n42145 = n42044 ^ n39423 ;
  assign n42146 = n42145 ^ n40653 ;
  assign n42147 = n42146 ^ n42044 ;
  assign n42148 = ~n42144 & ~n42147 ;
  assign n42149 = n42148 ^ n42145 ;
  assign n41078 = n40938 ^ n40896 ;
  assign n42156 = n41078 ^ n40570 ;
  assign n42157 = n40570 ^ n39430 ;
  assign n42158 = ~n42156 & n42157 ;
  assign n42159 = n42158 ^ n39430 ;
  assign n42060 = n41744 ^ n41704 ;
  assign n42160 = n42159 ^ n42060 ;
  assign n42166 = n41741 ^ n41709 ;
  assign n41088 = n40935 ^ n40903 ;
  assign n42161 = n41088 ^ n40560 ;
  assign n42162 = n40560 ^ n39437 ;
  assign n42163 = ~n42161 & ~n42162 ;
  assign n42164 = n42163 ^ n39437 ;
  assign n42167 = n42166 ^ n42164 ;
  assign n41930 = n41106 ^ n40460 ;
  assign n41931 = n41728 ^ n41718 ;
  assign n41932 = n41931 ^ n39789 ;
  assign n41933 = n41932 ^ n41106 ;
  assign n41934 = n41933 ^ n41931 ;
  assign n41935 = ~n41930 & ~n41934 ;
  assign n41936 = n41935 ^ n41932 ;
  assign n41096 = n40929 ^ n40913 ;
  assign n42007 = n41096 ^ n40454 ;
  assign n42008 = n40454 ^ n39793 ;
  assign n42009 = ~n42007 & n42008 ;
  assign n42010 = n42009 ^ n39793 ;
  assign n42011 = n42010 ^ n41931 ;
  assign n42012 = n42011 ^ n42010 ;
  assign n41887 = n41112 ^ n40466 ;
  assign n41888 = n40466 ^ n39784 ;
  assign n41889 = n41887 & ~n41888 ;
  assign n41890 = n41889 ^ n39784 ;
  assign n40999 = n40998 ^ n40995 ;
  assign n41891 = n41890 ^ n40999 ;
  assign n40452 = n40451 ^ n40450 ;
  assign n41000 = n40999 ^ n39774 ;
  assign n41001 = n41000 ^ n40450 ;
  assign n41002 = n41001 ^ n40999 ;
  assign n41003 = ~n40452 & ~n41002 ;
  assign n41004 = n41003 ^ n41000 ;
  assign n41602 = n39593 ^ n30900 ;
  assign n41603 = n41602 ^ n2657 ;
  assign n41604 = n41603 ^ n3221 ;
  assign n41839 = n41838 ^ n41604 ;
  assign n41834 = n38237 ^ n37248 ;
  assign n41832 = n40982 ^ n40816 ;
  assign n41588 = n40980 ^ n40839 ;
  assign n41831 = n41588 ^ n38932 ;
  assign n41833 = n41832 ^ n41831 ;
  assign n41835 = n41834 ^ n41833 ;
  assign n41840 = n41839 ^ n41835 ;
  assign n41011 = n40298 ^ n39662 ;
  assign n41016 = n40970 ^ n40847 ;
  assign n41012 = n39669 ^ n38832 ;
  assign n41013 = n40296 ^ n39669 ;
  assign n41014 = ~n41012 & n41013 ;
  assign n41015 = n41014 ^ n38832 ;
  assign n41017 = n41016 ^ n41015 ;
  assign n41023 = n40967 ^ n40852 ;
  assign n41018 = n39677 ^ n38783 ;
  assign n41020 = n41019 ^ n39677 ;
  assign n41021 = n41018 & ~n41020 ;
  assign n41022 = n41021 ^ n38783 ;
  assign n41024 = n41023 ^ n41022 ;
  assign n41026 = n41025 ^ n39678 ;
  assign n41027 = n40965 ^ n1674 ;
  assign n41028 = n41027 ^ n38748 ;
  assign n41029 = n41028 ^ n41025 ;
  assign n41030 = n41029 ^ n41027 ;
  assign n41031 = ~n41026 & n41030 ;
  assign n41032 = n41031 ^ n41028 ;
  assign n41034 = n40401 ^ n39381 ;
  assign n41036 = n41035 ^ n40401 ;
  assign n41037 = n41034 & n41036 ;
  assign n41038 = n41037 ^ n39381 ;
  assign n41033 = n40961 ^ n40859 ;
  assign n41039 = n41038 ^ n41033 ;
  assign n41042 = n41041 ^ n40323 ;
  assign n41043 = n40323 ^ n39389 ;
  assign n41044 = n41042 & ~n41043 ;
  assign n41045 = n41044 ^ n39389 ;
  assign n41351 = n41045 ^ n41038 ;
  assign n41040 = n40959 ^ n40862 ;
  assign n41046 = n41045 ^ n41040 ;
  assign n41048 = n40274 ^ n39484 ;
  assign n41049 = n40829 ^ n40274 ;
  assign n41050 = ~n41048 & ~n41049 ;
  assign n41051 = n41050 ^ n39484 ;
  assign n41052 = n41051 ^ n41047 ;
  assign n41053 = n39853 ^ n39394 ;
  assign n41054 = n40808 ^ n39853 ;
  assign n41055 = n41053 & ~n41054 ;
  assign n41056 = n41055 ^ n39394 ;
  assign n41058 = n41057 ^ n41056 ;
  assign n41059 = n39403 ^ n39368 ;
  assign n41060 = n40787 ^ n39368 ;
  assign n41061 = n41059 & n41060 ;
  assign n41062 = n41061 ^ n39403 ;
  assign n41064 = n41063 ^ n41062 ;
  assign n41065 = n39410 ^ n39385 ;
  assign n41066 = n40773 ^ n39385 ;
  assign n41067 = n41065 & n41066 ;
  assign n41068 = n41067 ^ n39410 ;
  assign n41070 = n41069 ^ n41068 ;
  assign n41075 = n40943 ^ n40886 ;
  assign n41071 = n39416 ^ n39387 ;
  assign n41072 = n40756 ^ n39387 ;
  assign n41073 = n41071 & ~n41072 ;
  assign n41074 = n41073 ^ n39416 ;
  assign n41076 = n41075 ^ n41074 ;
  assign n41077 = n40711 ^ n39396 ;
  assign n41079 = n41078 ^ n39431 ;
  assign n41080 = n41079 ^ n40711 ;
  assign n41081 = n41080 ^ n41078 ;
  assign n41082 = n41077 & ~n41081 ;
  assign n41083 = n41082 ^ n41079 ;
  assign n41084 = n39407 ^ n39356 ;
  assign n41085 = n40694 ^ n39407 ;
  assign n41086 = ~n41084 & n41085 ;
  assign n41087 = n41086 ^ n39356 ;
  assign n41089 = n41088 ^ n41087 ;
  assign n41091 = n40653 ^ n39414 ;
  assign n41092 = n39414 ^ n39067 ;
  assign n41093 = n41091 & n41092 ;
  assign n41094 = n41093 ^ n39067 ;
  assign n41090 = n40932 ^ n40908 ;
  assign n41095 = n41094 ^ n41090 ;
  assign n41097 = n40570 ^ n39421 ;
  assign n41098 = n39421 ^ n38851 ;
  assign n41099 = n41097 & n41098 ;
  assign n41100 = n41099 ^ n38851 ;
  assign n41101 = n41100 ^ n41096 ;
  assign n41309 = n41308 ^ n41105 ;
  assign n41310 = n41107 & n41309 ;
  assign n41311 = n41310 ^ n41106 ;
  assign n41312 = n41311 ^ n41096 ;
  assign n41313 = n41101 & n41312 ;
  assign n41314 = n41313 ^ n41100 ;
  assign n41315 = n41314 ^ n41090 ;
  assign n41316 = ~n41095 & ~n41315 ;
  assign n41317 = n41316 ^ n41094 ;
  assign n41318 = n41317 ^ n41087 ;
  assign n41319 = ~n41089 & n41318 ;
  assign n41320 = n41319 ^ n41088 ;
  assign n41321 = n41320 ^ n41078 ;
  assign n41322 = ~n41083 & n41321 ;
  assign n41323 = n41322 ^ n41078 ;
  assign n41325 = n41324 ^ n41323 ;
  assign n41326 = n40729 ^ n39840 ;
  assign n41327 = n41324 ^ n39424 ;
  assign n41328 = n41327 ^ n41324 ;
  assign n41329 = n41328 ^ n40729 ;
  assign n41330 = n41326 & ~n41329 ;
  assign n41331 = n41330 ^ n41327 ;
  assign n41332 = ~n41325 & n41331 ;
  assign n41333 = n41332 ^ n41324 ;
  assign n41334 = n41333 ^ n41074 ;
  assign n41335 = ~n41076 & n41334 ;
  assign n41336 = n41335 ^ n41075 ;
  assign n41337 = n41336 ^ n41068 ;
  assign n41338 = n41070 & n41337 ;
  assign n41339 = n41338 ^ n41069 ;
  assign n41340 = n41339 ^ n41062 ;
  assign n41341 = ~n41064 & ~n41340 ;
  assign n41342 = n41341 ^ n41063 ;
  assign n41343 = n41342 ^ n41056 ;
  assign n41344 = n41058 & ~n41343 ;
  assign n41345 = n41344 ^ n41057 ;
  assign n41346 = n41345 ^ n41047 ;
  assign n41347 = n41052 & ~n41346 ;
  assign n41348 = n41347 ^ n41051 ;
  assign n41349 = n41348 ^ n41040 ;
  assign n41350 = n41046 & n41349 ;
  assign n41352 = n41351 ^ n41350 ;
  assign n41353 = n41039 & ~n41352 ;
  assign n41354 = n41353 ^ n41038 ;
  assign n41355 = n41354 ^ n41027 ;
  assign n41356 = n41032 & ~n41355 ;
  assign n41357 = n41356 ^ n41027 ;
  assign n41358 = n41357 ^ n41022 ;
  assign n41359 = ~n41024 & ~n41358 ;
  assign n41360 = n41359 ^ n41023 ;
  assign n41361 = n41360 ^ n41015 ;
  assign n41362 = n41017 & ~n41361 ;
  assign n41363 = n41362 ^ n41016 ;
  assign n41364 = n41363 ^ n38969 ;
  assign n41365 = n41364 ^ n40298 ;
  assign n41366 = n41365 ^ n41363 ;
  assign n41367 = n41011 & ~n41366 ;
  assign n41368 = n41367 ^ n41364 ;
  assign n41374 = n40974 ^ n1231 ;
  assign n41369 = n39721 ^ n39003 ;
  assign n41370 = n40286 ^ n39721 ;
  assign n41371 = n41369 & ~n41370 ;
  assign n41372 = n41371 ^ n39003 ;
  assign n41375 = n41374 ^ n41372 ;
  assign n41373 = n41372 ^ n41363 ;
  assign n41376 = n41375 ^ n41373 ;
  assign n41377 = ~n41368 & n41376 ;
  assign n41378 = n41377 ^ n41375 ;
  assign n41590 = n41588 ^ n41372 ;
  assign n41379 = n40976 ^ n40843 ;
  assign n41589 = n41588 ^ n41379 ;
  assign n41591 = n41590 ^ n41589 ;
  assign n41592 = ~n41378 & ~n41591 ;
  assign n41593 = n41592 ^ n41590 ;
  assign n41594 = n39472 ^ n38935 ;
  assign n41595 = n40342 ^ n39472 ;
  assign n41596 = ~n41594 & n41595 ;
  assign n41597 = n41596 ^ n38935 ;
  assign n41829 = n41597 ^ n41588 ;
  assign n41830 = n41593 & n41829 ;
  assign n41841 = n41840 ^ n41830 ;
  assign n41598 = n41597 ^ n41593 ;
  assign n41599 = n41598 ^ n37248 ;
  assign n41382 = n41374 ^ n41368 ;
  assign n41383 = n41382 ^ n38157 ;
  assign n41385 = n41357 ^ n41024 ;
  assign n41386 = n41385 ^ n38166 ;
  assign n41387 = n41354 ^ n41032 ;
  assign n41388 = n41387 ^ n38167 ;
  assign n41390 = n41348 ^ n41046 ;
  assign n41391 = n41390 ^ n38951 ;
  assign n41393 = n41342 ^ n41058 ;
  assign n41394 = n41393 ^ n38777 ;
  assign n41395 = n41339 ^ n41064 ;
  assign n41396 = n41395 ^ n38735 ;
  assign n41398 = n41333 ^ n41076 ;
  assign n41399 = n41398 ^ n38336 ;
  assign n41477 = n41320 ^ n41083 ;
  assign n41401 = n41317 ^ n41089 ;
  assign n41402 = n41401 ^ n37788 ;
  assign n41403 = n41314 ^ n41095 ;
  assign n41404 = n41403 ^ n38312 ;
  assign n41405 = n41311 ^ n41101 ;
  assign n41406 = n41405 ^ n37798 ;
  assign n41465 = n41464 ^ n41407 ;
  assign n41466 = ~n41408 & ~n41465 ;
  assign n41467 = n41466 ^ n37811 ;
  assign n41468 = n41467 ^ n41405 ;
  assign n41469 = ~n41406 & ~n41468 ;
  assign n41470 = n41469 ^ n37798 ;
  assign n41471 = n41470 ^ n41403 ;
  assign n41472 = n41404 & n41471 ;
  assign n41473 = n41472 ^ n38312 ;
  assign n41474 = n41473 ^ n41401 ;
  assign n41475 = n41402 & n41474 ;
  assign n41476 = n41475 ^ n37788 ;
  assign n41478 = n41477 ^ n41476 ;
  assign n41479 = n41477 ^ n37786 ;
  assign n41480 = ~n41478 & n41479 ;
  assign n41481 = n41480 ^ n37786 ;
  assign n41400 = n41331 ^ n41323 ;
  assign n41482 = n41481 ^ n41400 ;
  assign n41483 = n41481 ^ n38331 ;
  assign n41484 = n41482 & n41483 ;
  assign n41485 = n41484 ^ n38331 ;
  assign n41486 = n41485 ^ n41398 ;
  assign n41487 = n41399 & n41486 ;
  assign n41488 = n41487 ^ n38336 ;
  assign n41397 = n41336 ^ n41070 ;
  assign n41489 = n41488 ^ n41397 ;
  assign n41490 = n41488 ^ n38476 ;
  assign n41491 = n41489 & ~n41490 ;
  assign n41492 = n41491 ^ n38476 ;
  assign n41493 = n41492 ^ n41395 ;
  assign n41494 = ~n41396 & ~n41493 ;
  assign n41495 = n41494 ^ n38735 ;
  assign n41496 = n41495 ^ n41393 ;
  assign n41497 = n41394 & n41496 ;
  assign n41498 = n41497 ^ n38777 ;
  assign n41392 = n41345 ^ n41052 ;
  assign n41499 = n41498 ^ n41392 ;
  assign n41500 = n41498 ^ n38817 ;
  assign n41501 = ~n41499 & ~n41500 ;
  assign n41502 = n41501 ^ n38817 ;
  assign n41503 = n41502 ^ n41390 ;
  assign n41504 = ~n41391 & n41503 ;
  assign n41505 = n41504 ^ n38951 ;
  assign n41389 = n41352 ^ n41033 ;
  assign n41506 = n41505 ^ n41389 ;
  assign n41507 = n41505 ^ n38986 ;
  assign n41508 = ~n41506 & ~n41507 ;
  assign n41509 = n41508 ^ n38986 ;
  assign n41510 = n41509 ^ n41387 ;
  assign n41511 = n41388 & ~n41510 ;
  assign n41512 = n41511 ^ n38167 ;
  assign n41513 = n41512 ^ n41385 ;
  assign n41514 = ~n41386 & ~n41513 ;
  assign n41515 = n41514 ^ n38166 ;
  assign n41384 = n41360 ^ n41017 ;
  assign n41516 = n41515 ^ n41384 ;
  assign n41517 = n41515 ^ n38160 ;
  assign n41518 = n41516 & n41517 ;
  assign n41519 = n41518 ^ n38160 ;
  assign n41520 = n41519 ^ n41382 ;
  assign n41521 = n41383 & n41520 ;
  assign n41522 = n41521 ^ n38157 ;
  assign n41380 = n41379 ^ n41378 ;
  assign n41584 = n41522 ^ n41380 ;
  assign n41585 = n41522 ^ n38213 ;
  assign n41586 = n41584 & ~n41585 ;
  assign n41587 = n41586 ^ n38213 ;
  assign n41827 = n41598 ^ n41587 ;
  assign n41828 = ~n41599 & ~n41827 ;
  assign n41842 = n41841 ^ n41828 ;
  assign n41824 = n39739 ^ n38932 ;
  assign n41825 = n40414 ^ n39739 ;
  assign n41826 = ~n41824 & n41825 ;
  assign n41843 = n41842 ^ n41826 ;
  assign n41381 = n41380 ^ n38213 ;
  assign n41523 = n41522 ^ n41381 ;
  assign n41524 = n41492 ^ n41396 ;
  assign n41525 = n41400 ^ n38331 ;
  assign n41526 = n41525 ^ n41481 ;
  assign n41527 = n41479 ^ n41476 ;
  assign n41549 = n41547 & n41548 ;
  assign n41550 = n41467 ^ n41406 ;
  assign n41551 = n41549 & ~n41550 ;
  assign n41552 = n41470 ^ n41404 ;
  assign n41553 = ~n41551 & n41552 ;
  assign n41554 = n41473 ^ n41402 ;
  assign n41555 = ~n41553 & n41554 ;
  assign n41556 = ~n41527 & n41555 ;
  assign n41557 = n41526 & n41556 ;
  assign n41558 = n41485 ^ n41399 ;
  assign n41559 = ~n41557 & n41558 ;
  assign n41560 = n41397 ^ n38476 ;
  assign n41561 = n41560 ^ n41488 ;
  assign n41562 = ~n41559 & n41561 ;
  assign n41563 = n41524 & n41562 ;
  assign n41564 = n41495 ^ n41394 ;
  assign n41565 = ~n41563 & ~n41564 ;
  assign n41566 = n41392 ^ n38817 ;
  assign n41567 = n41566 ^ n41498 ;
  assign n41568 = n41565 & ~n41567 ;
  assign n41569 = n41502 ^ n41391 ;
  assign n41570 = n41568 & n41569 ;
  assign n41571 = n41389 ^ n38986 ;
  assign n41572 = n41571 ^ n41505 ;
  assign n41573 = ~n41570 & ~n41572 ;
  assign n41574 = n41509 ^ n41388 ;
  assign n41575 = n41573 & ~n41574 ;
  assign n41576 = n41512 ^ n41386 ;
  assign n41577 = n41575 & n41576 ;
  assign n41578 = n41384 ^ n38160 ;
  assign n41579 = n41578 ^ n41515 ;
  assign n41580 = n41577 & ~n41579 ;
  assign n41581 = n41519 ^ n41383 ;
  assign n41582 = ~n41580 & ~n41581 ;
  assign n41583 = n41523 & n41582 ;
  assign n41600 = n41599 ^ n41587 ;
  assign n41823 = n41583 & n41600 ;
  assign n41844 = n41843 ^ n41823 ;
  assign n41601 = n41600 ^ n41583 ;
  assign n41605 = n41604 ^ n41601 ;
  assign n41609 = n41582 ^ n41523 ;
  assign n41606 = n39597 ^ n30857 ;
  assign n41607 = n41606 ^ n35773 ;
  assign n41608 = n41607 ^ n2597 ;
  assign n41610 = n41609 ^ n41608 ;
  assign n41612 = n39603 ^ n2651 ;
  assign n41613 = n41612 ^ n35731 ;
  assign n41614 = n41613 ^ n29378 ;
  assign n41611 = n41581 ^ n41580 ;
  assign n41615 = n41614 ^ n41611 ;
  assign n41616 = n39609 ^ n30639 ;
  assign n41617 = n41616 ^ n34061 ;
  assign n41618 = n41617 ^ n29469 ;
  assign n41814 = n41618 ^ n41611 ;
  assign n41619 = n41579 ^ n41577 ;
  assign n41620 = n41619 ^ n41618 ;
  assign n41621 = n41576 ^ n41575 ;
  assign n41622 = n41621 ^ n2858 ;
  assign n41626 = n41574 ^ n41573 ;
  assign n41623 = n30643 ^ n1436 ;
  assign n41624 = n41623 ^ n35529 ;
  assign n41625 = n41624 ^ n2842 ;
  assign n41627 = n41626 ^ n41625 ;
  assign n41632 = n41572 ^ n41570 ;
  assign n41628 = n1421 ^ n1332 ;
  assign n41629 = n41628 ^ n35534 ;
  assign n41630 = n41629 ^ n29387 ;
  assign n41633 = n41632 ^ n41630 ;
  assign n41634 = n41569 ^ n41568 ;
  assign n1742 = n1720 ^ n1314 ;
  assign n1743 = n1742 ^ n1739 ;
  assign n1747 = n1746 ^ n1743 ;
  assign n41635 = n41634 ^ n1747 ;
  assign n41636 = n41567 ^ n41565 ;
  assign n1724 = n1711 ^ n1299 ;
  assign n1731 = n1730 ^ n1724 ;
  assign n1732 = n1731 ^ n1070 ;
  assign n41637 = n41636 ^ n1732 ;
  assign n41641 = n41564 ^ n41563 ;
  assign n41638 = n39212 ^ n1694 ;
  assign n41639 = n41638 ^ n929 ;
  assign n41640 = n41639 ^ n1728 ;
  assign n41642 = n41641 ^ n41640 ;
  assign n41646 = n41562 ^ n41524 ;
  assign n41643 = n39217 ^ n1688 ;
  assign n41644 = n41643 ^ n35545 ;
  assign n41645 = n41644 ^ n921 ;
  assign n41647 = n41646 ^ n41645 ;
  assign n792 = n791 ^ n770 ;
  assign n820 = n819 ^ n792 ;
  assign n827 = n826 ^ n820 ;
  assign n41791 = n41646 ^ n827 ;
  assign n41648 = n41561 ^ n41559 ;
  assign n41649 = n41648 ^ n827 ;
  assign n41653 = n41558 ^ n41557 ;
  assign n41650 = n39224 ^ n2992 ;
  assign n41651 = n41650 ^ n35551 ;
  assign n41652 = n41651 ^ n811 ;
  assign n41654 = n41653 ^ n41652 ;
  assign n41658 = n41556 ^ n41526 ;
  assign n41659 = n41658 ^ n41657 ;
  assign n41663 = n41555 ^ n41527 ;
  assign n41664 = n41663 ^ n41662 ;
  assign n41669 = n41554 ^ n41553 ;
  assign n41665 = n39241 ^ n1535 ;
  assign n41666 = n41665 ^ n35558 ;
  assign n41667 = n41666 ^ n29411 ;
  assign n41670 = n41669 ^ n41667 ;
  assign n41672 = n39246 ^ n30670 ;
  assign n41673 = n41672 ^ n35568 ;
  assign n41674 = n41673 ^ n29416 ;
  assign n41671 = n41552 ^ n41551 ;
  assign n41675 = n41674 ^ n41671 ;
  assign n41677 = n39251 ^ n30674 ;
  assign n41678 = n41677 ^ n35657 ;
  assign n41679 = n41678 ^ n2939 ;
  assign n41774 = n41679 ^ n41671 ;
  assign n41676 = n41550 ^ n41549 ;
  assign n41680 = n41679 ^ n41676 ;
  assign n41685 = n41684 ^ n41681 ;
  assign n41770 = ~n41685 & n41769 ;
  assign n41771 = n41770 ^ n41684 ;
  assign n41772 = n41771 ^ n41679 ;
  assign n41773 = n41680 & n41772 ;
  assign n41775 = n41774 ^ n41773 ;
  assign n41776 = ~n41675 & n41775 ;
  assign n41777 = n41776 ^ n41674 ;
  assign n41778 = n41777 ^ n41667 ;
  assign n41779 = n41670 & n41778 ;
  assign n41668 = n41667 ^ n41662 ;
  assign n41780 = n41779 ^ n41668 ;
  assign n41781 = n41664 & ~n41780 ;
  assign n41782 = n41781 ^ n41663 ;
  assign n41783 = n41782 ^ n41657 ;
  assign n41784 = ~n41659 & ~n41783 ;
  assign n41785 = n41784 ^ n41658 ;
  assign n41786 = n41785 ^ n41652 ;
  assign n41787 = ~n41654 & n41786 ;
  assign n41788 = n41787 ^ n41653 ;
  assign n41789 = n41788 ^ n827 ;
  assign n41790 = n41649 & ~n41789 ;
  assign n41792 = n41791 ^ n41790 ;
  assign n41793 = ~n41647 & ~n41792 ;
  assign n41794 = n41793 ^ n41646 ;
  assign n41795 = n41794 ^ n41640 ;
  assign n41796 = n41642 & n41795 ;
  assign n41797 = n41796 ^ n41641 ;
  assign n41798 = n41797 ^ n41636 ;
  assign n41799 = ~n41637 & n41798 ;
  assign n41800 = n41799 ^ n1732 ;
  assign n41801 = n41800 ^ n1747 ;
  assign n41802 = n41635 & ~n41801 ;
  assign n41803 = n41802 ^ n41634 ;
  assign n41804 = n41803 ^ n41630 ;
  assign n41805 = ~n41633 & n41804 ;
  assign n41631 = n41630 ^ n41626 ;
  assign n41806 = n41805 ^ n41631 ;
  assign n41807 = n41627 & n41806 ;
  assign n41808 = n41807 ^ n41626 ;
  assign n41809 = n41808 ^ n2858 ;
  assign n41810 = ~n41622 & ~n41809 ;
  assign n41811 = n41810 ^ n41621 ;
  assign n41812 = n41811 ^ n41618 ;
  assign n41813 = n41620 & ~n41812 ;
  assign n41815 = n41814 ^ n41813 ;
  assign n41816 = n41615 & ~n41815 ;
  assign n41817 = n41816 ^ n41614 ;
  assign n41818 = n41817 ^ n41608 ;
  assign n41819 = n41610 & ~n41818 ;
  assign n41820 = n41819 ^ n41609 ;
  assign n41821 = n41820 ^ n41604 ;
  assign n41822 = n41605 & n41821 ;
  assign n41845 = n41844 ^ n41822 ;
  assign n41005 = n40478 ^ n39448 ;
  assign n41008 = n41007 ^ n40478 ;
  assign n41009 = ~n41005 & n41008 ;
  assign n41010 = n41009 ^ n39448 ;
  assign n41846 = n41845 ^ n41010 ;
  assign n41848 = n40488 ^ n39451 ;
  assign n41849 = n41125 ^ n40488 ;
  assign n41850 = ~n41848 & n41849 ;
  assign n41851 = n41850 ^ n39451 ;
  assign n41847 = n41820 ^ n41605 ;
  assign n41852 = n41851 ^ n41847 ;
  assign n41857 = n41817 ^ n41610 ;
  assign n41878 = n41857 ^ n41851 ;
  assign n41853 = n41132 ^ n39459 ;
  assign n41854 = n40522 ^ n39459 ;
  assign n41855 = n41853 & n41854 ;
  assign n41856 = n41855 ^ n40522 ;
  assign n41858 = n41857 ^ n41856 ;
  assign n41859 = n41138 ^ n40494 ;
  assign n41860 = n41811 ^ n41620 ;
  assign n41861 = n41145 ^ n38840 ;
  assign n41862 = n40514 ^ n38840 ;
  assign n41863 = ~n41861 & ~n41862 ;
  assign n41864 = n41863 ^ n40514 ;
  assign n41865 = ~n41860 & n41864 ;
  assign n41866 = n41865 ^ n39465 ;
  assign n41867 = n41866 ^ n41138 ;
  assign n41868 = n41867 ^ n41865 ;
  assign n41869 = ~n41859 & n41868 ;
  assign n41870 = n41869 ^ n41866 ;
  assign n41873 = n41865 ^ n41856 ;
  assign n41871 = n41815 ^ n41614 ;
  assign n41872 = n41871 ^ n41856 ;
  assign n41874 = n41873 ^ n41872 ;
  assign n41875 = ~n41870 & n41874 ;
  assign n41876 = n41875 ^ n41873 ;
  assign n41877 = ~n41858 & n41876 ;
  assign n41879 = n41878 ^ n41877 ;
  assign n41880 = ~n41852 & ~n41879 ;
  assign n41881 = n41880 ^ n41851 ;
  assign n41882 = n41881 ^ n41010 ;
  assign n41883 = n41846 & ~n41882 ;
  assign n41884 = n41883 ^ n41845 ;
  assign n41885 = n41884 ^ n40999 ;
  assign n41886 = ~n41004 & n41885 ;
  assign n41892 = n41891 ^ n41886 ;
  assign n41893 = n41725 ^ n41723 ;
  assign n41927 = n41893 ^ n41890 ;
  assign n41928 = ~n41892 & ~n41927 ;
  assign n41929 = n41928 ^ n41890 ;
  assign n42013 = n42012 ^ n41929 ;
  assign n42014 = n41936 & n42013 ;
  assign n42015 = n42014 ^ n42011 ;
  assign n42168 = n40550 ^ n39803 ;
  assign n42169 = n41090 ^ n40550 ;
  assign n42170 = n42168 & n42169 ;
  assign n42171 = n42170 ^ n39803 ;
  assign n42173 = n42171 ^ n42010 ;
  assign n42016 = n41731 ^ n41712 ;
  assign n42172 = n42171 ^ n42016 ;
  assign n42174 = n42173 ^ n42172 ;
  assign n42175 = n42015 & n42174 ;
  assign n42176 = n42175 ^ n42173 ;
  assign n42180 = n42171 ^ n42164 ;
  assign n42177 = n41738 ^ n41734 ;
  assign n42178 = n42177 ^ n41733 ;
  assign n42179 = n42178 ^ n42164 ;
  assign n42181 = n42180 ^ n42179 ;
  assign n42182 = ~n42176 & ~n42181 ;
  assign n42183 = n42182 ^ n42180 ;
  assign n42184 = n42167 & ~n42183 ;
  assign n42165 = n42164 ^ n42159 ;
  assign n42185 = n42184 ^ n42165 ;
  assign n42186 = ~n42160 & n42185 ;
  assign n42187 = n42186 ^ n42060 ;
  assign n42150 = n41075 ^ n40694 ;
  assign n42151 = n40694 ^ n39421 ;
  assign n42152 = ~n42150 & n42151 ;
  assign n42153 = n42152 ^ n39421 ;
  assign n42154 = n42153 ^ n42044 ;
  assign n42155 = n42154 ^ n42153 ;
  assign n42188 = n42187 ^ n42155 ;
  assign n42189 = n42149 & ~n42188 ;
  assign n42190 = n42189 ^ n42154 ;
  assign n42192 = n42153 ^ n42142 ;
  assign n42053 = n41757 ^ n2268 ;
  assign n42191 = n42142 ^ n42053 ;
  assign n42193 = n42192 ^ n42191 ;
  assign n42194 = ~n42190 & ~n42193 ;
  assign n42195 = n42194 ^ n42192 ;
  assign n42196 = n42143 & ~n42195 ;
  assign n42197 = n42196 ^ n42142 ;
  assign n42202 = n42201 ^ n42197 ;
  assign n42203 = n41762 ^ n41692 ;
  assign n42206 = n42203 ^ n42197 ;
  assign n42207 = ~n42202 & ~n42206 ;
  assign n42204 = n42203 ^ n42136 ;
  assign n42208 = n42207 ^ n42204 ;
  assign n42209 = ~n42137 & n42208 ;
  assign n42210 = n42209 ^ n42136 ;
  assign n42211 = n42210 ^ n42130 ;
  assign n42212 = ~n42131 & ~n42211 ;
  assign n42213 = n42212 ^ n42038 ;
  assign n42122 = n40787 ^ n39387 ;
  assign n42123 = n41040 ^ n40787 ;
  assign n42124 = ~n42122 & n42123 ;
  assign n42125 = n42124 ^ n39387 ;
  assign n42031 = n41771 ^ n41680 ;
  assign n42126 = n42125 ^ n42031 ;
  assign n42270 = n42213 ^ n42126 ;
  assign n42271 = n42270 ^ n39416 ;
  assign n42316 = n42210 ^ n42131 ;
  assign n42273 = n42203 ^ n42201 ;
  assign n42274 = n42273 ^ n42197 ;
  assign n42275 = n42274 ^ n39356 ;
  assign n42276 = n42190 ^ n42053 ;
  assign n42277 = n42276 ^ n38851 ;
  assign n42278 = n42187 ^ n42149 ;
  assign n42279 = n42278 ^ n38857 ;
  assign n42280 = n42185 ^ n42060 ;
  assign n42281 = n42280 ^ n38860 ;
  assign n42290 = n42183 ^ n42166 ;
  assign n42282 = n42178 ^ n42176 ;
  assign n42283 = n42282 ^ n38876 ;
  assign n42017 = n42016 ^ n42015 ;
  assign n42018 = n42017 ^ n38878 ;
  assign n41937 = n41936 ^ n41929 ;
  assign n41938 = n41937 ^ n38884 ;
  assign n41894 = n41893 ^ n41892 ;
  assign n41895 = n41894 ^ n38890 ;
  assign n41896 = n41884 ^ n41004 ;
  assign n41897 = n41896 ^ n38896 ;
  assign n41899 = n41879 ^ n41847 ;
  assign n41900 = n41899 ^ n38908 ;
  assign n41908 = n41876 ^ n41857 ;
  assign n41901 = n41864 ^ n41860 ;
  assign n41902 = ~n38922 & ~n41901 ;
  assign n41903 = n41902 ^ n38915 ;
  assign n41904 = n41871 ^ n41870 ;
  assign n41905 = n41904 ^ n41902 ;
  assign n41906 = ~n41903 & n41905 ;
  assign n41907 = n41906 ^ n38915 ;
  assign n41909 = n41908 ^ n41907 ;
  assign n41910 = n41908 ^ n38841 ;
  assign n41911 = ~n41909 & ~n41910 ;
  assign n41912 = n41911 ^ n38841 ;
  assign n41913 = n41912 ^ n41899 ;
  assign n41914 = ~n41900 & n41913 ;
  assign n41915 = n41914 ^ n38908 ;
  assign n41898 = n41881 ^ n41846 ;
  assign n41916 = n41915 ^ n41898 ;
  assign n41917 = n41896 ^ n38902 ;
  assign n41918 = n41917 ^ n41896 ;
  assign n41919 = n41918 ^ n41898 ;
  assign n41920 = n41916 & n41919 ;
  assign n41921 = n41920 ^ n41917 ;
  assign n41922 = n41897 & n41921 ;
  assign n41923 = n41922 ^ n38896 ;
  assign n41924 = n41923 ^ n41894 ;
  assign n41925 = ~n41895 & ~n41924 ;
  assign n41926 = n41925 ^ n38890 ;
  assign n42019 = n41937 ^ n41926 ;
  assign n42020 = ~n41938 & n42019 ;
  assign n42021 = n42020 ^ n38884 ;
  assign n42284 = n42021 ^ n42017 ;
  assign n42285 = ~n42018 & n42284 ;
  assign n42286 = n42285 ^ n38878 ;
  assign n42287 = n42286 ^ n42282 ;
  assign n42288 = ~n42283 & ~n42287 ;
  assign n42289 = n42288 ^ n38876 ;
  assign n42291 = n42290 ^ n42289 ;
  assign n42292 = n42290 ^ n38870 ;
  assign n42293 = n42291 & ~n42292 ;
  assign n42294 = n42293 ^ n38870 ;
  assign n42295 = n42294 ^ n42280 ;
  assign n42296 = n42281 & n42295 ;
  assign n42297 = n42296 ^ n38860 ;
  assign n42298 = n42297 ^ n42278 ;
  assign n42299 = ~n42279 & n42298 ;
  assign n42300 = n42299 ^ n38857 ;
  assign n42301 = n42300 ^ n42276 ;
  assign n42302 = n42277 & n42301 ;
  assign n42303 = n42302 ^ n38851 ;
  assign n42304 = n42303 ^ n39067 ;
  assign n42305 = n42195 ^ n42138 ;
  assign n42306 = n42305 ^ n42303 ;
  assign n42307 = ~n42304 & ~n42306 ;
  assign n42308 = n42307 ^ n39067 ;
  assign n42309 = n42308 ^ n42274 ;
  assign n42310 = n42275 & n42309 ;
  assign n42311 = n42310 ^ n39356 ;
  assign n42272 = n42208 ^ n42132 ;
  assign n42312 = n42311 ^ n42272 ;
  assign n42313 = n42311 ^ n39431 ;
  assign n42314 = n42312 & n42313 ;
  assign n42315 = n42314 ^ n39431 ;
  assign n42317 = n42316 ^ n42315 ;
  assign n42318 = n42316 ^ n39424 ;
  assign n42319 = n42317 & ~n42318 ;
  assign n42320 = n42319 ^ n39424 ;
  assign n42321 = n42320 ^ n42270 ;
  assign n42322 = ~n42271 & ~n42321 ;
  assign n42323 = n42322 ^ n39416 ;
  assign n42214 = n42213 ^ n42125 ;
  assign n42215 = ~n42126 & ~n42214 ;
  assign n42216 = n42215 ^ n42031 ;
  assign n42120 = n41775 ^ n41674 ;
  assign n42116 = n41033 ^ n40808 ;
  assign n42117 = n40808 ^ n39385 ;
  assign n42118 = ~n42116 & ~n42117 ;
  assign n42119 = n42118 ^ n39385 ;
  assign n42121 = n42120 ^ n42119 ;
  assign n42268 = n42216 ^ n42121 ;
  assign n42269 = n42268 ^ n39410 ;
  assign n42410 = n42323 ^ n42269 ;
  assign n42388 = n42318 ^ n42315 ;
  assign n42389 = n42300 ^ n42277 ;
  assign n42390 = n42292 ^ n42289 ;
  assign n42391 = n42286 ^ n42283 ;
  assign n41939 = n41938 ^ n41926 ;
  assign n41940 = n41910 ^ n41907 ;
  assign n41941 = n41912 ^ n41900 ;
  assign n41942 = ~n41940 & n41941 ;
  assign n41943 = n41898 ^ n38902 ;
  assign n41944 = n41943 ^ n41915 ;
  assign n41945 = n41942 & ~n41944 ;
  assign n41946 = n41921 ^ n38896 ;
  assign n41947 = ~n41945 & ~n41946 ;
  assign n41948 = n41923 ^ n41895 ;
  assign n41949 = ~n41947 & n41948 ;
  assign n42006 = ~n41939 & n41949 ;
  assign n42022 = n42021 ^ n42018 ;
  assign n42392 = ~n42006 & n42022 ;
  assign n42393 = n42391 & n42392 ;
  assign n42394 = n42390 & ~n42393 ;
  assign n42395 = n42294 ^ n42281 ;
  assign n42396 = n42394 & ~n42395 ;
  assign n42397 = n42297 ^ n42279 ;
  assign n42398 = n42396 & ~n42397 ;
  assign n42399 = n42389 & n42398 ;
  assign n42400 = n42305 ^ n42304 ;
  assign n42401 = ~n42399 & ~n42400 ;
  assign n42402 = n42308 ^ n42275 ;
  assign n42403 = ~n42401 & n42402 ;
  assign n42404 = n42272 ^ n39431 ;
  assign n42405 = n42404 ^ n42311 ;
  assign n42406 = n42403 & n42405 ;
  assign n42407 = n42388 & n42406 ;
  assign n42408 = n42320 ^ n42271 ;
  assign n42409 = ~n42407 & ~n42408 ;
  assign n42479 = n42410 ^ n42409 ;
  assign n42564 = n42483 ^ n42479 ;
  assign n42484 = n42408 ^ n42407 ;
  assign n42485 = n42484 ^ n42483 ;
  assign n42489 = n42406 ^ n42388 ;
  assign n42486 = n40106 ^ n1590 ;
  assign n42487 = n42486 ^ n36327 ;
  assign n42488 = n42487 ^ n2978 ;
  assign n42490 = n42489 ^ n42488 ;
  assign n42494 = n42405 ^ n42403 ;
  assign n42491 = n40111 ^ n31384 ;
  assign n42492 = n42491 ^ n2966 ;
  assign n42493 = n42492 ^ n29763 ;
  assign n42495 = n42494 ^ n42493 ;
  assign n42496 = n42402 ^ n42401 ;
  assign n42500 = n42499 ^ n42496 ;
  assign n42506 = n42400 ^ n42399 ;
  assign n42503 = n40122 ^ n2948 ;
  assign n42504 = n42503 ^ n36342 ;
  assign n42505 = n42504 ^ n29771 ;
  assign n42507 = n42506 ^ n42505 ;
  assign n42509 = n40126 ^ n31396 ;
  assign n42510 = n42509 ^ n36347 ;
  assign n42511 = n42510 ^ n29775 ;
  assign n42550 = n42511 ^ n42506 ;
  assign n42508 = n42398 ^ n42389 ;
  assign n42512 = n42511 ^ n42508 ;
  assign n42516 = n42397 ^ n42396 ;
  assign n42513 = n40131 ^ n31403 ;
  assign n42514 = n42513 ^ n36351 ;
  assign n42515 = n42514 ^ n29780 ;
  assign n42517 = n42516 ^ n42515 ;
  assign n42521 = n42395 ^ n42394 ;
  assign n42544 = n42521 ^ n42516 ;
  assign n42518 = n31461 ^ n2440 ;
  assign n42519 = n42518 ^ n36357 ;
  assign n42520 = n42519 ^ n29786 ;
  assign n42522 = n42521 ^ n42520 ;
  assign n42524 = n31407 ^ n2422 ;
  assign n42525 = n42524 ^ n36362 ;
  assign n42526 = n42525 ^ n29850 ;
  assign n42541 = n42526 ^ n42521 ;
  assign n42523 = n42393 ^ n42390 ;
  assign n42527 = n42526 ^ n42523 ;
  assign n42531 = n42392 ^ n42391 ;
  assign n42528 = n40141 ^ n2348 ;
  assign n42529 = n42528 ^ n36367 ;
  assign n42530 = n42529 ^ n29791 ;
  assign n42532 = n42531 ^ n42530 ;
  assign n42023 = n42022 ^ n42006 ;
  assign n41951 = n40151 ^ n31418 ;
  assign n41952 = n41951 ^ n36402 ;
  assign n41953 = n41952 ^ n29800 ;
  assign n42024 = n42023 ^ n41953 ;
  assign n41950 = n41949 ^ n41939 ;
  assign n41954 = n41953 ^ n41950 ;
  assign n41958 = n41948 ^ n41947 ;
  assign n41955 = n40155 ^ n31423 ;
  assign n41956 = n41955 ^ n36377 ;
  assign n41957 = n41956 ^ n2036 ;
  assign n41959 = n41958 ^ n41957 ;
  assign n41963 = n41946 ^ n41945 ;
  assign n41960 = n40161 ^ n31428 ;
  assign n41961 = n41960 ^ n1970 ;
  assign n41962 = n41961 ^ n29807 ;
  assign n41964 = n41963 ^ n41962 ;
  assign n41968 = n41944 ^ n41942 ;
  assign n41965 = n40185 ^ n31435 ;
  assign n41966 = n41965 ^ n36384 ;
  assign n41967 = n41966 ^ n1962 ;
  assign n41969 = n41968 ^ n41967 ;
  assign n41987 = n41941 ^ n41940 ;
  assign n41970 = n40169 ^ n30821 ;
  assign n41971 = n41970 ^ n3023 ;
  assign n41972 = n41971 ^ n29816 ;
  assign n41973 = n41972 ^ n41940 ;
  assign n2706 = n2705 ^ n2684 ;
  assign n2725 = n2724 ^ n2706 ;
  assign n2732 = n2731 ^ n2725 ;
  assign n41977 = n41901 ^ n38922 ;
  assign n41978 = n2732 & n41977 ;
  assign n41979 = n41978 ^ n41976 ;
  assign n41980 = n41904 ^ n41903 ;
  assign n41981 = n41980 ^ n41976 ;
  assign n41982 = n41979 & ~n41981 ;
  assign n41983 = n41982 ^ n41978 ;
  assign n41984 = n41983 ^ n41972 ;
  assign n41985 = ~n41973 & ~n41984 ;
  assign n41986 = n41985 ^ n41940 ;
  assign n41988 = n41987 ^ n41986 ;
  assign n41989 = n40165 ^ n1895 ;
  assign n41990 = n41989 ^ n35785 ;
  assign n41991 = n41990 ^ n3062 ;
  assign n41992 = n41991 ^ n41986 ;
  assign n41993 = ~n41988 & n41992 ;
  assign n41994 = n41993 ^ n41987 ;
  assign n41995 = n41994 ^ n41967 ;
  assign n41996 = n41969 & ~n41995 ;
  assign n41997 = n41996 ^ n41968 ;
  assign n41998 = n41997 ^ n41962 ;
  assign n41999 = n41964 & n41998 ;
  assign n42000 = n41999 ^ n41962 ;
  assign n42001 = n42000 ^ n41957 ;
  assign n42002 = n41959 & ~n42001 ;
  assign n42003 = n42002 ^ n41958 ;
  assign n42004 = n42003 ^ n41953 ;
  assign n42005 = n41954 & n42004 ;
  assign n42025 = n42024 ^ n42005 ;
  assign n42026 = n40146 ^ n2333 ;
  assign n42027 = n42026 ^ n36372 ;
  assign n42028 = n42027 ^ n29795 ;
  assign n42533 = n42028 ^ n42023 ;
  assign n42534 = n42025 & ~n42533 ;
  assign n42535 = n42534 ^ n42028 ;
  assign n42536 = n42535 ^ n42530 ;
  assign n42537 = n42532 & ~n42536 ;
  assign n42538 = n42537 ^ n42531 ;
  assign n42539 = n42538 ^ n42526 ;
  assign n42540 = n42527 & n42539 ;
  assign n42542 = n42541 ^ n42540 ;
  assign n42543 = n42522 & n42542 ;
  assign n42545 = n42544 ^ n42543 ;
  assign n42546 = n42517 & n42545 ;
  assign n42547 = n42546 ^ n42516 ;
  assign n42548 = n42547 ^ n42511 ;
  assign n42549 = ~n42512 & n42548 ;
  assign n42551 = n42550 ^ n42549 ;
  assign n42552 = n42507 & n42551 ;
  assign n42553 = n42552 ^ n42506 ;
  assign n42501 = n42499 ^ n42494 ;
  assign n42502 = n42501 ^ n42494 ;
  assign n42554 = n42553 ^ n42502 ;
  assign n42555 = n42500 & n42554 ;
  assign n42556 = n42555 ^ n42501 ;
  assign n42557 = ~n42495 & ~n42556 ;
  assign n42558 = n42557 ^ n42494 ;
  assign n42559 = n42558 ^ n42488 ;
  assign n42560 = ~n42490 & n42559 ;
  assign n42561 = n42560 ^ n42489 ;
  assign n42562 = n42561 ^ n42483 ;
  assign n42563 = n42485 & ~n42562 ;
  assign n42565 = n42564 ^ n42563 ;
  assign n43074 = n42565 ^ n1637 ;
  assign n42089 = n41788 ^ n41649 ;
  assign n44267 = n43074 ^ n42089 ;
  assign n42849 = n42542 ^ n42520 ;
  assign n42108 = n41780 ^ n41663 ;
  assign n42843 = n42108 ^ n41040 ;
  assign n42844 = n41040 ^ n40756 ;
  assign n42845 = n42843 & n42844 ;
  assign n42846 = n42845 ^ n40756 ;
  assign n42825 = n42538 ^ n42527 ;
  assign n42847 = n42846 ^ n42825 ;
  assign n42114 = n41777 ^ n41670 ;
  assign n42824 = n42114 ^ n41047 ;
  assign n42826 = n42825 ^ n40729 ;
  assign n42827 = n42826 ^ n42114 ;
  assign n42828 = n42827 ^ n42825 ;
  assign n42829 = ~n42824 & ~n42828 ;
  assign n42830 = n42829 ^ n42826 ;
  assign n42721 = n41057 ^ n40711 ;
  assign n42722 = n42120 ^ n41057 ;
  assign n42723 = ~n42721 & n42722 ;
  assign n42724 = n42723 ^ n40711 ;
  assign n42720 = n42535 ^ n42532 ;
  assign n42725 = n42724 ^ n42720 ;
  assign n42030 = n41063 ^ n40694 ;
  assign n42032 = n42031 ^ n41063 ;
  assign n42033 = n42030 & ~n42032 ;
  assign n42034 = n42033 ^ n40694 ;
  assign n42029 = n42028 ^ n42025 ;
  assign n42035 = n42034 ^ n42029 ;
  assign n42037 = n41069 ^ n40653 ;
  assign n42039 = n42038 ^ n41069 ;
  assign n42040 = ~n42037 & ~n42039 ;
  assign n42041 = n42040 ^ n40653 ;
  assign n42036 = n42003 ^ n41954 ;
  assign n42042 = n42041 ^ n42036 ;
  assign n42704 = n42132 ^ n41075 ;
  assign n42705 = n41075 ^ n40570 ;
  assign n42706 = n42704 & ~n42705 ;
  assign n42707 = n42706 ^ n40570 ;
  assign n42713 = n42707 ^ n42041 ;
  assign n42701 = n41997 ^ n41964 ;
  assign n42708 = n42707 ^ n42701 ;
  assign n42045 = n42044 ^ n41090 ;
  assign n42046 = n41983 ^ n41973 ;
  assign n42047 = n42046 ^ n40460 ;
  assign n42048 = n42047 ^ n41090 ;
  assign n42049 = n42048 ^ n42046 ;
  assign n42050 = n42045 & ~n42049 ;
  assign n42051 = n42050 ^ n42047 ;
  assign n42061 = n42060 ^ n41096 ;
  assign n42062 = n42060 ^ n40466 ;
  assign n42063 = ~n42061 & ~n42062 ;
  assign n42064 = n42063 ^ n40466 ;
  assign n42059 = n41980 ^ n41979 ;
  assign n42065 = n42064 ^ n42059 ;
  assign n42665 = n41977 ^ n2732 ;
  assign n42674 = n42665 ^ n42064 ;
  assign n42623 = n42178 ^ n41112 ;
  assign n42624 = n41112 ^ n40478 ;
  assign n42625 = ~n42623 & n42624 ;
  assign n42626 = n42625 ^ n40478 ;
  assign n42617 = n40509 ^ n39739 ;
  assign n42618 = n41247 ^ n40509 ;
  assign n42619 = ~n42617 & n42618 ;
  assign n42066 = n40989 ^ n40286 ;
  assign n42067 = n41797 ^ n41637 ;
  assign n42068 = n42067 ^ n39669 ;
  assign n42069 = n42068 ^ n40989 ;
  assign n42070 = n42069 ^ n42067 ;
  assign n42071 = n42066 & ~n42070 ;
  assign n42072 = n42071 ^ n42068 ;
  assign n42083 = n41794 ^ n41642 ;
  assign n42079 = n40298 ^ n39677 ;
  assign n42080 = n41832 ^ n40298 ;
  assign n42081 = n42079 & ~n42080 ;
  assign n42082 = n42081 ^ n39677 ;
  assign n42084 = n42083 ^ n42082 ;
  assign n42235 = n41792 ^ n41645 ;
  assign n42085 = n41019 ^ n40401 ;
  assign n42086 = n41379 ^ n41019 ;
  assign n42087 = ~n42085 & n42086 ;
  assign n42088 = n42087 ^ n40401 ;
  assign n42090 = n42089 ^ n42088 ;
  assign n42092 = n41785 ^ n41654 ;
  assign n42231 = n42092 ^ n42088 ;
  assign n42091 = n41374 ^ n41025 ;
  assign n42093 = n42092 ^ n40323 ;
  assign n42094 = n42093 ^ n41374 ;
  assign n42095 = n42094 ^ n42092 ;
  assign n42096 = n42091 & n42095 ;
  assign n42097 = n42096 ^ n42093 ;
  assign n42102 = n41782 ^ n41659 ;
  assign n42098 = n41035 ^ n40274 ;
  assign n42099 = n41035 ^ n41016 ;
  assign n42100 = n42098 & n42099 ;
  assign n42101 = n42100 ^ n40274 ;
  assign n42103 = n42102 ^ n42101 ;
  assign n42104 = n41041 ^ n39853 ;
  assign n42105 = n41041 ^ n41023 ;
  assign n42106 = ~n42104 & n42105 ;
  assign n42107 = n42106 ^ n39853 ;
  assign n42109 = n42108 ^ n42107 ;
  assign n42110 = n40829 ^ n39368 ;
  assign n42111 = n41027 ^ n40829 ;
  assign n42112 = n42110 & ~n42111 ;
  assign n42113 = n42112 ^ n39368 ;
  assign n42115 = n42114 ^ n42113 ;
  assign n42217 = n42216 ^ n42119 ;
  assign n42218 = n42121 & n42217 ;
  assign n42219 = n42218 ^ n42120 ;
  assign n42220 = n42219 ^ n42113 ;
  assign n42221 = ~n42115 & ~n42220 ;
  assign n42222 = n42221 ^ n42114 ;
  assign n42223 = n42222 ^ n42107 ;
  assign n42224 = n42109 & ~n42223 ;
  assign n42225 = n42224 ^ n42108 ;
  assign n42226 = n42225 ^ n42101 ;
  assign n42227 = n42103 & n42226 ;
  assign n42228 = n42227 ^ n42102 ;
  assign n42229 = n42228 ^ n42092 ;
  assign n42230 = n42097 & ~n42229 ;
  assign n42232 = n42231 ^ n42230 ;
  assign n42233 = ~n42090 & ~n42232 ;
  assign n42234 = n42233 ^ n42089 ;
  assign n42236 = n42235 ^ n42234 ;
  assign n42237 = n41588 ^ n40296 ;
  assign n42238 = n42235 ^ n39678 ;
  assign n42239 = n42238 ^ n41588 ;
  assign n42240 = n42239 ^ n42235 ;
  assign n42241 = n42237 & n42240 ;
  assign n42242 = n42241 ^ n42238 ;
  assign n42243 = n42236 & n42242 ;
  assign n42244 = n42243 ^ n42235 ;
  assign n42245 = n42244 ^ n42082 ;
  assign n42246 = n42084 & ~n42245 ;
  assign n42247 = n42246 ^ n42083 ;
  assign n42073 = n40342 ^ n39662 ;
  assign n42074 = n41260 ^ n40342 ;
  assign n42075 = ~n42073 & n42074 ;
  assign n42076 = n42075 ^ n39662 ;
  assign n42077 = n42076 ^ n42067 ;
  assign n42078 = n42077 ^ n42076 ;
  assign n42248 = n42247 ^ n42078 ;
  assign n42249 = n42072 & n42248 ;
  assign n42250 = n42249 ^ n42077 ;
  assign n42356 = n41803 ^ n41633 ;
  assign n42358 = n42356 ^ n42076 ;
  assign n42251 = n41800 ^ n41635 ;
  assign n42357 = n42356 ^ n42251 ;
  assign n42359 = n42358 ^ n42357 ;
  assign n42360 = ~n42250 & n42359 ;
  assign n42361 = n42360 ^ n42358 ;
  assign n42375 = n41806 ^ n41625 ;
  assign n42377 = n42375 ^ n42356 ;
  assign n42362 = n41270 ^ n40414 ;
  assign n42363 = n40414 ^ n39721 ;
  assign n42364 = ~n42362 & n42363 ;
  assign n42365 = n42364 ^ n39721 ;
  assign n42376 = n42375 ^ n42365 ;
  assign n42378 = n42377 ^ n42376 ;
  assign n42379 = ~n42361 & n42378 ;
  assign n42380 = n42379 ^ n42377 ;
  assign n42371 = n40432 ^ n39472 ;
  assign n42372 = n41257 ^ n39472 ;
  assign n42373 = ~n42371 & ~n42372 ;
  assign n42374 = n42373 ^ n40432 ;
  assign n42381 = n42380 ^ n42374 ;
  assign n42382 = n42381 ^ n38935 ;
  assign n42366 = n42365 ^ n42361 ;
  assign n42253 = n42247 ^ n42072 ;
  assign n42254 = n42253 ^ n38832 ;
  assign n42255 = n42244 ^ n42084 ;
  assign n42256 = n42255 ^ n38783 ;
  assign n42258 = n42232 ^ n42089 ;
  assign n42259 = n42258 ^ n39381 ;
  assign n42260 = n42228 ^ n42097 ;
  assign n42261 = n42260 ^ n39389 ;
  assign n42262 = n42225 ^ n42103 ;
  assign n42263 = n42262 ^ n39484 ;
  assign n42264 = n42222 ^ n42109 ;
  assign n42265 = n42264 ^ n39394 ;
  assign n42266 = n42219 ^ n42115 ;
  assign n42267 = n42266 ^ n39403 ;
  assign n42324 = n42323 ^ n42268 ;
  assign n42325 = ~n42269 & n42324 ;
  assign n42326 = n42325 ^ n39410 ;
  assign n42327 = n42326 ^ n42266 ;
  assign n42328 = ~n42267 & n42327 ;
  assign n42329 = n42328 ^ n39403 ;
  assign n42330 = n42329 ^ n42264 ;
  assign n42331 = n42265 & n42330 ;
  assign n42332 = n42331 ^ n39394 ;
  assign n42333 = n42332 ^ n42262 ;
  assign n42334 = n42263 & ~n42333 ;
  assign n42335 = n42334 ^ n39484 ;
  assign n42336 = n42335 ^ n42260 ;
  assign n42337 = n42261 & n42336 ;
  assign n42338 = n42337 ^ n39389 ;
  assign n42339 = n42338 ^ n42258 ;
  assign n42340 = ~n42259 & ~n42339 ;
  assign n42341 = n42340 ^ n39381 ;
  assign n42257 = n42242 ^ n42234 ;
  assign n42342 = n42341 ^ n42257 ;
  assign n42343 = n42341 ^ n38748 ;
  assign n42344 = n42342 & ~n42343 ;
  assign n42345 = n42344 ^ n38748 ;
  assign n42346 = n42345 ^ n42255 ;
  assign n42347 = n42256 & ~n42346 ;
  assign n42348 = n42347 ^ n38783 ;
  assign n42349 = n42348 ^ n42253 ;
  assign n42350 = ~n42254 & ~n42349 ;
  assign n42351 = n42350 ^ n38832 ;
  assign n42252 = n42251 ^ n42250 ;
  assign n42352 = n42351 ^ n42252 ;
  assign n42353 = n42351 ^ n38969 ;
  assign n42354 = n42352 & n42353 ;
  assign n42355 = n42354 ^ n38969 ;
  assign n42367 = n42366 ^ n42355 ;
  assign n42368 = n42366 ^ n39003 ;
  assign n42369 = ~n42367 & ~n42368 ;
  assign n42370 = n42369 ^ n39003 ;
  assign n42614 = n42381 ^ n42370 ;
  assign n42615 = ~n42382 & n42614 ;
  assign n42608 = n40340 ^ n3224 ;
  assign n42609 = n42608 ^ n36683 ;
  assign n42610 = n42609 ^ n2719 ;
  assign n42431 = n40284 ^ n2612 ;
  assign n42432 = n42431 ^ n36545 ;
  assign n42433 = n42432 ^ n30193 ;
  assign n42611 = n42610 ^ n42433 ;
  assign n42605 = n42375 ^ n39739 ;
  assign n42604 = n41808 ^ n41622 ;
  assign n42606 = n42605 ^ n42604 ;
  assign n42603 = n38935 ^ n38932 ;
  assign n42607 = n42606 ^ n42603 ;
  assign n42612 = n42611 ^ n42607 ;
  assign n42601 = n42375 ^ n42374 ;
  assign n42602 = ~n42380 & ~n42601 ;
  assign n42613 = n42612 ^ n42602 ;
  assign n42616 = n42615 ^ n42613 ;
  assign n42620 = n42619 ^ n42616 ;
  assign n42383 = n42382 ^ n42370 ;
  assign n42384 = n42368 ^ n42355 ;
  assign n42385 = n42348 ^ n42254 ;
  assign n42386 = n42257 ^ n38748 ;
  assign n42387 = n42386 ^ n42341 ;
  assign n42411 = ~n42409 & ~n42410 ;
  assign n42412 = n42326 ^ n42267 ;
  assign n42413 = n42411 & ~n42412 ;
  assign n42414 = n42329 ^ n42265 ;
  assign n42415 = ~n42413 & ~n42414 ;
  assign n42416 = n42332 ^ n42263 ;
  assign n42417 = n42415 & n42416 ;
  assign n42418 = n42335 ^ n42261 ;
  assign n42419 = n42417 & n42418 ;
  assign n42420 = n42338 ^ n42259 ;
  assign n42421 = ~n42419 & ~n42420 ;
  assign n42422 = ~n42387 & n42421 ;
  assign n42423 = n42345 ^ n42256 ;
  assign n42424 = n42422 & n42423 ;
  assign n42425 = ~n42385 & n42424 ;
  assign n42426 = n42252 ^ n38969 ;
  assign n42427 = n42426 ^ n42351 ;
  assign n42428 = ~n42425 & ~n42427 ;
  assign n42429 = ~n42384 & n42428 ;
  assign n42600 = n42383 & n42429 ;
  assign n42621 = n42620 ^ n42600 ;
  assign n42430 = n42429 ^ n42383 ;
  assign n42434 = n42433 ^ n42430 ;
  assign n42438 = n42428 ^ n42384 ;
  assign n42435 = n38845 ^ n31774 ;
  assign n42436 = n42435 ^ n36502 ;
  assign n42437 = n42436 ^ n3128 ;
  assign n42439 = n42438 ^ n42437 ;
  assign n42443 = n42427 ^ n42425 ;
  assign n42440 = n40060 ^ n31577 ;
  assign n42441 = n42440 ^ n36292 ;
  assign n42442 = n42441 ^ n30200 ;
  assign n42444 = n42443 ^ n42442 ;
  assign n42448 = n42424 ^ n42385 ;
  assign n42445 = n40065 ^ n2902 ;
  assign n42446 = n42445 ^ n36288 ;
  assign n42447 = n42446 ^ n30206 ;
  assign n42449 = n42448 ^ n42447 ;
  assign n42451 = n40070 ^ n2887 ;
  assign n42452 = n42451 ^ n36298 ;
  assign n42453 = n42452 ^ n30211 ;
  assign n42450 = n42423 ^ n42422 ;
  assign n42454 = n42453 ^ n42450 ;
  assign n42456 = n40075 ^ n31522 ;
  assign n42457 = n42456 ^ n1388 ;
  assign n42458 = n42457 ^ n30215 ;
  assign n42455 = n42421 ^ n42387 ;
  assign n42459 = n42458 ^ n42455 ;
  assign n42461 = n40079 ^ n1773 ;
  assign n42462 = n42461 ^ n36304 ;
  assign n42463 = n42462 ^ n1352 ;
  assign n42582 = n42463 ^ n42455 ;
  assign n42460 = n42420 ^ n42419 ;
  assign n42464 = n42463 ^ n42460 ;
  assign n42465 = n42418 ^ n42417 ;
  assign n1161 = n1160 ^ n1091 ;
  assign n1177 = n1176 ^ n1161 ;
  assign n1184 = n1183 ^ n1177 ;
  assign n42466 = n42465 ^ n1184 ;
  assign n42470 = n42416 ^ n42415 ;
  assign n42467 = n40086 ^ n1755 ;
  assign n42468 = n42467 ^ n1048 ;
  assign n42469 = n42468 ^ n1168 ;
  assign n42471 = n42470 ^ n42469 ;
  assign n42472 = n42414 ^ n42413 ;
  assign n1006 = n996 ^ n957 ;
  assign n1031 = n1030 ^ n1006 ;
  assign n1038 = n1037 ^ n1031 ;
  assign n42473 = n42472 ^ n1038 ;
  assign n42477 = n42412 ^ n42411 ;
  assign n42474 = n40093 ^ n892 ;
  assign n42475 = n42474 ^ n36317 ;
  assign n42476 = n42475 ^ n1022 ;
  assign n42478 = n42477 ^ n42476 ;
  assign n42480 = n42479 ^ n1637 ;
  assign n42566 = ~n42480 & ~n42565 ;
  assign n42567 = n42566 ^ n42479 ;
  assign n42568 = n42567 ^ n42476 ;
  assign n42569 = n42478 & n42568 ;
  assign n42570 = n42569 ^ n42477 ;
  assign n42571 = n42570 ^ n1038 ;
  assign n42572 = n42473 & ~n42571 ;
  assign n42573 = n42572 ^ n42472 ;
  assign n42574 = n42573 ^ n42469 ;
  assign n42575 = n42471 & ~n42574 ;
  assign n42576 = n42575 ^ n42470 ;
  assign n42577 = n42576 ^ n1184 ;
  assign n42578 = n42466 & ~n42577 ;
  assign n42579 = n42578 ^ n42465 ;
  assign n42580 = n42579 ^ n42463 ;
  assign n42581 = ~n42464 & n42580 ;
  assign n42583 = n42582 ^ n42581 ;
  assign n42584 = n42459 & ~n42583 ;
  assign n42585 = n42584 ^ n42458 ;
  assign n42586 = n42585 ^ n42450 ;
  assign n42587 = ~n42454 & n42586 ;
  assign n42588 = n42587 ^ n42453 ;
  assign n42589 = n42588 ^ n42447 ;
  assign n42590 = n42449 & ~n42589 ;
  assign n42591 = n42590 ^ n42448 ;
  assign n42592 = n42591 ^ n42442 ;
  assign n42593 = n42444 & ~n42592 ;
  assign n42594 = n42593 ^ n42443 ;
  assign n42595 = n42594 ^ n42437 ;
  assign n42596 = ~n42439 & ~n42595 ;
  assign n42597 = n42596 ^ n42438 ;
  assign n42598 = n42597 ^ n42433 ;
  assign n42599 = n42434 & ~n42598 ;
  assign n42622 = n42621 ^ n42599 ;
  assign n42627 = n42626 ^ n42622 ;
  assign n42632 = n42597 ^ n42434 ;
  assign n42628 = n42016 ^ n40450 ;
  assign n42629 = n40488 ^ n40450 ;
  assign n42630 = n42628 & ~n42629 ;
  assign n42631 = n42630 ^ n40488 ;
  assign n42633 = n42632 ^ n42631 ;
  assign n42635 = n41931 ^ n41007 ;
  assign n42636 = n41931 ^ n40522 ;
  assign n42637 = n42635 & ~n42636 ;
  assign n42638 = n42637 ^ n40522 ;
  assign n42658 = n42638 ^ n42631 ;
  assign n42634 = n42594 ^ n42439 ;
  assign n42639 = n42638 ^ n42634 ;
  assign n42641 = n42588 ^ n42449 ;
  assign n42642 = n41132 ^ n40514 ;
  assign n42643 = n41132 ^ n40999 ;
  assign n42644 = n42642 & n42643 ;
  assign n42645 = n42644 ^ n40514 ;
  assign n42646 = n42641 & n42645 ;
  assign n42640 = n42591 ^ n42444 ;
  assign n42647 = n42646 ^ n42640 ;
  assign n42648 = n41893 ^ n41125 ;
  assign n42649 = n42646 ^ n40494 ;
  assign n42650 = n42649 ^ n41125 ;
  assign n42651 = n42650 ^ n42646 ;
  assign n42652 = ~n42648 & n42651 ;
  assign n42653 = n42652 ^ n42649 ;
  assign n42654 = n42647 & ~n42653 ;
  assign n42655 = n42654 ^ n42646 ;
  assign n42656 = n42655 ^ n42634 ;
  assign n42657 = n42639 & n42656 ;
  assign n42659 = n42658 ^ n42657 ;
  assign n42660 = ~n42633 & n42659 ;
  assign n42661 = n42660 ^ n42632 ;
  assign n42662 = n42661 ^ n42622 ;
  assign n42663 = n42627 & n42662 ;
  assign n42664 = n42663 ^ n42626 ;
  assign n42666 = n42665 ^ n42664 ;
  assign n42667 = n42166 ^ n41106 ;
  assign n42668 = n42665 ^ n40451 ;
  assign n42669 = n42668 ^ n42166 ;
  assign n42670 = n42669 ^ n42665 ;
  assign n42671 = n42667 & ~n42670 ;
  assign n42672 = n42671 ^ n42668 ;
  assign n42673 = n42666 & ~n42672 ;
  assign n42675 = n42674 ^ n42673 ;
  assign n42676 = ~n42065 & ~n42675 ;
  assign n42677 = n42676 ^ n42064 ;
  assign n42052 = n41088 ^ n40454 ;
  assign n42054 = n42053 ^ n41088 ;
  assign n42055 = ~n42052 & ~n42054 ;
  assign n42056 = n42055 ^ n40454 ;
  assign n42057 = n42056 ^ n42046 ;
  assign n42058 = n42057 ^ n42056 ;
  assign n42678 = n42677 ^ n42058 ;
  assign n42679 = n42051 & n42678 ;
  assign n42680 = n42679 ^ n42057 ;
  assign n42686 = n41992 ^ n41987 ;
  assign n42681 = n41078 ^ n40550 ;
  assign n42682 = n42138 ^ n41078 ;
  assign n42683 = n42681 & ~n42682 ;
  assign n42684 = n42683 ^ n40550 ;
  assign n42687 = n42686 ^ n42684 ;
  assign n42685 = n42684 ^ n42056 ;
  assign n42688 = n42687 ^ n42685 ;
  assign n42689 = ~n42680 & ~n42688 ;
  assign n42690 = n42689 ^ n42685 ;
  assign n42696 = n41994 ^ n41969 ;
  assign n42691 = n41324 ^ n40560 ;
  assign n42692 = n42203 ^ n40560 ;
  assign n42693 = ~n42691 & n42692 ;
  assign n42694 = n42693 ^ n41324 ;
  assign n42695 = n42694 ^ n42684 ;
  assign n42697 = n42696 ^ n42695 ;
  assign n42698 = n42697 ^ n42694 ;
  assign n42699 = ~n42690 & ~n42698 ;
  assign n42700 = n42699 ^ n42695 ;
  assign n42702 = n42701 ^ n42694 ;
  assign n42703 = n42700 & n42702 ;
  assign n42709 = n42708 ^ n42703 ;
  assign n42710 = n42000 ^ n41959 ;
  assign n42711 = n42710 ^ n42707 ;
  assign n42712 = ~n42709 & ~n42711 ;
  assign n42714 = n42713 ^ n42712 ;
  assign n42715 = n42042 & ~n42714 ;
  assign n42716 = n42715 ^ n42041 ;
  assign n42717 = n42716 ^ n42029 ;
  assign n42718 = ~n42035 & n42717 ;
  assign n42719 = n42718 ^ n42034 ;
  assign n42831 = n42720 ^ n42719 ;
  assign n42832 = ~n42725 & ~n42831 ;
  assign n42833 = n42832 ^ n42724 ;
  assign n42841 = n42833 ^ n42825 ;
  assign n42842 = ~n42830 & ~n42841 ;
  assign n42848 = n42847 ^ n42842 ;
  assign n42850 = n42849 ^ n42848 ;
  assign n42851 = n42850 ^ n39396 ;
  assign n42834 = n42833 ^ n42830 ;
  assign n42835 = n42834 ^ n39407 ;
  assign n42728 = n42716 ^ n42035 ;
  assign n42729 = n42728 ^ n39421 ;
  assign n42730 = n42714 ^ n42036 ;
  assign n42731 = n42730 ^ n39423 ;
  assign n42732 = n42710 ^ n42709 ;
  assign n42733 = n42732 ^ n39430 ;
  assign n42734 = n42701 ^ n42700 ;
  assign n42735 = n42734 ^ n39437 ;
  assign n42778 = n42696 ^ n42690 ;
  assign n42736 = n42686 ^ n42680 ;
  assign n42737 = n42736 ^ n39793 ;
  assign n42738 = n42677 ^ n42051 ;
  assign n42739 = n42738 ^ n39789 ;
  assign n42767 = n42675 ^ n42059 ;
  assign n42740 = n42672 ^ n42664 ;
  assign n42741 = n42740 ^ n39774 ;
  assign n42742 = n42661 ^ n42627 ;
  assign n42743 = n42742 ^ n39448 ;
  assign n42744 = n42659 ^ n42632 ;
  assign n42745 = n42744 ^ n39451 ;
  assign n42753 = n42655 ^ n42639 ;
  assign n42746 = n42645 ^ n42641 ;
  assign n42747 = ~n38840 & n42746 ;
  assign n42748 = n42747 ^ n39465 ;
  assign n42749 = n42653 ^ n42640 ;
  assign n42750 = n42749 ^ n42747 ;
  assign n42751 = ~n42748 & n42750 ;
  assign n42752 = n42751 ^ n39465 ;
  assign n42754 = n42753 ^ n42752 ;
  assign n42755 = n42753 ^ n39459 ;
  assign n42756 = n42754 & ~n42755 ;
  assign n42757 = n42756 ^ n39459 ;
  assign n42758 = n42757 ^ n42744 ;
  assign n42759 = ~n42745 & n42758 ;
  assign n42760 = n42759 ^ n39451 ;
  assign n42761 = n42760 ^ n42742 ;
  assign n42762 = n42743 & ~n42761 ;
  assign n42763 = n42762 ^ n39448 ;
  assign n42764 = n42763 ^ n42740 ;
  assign n42765 = ~n42741 & ~n42764 ;
  assign n42766 = n42765 ^ n39774 ;
  assign n42768 = n42767 ^ n42766 ;
  assign n42769 = n42767 ^ n39784 ;
  assign n42770 = n42768 & ~n42769 ;
  assign n42771 = n42770 ^ n39784 ;
  assign n42772 = n42771 ^ n42738 ;
  assign n42773 = ~n42739 & n42772 ;
  assign n42774 = n42773 ^ n39789 ;
  assign n42775 = n42774 ^ n42736 ;
  assign n42776 = n42737 & ~n42775 ;
  assign n42777 = n42776 ^ n39793 ;
  assign n42779 = n42778 ^ n42777 ;
  assign n42780 = n42778 ^ n39803 ;
  assign n42781 = n42779 & n42780 ;
  assign n42782 = n42781 ^ n39803 ;
  assign n42783 = n42782 ^ n42734 ;
  assign n42784 = ~n42735 & ~n42783 ;
  assign n42785 = n42784 ^ n39437 ;
  assign n42786 = n42785 ^ n42732 ;
  assign n42787 = n42733 & n42786 ;
  assign n42788 = n42787 ^ n39430 ;
  assign n42789 = n42788 ^ n42730 ;
  assign n42790 = n42731 & ~n42789 ;
  assign n42791 = n42790 ^ n39423 ;
  assign n42792 = n42791 ^ n42728 ;
  assign n42793 = ~n42729 & ~n42792 ;
  assign n42794 = n42793 ^ n39421 ;
  assign n42726 = n42725 ^ n42719 ;
  assign n42820 = n42794 ^ n42726 ;
  assign n42821 = n42794 ^ n39414 ;
  assign n42822 = n42820 & ~n42821 ;
  assign n42823 = n42822 ^ n39414 ;
  assign n42838 = n42834 ^ n42823 ;
  assign n42839 = ~n42835 & n42838 ;
  assign n42840 = n42839 ^ n39407 ;
  assign n42852 = n42851 ^ n42840 ;
  assign n42727 = n42726 ^ n39414 ;
  assign n42795 = n42794 ^ n42727 ;
  assign n42796 = n42782 ^ n42735 ;
  assign n42797 = n42780 ^ n42777 ;
  assign n42798 = n42760 ^ n42743 ;
  assign n42799 = n42755 ^ n42752 ;
  assign n42800 = n42757 ^ n42745 ;
  assign n42801 = ~n42799 & ~n42800 ;
  assign n42802 = n42798 & n42801 ;
  assign n42803 = n42763 ^ n42741 ;
  assign n42804 = ~n42802 & n42803 ;
  assign n42805 = n42769 ^ n42766 ;
  assign n42806 = ~n42804 & n42805 ;
  assign n42807 = n42771 ^ n42739 ;
  assign n42808 = n42806 & n42807 ;
  assign n42809 = n42774 ^ n42737 ;
  assign n42810 = ~n42808 & n42809 ;
  assign n42811 = n42797 & n42810 ;
  assign n42812 = ~n42796 & ~n42811 ;
  assign n42813 = n42785 ^ n42733 ;
  assign n42814 = n42812 & ~n42813 ;
  assign n42815 = n42788 ^ n42731 ;
  assign n42816 = n42814 & n42815 ;
  assign n42817 = n42791 ^ n42729 ;
  assign n42818 = n42816 & ~n42817 ;
  assign n42819 = n42795 & ~n42818 ;
  assign n42836 = n42835 ^ n42823 ;
  assign n42837 = ~n42819 & ~n42836 ;
  assign n42895 = n42852 ^ n42837 ;
  assign n42892 = n40874 ^ n638 ;
  assign n42893 = n42892 ^ n37083 ;
  assign n42894 = n42893 ^ n30664 ;
  assign n42896 = n42895 ^ n42894 ;
  assign n42897 = n40879 ^ n31998 ;
  assign n42898 = n42897 ^ n37089 ;
  assign n42899 = n42898 ^ n1535 ;
  assign n43017 = n42899 ^ n42895 ;
  assign n42900 = n42836 ^ n42819 ;
  assign n42901 = n42900 ^ n42899 ;
  assign n42905 = n42818 ^ n42795 ;
  assign n42902 = n40884 ^ n32003 ;
  assign n42903 = n42902 ^ n37094 ;
  assign n42904 = n42903 ^ n30670 ;
  assign n42906 = n42905 ^ n42904 ;
  assign n42908 = n40889 ^ n32008 ;
  assign n42909 = n42908 ^ n37098 ;
  assign n42910 = n42909 ^ n30674 ;
  assign n42907 = n42817 ^ n42816 ;
  assign n42911 = n42910 ^ n42907 ;
  assign n42915 = n40895 ^ n32014 ;
  assign n42916 = n42915 ^ n37105 ;
  assign n42917 = n42916 ^ n30679 ;
  assign n42914 = n42815 ^ n42814 ;
  assign n42918 = n42917 ^ n42914 ;
  assign n42919 = n40902 ^ n32019 ;
  assign n42920 = n42919 ^ n37109 ;
  assign n42921 = n42920 ^ n30685 ;
  assign n43006 = n42921 ^ n42914 ;
  assign n42922 = n42813 ^ n42812 ;
  assign n42923 = n42922 ^ n42921 ;
  assign n42927 = n42811 ^ n42796 ;
  assign n42924 = n40906 ^ n32024 ;
  assign n42925 = n42924 ^ n37115 ;
  assign n42926 = n42925 ^ n2378 ;
  assign n42928 = n42927 ^ n42926 ;
  assign n42932 = n42810 ^ n42797 ;
  assign n42929 = n40911 ^ n32029 ;
  assign n42930 = n42929 ^ n2234 ;
  assign n42931 = n42930 ^ n30695 ;
  assign n42933 = n42932 ^ n42931 ;
  assign n42937 = n42809 ^ n42808 ;
  assign n42934 = n40916 ^ n32033 ;
  assign n42935 = n42934 ^ n37122 ;
  assign n42936 = n42935 ^ n2229 ;
  assign n42938 = n42937 ^ n42936 ;
  assign n42941 = n40448 ^ n32040 ;
  assign n42942 = n42941 ^ n37128 ;
  assign n42943 = n42942 ^ n2116 ;
  assign n42940 = n42805 ^ n42804 ;
  assign n42944 = n42943 ^ n42940 ;
  assign n42948 = n42803 ^ n42802 ;
  assign n42945 = n40424 ^ n2007 ;
  assign n42946 = n42945 ^ n37132 ;
  assign n42947 = n42946 ^ n30705 ;
  assign n42949 = n42948 ^ n42947 ;
  assign n42953 = n42801 ^ n42798 ;
  assign n42950 = n32048 ^ n3089 ;
  assign n42951 = n42950 ^ n37137 ;
  assign n42952 = n42951 ^ n30709 ;
  assign n42954 = n42953 ^ n42952 ;
  assign n42955 = n40363 ^ n32052 ;
  assign n42956 = n42955 ^ n36535 ;
  assign n42957 = n42956 ^ n30714 ;
  assign n42958 = n42957 ^ n42800 ;
  assign n42959 = n42958 ^ n42799 ;
  assign n42960 = n40372 ^ n3045 ;
  assign n42961 = n42960 ^ n36491 ;
  assign n42962 = n42961 ^ n30718 ;
  assign n42963 = n42962 ^ n42799 ;
  assign n42969 = n40367 ^ n2782 ;
  assign n42970 = n42969 ^ n35828 ;
  assign n42971 = n42970 ^ n30721 ;
  assign n42964 = n42746 ^ n38840 ;
  assign n42965 = n41244 ^ n2774 ;
  assign n42966 = n42965 ^ n3173 ;
  assign n42967 = n42966 ^ n31059 ;
  assign n42968 = ~n42964 & n42967 ;
  assign n42972 = n42971 ^ n42968 ;
  assign n42973 = n42749 ^ n42748 ;
  assign n42974 = n42973 ^ n42968 ;
  assign n42975 = n42972 & ~n42974 ;
  assign n42976 = n42975 ^ n42971 ;
  assign n42977 = n42976 ^ n42962 ;
  assign n42978 = ~n42963 & ~n42977 ;
  assign n42979 = n42978 ^ n42800 ;
  assign n42980 = ~n42959 & ~n42979 ;
  assign n42981 = n42980 ^ n42957 ;
  assign n42982 = n42981 ^ n42952 ;
  assign n42983 = ~n42954 & ~n42982 ;
  assign n42984 = n42983 ^ n42953 ;
  assign n42985 = n42984 ^ n42947 ;
  assign n42986 = ~n42949 & n42985 ;
  assign n42987 = n42986 ^ n42948 ;
  assign n42988 = n42987 ^ n42943 ;
  assign n42989 = n42944 & ~n42988 ;
  assign n42990 = n42989 ^ n42943 ;
  assign n42994 = n42990 ^ n42937 ;
  assign n42939 = n42807 ^ n42806 ;
  assign n42991 = n42990 ^ n42939 ;
  assign n2097 = n2096 ^ n2072 ;
  assign n2125 = n2124 ^ n2097 ;
  assign n2132 = n2131 ^ n2125 ;
  assign n42992 = n42939 ^ n2132 ;
  assign n42993 = ~n42991 & n42992 ;
  assign n42995 = n42994 ^ n42993 ;
  assign n42996 = ~n42938 & ~n42995 ;
  assign n42997 = n42996 ^ n42937 ;
  assign n42998 = n42997 ^ n42931 ;
  assign n42999 = n42933 & n42998 ;
  assign n43000 = n42999 ^ n42932 ;
  assign n43001 = n43000 ^ n42926 ;
  assign n43002 = ~n42928 & ~n43001 ;
  assign n43003 = n43002 ^ n42927 ;
  assign n43004 = n43003 ^ n42921 ;
  assign n43005 = n42923 & ~n43004 ;
  assign n43007 = n43006 ^ n43005 ;
  assign n43008 = ~n42918 & n43007 ;
  assign n43009 = n43008 ^ n42917 ;
  assign n42912 = n42910 ^ n42905 ;
  assign n42913 = n42912 ^ n42905 ;
  assign n43010 = n43009 ^ n42913 ;
  assign n43011 = n42911 & n43010 ;
  assign n43012 = n43011 ^ n42912 ;
  assign n43013 = ~n42906 & ~n43012 ;
  assign n43014 = n43013 ^ n42905 ;
  assign n43015 = n43014 ^ n42899 ;
  assign n43016 = ~n42901 & ~n43015 ;
  assign n43018 = n43017 ^ n43016 ;
  assign n43019 = n42896 & n43018 ;
  assign n43020 = n43019 ^ n42895 ;
  assign n42861 = n41033 ^ n40773 ;
  assign n42862 = n42102 ^ n41033 ;
  assign n42863 = n42861 & n42862 ;
  assign n42864 = n42863 ^ n40773 ;
  assign n42860 = n42545 ^ n42515 ;
  assign n42865 = n42864 ^ n42860 ;
  assign n42857 = n42849 ^ n42846 ;
  assign n42858 = ~n42848 & ~n42857 ;
  assign n42859 = n42858 ^ n42846 ;
  assign n42866 = n42865 ^ n42859 ;
  assign n42867 = n42866 ^ n39840 ;
  assign n42854 = n42850 ^ n42840 ;
  assign n42855 = ~n42851 & ~n42854 ;
  assign n42856 = n42855 ^ n39396 ;
  assign n42868 = n42867 ^ n42856 ;
  assign n42853 = n42837 & ~n42852 ;
  assign n42887 = n42868 ^ n42853 ;
  assign n42891 = n42890 ^ n42887 ;
  assign n43061 = n43020 ^ n42891 ;
  assign n44268 = n44267 ^ n43061 ;
  assign n43086 = n42556 ^ n42493 ;
  assign n44035 = n43086 ^ n42108 ;
  assign n43076 = n43012 ^ n42904 ;
  assign n44036 = n44035 ^ n43076 ;
  assign n43815 = n41752 ^ n2200 ;
  assign n43816 = n43815 ^ n37733 ;
  assign n43817 = n43816 ^ n2333 ;
  assign n43439 = n41931 ^ n41132 ;
  assign n43440 = n43439 ^ n42665 ;
  assign n43413 = n40815 ^ n32523 ;
  assign n43414 = n43413 ^ n37046 ;
  assign n43415 = n43414 ^ n30639 ;
  assign n43037 = n42089 ^ n41023 ;
  assign n43038 = n41023 ^ n40808 ;
  assign n43039 = n43037 & n43038 ;
  assign n43040 = n43039 ^ n40808 ;
  assign n43036 = n42551 ^ n42505 ;
  assign n43041 = n43040 ^ n43036 ;
  assign n42874 = n42092 ^ n41027 ;
  assign n42875 = n41027 ^ n40787 ;
  assign n42876 = n42874 & ~n42875 ;
  assign n42877 = n42876 ^ n40787 ;
  assign n42873 = n42547 ^ n42512 ;
  assign n42878 = n42877 ^ n42873 ;
  assign n42870 = n42860 ^ n42859 ;
  assign n42871 = n42865 & n42870 ;
  assign n42872 = n42871 ^ n42864 ;
  assign n43033 = n42873 ^ n42872 ;
  assign n43034 = ~n42878 & n43033 ;
  assign n43035 = n43034 ^ n42877 ;
  assign n43042 = n43041 ^ n43035 ;
  assign n43043 = n43042 ^ n39385 ;
  assign n42879 = n42878 ^ n42872 ;
  assign n42880 = n42879 ^ n39387 ;
  assign n42881 = n42866 ^ n42856 ;
  assign n42882 = ~n42867 & n42881 ;
  assign n42883 = n42882 ^ n39840 ;
  assign n43030 = n42883 ^ n42879 ;
  assign n43031 = n42880 & n43030 ;
  assign n43032 = n43031 ^ n39387 ;
  assign n43254 = n43042 ^ n43032 ;
  assign n43255 = ~n43043 & n43254 ;
  assign n43256 = n43255 ^ n39385 ;
  assign n43154 = n42235 ^ n41016 ;
  assign n43155 = n43036 ^ n43035 ;
  assign n43156 = n43041 & ~n43155 ;
  assign n43157 = n43156 ^ n43040 ;
  assign n43158 = n43157 ^ n40829 ;
  assign n43159 = n43158 ^ n42235 ;
  assign n43160 = n43159 ^ n43157 ;
  assign n43161 = n43154 & n43160 ;
  assign n43162 = n43161 ^ n43158 ;
  assign n43091 = n42553 ^ n42500 ;
  assign n43252 = n43162 ^ n43091 ;
  assign n43253 = n43252 ^ n39368 ;
  assign n43300 = n43256 ^ n43253 ;
  assign n43044 = n43043 ^ n43032 ;
  assign n42869 = n42853 & n42868 ;
  assign n42884 = n42883 ^ n42880 ;
  assign n43045 = ~n42869 & n42884 ;
  assign n43301 = ~n43044 & ~n43045 ;
  assign n43302 = n43300 & n43301 ;
  assign n43163 = n41374 ^ n41041 ;
  assign n43164 = n42083 ^ n41374 ;
  assign n43165 = ~n43163 & n43164 ;
  assign n43166 = n43165 ^ n41041 ;
  assign n43168 = n43166 ^ n43091 ;
  assign n43167 = n43166 ^ n43157 ;
  assign n43169 = n43168 ^ n43167 ;
  assign n43170 = n43162 & n43169 ;
  assign n43171 = n43170 ^ n43168 ;
  assign n43251 = n43171 ^ n43086 ;
  assign n43303 = n43251 ^ n39853 ;
  assign n43257 = n43256 ^ n43252 ;
  assign n43258 = n43253 & ~n43257 ;
  assign n43259 = n43258 ^ n39368 ;
  assign n43304 = n43303 ^ n43259 ;
  assign n43305 = ~n43302 & ~n43304 ;
  assign n43260 = n43259 ^ n43251 ;
  assign n43261 = n43259 ^ n39853 ;
  assign n43262 = n43260 & ~n43261 ;
  assign n43263 = n43262 ^ n39853 ;
  assign n43306 = n43263 ^ n40274 ;
  assign n43182 = n41379 ^ n41035 ;
  assign n43183 = n42067 ^ n41379 ;
  assign n43184 = ~n43182 & n43183 ;
  assign n43185 = n43184 ^ n41035 ;
  assign n43172 = n42558 ^ n42490 ;
  assign n43174 = n43172 ^ n43166 ;
  assign n43173 = n43172 ^ n43086 ;
  assign n43175 = n43174 ^ n43173 ;
  assign n43176 = n43171 & n43175 ;
  assign n43177 = n43176 ^ n43173 ;
  assign n43249 = n43185 ^ n43177 ;
  assign n43307 = n43306 ^ n43249 ;
  assign n43308 = n43305 & ~n43307 ;
  assign n43178 = n41588 ^ n41025 ;
  assign n43179 = n42251 ^ n41588 ;
  assign n43180 = n43178 & n43179 ;
  assign n43181 = n43180 ^ n41025 ;
  assign n43187 = n43181 ^ n43172 ;
  assign n43186 = n43185 ^ n43181 ;
  assign n43188 = n43187 ^ n43186 ;
  assign n43189 = ~n43177 & ~n43188 ;
  assign n43190 = n43189 ^ n43187 ;
  assign n43081 = n42561 ^ n42485 ;
  assign n43268 = n43190 ^ n43081 ;
  assign n43250 = n43249 ^ n40274 ;
  assign n43264 = n43263 ^ n43249 ;
  assign n43265 = ~n43250 & ~n43264 ;
  assign n43266 = n43265 ^ n40274 ;
  assign n43267 = n43266 ^ n40323 ;
  assign n43309 = n43268 ^ n43267 ;
  assign n43310 = n43308 & ~n43309 ;
  assign n43191 = n41832 ^ n41019 ;
  assign n43192 = n42356 ^ n41832 ;
  assign n43193 = n43191 & ~n43192 ;
  assign n43194 = n43193 ^ n41019 ;
  assign n43196 = n43194 ^ n43181 ;
  assign n43195 = n43194 ^ n43081 ;
  assign n43197 = n43196 ^ n43195 ;
  assign n43198 = ~n43190 & n43197 ;
  assign n43199 = n43198 ^ n43196 ;
  assign n43248 = n43199 ^ n43074 ;
  assign n43311 = n43248 ^ n40401 ;
  assign n43269 = n43268 ^ n43266 ;
  assign n43270 = ~n43267 & n43269 ;
  assign n43271 = n43270 ^ n40323 ;
  assign n43312 = n43311 ^ n43271 ;
  assign n43313 = ~n43310 & n43312 ;
  assign n43272 = n43271 ^ n43248 ;
  assign n43273 = n43271 ^ n40401 ;
  assign n43274 = n43272 & n43273 ;
  assign n43275 = n43274 ^ n40401 ;
  assign n43200 = n40989 ^ n40296 ;
  assign n43201 = n42375 ^ n40989 ;
  assign n43202 = n43200 & ~n43201 ;
  assign n43203 = n43202 ^ n40296 ;
  assign n43205 = n43203 ^ n43194 ;
  assign n43204 = n43203 ^ n43074 ;
  assign n43206 = n43205 ^ n43204 ;
  assign n43207 = n43199 & n43206 ;
  assign n43208 = n43207 ^ n43205 ;
  assign n43069 = n42567 ^ n42478 ;
  assign n43246 = n43208 ^ n43069 ;
  assign n43247 = n43246 ^ n39678 ;
  assign n43314 = n43275 ^ n43247 ;
  assign n43315 = n43313 & n43314 ;
  assign n43209 = n41260 ^ n40298 ;
  assign n43210 = n42604 ^ n41260 ;
  assign n43211 = ~n43209 & n43210 ;
  assign n43212 = n43211 ^ n40298 ;
  assign n43214 = n43212 ^ n43203 ;
  assign n43213 = n43212 ^ n43069 ;
  assign n43215 = n43214 ^ n43213 ;
  assign n43216 = ~n43208 & ~n43215 ;
  assign n43217 = n43216 ^ n43214 ;
  assign n43064 = n42570 ^ n42473 ;
  assign n43245 = n43217 ^ n43064 ;
  assign n43298 = n43245 ^ n39677 ;
  assign n43276 = n43275 ^ n43246 ;
  assign n43277 = ~n43247 & ~n43276 ;
  assign n43278 = n43277 ^ n39678 ;
  assign n43299 = n43298 ^ n43278 ;
  assign n43363 = n43315 ^ n43299 ;
  assign n43360 = n40839 ^ n32527 ;
  assign n43361 = n43360 ^ n37055 ;
  assign n43362 = n43361 ^ n2828 ;
  assign n43364 = n43363 ^ n43362 ;
  assign n43368 = n43314 ^ n43313 ;
  assign n43372 = n43371 ^ n43368 ;
  assign n43374 = n43312 ^ n43310 ;
  assign n1325 = n1285 ^ n1231 ;
  assign n1326 = n1325 ^ n1322 ;
  assign n1333 = n1332 ^ n1326 ;
  assign n43375 = n43374 ^ n1333 ;
  assign n43376 = n43309 ^ n43308 ;
  assign n1289 = n1270 ^ n1213 ;
  assign n1308 = n1307 ^ n1289 ;
  assign n1315 = n1314 ^ n1308 ;
  assign n43377 = n43376 ^ n1315 ;
  assign n43379 = n40851 ^ n1124 ;
  assign n43380 = n43379 ^ n1699 ;
  assign n43381 = n43380 ^ n1299 ;
  assign n43378 = n43307 ^ n43305 ;
  assign n43382 = n43381 ^ n43378 ;
  assign n43383 = n43304 ^ n43302 ;
  assign n1681 = n1674 ^ n1116 ;
  assign n1691 = n1690 ^ n1681 ;
  assign n1695 = n1694 ^ n1691 ;
  assign n43384 = n43383 ^ n1695 ;
  assign n43388 = n43301 ^ n43300 ;
  assign n43385 = n40857 ^ n1657 ;
  assign n43386 = n43385 ^ n37071 ;
  assign n43387 = n43386 ^ n1688 ;
  assign n43389 = n43388 ^ n43387 ;
  assign n43046 = n43045 ^ n43044 ;
  assign n43027 = n40862 ^ n1648 ;
  assign n43028 = n43027 ^ n37067 ;
  assign n43029 = n43028 ^ n791 ;
  assign n43047 = n43046 ^ n43029 ;
  assign n42885 = n42884 ^ n42869 ;
  assign n2988 = n2987 ^ n2984 ;
  assign n2989 = n2988 ^ n722 ;
  assign n2993 = n2992 ^ n2989 ;
  assign n42886 = n42885 ^ n2993 ;
  assign n43023 = n42890 ^ n42885 ;
  assign n43021 = n43020 ^ n42890 ;
  assign n43022 = ~n42891 & n43021 ;
  assign n43024 = n43023 ^ n43022 ;
  assign n43025 = ~n42886 & ~n43024 ;
  assign n43026 = n43025 ^ n42885 ;
  assign n43390 = n43029 ^ n43026 ;
  assign n43391 = ~n43047 & n43390 ;
  assign n43392 = n43391 ^ n43046 ;
  assign n43393 = n43392 ^ n43387 ;
  assign n43394 = ~n43389 & n43393 ;
  assign n43395 = n43394 ^ n43388 ;
  assign n43396 = n43395 ^ n1695 ;
  assign n43397 = n43384 & n43396 ;
  assign n43398 = n43397 ^ n43383 ;
  assign n43399 = n43398 ^ n43381 ;
  assign n43400 = ~n43382 & n43399 ;
  assign n43401 = n43400 ^ n43381 ;
  assign n43402 = n43401 ^ n1315 ;
  assign n43403 = ~n43377 & ~n43402 ;
  assign n43404 = n43403 ^ n43376 ;
  assign n43405 = n43404 ^ n1333 ;
  assign n43406 = n43375 & ~n43405 ;
  assign n43373 = n43368 ^ n1333 ;
  assign n43407 = n43406 ^ n43373 ;
  assign n43408 = ~n43372 & n43407 ;
  assign n43409 = n43408 ^ n43371 ;
  assign n43316 = n43299 & n43315 ;
  assign n43279 = n43278 ^ n43245 ;
  assign n43280 = n43278 ^ n39677 ;
  assign n43281 = ~n43279 & n43280 ;
  assign n43282 = n43281 ^ n39677 ;
  assign n43218 = n41270 ^ n40286 ;
  assign n43219 = n41860 ^ n41270 ;
  assign n43220 = n43218 & ~n43219 ;
  assign n43221 = n43220 ^ n40286 ;
  assign n43223 = n43221 ^ n43212 ;
  assign n43222 = n43221 ^ n43064 ;
  assign n43224 = n43223 ^ n43222 ;
  assign n43225 = ~n43217 & ~n43224 ;
  assign n43226 = n43225 ^ n43223 ;
  assign n43059 = n42573 ^ n42471 ;
  assign n43243 = n43226 ^ n43059 ;
  assign n43244 = n43243 ^ n39669 ;
  assign n43297 = n43282 ^ n43244 ;
  assign n43365 = n43316 ^ n43297 ;
  assign n43366 = n43365 ^ n43362 ;
  assign n43367 = n43366 ^ n43365 ;
  assign n43410 = n43409 ^ n43367 ;
  assign n43411 = ~n43364 & n43410 ;
  assign n43412 = n43411 ^ n43366 ;
  assign n43438 = n43415 ^ n43412 ;
  assign n43561 = n43440 ^ n43438 ;
  assign n43562 = n40514 & n43561 ;
  assign n43685 = n43562 ^ n40494 ;
  assign n43149 = n41257 ^ n40342 ;
  assign n43150 = n41871 ^ n41257 ;
  assign n43151 = ~n43149 & ~n43150 ;
  assign n43152 = n43151 ^ n40342 ;
  assign n43229 = n43221 ^ n43152 ;
  assign n43227 = n43221 ^ n43059 ;
  assign n43228 = n43226 & ~n43227 ;
  assign n43230 = n43229 ^ n43228 ;
  assign n43054 = n42576 ^ n42466 ;
  assign n43242 = n43230 ^ n43054 ;
  assign n43318 = n43242 ^ n39662 ;
  assign n43283 = n43282 ^ n43243 ;
  assign n43284 = ~n43244 & n43283 ;
  assign n43285 = n43284 ^ n39669 ;
  assign n43319 = n43318 ^ n43285 ;
  assign n43317 = ~n43297 & n43316 ;
  assign n43358 = n43319 ^ n43317 ;
  assign n43417 = n43365 ^ n43358 ;
  assign n43416 = n43415 ^ n43358 ;
  assign n43418 = n43417 ^ n43416 ;
  assign n43419 = ~n43412 & n43418 ;
  assign n43420 = n43419 ^ n43416 ;
  assign n43355 = n40988 ^ n32518 ;
  assign n43356 = n43355 ^ n37050 ;
  assign n43357 = n43356 ^ n2651 ;
  assign n43446 = n43420 ^ n43357 ;
  assign n43443 = n42016 ^ n41125 ;
  assign n43444 = n43443 ^ n42059 ;
  assign n43441 = n43438 & n43440 ;
  assign n43445 = n43444 ^ n43441 ;
  assign n43563 = n43446 ^ n43445 ;
  assign n43686 = n43685 ^ n43563 ;
  assign n43564 = n43563 ^ n43562 ;
  assign n43565 = n43563 ^ n40494 ;
  assign n43566 = n43564 & n43565 ;
  assign n43567 = n43566 ^ n40494 ;
  assign n43447 = n43446 ^ n43441 ;
  assign n43448 = ~n43445 & n43447 ;
  assign n43359 = n43358 ^ n43357 ;
  assign n43421 = n43359 & n43420 ;
  assign n43422 = n43421 ^ n43358 ;
  assign n43351 = n41212 ^ n32512 ;
  assign n43352 = n43351 ^ n37392 ;
  assign n43353 = n43352 ^ n30857 ;
  assign n43320 = ~n43317 & ~n43319 ;
  assign n43153 = n43152 ^ n43054 ;
  assign n43231 = ~n43153 & ~n43230 ;
  assign n43232 = n43231 ^ n43054 ;
  assign n43140 = n41857 ^ n41247 ;
  assign n43050 = n42579 ^ n42464 ;
  assign n43141 = n43050 ^ n40414 ;
  assign n43142 = n43141 ^ n41857 ;
  assign n43143 = n43142 ^ n43050 ;
  assign n43144 = ~n43140 & ~n43143 ;
  assign n43145 = n43144 ^ n43141 ;
  assign n43290 = n43232 ^ n43145 ;
  assign n43292 = n43290 ^ n39721 ;
  assign n43286 = n43285 ^ n43242 ;
  assign n43287 = n43285 ^ n39662 ;
  assign n43288 = n43286 & ~n43287 ;
  assign n43289 = n43288 ^ n39662 ;
  assign n43296 = n43292 ^ n43289 ;
  assign n43350 = n43320 ^ n43296 ;
  assign n43354 = n43353 ^ n43350 ;
  assign n43436 = n43422 ^ n43354 ;
  assign n43442 = n43441 ^ n43436 ;
  assign n43449 = n43448 ^ n43442 ;
  assign n43434 = n42178 ^ n41007 ;
  assign n43435 = n43434 ^ n42046 ;
  assign n43559 = n43449 ^ n43435 ;
  assign n43560 = n43559 ^ n40522 ;
  assign n43687 = n43567 ^ n43560 ;
  assign n43688 = ~n43686 & n43687 ;
  assign n43568 = n43567 ^ n43559 ;
  assign n43569 = n43560 & ~n43568 ;
  assign n43570 = n43569 ^ n40522 ;
  assign n43437 = n43436 ^ n43435 ;
  assign n43450 = ~n43437 & ~n43449 ;
  assign n43451 = n43450 ^ n43436 ;
  assign n43431 = n42166 ^ n40450 ;
  assign n43432 = n43431 ^ n42686 ;
  assign n43423 = n43422 ^ n43353 ;
  assign n43424 = ~n43354 & n43423 ;
  assign n43425 = n43424 ^ n43353 ;
  assign n43321 = ~n43296 & n43320 ;
  assign n43291 = n43290 ^ n43289 ;
  assign n43293 = ~n43291 & ~n43292 ;
  assign n43294 = n43293 ^ n39721 ;
  assign n43236 = n41145 ^ n40432 ;
  assign n43237 = n41847 ^ n41145 ;
  assign n43238 = n43236 & n43237 ;
  assign n43239 = n43238 ^ n40432 ;
  assign n43146 = n42583 ^ n42458 ;
  assign n43147 = n43146 ^ n43050 ;
  assign n43148 = n43147 ^ n43146 ;
  assign n43233 = n43232 ^ n43148 ;
  assign n43234 = n43145 & ~n43233 ;
  assign n43235 = n43234 ^ n43147 ;
  assign n43240 = n43239 ^ n43235 ;
  assign n43241 = n43240 ^ n39472 ;
  assign n43295 = n43294 ^ n43241 ;
  assign n43348 = n43321 ^ n43295 ;
  assign n43336 = n41206 ^ n3143 ;
  assign n43337 = n43336 ^ n37387 ;
  assign n43338 = n43337 ^ n30900 ;
  assign n43349 = n43348 ^ n43338 ;
  assign n43430 = n43425 ^ n43349 ;
  assign n43433 = n43432 ^ n43430 ;
  assign n43557 = n43451 ^ n43433 ;
  assign n43558 = n43557 ^ n40488 ;
  assign n43689 = n43570 ^ n43558 ;
  assign n43690 = ~n43688 & ~n43689 ;
  assign n43571 = n43570 ^ n43557 ;
  assign n43572 = n43558 & n43571 ;
  assign n43573 = n43572 ^ n40488 ;
  assign n43426 = n43425 ^ n43338 ;
  assign n43427 = ~n43349 & n43426 ;
  assign n43343 = n41138 ^ n40509 ;
  assign n43344 = n41845 ^ n41138 ;
  assign n43345 = n43343 & ~n43344 ;
  assign n43333 = n41153 ^ n32501 ;
  assign n43334 = n43333 ^ n37373 ;
  assign n43335 = n43334 ^ n3171 ;
  assign n43339 = n43338 ^ n43335 ;
  assign n43331 = n39739 ^ n39472 ;
  assign n43328 = n42585 ^ n42454 ;
  assign n43329 = n43328 ^ n40509 ;
  assign n43330 = n43329 ^ n43146 ;
  assign n43332 = n43331 ^ n43330 ;
  assign n43340 = n43339 ^ n43332 ;
  assign n43326 = n43239 ^ n43146 ;
  assign n43327 = ~n43235 & ~n43326 ;
  assign n43341 = n43340 ^ n43327 ;
  assign n43323 = n43294 ^ n43240 ;
  assign n43324 = n43294 ^ n39472 ;
  assign n43325 = n43323 & ~n43324 ;
  assign n43342 = n43341 ^ n43325 ;
  assign n43346 = n43345 ^ n43342 ;
  assign n43322 = ~n43295 & n43321 ;
  assign n43347 = n43346 ^ n43322 ;
  assign n43428 = n43427 ^ n43347 ;
  assign n43454 = n43430 ^ n43428 ;
  assign n43452 = n43451 ^ n43430 ;
  assign n43453 = ~n43433 & n43452 ;
  assign n43455 = n43454 ^ n43453 ;
  assign n43138 = n42060 ^ n41112 ;
  assign n43139 = n43138 ^ n42696 ;
  assign n43555 = n43455 ^ n43139 ;
  assign n43556 = n43555 ^ n40478 ;
  assign n43691 = n43573 ^ n43556 ;
  assign n43692 = ~n43690 & ~n43691 ;
  assign n43429 = n43428 ^ n43139 ;
  assign n43456 = ~n43429 & n43455 ;
  assign n43457 = n43456 ^ n43428 ;
  assign n43136 = n42967 ^ n42964 ;
  assign n43134 = n42044 ^ n41106 ;
  assign n43135 = n43134 ^ n42701 ;
  assign n43137 = n43136 ^ n43135 ;
  assign n43554 = n43457 ^ n43137 ;
  assign n43693 = n43554 ^ n40451 ;
  assign n43574 = n43573 ^ n43555 ;
  assign n43575 = n43556 & ~n43574 ;
  assign n43576 = n43575 ^ n40478 ;
  assign n43694 = n43693 ^ n43576 ;
  assign n43695 = ~n43692 & ~n43694 ;
  assign n43577 = n43576 ^ n43554 ;
  assign n43578 = n43576 ^ n40451 ;
  assign n43579 = ~n43577 & ~n43578 ;
  assign n43580 = n43579 ^ n40451 ;
  assign n43458 = n43457 ^ n43136 ;
  assign n43459 = ~n43137 & n43458 ;
  assign n43460 = n43459 ^ n43136 ;
  assign n43132 = n42973 ^ n42972 ;
  assign n43130 = n42710 ^ n42053 ;
  assign n43131 = n43130 ^ n41096 ;
  assign n43133 = n43132 ^ n43131 ;
  assign n43552 = n43460 ^ n43133 ;
  assign n43553 = n43552 ^ n40466 ;
  assign n43696 = n43580 ^ n43553 ;
  assign n43697 = ~n43695 & ~n43696 ;
  assign n43461 = n43460 ^ n43131 ;
  assign n43462 = ~n43133 & ~n43461 ;
  assign n43463 = n43462 ^ n43132 ;
  assign n43127 = n42138 ^ n41090 ;
  assign n43128 = n43127 ^ n42036 ;
  assign n43126 = n42976 ^ n42963 ;
  assign n43129 = n43128 ^ n43126 ;
  assign n43584 = n43463 ^ n43129 ;
  assign n43698 = n43584 ^ n40460 ;
  assign n43581 = n43580 ^ n43552 ;
  assign n43582 = ~n43553 & n43581 ;
  assign n43583 = n43582 ^ n40466 ;
  assign n43699 = n43698 ^ n43583 ;
  assign n43700 = n43697 & ~n43699 ;
  assign n43585 = n43584 ^ n43583 ;
  assign n43464 = n43463 ^ n43126 ;
  assign n43465 = n43129 & n43464 ;
  assign n43466 = n43465 ^ n43128 ;
  assign n43121 = n42203 ^ n41088 ;
  assign n43122 = n43121 ^ n42029 ;
  assign n43120 = n42979 ^ n42957 ;
  assign n43123 = n43122 ^ n43120 ;
  assign n43550 = n43466 ^ n43123 ;
  assign n43586 = n43550 ^ n40460 ;
  assign n43587 = n43586 ^ n43583 ;
  assign n43588 = n43587 ^ n43550 ;
  assign n43589 = n43585 & n43588 ;
  assign n43590 = n43589 ^ n43586 ;
  assign n43684 = n43590 ^ n40454 ;
  assign n43814 = n43700 ^ n43684 ;
  assign n43818 = n43817 ^ n43814 ;
  assign n43824 = n43699 ^ n43697 ;
  assign n43821 = n41702 ^ n2185 ;
  assign n43822 = n43821 ^ n37686 ;
  assign n43823 = n43822 ^ n31418 ;
  assign n43825 = n43824 ^ n43823 ;
  assign n43826 = n41708 ^ n33124 ;
  assign n43827 = n43826 ^ n37691 ;
  assign n43828 = n43827 ^ n31423 ;
  assign n43878 = n43828 ^ n43824 ;
  assign n43829 = n43696 ^ n43695 ;
  assign n43830 = n43829 ^ n43828 ;
  assign n43834 = n43694 ^ n43692 ;
  assign n43831 = n41738 ^ n33128 ;
  assign n43832 = n43831 ^ n37720 ;
  assign n43833 = n43832 ^ n31428 ;
  assign n43835 = n43834 ^ n43833 ;
  assign n43837 = n41712 ^ n33134 ;
  assign n43838 = n43837 ^ n37695 ;
  assign n43839 = n43838 ^ n31435 ;
  assign n43872 = n43839 ^ n43834 ;
  assign n43836 = n43691 ^ n43690 ;
  assign n43840 = n43839 ^ n43836 ;
  assign n43844 = n43689 ^ n43688 ;
  assign n43841 = n41717 ^ n33138 ;
  assign n43842 = n43841 ^ n37700 ;
  assign n43843 = n43842 ^ n1895 ;
  assign n43845 = n43844 ^ n43843 ;
  assign n43847 = n41721 ^ n33147 ;
  assign n43848 = n43847 ^ n37704 ;
  assign n43849 = n43848 ^ n30821 ;
  assign n43846 = n43687 ^ n43686 ;
  assign n43850 = n43849 ^ n43846 ;
  assign n43857 = n43561 ^ n40514 ;
  assign n43858 = n43856 & n43857 ;
  assign n43851 = n40998 ^ n33142 ;
  assign n43852 = n43851 ^ n37247 ;
  assign n43853 = n43852 ^ n3236 ;
  assign n43859 = n43858 ^ n43853 ;
  assign n44055 = n43853 ^ n43686 ;
  assign n43863 = ~n43859 & ~n44055 ;
  assign n43860 = n43849 ^ n43686 ;
  assign n43864 = n43863 ^ n43860 ;
  assign n43865 = n43850 & ~n43864 ;
  assign n43866 = n43865 ^ n43849 ;
  assign n43867 = n43866 ^ n43843 ;
  assign n43868 = n43845 & ~n43867 ;
  assign n43869 = n43868 ^ n43844 ;
  assign n43870 = n43869 ^ n43839 ;
  assign n43871 = ~n43840 & n43870 ;
  assign n43873 = n43872 ^ n43871 ;
  assign n43874 = n43835 & n43873 ;
  assign n43875 = n43874 ^ n43834 ;
  assign n43876 = n43875 ^ n43828 ;
  assign n43877 = ~n43830 & n43876 ;
  assign n43879 = n43878 ^ n43877 ;
  assign n43880 = n43825 & n43879 ;
  assign n43881 = n43880 ^ n43824 ;
  assign n43882 = n43881 ^ n43817 ;
  assign n43883 = n43818 & n43882 ;
  assign n43467 = n43466 ^ n43120 ;
  assign n43468 = n43123 & ~n43467 ;
  assign n43118 = n42981 ^ n42954 ;
  assign n43124 = n43120 ^ n43118 ;
  assign n43469 = n43468 ^ n43124 ;
  assign n43116 = n42132 ^ n41078 ;
  assign n43117 = n43116 ^ n42720 ;
  assign n43549 = n43469 ^ n43117 ;
  assign n43702 = n43549 ^ n40550 ;
  assign n43551 = n43550 ^ n40454 ;
  assign n43591 = ~n43551 & ~n43590 ;
  assign n43592 = n43591 ^ n40454 ;
  assign n43703 = n43702 ^ n43592 ;
  assign n43701 = ~n43684 & n43700 ;
  assign n43812 = n43703 ^ n43701 ;
  assign n43819 = n43817 ^ n43812 ;
  assign n43884 = n43883 ^ n43819 ;
  assign n2317 = n2310 ^ n2268 ;
  assign n2342 = n2341 ^ n2317 ;
  assign n2349 = n2348 ^ n2342 ;
  assign n44034 = n43884 ^ n2349 ;
  assign n44037 = n44036 ^ n44034 ;
  assign n44043 = n43881 ^ n43818 ;
  assign n44041 = n43091 ^ n42114 ;
  assign n43083 = n43009 ^ n42911 ;
  assign n44042 = n44041 ^ n43083 ;
  assign n44044 = n44043 ^ n44042 ;
  assign n44047 = n43879 ^ n43823 ;
  assign n44045 = n43036 ^ n42120 ;
  assign n43495 = n43007 ^ n42917 ;
  assign n44046 = n44045 ^ n43495 ;
  assign n44048 = n44047 ^ n44046 ;
  assign n44050 = n42873 ^ n42031 ;
  assign n43088 = n43003 ^ n42923 ;
  assign n44051 = n44050 ^ n43088 ;
  assign n44049 = n43875 ^ n43830 ;
  assign n44052 = n44051 ^ n44049 ;
  assign n44152 = n43873 ^ n43833 ;
  assign n44162 = n44152 ^ n44049 ;
  assign n44056 = n44055 ^ n43858 ;
  assign n44053 = n42053 ^ n42029 ;
  assign n43110 = n42987 ^ n42944 ;
  assign n44054 = n44053 ^ n43110 ;
  assign n44057 = n44056 ^ n44054 ;
  assign n44063 = n43857 ^ n43856 ;
  assign n44061 = n42044 ^ n42036 ;
  assign n43114 = n42984 ^ n42949 ;
  assign n44062 = n44061 ^ n43114 ;
  assign n44064 = n44063 ^ n44062 ;
  assign n44077 = n41145 ^ n40999 ;
  assign n44078 = n44077 ^ n42632 ;
  assign n43521 = n43392 ^ n43389 ;
  assign n43519 = n41860 ^ n40989 ;
  assign n43520 = n43519 ^ n43146 ;
  assign n43522 = n43521 ^ n43520 ;
  assign n43652 = n43395 ^ n43384 ;
  assign n43653 = n43652 ^ n43521 ;
  assign n43654 = n43653 ^ n43652 ;
  assign n43049 = n42604 ^ n41832 ;
  assign n43051 = n43050 ^ n43049 ;
  assign n43048 = n43047 ^ n43026 ;
  assign n43052 = n43051 ^ n43048 ;
  assign n43056 = n43024 ^ n2993 ;
  assign n43053 = n42375 ^ n41588 ;
  assign n43055 = n43054 ^ n43053 ;
  assign n43057 = n43056 ^ n43055 ;
  assign n43512 = n43061 ^ n43056 ;
  assign n43058 = n42356 ^ n41379 ;
  assign n43060 = n43059 ^ n43058 ;
  assign n43062 = n43061 ^ n43060 ;
  assign n43066 = n43018 ^ n42894 ;
  assign n43063 = n42251 ^ n41374 ;
  assign n43065 = n43064 ^ n43063 ;
  assign n43067 = n43066 ^ n43065 ;
  assign n43071 = n43014 ^ n42901 ;
  assign n43506 = n43071 ^ n43066 ;
  assign n43068 = n42067 ^ n41016 ;
  assign n43070 = n43069 ^ n43068 ;
  assign n43072 = n43071 ^ n43070 ;
  assign n43073 = n42083 ^ n41023 ;
  assign n43075 = n43074 ^ n43073 ;
  assign n43077 = n43076 ^ n43075 ;
  assign n43080 = n42235 ^ n41027 ;
  assign n43082 = n43081 ^ n43080 ;
  assign n43084 = n43083 ^ n43082 ;
  assign n43498 = n43495 ^ n43083 ;
  assign n43492 = n42089 ^ n41033 ;
  assign n43493 = n43492 ^ n43172 ;
  assign n43085 = n42092 ^ n41040 ;
  assign n43087 = n43086 ^ n43085 ;
  assign n43089 = n43088 ^ n43087 ;
  assign n43093 = n43000 ^ n42928 ;
  assign n43090 = n42102 ^ n41047 ;
  assign n43092 = n43091 ^ n43090 ;
  assign n43094 = n43093 ^ n43092 ;
  assign n43097 = n42108 ^ n41057 ;
  assign n43098 = n43097 ^ n43036 ;
  assign n43095 = n42997 ^ n42933 ;
  assign n43099 = n43098 ^ n43095 ;
  assign n43102 = n42995 ^ n42936 ;
  assign n43100 = n42114 ^ n41063 ;
  assign n43101 = n43100 ^ n42873 ;
  assign n43103 = n43102 ^ n43101 ;
  assign n43106 = n42992 ^ n42990 ;
  assign n43480 = n43106 ^ n43102 ;
  assign n43104 = n42120 ^ n41069 ;
  assign n43105 = n43104 ^ n42860 ;
  assign n43107 = n43106 ^ n43105 ;
  assign n43108 = n42031 ^ n41075 ;
  assign n43109 = n43108 ^ n42849 ;
  assign n43111 = n43110 ^ n43109 ;
  assign n43112 = n42038 ^ n41324 ;
  assign n43113 = n43112 ^ n42825 ;
  assign n43115 = n43114 ^ n43113 ;
  assign n43119 = n43118 ^ n43117 ;
  assign n43470 = ~n43119 & ~n43469 ;
  assign n43471 = n43470 ^ n43118 ;
  assign n43472 = n43471 ^ n43113 ;
  assign n43473 = ~n43115 & ~n43472 ;
  assign n43474 = n43473 ^ n43114 ;
  assign n43475 = n43474 ^ n43109 ;
  assign n43476 = ~n43111 & ~n43475 ;
  assign n43477 = n43476 ^ n43110 ;
  assign n43478 = n43477 ^ n43106 ;
  assign n43479 = ~n43107 & n43478 ;
  assign n43481 = n43480 ^ n43479 ;
  assign n43482 = n43103 & n43481 ;
  assign n43483 = n43482 ^ n43102 ;
  assign n43484 = n43483 ^ n43095 ;
  assign n43485 = ~n43099 & n43484 ;
  assign n43096 = n43095 ^ n43093 ;
  assign n43486 = n43485 ^ n43096 ;
  assign n43487 = n43094 & n43486 ;
  assign n43488 = n43487 ^ n43093 ;
  assign n43489 = n43488 ^ n43087 ;
  assign n43490 = ~n43089 & n43489 ;
  assign n43491 = n43490 ^ n43088 ;
  assign n43494 = n43493 ^ n43491 ;
  assign n43496 = n43495 ^ n43493 ;
  assign n43497 = ~n43494 & n43496 ;
  assign n43499 = n43498 ^ n43497 ;
  assign n43500 = ~n43084 & ~n43499 ;
  assign n43501 = n43500 ^ n43083 ;
  assign n43502 = n43501 ^ n43076 ;
  assign n43503 = ~n43077 & ~n43502 ;
  assign n43078 = n43076 ^ n43071 ;
  assign n43504 = n43503 ^ n43078 ;
  assign n43505 = n43072 & ~n43504 ;
  assign n43507 = n43506 ^ n43505 ;
  assign n43508 = n43067 & n43507 ;
  assign n43509 = n43508 ^ n43066 ;
  assign n43510 = n43509 ^ n43060 ;
  assign n43511 = n43062 & n43510 ;
  assign n43513 = n43512 ^ n43511 ;
  assign n43514 = n43057 & n43513 ;
  assign n43515 = n43514 ^ n43056 ;
  assign n43516 = n43515 ^ n43048 ;
  assign n43517 = ~n43052 & n43516 ;
  assign n43518 = n43517 ^ n43051 ;
  assign n43655 = n43654 ^ n43518 ;
  assign n43656 = ~n43522 & ~n43655 ;
  assign n43657 = n43656 ^ n43653 ;
  assign n43665 = n43398 ^ n43382 ;
  assign n43667 = n43665 ^ n43652 ;
  assign n43658 = n41871 ^ n41260 ;
  assign n43659 = n43658 ^ n43328 ;
  assign n43666 = n43665 ^ n43659 ;
  assign n43668 = n43667 ^ n43666 ;
  assign n43669 = ~n43657 & n43668 ;
  assign n43670 = n43669 ^ n43667 ;
  assign n43946 = n43401 ^ n43377 ;
  assign n43948 = n43946 ^ n43665 ;
  assign n43671 = n41857 ^ n41270 ;
  assign n43672 = n43671 ^ n42641 ;
  assign n43947 = n43946 ^ n43672 ;
  assign n43949 = n43948 ^ n43947 ;
  assign n43950 = n43670 & n43949 ;
  assign n43951 = n43950 ^ n43948 ;
  assign n43992 = n43404 ^ n43375 ;
  assign n43994 = n43992 ^ n43946 ;
  assign n43952 = n41847 ^ n41257 ;
  assign n43953 = n43952 ^ n42640 ;
  assign n43993 = n43992 ^ n43953 ;
  assign n43995 = n43994 ^ n43993 ;
  assign n43996 = n43951 & ~n43995 ;
  assign n43997 = n43996 ^ n43994 ;
  assign n44071 = n43407 ^ n43371 ;
  assign n44073 = n44071 ^ n43992 ;
  assign n43998 = n41845 ^ n41247 ;
  assign n43999 = n43998 ^ n42634 ;
  assign n44072 = n44071 ^ n43999 ;
  assign n44074 = n44073 ^ n44072 ;
  assign n44075 = n43997 & ~n44074 ;
  assign n44076 = n44075 ^ n44073 ;
  assign n44079 = n44078 ^ n44076 ;
  assign n44080 = n44079 ^ n40432 ;
  assign n43954 = n43953 ^ n43951 ;
  assign n43955 = n43954 ^ n40342 ;
  assign n43673 = n43672 ^ n43670 ;
  assign n43674 = n43673 ^ n40286 ;
  assign n43660 = n43659 ^ n43657 ;
  assign n43523 = n43522 ^ n43518 ;
  assign n43524 = n43523 ^ n40296 ;
  assign n43525 = n43515 ^ n43052 ;
  assign n43526 = n43525 ^ n41019 ;
  assign n43527 = n43513 ^ n43055 ;
  assign n43528 = n43527 ^ n41025 ;
  assign n43529 = n43509 ^ n43062 ;
  assign n43530 = n43529 ^ n41035 ;
  assign n43531 = n43507 ^ n43065 ;
  assign n43532 = n43531 ^ n41041 ;
  assign n43534 = n43501 ^ n43077 ;
  assign n43535 = n43534 ^ n40808 ;
  assign n43536 = n43499 ^ n43082 ;
  assign n43537 = n43536 ^ n40787 ;
  assign n43538 = n43496 ^ n43491 ;
  assign n43539 = n43538 ^ n40773 ;
  assign n43618 = n43488 ^ n43089 ;
  assign n43540 = n43486 ^ n43092 ;
  assign n43541 = n43540 ^ n40729 ;
  assign n43543 = n43481 ^ n43101 ;
  assign n43544 = n43543 ^ n40694 ;
  assign n43545 = n43477 ^ n43107 ;
  assign n43546 = n43545 ^ n40653 ;
  assign n43600 = n43474 ^ n43111 ;
  assign n43547 = n43471 ^ n43115 ;
  assign n43548 = n43547 ^ n40560 ;
  assign n43593 = n43592 ^ n43549 ;
  assign n43594 = n43592 ^ n40550 ;
  assign n43595 = n43593 & ~n43594 ;
  assign n43596 = n43595 ^ n40550 ;
  assign n43597 = n43596 ^ n43547 ;
  assign n43598 = ~n43548 & n43597 ;
  assign n43599 = n43598 ^ n40560 ;
  assign n43601 = n43600 ^ n43599 ;
  assign n43602 = n43600 ^ n40570 ;
  assign n43603 = ~n43601 & n43602 ;
  assign n43604 = n43603 ^ n40570 ;
  assign n43605 = n43604 ^ n43545 ;
  assign n43606 = n43546 & n43605 ;
  assign n43607 = n43606 ^ n40653 ;
  assign n43608 = n43607 ^ n43543 ;
  assign n43609 = ~n43544 & n43608 ;
  assign n43610 = n43609 ^ n40694 ;
  assign n43542 = n43483 ^ n43099 ;
  assign n43611 = n43610 ^ n43542 ;
  assign n43612 = n43610 ^ n40711 ;
  assign n43613 = ~n43611 & ~n43612 ;
  assign n43614 = n43613 ^ n40711 ;
  assign n43615 = n43614 ^ n43540 ;
  assign n43616 = n43541 & ~n43615 ;
  assign n43617 = n43616 ^ n40729 ;
  assign n43619 = n43618 ^ n43617 ;
  assign n43620 = n43618 ^ n40756 ;
  assign n43621 = n43619 & ~n43620 ;
  assign n43622 = n43621 ^ n40756 ;
  assign n43623 = n43622 ^ n43538 ;
  assign n43624 = ~n43539 & ~n43623 ;
  assign n43625 = n43624 ^ n40773 ;
  assign n43626 = n43625 ^ n43536 ;
  assign n43627 = n43537 & ~n43626 ;
  assign n43628 = n43627 ^ n40787 ;
  assign n43629 = n43628 ^ n43534 ;
  assign n43630 = ~n43535 & n43629 ;
  assign n43631 = n43630 ^ n40808 ;
  assign n43533 = n43504 ^ n43070 ;
  assign n43632 = n43631 ^ n43533 ;
  assign n43633 = n43531 ^ n40829 ;
  assign n43634 = n43633 ^ n43531 ;
  assign n43635 = n43634 ^ n43533 ;
  assign n43636 = n43632 & n43635 ;
  assign n43637 = n43636 ^ n43633 ;
  assign n43638 = ~n43532 & n43637 ;
  assign n43639 = n43638 ^ n41041 ;
  assign n43640 = n43639 ^ n43529 ;
  assign n43641 = ~n43530 & n43640 ;
  assign n43642 = n43641 ^ n41035 ;
  assign n43643 = n43642 ^ n43527 ;
  assign n43644 = n43528 & ~n43643 ;
  assign n43645 = n43644 ^ n41025 ;
  assign n43646 = n43645 ^ n43525 ;
  assign n43647 = ~n43526 & n43646 ;
  assign n43648 = n43647 ^ n41019 ;
  assign n43649 = n43648 ^ n43523 ;
  assign n43650 = n43524 & n43649 ;
  assign n43651 = n43650 ^ n40296 ;
  assign n43661 = n43660 ^ n43651 ;
  assign n43662 = n43660 ^ n40298 ;
  assign n43663 = ~n43661 & ~n43662 ;
  assign n43664 = n43663 ^ n40298 ;
  assign n43943 = n43673 ^ n43664 ;
  assign n43944 = n43674 & ~n43943 ;
  assign n43945 = n43944 ^ n40286 ;
  assign n44002 = n43954 ^ n43945 ;
  assign n44003 = ~n43955 & n44002 ;
  assign n44004 = n44003 ^ n40342 ;
  assign n44000 = n43999 ^ n43997 ;
  assign n44067 = n44004 ^ n44000 ;
  assign n44068 = n44004 ^ n40414 ;
  assign n44069 = n44067 & n44068 ;
  assign n44070 = n44069 ^ n40414 ;
  assign n44081 = n44080 ^ n44070 ;
  assign n43956 = n43955 ^ n43945 ;
  assign n43675 = n43674 ^ n43664 ;
  assign n43676 = n43662 ^ n43651 ;
  assign n43677 = n43625 ^ n43537 ;
  assign n43678 = n43620 ^ n43617 ;
  assign n43679 = n43614 ^ n43541 ;
  assign n43680 = n43542 ^ n40711 ;
  assign n43681 = n43680 ^ n43610 ;
  assign n43682 = n43604 ^ n43546 ;
  assign n43683 = n43602 ^ n43599 ;
  assign n43704 = ~n43701 & n43703 ;
  assign n43705 = n43596 ^ n43548 ;
  assign n43706 = n43704 & n43705 ;
  assign n43707 = ~n43683 & n43706 ;
  assign n43708 = ~n43682 & n43707 ;
  assign n43709 = n43607 ^ n43544 ;
  assign n43710 = n43708 & ~n43709 ;
  assign n43711 = n43681 & ~n43710 ;
  assign n43712 = n43679 & n43711 ;
  assign n43713 = n43678 & ~n43712 ;
  assign n43714 = n43622 ^ n43539 ;
  assign n43715 = ~n43713 & ~n43714 ;
  assign n43716 = n43677 & ~n43715 ;
  assign n43717 = n43628 ^ n43535 ;
  assign n43718 = n43716 & ~n43717 ;
  assign n43719 = n43533 ^ n40829 ;
  assign n43720 = n43719 ^ n43631 ;
  assign n43721 = n43718 & n43720 ;
  assign n43722 = n43637 ^ n41041 ;
  assign n43723 = ~n43721 & ~n43722 ;
  assign n43724 = n43639 ^ n43530 ;
  assign n43725 = n43723 & ~n43724 ;
  assign n43726 = n43642 ^ n43528 ;
  assign n43727 = ~n43725 & ~n43726 ;
  assign n43728 = n43645 ^ n43526 ;
  assign n43729 = n43727 & n43728 ;
  assign n43730 = n43648 ^ n43524 ;
  assign n43731 = ~n43729 & n43730 ;
  assign n43732 = ~n43676 & ~n43731 ;
  assign n43957 = n43675 & ~n43732 ;
  assign n43991 = n43956 & ~n43957 ;
  assign n44001 = n44000 ^ n40414 ;
  assign n44005 = n44004 ^ n44001 ;
  assign n44082 = n43991 & n44005 ;
  assign n44111 = n44081 & ~n44082 ;
  assign n44104 = n41604 ^ n33445 ;
  assign n44105 = n44104 ^ n2660 ;
  assign n44106 = n44105 ^ n3224 ;
  assign n44102 = n40509 ^ n40432 ;
  assign n44098 = n41893 ^ n41138 ;
  assign n44099 = n44098 ^ n42622 ;
  assign n44028 = n43409 ^ n43364 ;
  assign n44100 = n44099 ^ n44028 ;
  assign n44101 = n44100 ^ n44078 ;
  assign n44103 = n44102 ^ n44101 ;
  assign n44107 = n44106 ^ n44103 ;
  assign n44084 = n41608 ^ n33310 ;
  assign n44085 = n44084 ^ n38064 ;
  assign n44086 = n44085 ^ n2612 ;
  assign n44108 = n44107 ^ n44086 ;
  assign n44096 = n44079 ^ n44070 ;
  assign n44097 = n44080 & ~n44096 ;
  assign n44109 = n44108 ^ n44097 ;
  assign n44094 = n44078 ^ n44071 ;
  assign n44095 = ~n44076 & n44094 ;
  assign n44110 = n44109 ^ n44095 ;
  assign n44112 = n44111 ^ n44110 ;
  assign n44083 = n44082 ^ n44081 ;
  assign n44087 = n44086 ^ n44083 ;
  assign n44007 = n41614 ^ n2654 ;
  assign n44008 = n44007 ^ n38069 ;
  assign n44009 = n44008 ^ n31774 ;
  assign n44006 = n44005 ^ n43991 ;
  assign n44010 = n44009 ^ n44006 ;
  assign n44088 = n44083 ^ n44009 ;
  assign n44089 = n44088 ^ n44083 ;
  assign n43958 = n43957 ^ n43956 ;
  assign n43940 = n41618 ^ n33006 ;
  assign n43941 = n43940 ^ n38073 ;
  assign n43942 = n43941 ^ n31577 ;
  assign n43959 = n43958 ^ n43942 ;
  assign n43733 = n43732 ^ n43675 ;
  assign n2874 = n2873 ^ n2858 ;
  assign n2896 = n2895 ^ n2874 ;
  assign n2903 = n2902 ^ n2896 ;
  assign n43734 = n43733 ^ n2903 ;
  assign n43736 = n41625 ^ n32973 ;
  assign n43737 = n43736 ^ n38083 ;
  assign n43738 = n43737 ^ n2887 ;
  assign n43936 = n43738 ^ n43733 ;
  assign n43735 = n43731 ^ n43676 ;
  assign n43739 = n43738 ^ n43735 ;
  assign n43741 = n41630 ^ n1446 ;
  assign n43742 = n43741 ^ n38088 ;
  assign n43743 = n43742 ^ n31522 ;
  assign n43740 = n43730 ^ n43729 ;
  assign n43744 = n43743 ^ n43740 ;
  assign n43745 = n43728 ^ n43727 ;
  assign n1769 = n1747 ^ n1428 ;
  assign n1770 = n1769 ^ n1766 ;
  assign n1774 = n1773 ^ n1770 ;
  assign n43746 = n43745 ^ n1774 ;
  assign n1751 = n1732 ^ n1420 ;
  assign n1758 = n1757 ^ n1751 ;
  assign n1759 = n1758 ^ n1160 ;
  assign n43927 = n43745 ^ n1759 ;
  assign n43747 = n43726 ^ n43725 ;
  assign n43748 = n43747 ^ n1759 ;
  assign n43752 = n43724 ^ n43723 ;
  assign n43749 = n41640 ^ n1715 ;
  assign n43750 = n43749 ^ n1004 ;
  assign n43751 = n43750 ^ n1755 ;
  assign n43753 = n43752 ^ n43751 ;
  assign n43755 = n41645 ^ n1709 ;
  assign n43756 = n43755 ^ n38098 ;
  assign n43757 = n43756 ^ n996 ;
  assign n43921 = n43757 ^ n43752 ;
  assign n43754 = n43722 ^ n43721 ;
  assign n43758 = n43757 ^ n43754 ;
  assign n43759 = n43720 ^ n43718 ;
  assign n858 = n857 ^ n827 ;
  assign n886 = n885 ^ n858 ;
  assign n893 = n892 ^ n886 ;
  assign n43760 = n43759 ^ n893 ;
  assign n43764 = n43717 ^ n43716 ;
  assign n43761 = n41652 ^ n33051 ;
  assign n43762 = n43761 ^ n37767 ;
  assign n43763 = n43762 ^ n877 ;
  assign n43765 = n43764 ^ n43763 ;
  assign n43769 = n43715 ^ n43677 ;
  assign n43770 = n43769 ^ n43768 ;
  assign n43774 = n43714 ^ n43713 ;
  assign n43775 = n43774 ^ n43773 ;
  assign n43779 = n43712 ^ n43678 ;
  assign n43776 = n41667 ^ n1553 ;
  assign n43777 = n43776 ^ n37647 ;
  assign n43778 = n43777 ^ n31384 ;
  assign n43780 = n43779 ^ n43778 ;
  assign n43785 = n43711 ^ n43679 ;
  assign n43781 = n41674 ^ n33087 ;
  assign n43782 = n43781 ^ n37652 ;
  assign n43783 = n43782 ^ n31390 ;
  assign n43786 = n43785 ^ n43783 ;
  assign n43788 = n41679 ^ n33092 ;
  assign n43789 = n43788 ^ n37658 ;
  assign n43790 = n43789 ^ n2948 ;
  assign n43787 = n43710 ^ n43681 ;
  assign n43791 = n43790 ^ n43787 ;
  assign n43793 = n41684 ^ n33097 ;
  assign n43794 = n43793 ^ n37665 ;
  assign n43795 = n43794 ^ n31396 ;
  assign n43792 = n43709 ^ n43708 ;
  assign n43796 = n43795 ^ n43792 ;
  assign n43800 = n43707 ^ n43682 ;
  assign n43797 = n41689 ^ n33103 ;
  assign n43798 = n43797 ^ n37669 ;
  assign n43799 = n43798 ^ n31403 ;
  assign n43801 = n43800 ^ n43799 ;
  assign n43805 = n43706 ^ n43683 ;
  assign n43802 = n33107 ^ n2396 ;
  assign n43803 = n43802 ^ n37675 ;
  assign n43804 = n43803 ^ n31461 ;
  assign n43806 = n43805 ^ n43804 ;
  assign n43810 = n43705 ^ n43704 ;
  assign n43807 = n41695 ^ n33112 ;
  assign n43808 = n43807 ^ n2359 ;
  assign n43809 = n43808 ^ n31407 ;
  assign n43811 = n43810 ^ n43809 ;
  assign n43813 = n43812 ^ n2349 ;
  assign n43885 = ~n43813 & ~n43884 ;
  assign n43886 = n43885 ^ n43812 ;
  assign n43887 = n43886 ^ n43809 ;
  assign n43888 = n43811 & n43887 ;
  assign n43889 = n43888 ^ n43810 ;
  assign n43890 = n43889 ^ n43804 ;
  assign n43891 = ~n43806 & ~n43890 ;
  assign n43892 = n43891 ^ n43805 ;
  assign n43893 = n43892 ^ n43799 ;
  assign n43894 = ~n43801 & n43893 ;
  assign n43895 = n43894 ^ n43800 ;
  assign n43896 = n43895 ^ n43792 ;
  assign n43897 = ~n43796 & ~n43896 ;
  assign n43898 = n43897 ^ n43795 ;
  assign n43899 = n43898 ^ n43787 ;
  assign n43900 = n43791 & ~n43899 ;
  assign n43901 = n43900 ^ n43790 ;
  assign n43902 = n43901 ^ n43783 ;
  assign n43903 = ~n43786 & n43902 ;
  assign n43784 = n43783 ^ n43779 ;
  assign n43904 = n43903 ^ n43784 ;
  assign n43905 = ~n43780 & ~n43904 ;
  assign n43906 = n43905 ^ n43779 ;
  assign n43907 = n43906 ^ n43773 ;
  assign n43908 = ~n43775 & n43907 ;
  assign n43909 = n43908 ^ n43774 ;
  assign n43910 = n43909 ^ n43768 ;
  assign n43911 = ~n43770 & n43910 ;
  assign n43912 = n43911 ^ n43769 ;
  assign n43913 = n43912 ^ n43763 ;
  assign n43914 = ~n43765 & n43913 ;
  assign n43915 = n43914 ^ n43764 ;
  assign n43916 = n43915 ^ n893 ;
  assign n43917 = n43760 & n43916 ;
  assign n43918 = n43917 ^ n43759 ;
  assign n43919 = n43918 ^ n43757 ;
  assign n43920 = ~n43758 & n43919 ;
  assign n43922 = n43921 ^ n43920 ;
  assign n43923 = n43753 & n43922 ;
  assign n43924 = n43923 ^ n43752 ;
  assign n43925 = n43924 ^ n1759 ;
  assign n43926 = n43748 & n43925 ;
  assign n43928 = n43927 ^ n43926 ;
  assign n43929 = n43746 & ~n43928 ;
  assign n43930 = n43929 ^ n1774 ;
  assign n43931 = n43930 ^ n43740 ;
  assign n43932 = n43744 & ~n43931 ;
  assign n43933 = n43932 ^ n43743 ;
  assign n43934 = n43933 ^ n43738 ;
  assign n43935 = n43739 & n43934 ;
  assign n43937 = n43936 ^ n43935 ;
  assign n43938 = n43734 & n43937 ;
  assign n43939 = n43938 ^ n43733 ;
  assign n43988 = n43942 ^ n43939 ;
  assign n43989 = ~n43959 & ~n43988 ;
  assign n43990 = n43989 ^ n43958 ;
  assign n44090 = n44089 ^ n43990 ;
  assign n44091 = n44010 & ~n44090 ;
  assign n44092 = n44091 ^ n44088 ;
  assign n44093 = n44087 & ~n44092 ;
  assign n44113 = n44112 ^ n44093 ;
  assign n44065 = n42710 ^ n42060 ;
  assign n44066 = n44065 ^ n43118 ;
  assign n44114 = n44113 ^ n44066 ;
  assign n44117 = n44092 ^ n44086 ;
  assign n44124 = n44117 ^ n44113 ;
  assign n44115 = n42701 ^ n42166 ;
  assign n44116 = n44115 ^ n43120 ;
  assign n44118 = n44117 ^ n44116 ;
  assign n43965 = n42686 ^ n42016 ;
  assign n43966 = n43965 ^ n43132 ;
  assign n43961 = n43937 ^ n2903 ;
  assign n43962 = n42046 ^ n41931 ;
  assign n43963 = n43962 ^ n43136 ;
  assign n43964 = n43961 & n43963 ;
  assign n43967 = n43966 ^ n43964 ;
  assign n43960 = n43959 ^ n43939 ;
  assign n44013 = n43964 ^ n43960 ;
  assign n44014 = ~n43967 & ~n44013 ;
  assign n44011 = n44010 ^ n43990 ;
  assign n44012 = n44011 ^ n43964 ;
  assign n44015 = n44014 ^ n44012 ;
  assign n44016 = n42696 ^ n42178 ;
  assign n44017 = n44016 ^ n43126 ;
  assign n44119 = n44017 ^ n44011 ;
  assign n44120 = ~n44015 & n44119 ;
  assign n44121 = n44120 ^ n44011 ;
  assign n44122 = n44121 ^ n44117 ;
  assign n44123 = n44118 & ~n44122 ;
  assign n44125 = n44124 ^ n44123 ;
  assign n44126 = ~n44114 & n44125 ;
  assign n44127 = n44126 ^ n44113 ;
  assign n44128 = n44127 ^ n44062 ;
  assign n44129 = ~n44064 & n44128 ;
  assign n44130 = n44129 ^ n44063 ;
  assign n44058 = n43864 ^ n43846 ;
  assign n44059 = n44058 ^ n44056 ;
  assign n44060 = n44059 ^ n44058 ;
  assign n44131 = n44130 ^ n44060 ;
  assign n44132 = n44057 & ~n44131 ;
  assign n44133 = n44132 ^ n44059 ;
  assign n44134 = n43866 ^ n43845 ;
  assign n44138 = n44134 ^ n44058 ;
  assign n44135 = n42720 ^ n42138 ;
  assign n44136 = n44135 ^ n43106 ;
  assign n44137 = n44136 ^ n44134 ;
  assign n44139 = n44138 ^ n44137 ;
  assign n44140 = n44133 & ~n44139 ;
  assign n44141 = n44140 ^ n44138 ;
  assign n44144 = n43869 ^ n43840 ;
  assign n44146 = n44144 ^ n44134 ;
  assign n44142 = n42825 ^ n42203 ;
  assign n44143 = n44142 ^ n43102 ;
  assign n44145 = n44144 ^ n44143 ;
  assign n44147 = n44146 ^ n44145 ;
  assign n44148 = ~n44141 & ~n44147 ;
  assign n44149 = n44148 ^ n44146 ;
  assign n44154 = n44152 ^ n44144 ;
  assign n44150 = n42849 ^ n42132 ;
  assign n44151 = n44150 ^ n43095 ;
  assign n44153 = n44152 ^ n44151 ;
  assign n44155 = n44154 ^ n44153 ;
  assign n44156 = ~n44149 & ~n44155 ;
  assign n44157 = n44156 ^ n44154 ;
  assign n44158 = n42860 ^ n42038 ;
  assign n44159 = n44158 ^ n43093 ;
  assign n44160 = n44159 ^ n44152 ;
  assign n44161 = ~n44157 & n44160 ;
  assign n44163 = n44162 ^ n44161 ;
  assign n44164 = ~n44052 & n44163 ;
  assign n44165 = n44164 ^ n44051 ;
  assign n44166 = n44165 ^ n44046 ;
  assign n44167 = n44048 & ~n44166 ;
  assign n44168 = n44167 ^ n44047 ;
  assign n44169 = n44168 ^ n44042 ;
  assign n44170 = n44044 & ~n44169 ;
  assign n44171 = n44170 ^ n44043 ;
  assign n44038 = n43886 ^ n43811 ;
  assign n44039 = n44038 ^ n44034 ;
  assign n44040 = n44039 ^ n44038 ;
  assign n44172 = n44171 ^ n44040 ;
  assign n44173 = ~n44037 & ~n44172 ;
  assign n44174 = n44173 ^ n44039 ;
  assign n44175 = n43889 ^ n43806 ;
  assign n44179 = n44175 ^ n44038 ;
  assign n44176 = n43172 ^ n42102 ;
  assign n44177 = n44176 ^ n43071 ;
  assign n44178 = n44177 ^ n44175 ;
  assign n44180 = n44179 ^ n44178 ;
  assign n44181 = n44174 & n44180 ;
  assign n44182 = n44181 ^ n44179 ;
  assign n44261 = n43892 ^ n43801 ;
  assign n44263 = n44261 ^ n44175 ;
  assign n44183 = n43081 ^ n42092 ;
  assign n44184 = n44183 ^ n43066 ;
  assign n44262 = n44261 ^ n44184 ;
  assign n44264 = n44263 ^ n44262 ;
  assign n44265 = n44182 & n44264 ;
  assign n44266 = n44265 ^ n44263 ;
  assign n44269 = n44268 ^ n44266 ;
  assign n44270 = n44269 ^ n41033 ;
  assign n44185 = n44184 ^ n44182 ;
  assign n44186 = n44185 ^ n41040 ;
  assign n44187 = n44177 ^ n44174 ;
  assign n44188 = n44187 ^ n41047 ;
  assign n44189 = n44171 ^ n44037 ;
  assign n44190 = n44189 ^ n41057 ;
  assign n44191 = n44168 ^ n44044 ;
  assign n44192 = n44191 ^ n41063 ;
  assign n44244 = n44165 ^ n44048 ;
  assign n44193 = n44163 ^ n44051 ;
  assign n44194 = n44193 ^ n41075 ;
  assign n44196 = n44151 ^ n44149 ;
  assign n44197 = n44196 ^ n41078 ;
  assign n44199 = n44136 ^ n44133 ;
  assign n44200 = n44199 ^ n41090 ;
  assign n44201 = n44130 ^ n44057 ;
  assign n44202 = n44201 ^ n41096 ;
  assign n44203 = n44127 ^ n44064 ;
  assign n44204 = n44203 ^ n41106 ;
  assign n44213 = n44125 ^ n44066 ;
  assign n44018 = n44017 ^ n44015 ;
  assign n44019 = n44018 ^ n41007 ;
  assign n43969 = n43963 ^ n43961 ;
  assign n43970 = n41132 & n43969 ;
  assign n43971 = n43970 ^ n41125 ;
  assign n43968 = n43967 ^ n43960 ;
  assign n43985 = n43970 ^ n43968 ;
  assign n43986 = ~n43971 & ~n43985 ;
  assign n43987 = n43986 ^ n41125 ;
  assign n44205 = n44018 ^ n43987 ;
  assign n44206 = ~n44019 & n44205 ;
  assign n44207 = n44206 ^ n41007 ;
  assign n44208 = n44207 ^ n40450 ;
  assign n44209 = n44121 ^ n44118 ;
  assign n44210 = n44209 ^ n44207 ;
  assign n44211 = n44208 & ~n44210 ;
  assign n44212 = n44211 ^ n40450 ;
  assign n44214 = n44213 ^ n44212 ;
  assign n44215 = n44203 ^ n41112 ;
  assign n44216 = n44215 ^ n44203 ;
  assign n44217 = n44216 ^ n44212 ;
  assign n44218 = ~n44214 & ~n44217 ;
  assign n44219 = n44218 ^ n44215 ;
  assign n44220 = n44204 & n44219 ;
  assign n44221 = n44220 ^ n41106 ;
  assign n44222 = n44221 ^ n44201 ;
  assign n44223 = n44202 & n44222 ;
  assign n44224 = n44223 ^ n41096 ;
  assign n44225 = n44224 ^ n44199 ;
  assign n44226 = n44200 & ~n44225 ;
  assign n44227 = n44226 ^ n41090 ;
  assign n44198 = n44143 ^ n44141 ;
  assign n44228 = n44227 ^ n44198 ;
  assign n44229 = n44196 ^ n41088 ;
  assign n44230 = n44229 ^ n44196 ;
  assign n44231 = n44230 ^ n44198 ;
  assign n44232 = ~n44228 & ~n44231 ;
  assign n44233 = n44232 ^ n44229 ;
  assign n44234 = n44197 & ~n44233 ;
  assign n44235 = n44234 ^ n41078 ;
  assign n44195 = n44159 ^ n44157 ;
  assign n44236 = n44235 ^ n44195 ;
  assign n44237 = n44193 ^ n41324 ;
  assign n44238 = n44237 ^ n44193 ;
  assign n44239 = n44238 ^ n44195 ;
  assign n44240 = ~n44236 & ~n44239 ;
  assign n44241 = n44240 ^ n44237 ;
  assign n44242 = ~n44194 & n44241 ;
  assign n44243 = n44242 ^ n41075 ;
  assign n44245 = n44244 ^ n44243 ;
  assign n44246 = n44244 ^ n41069 ;
  assign n44247 = ~n44245 & ~n44246 ;
  assign n44248 = n44247 ^ n41069 ;
  assign n44249 = n44248 ^ n44191 ;
  assign n44250 = n44192 & n44249 ;
  assign n44251 = n44250 ^ n41063 ;
  assign n44252 = n44251 ^ n44189 ;
  assign n44253 = ~n44190 & n44252 ;
  assign n44254 = n44253 ^ n41057 ;
  assign n44255 = n44254 ^ n44187 ;
  assign n44256 = ~n44188 & n44255 ;
  assign n44257 = n44256 ^ n41047 ;
  assign n44258 = n44257 ^ n44185 ;
  assign n44259 = n44186 & n44258 ;
  assign n44260 = n44259 ^ n41040 ;
  assign n44271 = n44270 ^ n44260 ;
  assign n44272 = n44248 ^ n44192 ;
  assign n44273 = n44246 ^ n44243 ;
  assign n44274 = n44241 ^ n41075 ;
  assign n44275 = n44195 ^ n41324 ;
  assign n44276 = n44275 ^ n44235 ;
  assign n44277 = n44233 ^ n41078 ;
  assign n44278 = n44209 ^ n44208 ;
  assign n43972 = n43971 ^ n43968 ;
  assign n44020 = n44019 ^ n43987 ;
  assign n44279 = n43972 & ~n44020 ;
  assign n44280 = ~n44278 & ~n44279 ;
  assign n44281 = n44213 ^ n41112 ;
  assign n44282 = n44281 ^ n44212 ;
  assign n44283 = ~n44280 & ~n44282 ;
  assign n44284 = n44219 ^ n41106 ;
  assign n44285 = ~n44283 & n44284 ;
  assign n44286 = n44221 ^ n44202 ;
  assign n44287 = ~n44285 & n44286 ;
  assign n44288 = n44224 ^ n44200 ;
  assign n44289 = n44287 & ~n44288 ;
  assign n44290 = n44198 ^ n41088 ;
  assign n44291 = n44290 ^ n44227 ;
  assign n44292 = n44289 & n44291 ;
  assign n44293 = ~n44277 & ~n44292 ;
  assign n44294 = n44276 & n44293 ;
  assign n44295 = ~n44274 & n44294 ;
  assign n44296 = ~n44273 & n44295 ;
  assign n44297 = ~n44272 & n44296 ;
  assign n44298 = n44251 ^ n44190 ;
  assign n44299 = ~n44297 & n44298 ;
  assign n44300 = n44254 ^ n44188 ;
  assign n44301 = n44299 & n44300 ;
  assign n44302 = n44257 ^ n44186 ;
  assign n44303 = ~n44301 & n44302 ;
  assign n44304 = n44271 & ~n44303 ;
  assign n44314 = n43069 ^ n42235 ;
  assign n44315 = n44314 ^ n43056 ;
  assign n44308 = n43895 ^ n43796 ;
  assign n44310 = n44308 ^ n44261 ;
  assign n44309 = n44308 ^ n44268 ;
  assign n44311 = n44310 ^ n44309 ;
  assign n44312 = ~n44266 & ~n44311 ;
  assign n44313 = n44312 ^ n44310 ;
  assign n44316 = n44315 ^ n44313 ;
  assign n44317 = n44316 ^ n41027 ;
  assign n44305 = n44269 ^ n44260 ;
  assign n44306 = n44270 & n44305 ;
  assign n44307 = n44306 ^ n41033 ;
  assign n44318 = n44317 ^ n44307 ;
  assign n44451 = ~n44304 & n44318 ;
  assign n44462 = n44316 ^ n44307 ;
  assign n44463 = n44317 & n44462 ;
  assign n44464 = n44463 ^ n41027 ;
  assign n44458 = n43064 ^ n42083 ;
  assign n44459 = n44458 ^ n43048 ;
  assign n44452 = n43898 ^ n43791 ;
  assign n44454 = n44452 ^ n44308 ;
  assign n44453 = n44452 ^ n44315 ;
  assign n44455 = n44454 ^ n44453 ;
  assign n44456 = n44313 & ~n44455 ;
  assign n44457 = n44456 ^ n44454 ;
  assign n44460 = n44459 ^ n44457 ;
  assign n44461 = n44460 ^ n41023 ;
  assign n44465 = n44464 ^ n44461 ;
  assign n44629 = n44451 & n44465 ;
  assign n44512 = n43901 ^ n43786 ;
  assign n44566 = n44512 ^ n44452 ;
  assign n44565 = n44512 ^ n44459 ;
  assign n44567 = n44566 ^ n44565 ;
  assign n44568 = n44457 & ~n44567 ;
  assign n44569 = n44568 ^ n44566 ;
  assign n44562 = n43059 ^ n42067 ;
  assign n44563 = n44562 ^ n43521 ;
  assign n44596 = n44569 ^ n44563 ;
  assign n44598 = n44596 ^ n41016 ;
  assign n44592 = n44464 ^ n44460 ;
  assign n44593 = n44464 ^ n41023 ;
  assign n44594 = ~n44592 & ~n44593 ;
  assign n44595 = n44594 ^ n41023 ;
  assign n44628 = n44598 ^ n44595 ;
  assign n44675 = n44629 ^ n44628 ;
  assign n44676 = n44675 ^ n1658 ;
  assign n44466 = n44465 ^ n44451 ;
  assign n44467 = n44466 ^ n44450 ;
  assign n44319 = n44318 ^ n44304 ;
  assign n44031 = n42488 ^ n1611 ;
  assign n44032 = n44031 ^ n38571 ;
  assign n44033 = n44032 ^ n2987 ;
  assign n44320 = n44319 ^ n44033 ;
  assign n44324 = n44303 ^ n44271 ;
  assign n44321 = n42493 ^ n33880 ;
  assign n44322 = n44321 ^ n2975 ;
  assign n44323 = n44322 ^ n31991 ;
  assign n44325 = n44324 ^ n44323 ;
  assign n44329 = n44302 ^ n44301 ;
  assign n44441 = n44329 ^ n44324 ;
  assign n44330 = n44329 ^ n44328 ;
  assign n44332 = n42505 ^ n2957 ;
  assign n44333 = n44332 ^ n38583 ;
  assign n44334 = n44333 ^ n31998 ;
  assign n44438 = n44334 ^ n44329 ;
  assign n44331 = n44300 ^ n44299 ;
  assign n44335 = n44334 ^ n44331 ;
  assign n44339 = n44298 ^ n44297 ;
  assign n44336 = n42511 ^ n33917 ;
  assign n44337 = n44336 ^ n38589 ;
  assign n44338 = n44337 ^ n32003 ;
  assign n44340 = n44339 ^ n44338 ;
  assign n44344 = n44296 ^ n44272 ;
  assign n44341 = n42515 ^ n33922 ;
  assign n44342 = n44341 ^ n38593 ;
  assign n44343 = n44342 ^ n32008 ;
  assign n44345 = n44344 ^ n44343 ;
  assign n44349 = n44295 ^ n44273 ;
  assign n44346 = n42520 ^ n33926 ;
  assign n44347 = n44346 ^ n38599 ;
  assign n44348 = n44347 ^ n32014 ;
  assign n44350 = n44349 ^ n44348 ;
  assign n44354 = n44294 ^ n44274 ;
  assign n44351 = n42526 ^ n33931 ;
  assign n44352 = n44351 ^ n38604 ;
  assign n44353 = n44352 ^ n32019 ;
  assign n44355 = n44354 ^ n44353 ;
  assign n44357 = n42530 ^ n2429 ;
  assign n44358 = n44357 ^ n38608 ;
  assign n44359 = n44358 ^ n32024 ;
  assign n44356 = n44293 ^ n44276 ;
  assign n44360 = n44359 ^ n44356 ;
  assign n44366 = n44292 ^ n44277 ;
  assign n44420 = n44366 ^ n44356 ;
  assign n44362 = n38620 ^ n33941 ;
  assign n44363 = n44362 ^ n41953 ;
  assign n44364 = n44363 ^ n32033 ;
  assign n44361 = n44291 ^ n44289 ;
  assign n44365 = n44364 ^ n44361 ;
  assign n44404 = n44288 ^ n44287 ;
  assign n44372 = n44286 ^ n44285 ;
  assign n44369 = n41962 ^ n33951 ;
  assign n44370 = n44369 ^ n2015 ;
  assign n44371 = n44370 ^ n32040 ;
  assign n44373 = n44372 ^ n44371 ;
  assign n44377 = n44284 ^ n44283 ;
  assign n44374 = n41967 ^ n33955 ;
  assign n44375 = n44374 ^ n38632 ;
  assign n44376 = n44375 ^ n2007 ;
  assign n44378 = n44377 ^ n44376 ;
  assign n44383 = n44282 ^ n44280 ;
  assign n44379 = n41991 ^ n1928 ;
  assign n44380 = n44379 ^ n38636 ;
  assign n44381 = n44380 ^ n32048 ;
  assign n44384 = n44383 ^ n44381 ;
  assign n44388 = n44279 ^ n44278 ;
  assign n44385 = n41972 ^ n33281 ;
  assign n44386 = n44385 ^ n3053 ;
  assign n44387 = n44386 ^ n32052 ;
  assign n44389 = n44388 ^ n44387 ;
  assign n44021 = n44020 ^ n43972 ;
  assign n43982 = n41976 ^ n3242 ;
  assign n43983 = n43982 ^ n38644 ;
  assign n43984 = n43983 ^ n3045 ;
  assign n44022 = n44021 ^ n43984 ;
  assign n2757 = n2756 ^ n2732 ;
  assign n2776 = n2775 ^ n2757 ;
  assign n2783 = n2782 ^ n2776 ;
  assign n43973 = n43972 ^ n2783 ;
  assign n43974 = n42610 ^ n3227 ;
  assign n43975 = n43974 ^ n38993 ;
  assign n43976 = n43975 ^ n2774 ;
  assign n43977 = n43969 ^ n41132 ;
  assign n43978 = n43976 & n43977 ;
  assign n43979 = n43978 ^ n2783 ;
  assign n43980 = n43973 & ~n43979 ;
  assign n43981 = n43980 ^ n43972 ;
  assign n44390 = n43984 ^ n43981 ;
  assign n44391 = n44022 & n44390 ;
  assign n44392 = n44391 ^ n43984 ;
  assign n44393 = n44392 ^ n44387 ;
  assign n44394 = n44389 & ~n44393 ;
  assign n44395 = n44394 ^ n44388 ;
  assign n44396 = n44395 ^ n44381 ;
  assign n44397 = ~n44384 & n44396 ;
  assign n44382 = n44381 ^ n44377 ;
  assign n44398 = n44397 ^ n44382 ;
  assign n44399 = ~n44378 & ~n44398 ;
  assign n44400 = n44399 ^ n44377 ;
  assign n44401 = n44400 ^ n44371 ;
  assign n44402 = n44373 & n44401 ;
  assign n44403 = n44402 ^ n44372 ;
  assign n44405 = n44404 ^ n44403 ;
  assign n44406 = n41957 ^ n33946 ;
  assign n44407 = n44406 ^ n38624 ;
  assign n44408 = n44407 ^ n2096 ;
  assign n44409 = n44408 ^ n44403 ;
  assign n44410 = ~n44405 & n44409 ;
  assign n44411 = n44410 ^ n44408 ;
  assign n44367 = n44366 ^ n44364 ;
  assign n44368 = n44367 ^ n44366 ;
  assign n44412 = n44411 ^ n44368 ;
  assign n44413 = ~n44365 & n44412 ;
  assign n44414 = n44413 ^ n44367 ;
  assign n44415 = n42028 ^ n2414 ;
  assign n44416 = n44415 ^ n38614 ;
  assign n44417 = n44416 ^ n32029 ;
  assign n44418 = n44417 ^ n44366 ;
  assign n44419 = n44414 & n44418 ;
  assign n44421 = n44420 ^ n44419 ;
  assign n44422 = n44360 & ~n44421 ;
  assign n44423 = n44422 ^ n44359 ;
  assign n44424 = n44423 ^ n44353 ;
  assign n44425 = ~n44355 & ~n44424 ;
  assign n44426 = n44425 ^ n44354 ;
  assign n44427 = n44426 ^ n44348 ;
  assign n44428 = ~n44350 & n44427 ;
  assign n44429 = n44428 ^ n44349 ;
  assign n44430 = n44429 ^ n44343 ;
  assign n44431 = ~n44345 & n44430 ;
  assign n44432 = n44431 ^ n44344 ;
  assign n44433 = n44432 ^ n44338 ;
  assign n44434 = n44340 & n44433 ;
  assign n44435 = n44434 ^ n44339 ;
  assign n44436 = n44435 ^ n44334 ;
  assign n44437 = ~n44335 & n44436 ;
  assign n44439 = n44438 ^ n44437 ;
  assign n44440 = ~n44330 & ~n44439 ;
  assign n44442 = n44441 ^ n44440 ;
  assign n44443 = n44325 & ~n44442 ;
  assign n44444 = n44443 ^ n44324 ;
  assign n44445 = n44444 ^ n44033 ;
  assign n44446 = ~n44320 & ~n44445 ;
  assign n44447 = n44446 ^ n44319 ;
  assign n44677 = n44450 ^ n44447 ;
  assign n44678 = n44467 & n44677 ;
  assign n44679 = n44678 ^ n44466 ;
  assign n44680 = n44679 ^ n1658 ;
  assign n44681 = n44676 & ~n44680 ;
  assign n44682 = n44681 ^ n44675 ;
  assign n44630 = n44628 & n44629 ;
  assign n44564 = n44563 ^ n44512 ;
  assign n44570 = n44564 & ~n44569 ;
  assign n44571 = n44570 ^ n44512 ;
  assign n44560 = n43054 ^ n42251 ;
  assign n44561 = n44560 ^ n43652 ;
  assign n44572 = n44571 ^ n44561 ;
  assign n44506 = n43904 ^ n43778 ;
  assign n44591 = n44572 ^ n44506 ;
  assign n44626 = n44591 ^ n41374 ;
  assign n44597 = n44596 ^ n44595 ;
  assign n44599 = ~n44597 & n44598 ;
  assign n44600 = n44599 ^ n41016 ;
  assign n44627 = n44626 ^ n44600 ;
  assign n44673 = n44630 ^ n44627 ;
  assign n44670 = n42476 ^ n964 ;
  assign n44671 = n44670 ^ n38559 ;
  assign n44672 = n44671 ^ n1116 ;
  assign n44674 = n44673 ^ n44672 ;
  assign n45277 = n44682 ^ n44674 ;
  assign n44481 = n43918 ^ n43758 ;
  assign n46527 = n45277 ^ n44481 ;
  assign n45109 = n42890 ^ n34522 ;
  assign n45110 = n45109 ^ n39224 ;
  assign n45111 = n45110 ^ n762 ;
  assign n44497 = n43521 ^ n43069 ;
  assign n44496 = n43909 ^ n43770 ;
  assign n44498 = n44497 ^ n44496 ;
  assign n44495 = n44429 ^ n44345 ;
  assign n44499 = n44498 ^ n44495 ;
  assign n44503 = n43074 ^ n43048 ;
  assign n44502 = n43906 ^ n43775 ;
  assign n44504 = n44503 ^ n44502 ;
  assign n44500 = n44426 ^ n44350 ;
  assign n44505 = n44504 ^ n44500 ;
  assign n44509 = n44423 ^ n44355 ;
  assign n44507 = n44506 ^ n43081 ;
  assign n44508 = n44507 ^ n43056 ;
  assign n44510 = n44509 ^ n44508 ;
  assign n44513 = n43172 ^ n43061 ;
  assign n44514 = n44513 ^ n44512 ;
  assign n44511 = n44421 ^ n44359 ;
  assign n44515 = n44514 ^ n44511 ;
  assign n44518 = n44417 ^ n44414 ;
  assign n44875 = n44518 ^ n44511 ;
  assign n44516 = n43086 ^ n43066 ;
  assign n44517 = n44516 ^ n44452 ;
  assign n44519 = n44518 ^ n44517 ;
  assign n44521 = n43091 ^ n43071 ;
  assign n44522 = n44521 ^ n44308 ;
  assign n44520 = n44411 ^ n44365 ;
  assign n44523 = n44522 ^ n44520 ;
  assign n44525 = n43076 ^ n43036 ;
  assign n44526 = n44525 ^ n44261 ;
  assign n44524 = n44408 ^ n44405 ;
  assign n44527 = n44526 ^ n44524 ;
  assign n44529 = n43083 ^ n42873 ;
  assign n44530 = n44529 ^ n44175 ;
  assign n44528 = n44400 ^ n44373 ;
  assign n44531 = n44530 ^ n44528 ;
  assign n44534 = n44398 ^ n44376 ;
  assign n44863 = n44534 ^ n44528 ;
  assign n44532 = n43495 ^ n42860 ;
  assign n44533 = n44532 ^ n44038 ;
  assign n44535 = n44534 ^ n44533 ;
  assign n44537 = n43088 ^ n42849 ;
  assign n44538 = n44537 ^ n44034 ;
  assign n44536 = n44395 ^ n44384 ;
  assign n44539 = n44538 ^ n44536 ;
  assign n44542 = n44392 ^ n44389 ;
  assign n44857 = n44542 ^ n44536 ;
  assign n44540 = n43093 ^ n42825 ;
  assign n44541 = n44540 ^ n44043 ;
  assign n44543 = n44542 ^ n44541 ;
  assign n44544 = n43095 ^ n42720 ;
  assign n44545 = n44544 ^ n44047 ;
  assign n44023 = n44022 ^ n43981 ;
  assign n44546 = n44545 ^ n44023 ;
  assign n44549 = n43978 ^ n43973 ;
  assign n44851 = n44549 ^ n44023 ;
  assign n44547 = n43102 ^ n42029 ;
  assign n44548 = n44547 ^ n44049 ;
  assign n44550 = n44549 ^ n44548 ;
  assign n44553 = n43977 ^ n43976 ;
  assign n44551 = n43106 ^ n42036 ;
  assign n44552 = n44551 ^ n44152 ;
  assign n44554 = n44553 ^ n44552 ;
  assign n44471 = n43924 ^ n43748 ;
  assign n44027 = n43928 ^ n1774 ;
  assign n44763 = n44471 ^ n44027 ;
  assign n44475 = n43922 ^ n43751 ;
  assign n44740 = n44475 ^ n44471 ;
  assign n44707 = n44481 ^ n44475 ;
  assign n44485 = n43915 ^ n43760 ;
  assign n44649 = n44485 ^ n44481 ;
  assign n44490 = n43912 ^ n43765 ;
  assign n44621 = n44490 ^ n44485 ;
  assign n44586 = n44496 ^ n44490 ;
  assign n44580 = n44502 ^ n44496 ;
  assign n44573 = n44571 ^ n44506 ;
  assign n44574 = ~n44572 & n44573 ;
  assign n44559 = n44506 ^ n44502 ;
  assign n44575 = n44574 ^ n44559 ;
  assign n44576 = n43050 ^ n42356 ;
  assign n44577 = n44576 ^ n43665 ;
  assign n44578 = n44577 ^ n44502 ;
  assign n44579 = ~n44575 & ~n44578 ;
  assign n44581 = n44580 ^ n44579 ;
  assign n44582 = n43146 ^ n42375 ;
  assign n44583 = n44582 ^ n43946 ;
  assign n44584 = n44583 ^ n44496 ;
  assign n44585 = n44581 & ~n44584 ;
  assign n44587 = n44586 ^ n44585 ;
  assign n44557 = n43328 ^ n42604 ;
  assign n44558 = n44557 ^ n43992 ;
  assign n44619 = n44558 ^ n44490 ;
  assign n44620 = n44587 & ~n44619 ;
  assign n44622 = n44621 ^ n44620 ;
  assign n44617 = n42641 ^ n41860 ;
  assign n44618 = n44617 ^ n44071 ;
  assign n44647 = n44618 ^ n44485 ;
  assign n44648 = ~n44622 & ~n44647 ;
  assign n44650 = n44649 ^ n44648 ;
  assign n44645 = n42640 ^ n41871 ;
  assign n44646 = n44645 ^ n44028 ;
  assign n44705 = n44646 ^ n44481 ;
  assign n44706 = n44650 & n44705 ;
  assign n44708 = n44707 ^ n44706 ;
  assign n44703 = n42634 ^ n41857 ;
  assign n44704 = n44703 ^ n43438 ;
  assign n44738 = n44704 ^ n44475 ;
  assign n44739 = ~n44708 & ~n44738 ;
  assign n44741 = n44740 ^ n44739 ;
  assign n44736 = n42632 ^ n41847 ;
  assign n44737 = n44736 ^ n43446 ;
  assign n44761 = n44737 ^ n44471 ;
  assign n44762 = n44741 & ~n44761 ;
  assign n44764 = n44763 ^ n44762 ;
  assign n44759 = n42622 ^ n41845 ;
  assign n44760 = n44759 ^ n43436 ;
  assign n44765 = n44764 ^ n44760 ;
  assign n44766 = n44765 ^ n41247 ;
  assign n44790 = n42665 ^ n40999 ;
  assign n44791 = n44790 ^ n43430 ;
  assign n44784 = n43930 ^ n43744 ;
  assign n44785 = n44784 ^ n44027 ;
  assign n44786 = n44785 ^ n44760 ;
  assign n44787 = n44786 ^ n44784 ;
  assign n44788 = n44764 & n44787 ;
  assign n44789 = n44788 ^ n44785 ;
  assign n44792 = n44791 ^ n44789 ;
  assign n44793 = n44792 ^ n41247 ;
  assign n44742 = n44741 ^ n44737 ;
  assign n44743 = n44742 ^ n41257 ;
  assign n44709 = n44708 ^ n44704 ;
  assign n44710 = n44709 ^ n41270 ;
  assign n44623 = n44622 ^ n44618 ;
  assign n44624 = n44623 ^ n40989 ;
  assign n44589 = n44577 ^ n44575 ;
  assign n44590 = n44589 ^ n41379 ;
  assign n44601 = n44600 ^ n44591 ;
  assign n44602 = n44600 ^ n41374 ;
  assign n44603 = n44601 & n44602 ;
  assign n44604 = n44603 ^ n41374 ;
  assign n44605 = n44604 ^ n44589 ;
  assign n44606 = n44590 & ~n44605 ;
  assign n44607 = n44606 ^ n41379 ;
  assign n44608 = n44607 ^ n41588 ;
  assign n44609 = n44583 ^ n44581 ;
  assign n44610 = n44609 ^ n44607 ;
  assign n44611 = ~n44608 & n44610 ;
  assign n44612 = n44611 ^ n41588 ;
  assign n44588 = n44587 ^ n44558 ;
  assign n44613 = n44612 ^ n44588 ;
  assign n44614 = n44612 ^ n41832 ;
  assign n44615 = ~n44613 & n44614 ;
  assign n44616 = n44615 ^ n41832 ;
  assign n44653 = n44623 ^ n44616 ;
  assign n44654 = ~n44624 & ~n44653 ;
  assign n44655 = n44654 ^ n40989 ;
  assign n44651 = n44650 ^ n44646 ;
  assign n44699 = n44655 ^ n44651 ;
  assign n44700 = n44655 ^ n41260 ;
  assign n44701 = n44699 & n44700 ;
  assign n44702 = n44701 ^ n41260 ;
  assign n44733 = n44709 ^ n44702 ;
  assign n44734 = ~n44710 & ~n44733 ;
  assign n44735 = n44734 ^ n41270 ;
  assign n44756 = n44742 ^ n44735 ;
  assign n44757 = ~n44743 & ~n44756 ;
  assign n44758 = n44757 ^ n41257 ;
  assign n44794 = n44793 ^ n44758 ;
  assign n44795 = n44794 ^ n44792 ;
  assign n44796 = n44766 & n44795 ;
  assign n44797 = n44796 ^ n44793 ;
  assign n44767 = n44766 ^ n44758 ;
  assign n44652 = n44651 ^ n41260 ;
  assign n44656 = n44655 ^ n44652 ;
  assign n44625 = n44624 ^ n44616 ;
  assign n44631 = n44627 & ~n44630 ;
  assign n44632 = n44604 ^ n41379 ;
  assign n44633 = n44632 ^ n44589 ;
  assign n44634 = n44631 & ~n44633 ;
  assign n44635 = n44609 ^ n44608 ;
  assign n44636 = ~n44634 & n44635 ;
  assign n44637 = n44588 ^ n41832 ;
  assign n44638 = n44637 ^ n44612 ;
  assign n44639 = n44636 & ~n44638 ;
  assign n44657 = ~n44625 & ~n44639 ;
  assign n44698 = ~n44656 & ~n44657 ;
  assign n44711 = n44710 ^ n44702 ;
  assign n44732 = ~n44698 & n44711 ;
  assign n44744 = n44743 ^ n44735 ;
  assign n44768 = ~n44732 & n44744 ;
  assign n44799 = n44767 & n44768 ;
  assign n44830 = n44799 ^ n44792 ;
  assign n44831 = ~n44797 & ~n44830 ;
  assign n44824 = n41145 ^ n41138 ;
  assign n44820 = n42059 ^ n41893 ;
  assign n44821 = n44820 ^ n44791 ;
  assign n44822 = n44821 ^ n43428 ;
  assign n44819 = n43933 ^ n43739 ;
  assign n44823 = n44822 ^ n44819 ;
  assign n44825 = n44824 ^ n44823 ;
  assign n44816 = n42433 ^ n2676 ;
  assign n44817 = n44816 ^ n38949 ;
  assign n44818 = n44817 ^ n32501 ;
  assign n44826 = n44825 ^ n44818 ;
  assign n44781 = n42437 ^ n34215 ;
  assign n44782 = n44781 ^ n38812 ;
  assign n44783 = n44782 ^ n3143 ;
  assign n44827 = n44826 ^ n44783 ;
  assign n44814 = n44791 ^ n44784 ;
  assign n44815 = ~n44789 & n44814 ;
  assign n44828 = n44827 ^ n44815 ;
  assign n44812 = n44799 ^ n44797 ;
  assign n44813 = ~n41145 & n44812 ;
  assign n44829 = n44828 ^ n44813 ;
  assign n44832 = n44831 ^ n44829 ;
  assign n44798 = n44797 ^ n41145 ;
  assign n44800 = n44799 ^ n44798 ;
  assign n44801 = n44800 ^ n44783 ;
  assign n44769 = n44768 ^ n44767 ;
  assign n44753 = n42442 ^ n34204 ;
  assign n44754 = n44753 ^ n38763 ;
  assign n44755 = n44754 ^ n32512 ;
  assign n44770 = n44769 ^ n44755 ;
  assign n44745 = n44744 ^ n44732 ;
  assign n44729 = n42447 ^ n34021 ;
  assign n44730 = n44729 ^ n38746 ;
  assign n44731 = n44730 ^ n32518 ;
  assign n44746 = n44745 ^ n44731 ;
  assign n44641 = n42463 ^ n33838 ;
  assign n44642 = n44641 ^ n38548 ;
  assign n44643 = n44642 ^ n32533 ;
  assign n44640 = n44639 ^ n44625 ;
  assign n44644 = n44643 ^ n44640 ;
  assign n44661 = n44638 ^ n44636 ;
  assign n1263 = n1262 ^ n1184 ;
  assign n1279 = n1278 ^ n1263 ;
  assign n1286 = n1285 ^ n1279 ;
  assign n44662 = n44661 ^ n1286 ;
  assign n44666 = n44635 ^ n44634 ;
  assign n44663 = n42469 ^ n33845 ;
  assign n44664 = n44663 ^ n1135 ;
  assign n44665 = n44664 ^ n1270 ;
  assign n44667 = n44666 ^ n44665 ;
  assign n44668 = n44633 ^ n44631 ;
  assign n1093 = n1083 ^ n1038 ;
  assign n1118 = n1117 ^ n1093 ;
  assign n1125 = n1124 ^ n1118 ;
  assign n44669 = n44668 ^ n1125 ;
  assign n44685 = n44672 ^ n44668 ;
  assign n44683 = n44682 ^ n44672 ;
  assign n44684 = n44674 & n44683 ;
  assign n44686 = n44685 ^ n44684 ;
  assign n44687 = n44669 & n44686 ;
  assign n44688 = n44687 ^ n44668 ;
  assign n44689 = n44688 ^ n44665 ;
  assign n44690 = ~n44667 & ~n44689 ;
  assign n44691 = n44690 ^ n44666 ;
  assign n44692 = n44691 ^ n1286 ;
  assign n44693 = ~n44662 & n44692 ;
  assign n44694 = n44693 ^ n44661 ;
  assign n44658 = n44657 ^ n44656 ;
  assign n44659 = n44658 ^ n44643 ;
  assign n44660 = n44659 ^ n44658 ;
  assign n44695 = n44694 ^ n44660 ;
  assign n44696 = ~n44644 & ~n44695 ;
  assign n44697 = n44696 ^ n44659 ;
  assign n44712 = n44711 ^ n44698 ;
  assign n44717 = n44712 ^ n44658 ;
  assign n44713 = n42458 ^ n33833 ;
  assign n44714 = n44713 ^ n38544 ;
  assign n44715 = n44714 ^ n32527 ;
  assign n44716 = n44715 ^ n44712 ;
  assign n44718 = n44717 ^ n44716 ;
  assign n44719 = n44697 & n44718 ;
  assign n44720 = n44719 ^ n44717 ;
  assign n44721 = n42453 ^ n33828 ;
  assign n44722 = n44721 ^ n38539 ;
  assign n44723 = n44722 ^ n32523 ;
  assign n44747 = n44723 ^ n44712 ;
  assign n44748 = n44720 & n44747 ;
  assign n44749 = n44748 ^ n44712 ;
  assign n44750 = n44749 ^ n44731 ;
  assign n44751 = ~n44746 & ~n44750 ;
  assign n44752 = n44751 ^ n44745 ;
  assign n44778 = n44755 ^ n44752 ;
  assign n44779 = n44770 & n44778 ;
  assign n44780 = n44779 ^ n44769 ;
  assign n44810 = n44783 ^ n44780 ;
  assign n44811 = n44801 & n44810 ;
  assign n44833 = n44832 ^ n44811 ;
  assign n44845 = n44833 ^ n44552 ;
  assign n44724 = n44723 ^ n44720 ;
  assign n44725 = n43126 ^ n42046 ;
  assign n44726 = n44725 ^ n44063 ;
  assign n44727 = n44724 & n44726 ;
  assign n44555 = n43120 ^ n42686 ;
  assign n44556 = n44555 ^ n44056 ;
  assign n44728 = n44727 ^ n44556 ;
  assign n44774 = n44749 ^ n44746 ;
  assign n44771 = n44770 ^ n44752 ;
  assign n44772 = n44771 ^ n44556 ;
  assign n44773 = n44772 ^ n44771 ;
  assign n44775 = n44774 ^ n44773 ;
  assign n44776 = n44728 & ~n44775 ;
  assign n44777 = n44776 ^ n44772 ;
  assign n44802 = n44801 ^ n44780 ;
  assign n44806 = n44802 ^ n44771 ;
  assign n44803 = n43118 ^ n42696 ;
  assign n44804 = n44803 ^ n44058 ;
  assign n44805 = n44804 ^ n44802 ;
  assign n44807 = n44806 ^ n44805 ;
  assign n44808 = ~n44777 & ~n44807 ;
  assign n44809 = n44808 ^ n44806 ;
  assign n44835 = n43114 ^ n42701 ;
  assign n44836 = n44835 ^ n44134 ;
  assign n44837 = n44836 ^ n44833 ;
  assign n44834 = n44833 ^ n44802 ;
  assign n44838 = n44837 ^ n44834 ;
  assign n44839 = ~n44809 & n44838 ;
  assign n44840 = n44839 ^ n44834 ;
  assign n44841 = n43110 ^ n42710 ;
  assign n44842 = n44841 ^ n44144 ;
  assign n44843 = n44842 ^ n44833 ;
  assign n44844 = n44840 & n44843 ;
  assign n44846 = n44845 ^ n44844 ;
  assign n44847 = ~n44554 & n44846 ;
  assign n44848 = n44847 ^ n44553 ;
  assign n44849 = n44848 ^ n44548 ;
  assign n44850 = ~n44550 & n44849 ;
  assign n44852 = n44851 ^ n44850 ;
  assign n44853 = ~n44546 & n44852 ;
  assign n44854 = n44853 ^ n44023 ;
  assign n44855 = n44854 ^ n44542 ;
  assign n44856 = ~n44543 & n44855 ;
  assign n44858 = n44857 ^ n44856 ;
  assign n44859 = ~n44539 & n44858 ;
  assign n44860 = n44859 ^ n44538 ;
  assign n44861 = n44860 ^ n44533 ;
  assign n44862 = ~n44535 & ~n44861 ;
  assign n44864 = n44863 ^ n44862 ;
  assign n44865 = ~n44531 & ~n44864 ;
  assign n44866 = n44865 ^ n44530 ;
  assign n44867 = n44866 ^ n44524 ;
  assign n44868 = ~n44527 & ~n44867 ;
  assign n44869 = n44868 ^ n44526 ;
  assign n44870 = n44869 ^ n44520 ;
  assign n44871 = ~n44523 & ~n44870 ;
  assign n44872 = n44871 ^ n44522 ;
  assign n44873 = n44872 ^ n44517 ;
  assign n44874 = ~n44519 & n44873 ;
  assign n44876 = n44875 ^ n44874 ;
  assign n44877 = n44515 & ~n44876 ;
  assign n44878 = n44877 ^ n44514 ;
  assign n44879 = n44878 ^ n44508 ;
  assign n44880 = n44510 & n44879 ;
  assign n44881 = n44880 ^ n44509 ;
  assign n44882 = n44881 ^ n44500 ;
  assign n44883 = ~n44505 & ~n44882 ;
  assign n44501 = n44500 ^ n44495 ;
  assign n44884 = n44883 ^ n44501 ;
  assign n44885 = ~n44499 & ~n44884 ;
  assign n44886 = n44885 ^ n44498 ;
  assign n44493 = n44432 ^ n44340 ;
  assign n44491 = n43652 ^ n43064 ;
  assign n44492 = n44491 ^ n44490 ;
  assign n44494 = n44493 ^ n44492 ;
  assign n45010 = n44886 ^ n44494 ;
  assign n45012 = n45010 ^ n42083 ;
  assign n44917 = n44884 ^ n44498 ;
  assign n44918 = n44917 ^ n42235 ;
  assign n44919 = n44881 ^ n44505 ;
  assign n44920 = n44919 ^ n42089 ;
  assign n44921 = n44878 ^ n44510 ;
  assign n44922 = n44921 ^ n42092 ;
  assign n44996 = n44876 ^ n44514 ;
  assign n44923 = n44872 ^ n44519 ;
  assign n44924 = n44923 ^ n42108 ;
  assign n44925 = n44869 ^ n44523 ;
  assign n44926 = n44925 ^ n42114 ;
  assign n44927 = n44866 ^ n44527 ;
  assign n44928 = n44927 ^ n42120 ;
  assign n44929 = n44864 ^ n44530 ;
  assign n44930 = n44929 ^ n42031 ;
  assign n44931 = n44860 ^ n44535 ;
  assign n44932 = n44931 ^ n42038 ;
  assign n44933 = n44858 ^ n44538 ;
  assign n44934 = n44933 ^ n42132 ;
  assign n44935 = n44854 ^ n44543 ;
  assign n44936 = n44935 ^ n42203 ;
  assign n44937 = n44852 ^ n44545 ;
  assign n44938 = n44937 ^ n42138 ;
  assign n44962 = n44846 ^ n44553 ;
  assign n44940 = n44842 ^ n44840 ;
  assign n44941 = n44940 ^ n42060 ;
  assign n44942 = n44836 ^ n44809 ;
  assign n44943 = n44942 ^ n42166 ;
  assign n44944 = n44804 ^ n44777 ;
  assign n44945 = n44944 ^ n42178 ;
  assign n44946 = n44726 ^ n44724 ;
  assign n44947 = n41931 & n44946 ;
  assign n44948 = n44947 ^ n42016 ;
  assign n44949 = n44774 ^ n44728 ;
  assign n44950 = n44949 ^ n44947 ;
  assign n44951 = n44948 & n44950 ;
  assign n44952 = n44951 ^ n42016 ;
  assign n44953 = n44952 ^ n44944 ;
  assign n44954 = ~n44945 & n44953 ;
  assign n44955 = n44954 ^ n42178 ;
  assign n44956 = n44955 ^ n44942 ;
  assign n44957 = ~n44943 & n44956 ;
  assign n44958 = n44957 ^ n42166 ;
  assign n44959 = n44958 ^ n44940 ;
  assign n44960 = n44941 & ~n44959 ;
  assign n44961 = n44960 ^ n42060 ;
  assign n44963 = n44962 ^ n44961 ;
  assign n44964 = n44962 ^ n42044 ;
  assign n44965 = n44963 & n44964 ;
  assign n44966 = n44965 ^ n42044 ;
  assign n44939 = n44848 ^ n44550 ;
  assign n44967 = n44966 ^ n44939 ;
  assign n44968 = n44937 ^ n42053 ;
  assign n44969 = n44968 ^ n44937 ;
  assign n44970 = n44969 ^ n44939 ;
  assign n44971 = ~n44967 & n44970 ;
  assign n44972 = n44971 ^ n44968 ;
  assign n44973 = n44938 & ~n44972 ;
  assign n44974 = n44973 ^ n42138 ;
  assign n44975 = n44974 ^ n44935 ;
  assign n44976 = ~n44936 & ~n44975 ;
  assign n44977 = n44976 ^ n42203 ;
  assign n44978 = n44977 ^ n44933 ;
  assign n44979 = n44934 & n44978 ;
  assign n44980 = n44979 ^ n42132 ;
  assign n44981 = n44980 ^ n44931 ;
  assign n44982 = n44932 & ~n44981 ;
  assign n44983 = n44982 ^ n42038 ;
  assign n44984 = n44983 ^ n44929 ;
  assign n44985 = n44930 & n44984 ;
  assign n44986 = n44985 ^ n42031 ;
  assign n44987 = n44986 ^ n44927 ;
  assign n44988 = n44928 & n44987 ;
  assign n44989 = n44988 ^ n42120 ;
  assign n44990 = n44989 ^ n44925 ;
  assign n44991 = n44926 & n44990 ;
  assign n44992 = n44991 ^ n42114 ;
  assign n44993 = n44992 ^ n44923 ;
  assign n44994 = ~n44924 & n44993 ;
  assign n44995 = n44994 ^ n42108 ;
  assign n44997 = n44996 ^ n44995 ;
  assign n44998 = n44996 ^ n42102 ;
  assign n44999 = ~n44997 & ~n44998 ;
  assign n45000 = n44999 ^ n42102 ;
  assign n45001 = n45000 ^ n44921 ;
  assign n45002 = n44922 & n45001 ;
  assign n45003 = n45002 ^ n42092 ;
  assign n45004 = n45003 ^ n44919 ;
  assign n45005 = ~n44920 & ~n45004 ;
  assign n45006 = n45005 ^ n42089 ;
  assign n45007 = n45006 ^ n44917 ;
  assign n45008 = n44918 & ~n45007 ;
  assign n45009 = n45008 ^ n42235 ;
  assign n45071 = n45012 ^ n45009 ;
  assign n45035 = n45006 ^ n44918 ;
  assign n45036 = n45000 ^ n44922 ;
  assign n45037 = n44998 ^ n44995 ;
  assign n45038 = n44939 ^ n42053 ;
  assign n45039 = n45038 ^ n44966 ;
  assign n45040 = n44964 ^ n44961 ;
  assign n45041 = n44958 ^ n44941 ;
  assign n45042 = n44949 ^ n44948 ;
  assign n45043 = n44952 ^ n44945 ;
  assign n45044 = n45042 & n45043 ;
  assign n45045 = n44955 ^ n44943 ;
  assign n45046 = ~n45044 & ~n45045 ;
  assign n45047 = ~n45041 & ~n45046 ;
  assign n45048 = n45040 & ~n45047 ;
  assign n45049 = n45039 & ~n45048 ;
  assign n45050 = n44972 ^ n42138 ;
  assign n45051 = n45049 & n45050 ;
  assign n45052 = n44974 ^ n44936 ;
  assign n45053 = n45051 & ~n45052 ;
  assign n45054 = n44977 ^ n44934 ;
  assign n45055 = ~n45053 & n45054 ;
  assign n45056 = n44980 ^ n44932 ;
  assign n45057 = n45055 & ~n45056 ;
  assign n45058 = n44983 ^ n44930 ;
  assign n45059 = n45057 & ~n45058 ;
  assign n45060 = n44986 ^ n44928 ;
  assign n45061 = n45059 & n45060 ;
  assign n45062 = n44989 ^ n44926 ;
  assign n45063 = n45061 & ~n45062 ;
  assign n45064 = n44992 ^ n44924 ;
  assign n45065 = ~n45063 & n45064 ;
  assign n45066 = n45037 & n45065 ;
  assign n45067 = ~n45036 & ~n45066 ;
  assign n45068 = n45003 ^ n44920 ;
  assign n45069 = ~n45067 & n45068 ;
  assign n45070 = ~n45035 & ~n45069 ;
  assign n45107 = n45071 ^ n45070 ;
  assign n45254 = n45111 ^ n45107 ;
  assign n45112 = n45069 ^ n45035 ;
  assign n45113 = n45112 ^ n45111 ;
  assign n45117 = n45068 ^ n45067 ;
  assign n45114 = n42894 ^ n680 ;
  assign n45115 = n45114 ^ n39229 ;
  assign n45116 = n45115 ^ n33055 ;
  assign n45118 = n45117 ^ n45116 ;
  assign n45122 = n45066 ^ n45036 ;
  assign n45119 = n42899 ^ n34553 ;
  assign n45120 = n45119 ^ n39234 ;
  assign n45121 = n45120 ^ n1553 ;
  assign n45123 = n45122 ^ n45121 ;
  assign n45127 = n45065 ^ n45037 ;
  assign n45124 = n42904 ^ n34558 ;
  assign n45125 = n45124 ^ n39241 ;
  assign n45126 = n45125 ^ n33087 ;
  assign n45128 = n45127 ^ n45126 ;
  assign n45132 = n45064 ^ n45063 ;
  assign n45129 = n42910 ^ n34563 ;
  assign n45130 = n45129 ^ n39246 ;
  assign n45131 = n45130 ^ n33092 ;
  assign n45133 = n45132 ^ n45131 ;
  assign n45135 = n42917 ^ n34569 ;
  assign n45136 = n45135 ^ n39251 ;
  assign n45137 = n45136 ^ n33097 ;
  assign n45134 = n45062 ^ n45061 ;
  assign n45138 = n45137 ^ n45134 ;
  assign n45140 = n42921 ^ n34574 ;
  assign n45141 = n45140 ^ n39255 ;
  assign n45142 = n45141 ^ n33103 ;
  assign n45139 = n45060 ^ n45059 ;
  assign n45143 = n45142 ^ n45139 ;
  assign n45147 = n45058 ^ n45057 ;
  assign n45144 = n42926 ^ n34580 ;
  assign n45145 = n45144 ^ n39261 ;
  assign n45146 = n45145 ^ n33107 ;
  assign n45148 = n45147 ^ n45146 ;
  assign n45152 = n45056 ^ n45055 ;
  assign n45149 = n42931 ^ n34591 ;
  assign n45150 = n45149 ^ n2315 ;
  assign n45151 = n45150 ^ n33112 ;
  assign n45153 = n45152 ^ n45151 ;
  assign n45157 = n45054 ^ n45053 ;
  assign n45154 = n42936 ^ n34586 ;
  assign n45155 = n45154 ^ n39268 ;
  assign n45156 = n45155 ^ n2310 ;
  assign n45158 = n45157 ^ n45156 ;
  assign n45159 = n45052 ^ n45051 ;
  assign n45224 = n45159 ^ n45157 ;
  assign n2166 = n2165 ^ n2132 ;
  assign n2194 = n2193 ^ n2166 ;
  assign n2201 = n2200 ^ n2194 ;
  assign n45160 = n45159 ^ n2201 ;
  assign n45163 = n42943 ^ n34613 ;
  assign n45164 = n45163 ^ n39274 ;
  assign n45165 = n45164 ^ n2185 ;
  assign n45161 = n45050 ^ n45049 ;
  assign n45166 = n45165 ^ n45161 ;
  assign n45170 = n45048 ^ n45039 ;
  assign n45167 = n42947 ^ n2064 ;
  assign n45168 = n45167 ^ n39279 ;
  assign n45169 = n45168 ^ n33124 ;
  assign n45171 = n45170 ^ n45169 ;
  assign n45175 = n42952 ^ n34621 ;
  assign n45176 = n45175 ^ n39296 ;
  assign n45177 = n45176 ^ n33128 ;
  assign n45174 = n45047 ^ n45040 ;
  assign n45178 = n45177 ^ n45174 ;
  assign n45179 = n42957 ^ n34625 ;
  assign n45180 = n45179 ^ n39284 ;
  assign n45181 = n45180 ^ n33134 ;
  assign n45214 = n45181 ^ n45174 ;
  assign n45182 = n45046 ^ n45041 ;
  assign n45183 = n45182 ^ n45181 ;
  assign n45187 = n45045 ^ n45044 ;
  assign n45184 = n42962 ^ n3081 ;
  assign n45185 = n45184 ^ n38797 ;
  assign n45186 = n45185 ^ n33138 ;
  assign n45188 = n45187 ^ n45186 ;
  assign n45190 = n42971 ^ n34632 ;
  assign n45191 = n45190 ^ n38754 ;
  assign n45192 = n45191 ^ n33147 ;
  assign n45189 = n45043 ^ n45042 ;
  assign n45193 = n45192 ^ n45189 ;
  assign n45194 = n42967 ^ n34054 ;
  assign n45195 = n45194 ^ n3194 ;
  assign n45196 = n45195 ^ n33142 ;
  assign n45197 = n45196 ^ n45042 ;
  assign n45198 = n43335 ^ n35198 ;
  assign n45199 = n45198 ^ n39714 ;
  assign n45200 = n45199 ^ n3193 ;
  assign n45201 = n44946 ^ n41931 ;
  assign n45202 = n45200 & n45201 ;
  assign n45203 = n45202 ^ n45196 ;
  assign n45204 = n45197 & ~n45203 ;
  assign n45205 = n45204 ^ n45042 ;
  assign n45206 = n45205 ^ n45192 ;
  assign n45207 = ~n45193 & n45206 ;
  assign n45208 = n45207 ^ n45192 ;
  assign n45209 = n45208 ^ n45186 ;
  assign n45210 = n45188 & ~n45209 ;
  assign n45211 = n45210 ^ n45187 ;
  assign n45212 = n45211 ^ n45181 ;
  assign n45213 = ~n45183 & n45212 ;
  assign n45215 = n45214 ^ n45213 ;
  assign n45216 = ~n45178 & n45215 ;
  assign n45217 = n45216 ^ n45177 ;
  assign n45172 = n45169 ^ n45161 ;
  assign n45173 = n45172 ^ n45161 ;
  assign n45218 = n45217 ^ n45173 ;
  assign n45219 = n45171 & n45218 ;
  assign n45220 = n45219 ^ n45172 ;
  assign n45221 = ~n45166 & ~n45220 ;
  assign n45162 = n45161 ^ n45159 ;
  assign n45222 = n45221 ^ n45162 ;
  assign n45223 = n45160 & ~n45222 ;
  assign n45225 = n45224 ^ n45223 ;
  assign n45226 = ~n45158 & ~n45225 ;
  assign n45227 = n45226 ^ n45157 ;
  assign n45228 = n45227 ^ n45151 ;
  assign n45229 = ~n45153 & n45228 ;
  assign n45230 = n45229 ^ n45152 ;
  assign n45231 = n45230 ^ n45146 ;
  assign n45232 = ~n45148 & n45231 ;
  assign n45233 = n45232 ^ n45147 ;
  assign n45234 = n45233 ^ n45139 ;
  assign n45235 = n45143 & n45234 ;
  assign n45236 = n45235 ^ n45142 ;
  assign n45237 = n45236 ^ n45134 ;
  assign n45238 = ~n45138 & n45237 ;
  assign n45239 = n45238 ^ n45137 ;
  assign n45240 = n45239 ^ n45131 ;
  assign n45241 = n45133 & ~n45240 ;
  assign n45242 = n45241 ^ n45132 ;
  assign n45243 = n45242 ^ n45126 ;
  assign n45244 = ~n45128 & ~n45243 ;
  assign n45245 = n45244 ^ n45127 ;
  assign n45246 = n45245 ^ n45121 ;
  assign n45247 = n45123 & n45246 ;
  assign n45248 = n45247 ^ n45122 ;
  assign n45249 = n45248 ^ n45116 ;
  assign n45250 = n45118 & ~n45249 ;
  assign n45251 = n45250 ^ n45117 ;
  assign n45252 = n45251 ^ n45111 ;
  assign n45253 = n45113 & n45252 ;
  assign n45255 = n45254 ^ n45253 ;
  assign n45104 = n34517 ^ n2993 ;
  assign n45105 = n45104 ^ n770 ;
  assign n45106 = n45105 ^ n33051 ;
  assign n45930 = n45255 ^ n45106 ;
  assign n46528 = n46527 ^ n45930 ;
  assign n45514 = n44452 ^ n43076 ;
  assign n45515 = n45514 ^ n44500 ;
  assign n45503 = n45217 ^ n45171 ;
  assign n45319 = n45215 ^ n45177 ;
  assign n45504 = n45503 ^ n45319 ;
  assign n45317 = n44261 ^ n43495 ;
  assign n45318 = n45317 ^ n44511 ;
  assign n45320 = n45319 ^ n45318 ;
  assign n45322 = n44175 ^ n43088 ;
  assign n45323 = n45322 ^ n44518 ;
  assign n45321 = n45211 ^ n45183 ;
  assign n45324 = n45323 ^ n45321 ;
  assign n45327 = n45208 ^ n45188 ;
  assign n45497 = n45327 ^ n45321 ;
  assign n45325 = n44038 ^ n43093 ;
  assign n45326 = n45325 ^ n44520 ;
  assign n45328 = n45327 ^ n45326 ;
  assign n45331 = n45205 ^ n45193 ;
  assign n45329 = n44034 ^ n43095 ;
  assign n45330 = n45329 ^ n44524 ;
  assign n45332 = n45331 ^ n45330 ;
  assign n45333 = n45202 ^ n45197 ;
  assign n45491 = n45333 ^ n45331 ;
  assign n45334 = n44043 ^ n43102 ;
  assign n45335 = n45334 ^ n44528 ;
  assign n45336 = n45335 ^ n45333 ;
  assign n45339 = n45201 ^ n45200 ;
  assign n45337 = n44047 ^ n43106 ;
  assign n45338 = n45337 ^ n44534 ;
  assign n45340 = n45339 ^ n45338 ;
  assign n45371 = n44694 ^ n44644 ;
  assign n45369 = n43136 ^ n42665 ;
  assign n45370 = n45369 ^ n44117 ;
  assign n45372 = n45371 ^ n45370 ;
  assign n45345 = n44691 ^ n44662 ;
  assign n45343 = n43428 ^ n42622 ;
  assign n45344 = n45343 ^ n44011 ;
  assign n45346 = n45345 ^ n45344 ;
  assign n45349 = n44688 ^ n44667 ;
  assign n45347 = n43430 ^ n42632 ;
  assign n45348 = n45347 ^ n43960 ;
  assign n45350 = n45349 ^ n45348 ;
  assign n45354 = n44686 ^ n1125 ;
  assign n45352 = n43961 ^ n43436 ;
  assign n45353 = n45352 ^ n42634 ;
  assign n45355 = n45354 ^ n45353 ;
  assign n44907 = n44679 ^ n44676 ;
  assign n44905 = n43438 ^ n42641 ;
  assign n44906 = n44905 ^ n44784 ;
  assign n44908 = n44907 ^ n44906 ;
  assign n45278 = n45277 ^ n44907 ;
  assign n45279 = n45278 ^ n45277 ;
  assign n44468 = n44467 ^ n44447 ;
  assign n44029 = n44028 ^ n43328 ;
  assign n44030 = n44029 ^ n44027 ;
  assign n44469 = n44468 ^ n44030 ;
  assign n44472 = n44071 ^ n43146 ;
  assign n44473 = n44472 ^ n44471 ;
  assign n44470 = n44444 ^ n44320 ;
  assign n44474 = n44473 ^ n44470 ;
  assign n44478 = n44442 ^ n44323 ;
  assign n44898 = n44478 ^ n44470 ;
  assign n44476 = n43992 ^ n43050 ;
  assign n44477 = n44476 ^ n44475 ;
  assign n44479 = n44478 ^ n44477 ;
  assign n44482 = n43946 ^ n43054 ;
  assign n44483 = n44482 ^ n44481 ;
  assign n44480 = n44439 ^ n44328 ;
  assign n44484 = n44483 ^ n44480 ;
  assign n44488 = n44435 ^ n44335 ;
  assign n44892 = n44488 ^ n44480 ;
  assign n44486 = n44485 ^ n43059 ;
  assign n44487 = n44486 ^ n43665 ;
  assign n44489 = n44488 ^ n44487 ;
  assign n44889 = n44493 ^ n44488 ;
  assign n44887 = n44886 ^ n44493 ;
  assign n44888 = n44494 & n44887 ;
  assign n44890 = n44889 ^ n44888 ;
  assign n44891 = ~n44489 & n44890 ;
  assign n44893 = n44892 ^ n44891 ;
  assign n44894 = ~n44484 & ~n44893 ;
  assign n44895 = n44894 ^ n44483 ;
  assign n44896 = n44895 ^ n44478 ;
  assign n44897 = ~n44479 & ~n44896 ;
  assign n44899 = n44898 ^ n44897 ;
  assign n44900 = n44474 & ~n44899 ;
  assign n44901 = n44900 ^ n44473 ;
  assign n44902 = n44901 ^ n44030 ;
  assign n44903 = ~n44469 & n44902 ;
  assign n44904 = n44903 ^ n44468 ;
  assign n45280 = n45279 ^ n44904 ;
  assign n45281 = n44908 & ~n45280 ;
  assign n45282 = n45281 ^ n45278 ;
  assign n45357 = n45354 ^ n45277 ;
  assign n45283 = n44819 ^ n42640 ;
  assign n45284 = n45283 ^ n43446 ;
  assign n45356 = n45354 ^ n45284 ;
  assign n45358 = n45357 ^ n45356 ;
  assign n45359 = n45282 & n45358 ;
  assign n45360 = n45359 ^ n45357 ;
  assign n45361 = n45355 & n45360 ;
  assign n45362 = n45361 ^ n45354 ;
  assign n45351 = n45349 ^ n45345 ;
  assign n45363 = n45362 ^ n45351 ;
  assign n45364 = n45363 ^ n45345 ;
  assign n45365 = n45350 & ~n45364 ;
  assign n45366 = n45365 ^ n45351 ;
  assign n45367 = n45346 & ~n45366 ;
  assign n45368 = n45367 ^ n45345 ;
  assign n45373 = n45372 ^ n45368 ;
  assign n45403 = n45373 ^ n40999 ;
  assign n45374 = n45366 ^ n45344 ;
  assign n45375 = n45374 ^ n41845 ;
  assign n45376 = n45362 ^ n45350 ;
  assign n45377 = n45376 ^ n41847 ;
  assign n45378 = n45360 ^ n45353 ;
  assign n45379 = n45378 ^ n41857 ;
  assign n44909 = n44908 ^ n44904 ;
  assign n44910 = n44909 ^ n41860 ;
  assign n44911 = n44901 ^ n44469 ;
  assign n44912 = n44911 ^ n42604 ;
  assign n45026 = n44899 ^ n44473 ;
  assign n44913 = n44895 ^ n44479 ;
  assign n44914 = n44913 ^ n42356 ;
  assign n45018 = n44893 ^ n44483 ;
  assign n44915 = n44890 ^ n44487 ;
  assign n44916 = n44915 ^ n42067 ;
  assign n45011 = n45010 ^ n45009 ;
  assign n45013 = ~n45011 & n45012 ;
  assign n45014 = n45013 ^ n42083 ;
  assign n45015 = n45014 ^ n44915 ;
  assign n45016 = ~n44916 & n45015 ;
  assign n45017 = n45016 ^ n42067 ;
  assign n45019 = n45018 ^ n45017 ;
  assign n45020 = n45018 ^ n42251 ;
  assign n45021 = n45019 & n45020 ;
  assign n45022 = n45021 ^ n42251 ;
  assign n45023 = n45022 ^ n44913 ;
  assign n45024 = n44914 & n45023 ;
  assign n45025 = n45024 ^ n42356 ;
  assign n45027 = n45026 ^ n45025 ;
  assign n45028 = n45026 ^ n42375 ;
  assign n45029 = ~n45027 & ~n45028 ;
  assign n45030 = n45029 ^ n42375 ;
  assign n45031 = n45030 ^ n44911 ;
  assign n45032 = ~n44912 & ~n45031 ;
  assign n45033 = n45032 ^ n42604 ;
  assign n45287 = n45033 ^ n44909 ;
  assign n45288 = n44910 & ~n45287 ;
  assign n45289 = n45288 ^ n41860 ;
  assign n45285 = n45284 ^ n45282 ;
  assign n45380 = n45289 ^ n45285 ;
  assign n45381 = n45289 ^ n41871 ;
  assign n45382 = n45380 & ~n45381 ;
  assign n45383 = n45382 ^ n41871 ;
  assign n45384 = n45383 ^ n45378 ;
  assign n45385 = n45379 & ~n45384 ;
  assign n45386 = n45385 ^ n41857 ;
  assign n45387 = n45386 ^ n45376 ;
  assign n45388 = n45377 & ~n45387 ;
  assign n45389 = n45388 ^ n41847 ;
  assign n45390 = n45389 ^ n41845 ;
  assign n45391 = n45375 & ~n45390 ;
  assign n45392 = n45391 ^ n41845 ;
  assign n45404 = n45403 ^ n45392 ;
  assign n45396 = n45383 ^ n45379 ;
  assign n45034 = n45033 ^ n44910 ;
  assign n45072 = n45070 & ~n45071 ;
  assign n45073 = n45014 ^ n44916 ;
  assign n45074 = n45072 & n45073 ;
  assign n45075 = n45020 ^ n45017 ;
  assign n45076 = ~n45074 & n45075 ;
  assign n45077 = n45022 ^ n44914 ;
  assign n45078 = n45076 & ~n45077 ;
  assign n45079 = n45028 ^ n45025 ;
  assign n45080 = ~n45078 & n45079 ;
  assign n45081 = n45030 ^ n44912 ;
  assign n45082 = n45080 & ~n45081 ;
  assign n45276 = n45034 & ~n45082 ;
  assign n45286 = n45285 ^ n41871 ;
  assign n45290 = n45289 ^ n45286 ;
  assign n45397 = ~n45276 & ~n45290 ;
  assign n45398 = ~n45396 & ~n45397 ;
  assign n45399 = n45386 ^ n45377 ;
  assign n45400 = ~n45398 & n45399 ;
  assign n45401 = n45389 ^ n45375 ;
  assign n45402 = n45400 & n45401 ;
  assign n45424 = n45404 ^ n45402 ;
  assign n45406 = n43353 ^ n35042 ;
  assign n45407 = n45406 ^ n39593 ;
  assign n45408 = n45407 ^ n33310 ;
  assign n45425 = n45424 ^ n45408 ;
  assign n45427 = n43357 ^ n35115 ;
  assign n45428 = n45427 ^ n39597 ;
  assign n45429 = n45428 ^ n2654 ;
  assign n45453 = n45429 ^ n45424 ;
  assign n45426 = n45401 ^ n45400 ;
  assign n45430 = n45429 ^ n45426 ;
  assign n45432 = n43415 ^ n35047 ;
  assign n45433 = n45432 ^ n39603 ;
  assign n45434 = n45433 ^ n33006 ;
  assign n45431 = n45399 ^ n45398 ;
  assign n45435 = n45434 ^ n45431 ;
  assign n45441 = n45397 ^ n45396 ;
  assign n45438 = n43362 ^ n35051 ;
  assign n45439 = n45438 ^ n39609 ;
  assign n45440 = n45439 ^ n2873 ;
  assign n45442 = n45441 ^ n45440 ;
  assign n45291 = n45290 ^ n45276 ;
  assign n45295 = n45294 ^ n45291 ;
  assign n45083 = n45082 ^ n45034 ;
  assign n1439 = n1399 ^ n1333 ;
  assign n1440 = n1439 ^ n1436 ;
  assign n1447 = n1446 ^ n1440 ;
  assign n45084 = n45083 ^ n1447 ;
  assign n1403 = n1362 ^ n1315 ;
  assign n1422 = n1421 ^ n1403 ;
  assign n1429 = n1428 ^ n1422 ;
  assign n45272 = n45083 ^ n1429 ;
  assign n45085 = n45081 ^ n45080 ;
  assign n45086 = n45085 ^ n1429 ;
  assign n45088 = n1720 ^ n1220 ;
  assign n45089 = n45088 ^ n43381 ;
  assign n45090 = n45089 ^ n1420 ;
  assign n45087 = n45079 ^ n45078 ;
  assign n45091 = n45090 ^ n45087 ;
  assign n45092 = n45077 ^ n45076 ;
  assign n1702 = n1695 ^ n1205 ;
  assign n1712 = n1711 ^ n1702 ;
  assign n1716 = n1715 ^ n1712 ;
  assign n45093 = n45092 ^ n1716 ;
  assign n45097 = n45075 ^ n45074 ;
  assign n45094 = n43387 ^ n1678 ;
  assign n45095 = n45094 ^ n39212 ;
  assign n45096 = n45095 ^ n1709 ;
  assign n45098 = n45097 ^ n45096 ;
  assign n45102 = n45073 ^ n45072 ;
  assign n45099 = n43029 ^ n1669 ;
  assign n45100 = n45099 ^ n39217 ;
  assign n45101 = n45100 ^ n857 ;
  assign n45103 = n45102 ^ n45101 ;
  assign n45108 = n45107 ^ n45106 ;
  assign n45256 = ~n45108 & ~n45255 ;
  assign n45257 = n45256 ^ n45107 ;
  assign n45258 = n45257 ^ n45101 ;
  assign n45259 = n45103 & n45258 ;
  assign n45260 = n45259 ^ n45102 ;
  assign n45261 = n45260 ^ n45096 ;
  assign n45262 = n45098 & ~n45261 ;
  assign n45263 = n45262 ^ n45097 ;
  assign n45264 = n45263 ^ n1716 ;
  assign n45265 = n45093 & ~n45264 ;
  assign n45266 = n45265 ^ n45092 ;
  assign n45267 = n45266 ^ n45087 ;
  assign n45268 = ~n45091 & n45267 ;
  assign n45269 = n45268 ^ n45090 ;
  assign n45270 = n45269 ^ n1429 ;
  assign n45271 = ~n45086 & n45270 ;
  assign n45273 = n45272 ^ n45271 ;
  assign n45274 = n45084 & n45273 ;
  assign n45275 = n45274 ^ n45083 ;
  assign n45443 = n45291 ^ n45275 ;
  assign n45444 = n45295 & ~n45443 ;
  assign n45445 = n45444 ^ n45294 ;
  assign n45446 = n45445 ^ n45440 ;
  assign n45447 = ~n45442 & ~n45446 ;
  assign n45448 = n45447 ^ n45441 ;
  assign n45449 = n45448 ^ n45434 ;
  assign n45450 = ~n45435 & ~n45449 ;
  assign n45436 = n45434 ^ n45429 ;
  assign n45451 = n45450 ^ n45436 ;
  assign n45452 = n45430 & n45451 ;
  assign n45454 = n45453 ^ n45452 ;
  assign n45455 = n45425 & ~n45454 ;
  assign n45420 = n45370 ^ n45368 ;
  assign n45421 = ~n45372 & ~n45420 ;
  assign n45410 = n43338 ^ n3158 ;
  assign n45411 = n45410 ^ n39660 ;
  assign n45412 = n45411 ^ n33445 ;
  assign n45413 = n45412 ^ n44820 ;
  assign n45297 = n44715 ^ n44697 ;
  assign n45414 = n45413 ^ n45297 ;
  assign n45415 = n45414 ^ n43132 ;
  assign n45416 = n45415 ^ n45370 ;
  assign n45409 = n44113 ^ n40999 ;
  assign n45417 = n45416 ^ n45409 ;
  assign n45418 = n45417 ^ n45408 ;
  assign n45405 = ~n45402 & n45404 ;
  assign n45419 = n45418 ^ n45405 ;
  assign n45422 = n45421 ^ n45419 ;
  assign n45393 = n45392 ^ n45373 ;
  assign n45394 = n45392 ^ n40999 ;
  assign n45395 = ~n45393 & n45394 ;
  assign n45423 = n45422 ^ n45395 ;
  assign n45456 = n45455 ^ n45423 ;
  assign n45341 = n44049 ^ n43110 ;
  assign n45342 = n45341 ^ n44536 ;
  assign n45457 = n45456 ^ n45342 ;
  assign n45460 = n45454 ^ n45408 ;
  assign n45482 = n45460 ^ n45456 ;
  assign n45458 = n44152 ^ n43114 ;
  assign n45459 = n45458 ^ n44542 ;
  assign n45461 = n45460 ^ n45459 ;
  assign n45464 = n45451 ^ n45426 ;
  assign n45462 = n44144 ^ n44023 ;
  assign n45463 = n45462 ^ n43118 ;
  assign n45465 = n45464 ^ n45463 ;
  assign n45468 = n44058 ^ n43126 ;
  assign n45469 = n45468 ^ n44553 ;
  assign n45470 = n45445 ^ n45442 ;
  assign n45471 = n45469 & ~n45470 ;
  assign n45466 = n44134 ^ n43120 ;
  assign n45467 = n45466 ^ n44549 ;
  assign n45472 = n45471 ^ n45467 ;
  assign n45473 = n45448 ^ n45435 ;
  assign n45474 = n45473 ^ n45467 ;
  assign n45475 = ~n45472 & n45474 ;
  assign n45476 = n45475 ^ n45473 ;
  assign n45477 = n45476 ^ n45463 ;
  assign n45478 = n45465 & ~n45477 ;
  assign n45479 = n45478 ^ n45464 ;
  assign n45480 = n45479 ^ n45459 ;
  assign n45481 = n45461 & ~n45480 ;
  assign n45483 = n45482 ^ n45481 ;
  assign n45484 = n45457 & ~n45483 ;
  assign n45485 = n45484 ^ n45456 ;
  assign n45486 = n45485 ^ n45338 ;
  assign n45487 = n45340 & n45486 ;
  assign n45488 = n45487 ^ n45339 ;
  assign n45489 = n45488 ^ n45333 ;
  assign n45490 = n45336 & n45489 ;
  assign n45492 = n45491 ^ n45490 ;
  assign n45493 = ~n45332 & ~n45492 ;
  assign n45494 = n45493 ^ n45331 ;
  assign n45495 = n45494 ^ n45326 ;
  assign n45496 = ~n45328 & ~n45495 ;
  assign n45498 = n45497 ^ n45496 ;
  assign n45499 = ~n45324 & n45498 ;
  assign n45500 = n45499 ^ n45323 ;
  assign n45501 = n45500 ^ n45319 ;
  assign n45502 = n45320 & ~n45501 ;
  assign n45505 = n45504 ^ n45502 ;
  assign n45509 = n44308 ^ n43083 ;
  assign n45510 = n45509 ^ n44509 ;
  assign n45506 = n45220 ^ n45165 ;
  assign n45507 = n45506 ^ n45503 ;
  assign n45508 = n45507 ^ n45506 ;
  assign n45511 = n45510 ^ n45508 ;
  assign n45512 = ~n45505 & ~n45511 ;
  assign n45513 = n45512 ^ n45507 ;
  assign n45621 = n45515 ^ n45513 ;
  assign n45623 = n45621 ^ n43036 ;
  assign n45564 = n45510 ^ n45505 ;
  assign n45565 = n45564 ^ n42873 ;
  assign n45566 = n45500 ^ n45320 ;
  assign n45567 = n45566 ^ n42860 ;
  assign n45568 = n45498 ^ n45323 ;
  assign n45569 = n45568 ^ n42849 ;
  assign n45570 = n45494 ^ n45328 ;
  assign n45571 = n45570 ^ n42825 ;
  assign n45604 = n45492 ^ n45330 ;
  assign n45572 = n45488 ^ n45336 ;
  assign n45573 = n45572 ^ n42029 ;
  assign n45574 = n45485 ^ n45340 ;
  assign n45575 = n45574 ^ n42036 ;
  assign n45593 = n45483 ^ n45342 ;
  assign n45576 = n45479 ^ n45461 ;
  assign n45577 = n45576 ^ n42701 ;
  assign n45585 = n45476 ^ n45465 ;
  assign n45580 = n45473 ^ n45472 ;
  assign n45578 = n45470 ^ n45469 ;
  assign n45579 = ~n42046 & ~n45578 ;
  assign n45581 = n45580 ^ n45579 ;
  assign n45582 = n45580 ^ n42686 ;
  assign n45583 = ~n45581 & ~n45582 ;
  assign n45584 = n45583 ^ n42686 ;
  assign n45586 = n45585 ^ n45584 ;
  assign n45587 = n45585 ^ n42696 ;
  assign n45588 = n45586 & n45587 ;
  assign n45589 = n45588 ^ n42696 ;
  assign n45590 = n45589 ^ n45576 ;
  assign n45591 = n45577 & ~n45590 ;
  assign n45592 = n45591 ^ n42701 ;
  assign n45594 = n45593 ^ n45592 ;
  assign n45595 = n45593 ^ n42710 ;
  assign n45596 = ~n45594 & n45595 ;
  assign n45597 = n45596 ^ n42710 ;
  assign n45598 = n45597 ^ n45574 ;
  assign n45599 = ~n45575 & n45598 ;
  assign n45600 = n45599 ^ n42036 ;
  assign n45601 = n45600 ^ n45572 ;
  assign n45602 = ~n45573 & ~n45601 ;
  assign n45603 = n45602 ^ n42029 ;
  assign n45605 = n45604 ^ n45603 ;
  assign n45606 = n45604 ^ n42720 ;
  assign n45607 = ~n45605 & ~n45606 ;
  assign n45608 = n45607 ^ n42720 ;
  assign n45609 = n45608 ^ n45570 ;
  assign n45610 = n45571 & ~n45609 ;
  assign n45611 = n45610 ^ n42825 ;
  assign n45612 = n45611 ^ n45568 ;
  assign n45613 = ~n45569 & n45612 ;
  assign n45614 = n45613 ^ n42849 ;
  assign n45615 = n45614 ^ n45566 ;
  assign n45616 = n45567 & ~n45615 ;
  assign n45617 = n45616 ^ n42860 ;
  assign n45618 = n45617 ^ n45564 ;
  assign n45619 = ~n45565 & ~n45618 ;
  assign n45620 = n45619 ^ n42873 ;
  assign n45676 = n45623 ^ n45620 ;
  assign n45654 = n45617 ^ n45565 ;
  assign n45655 = n45614 ^ n45567 ;
  assign n45656 = n45579 ^ n42686 ;
  assign n45657 = n45656 ^ n45580 ;
  assign n45658 = n45587 ^ n45584 ;
  assign n45659 = n45657 & n45658 ;
  assign n45660 = n45589 ^ n45577 ;
  assign n45661 = ~n45659 & n45660 ;
  assign n45662 = n45595 ^ n45592 ;
  assign n45663 = ~n45661 & ~n45662 ;
  assign n45664 = n45597 ^ n45575 ;
  assign n45665 = ~n45663 & ~n45664 ;
  assign n45666 = n45600 ^ n45573 ;
  assign n45667 = ~n45665 & n45666 ;
  assign n45668 = n45606 ^ n45603 ;
  assign n45669 = n45667 & ~n45668 ;
  assign n45670 = n45608 ^ n45571 ;
  assign n45671 = n45669 & ~n45670 ;
  assign n45672 = n45611 ^ n45569 ;
  assign n45673 = ~n45671 & ~n45672 ;
  assign n45674 = n45655 & n45673 ;
  assign n45675 = ~n45654 & n45674 ;
  assign n45797 = n45676 ^ n45675 ;
  assign n45794 = n43804 ^ n35573 ;
  assign n45795 = n45794 ^ n40131 ;
  assign n45796 = n45795 ^ n33926 ;
  assign n45798 = n45797 ^ n45796 ;
  assign n45802 = n45674 ^ n45654 ;
  assign n45799 = n43809 ^ n35578 ;
  assign n45800 = n45799 ^ n2440 ;
  assign n45801 = n45800 ^ n33931 ;
  assign n45803 = n45802 ^ n45801 ;
  assign n45804 = n45673 ^ n45655 ;
  assign n2398 = n2391 ^ n2349 ;
  assign n2423 = n2422 ^ n2398 ;
  assign n2430 = n2429 ^ n2423 ;
  assign n45805 = n45804 ^ n2430 ;
  assign n45807 = n43817 ^ n2278 ;
  assign n45808 = n45807 ^ n40141 ;
  assign n45809 = n45808 ^ n2414 ;
  assign n45806 = n45672 ^ n45671 ;
  assign n45810 = n45809 ^ n45806 ;
  assign n45811 = n43823 ^ n2260 ;
  assign n45812 = n45811 ^ n40146 ;
  assign n45813 = n45812 ^ n33941 ;
  assign n45878 = n45813 ^ n45806 ;
  assign n45814 = n45670 ^ n45669 ;
  assign n45815 = n45814 ^ n45813 ;
  assign n45817 = n43828 ^ n35590 ;
  assign n45818 = n45817 ^ n40151 ;
  assign n45819 = n45818 ^ n33946 ;
  assign n45816 = n45668 ^ n45667 ;
  assign n45820 = n45819 ^ n45816 ;
  assign n45822 = n43833 ^ n35594 ;
  assign n45823 = n45822 ^ n40155 ;
  assign n45824 = n45823 ^ n33951 ;
  assign n45872 = n45824 ^ n45816 ;
  assign n45821 = n45666 ^ n45665 ;
  assign n45825 = n45824 ^ n45821 ;
  assign n45829 = n45664 ^ n45663 ;
  assign n45826 = n43839 ^ n35624 ;
  assign n45827 = n45826 ^ n40161 ;
  assign n45828 = n45827 ^ n33955 ;
  assign n45830 = n45829 ^ n45828 ;
  assign n45831 = n43843 ^ n35616 ;
  assign n45832 = n45831 ^ n40185 ;
  assign n45833 = n45832 ^ n1928 ;
  assign n45866 = n45833 ^ n45829 ;
  assign n45834 = n45662 ^ n45661 ;
  assign n45835 = n45834 ^ n45833 ;
  assign n45839 = n45660 ^ n45659 ;
  assign n45836 = n43849 ^ n35612 ;
  assign n45837 = n45836 ^ n40165 ;
  assign n45838 = n45837 ^ n33281 ;
  assign n45840 = n45839 ^ n45838 ;
  assign n45842 = n43853 ^ n35599 ;
  assign n45843 = n45842 ^ n40169 ;
  assign n45844 = n45843 ^ n3242 ;
  assign n45841 = n45658 ^ n45657 ;
  assign n45845 = n45844 ^ n45841 ;
  assign n45849 = n45848 ^ n45657 ;
  assign n45850 = n44106 ^ n35958 ;
  assign n45851 = n45850 ^ n2684 ;
  assign n45852 = n45851 ^ n3227 ;
  assign n45853 = n45578 ^ n42046 ;
  assign n45854 = n45852 & n45853 ;
  assign n45855 = n45854 ^ n45657 ;
  assign n45856 = n45849 & ~n45855 ;
  assign n45857 = n45856 ^ n45848 ;
  assign n45858 = n45857 ^ n45844 ;
  assign n45859 = ~n45845 & n45858 ;
  assign n45860 = n45859 ^ n45844 ;
  assign n45861 = n45860 ^ n45838 ;
  assign n45862 = ~n45840 & ~n45861 ;
  assign n45863 = n45862 ^ n45839 ;
  assign n45864 = n45863 ^ n45833 ;
  assign n45865 = ~n45835 & ~n45864 ;
  assign n45867 = n45866 ^ n45865 ;
  assign n45868 = n45830 & n45867 ;
  assign n45869 = n45868 ^ n45829 ;
  assign n45870 = n45869 ^ n45824 ;
  assign n45871 = n45825 & n45870 ;
  assign n45873 = n45872 ^ n45871 ;
  assign n45874 = n45820 & ~n45873 ;
  assign n45875 = n45874 ^ n45819 ;
  assign n45876 = n45875 ^ n45813 ;
  assign n45877 = n45815 & n45876 ;
  assign n45879 = n45878 ^ n45877 ;
  assign n45880 = n45810 & ~n45879 ;
  assign n45881 = n45880 ^ n45809 ;
  assign n45882 = n45881 ^ n2430 ;
  assign n45883 = n45805 & ~n45882 ;
  assign n45884 = n45883 ^ n45804 ;
  assign n45885 = n45884 ^ n45801 ;
  assign n45886 = ~n45803 & ~n45885 ;
  assign n45887 = n45886 ^ n45802 ;
  assign n45888 = n45887 ^ n45796 ;
  assign n45889 = ~n45798 & n45888 ;
  assign n45890 = n45889 ^ n45797 ;
  assign n45677 = n45675 & ~n45676 ;
  assign n45622 = n45621 ^ n45620 ;
  assign n45624 = n45622 & n45623 ;
  assign n45625 = n45624 ^ n43036 ;
  assign n45522 = n44512 ^ n43071 ;
  assign n45523 = n45522 ^ n44495 ;
  assign n45516 = n45222 ^ n2201 ;
  assign n45518 = n45516 ^ n45506 ;
  assign n45517 = n45516 ^ n45515 ;
  assign n45519 = n45518 ^ n45517 ;
  assign n45520 = ~n45513 & n45519 ;
  assign n45521 = n45520 ^ n45518 ;
  assign n45562 = n45523 ^ n45521 ;
  assign n45563 = n45562 ^ n43091 ;
  assign n45653 = n45625 ^ n45563 ;
  assign n45792 = n45677 ^ n45653 ;
  assign n45789 = n43799 ^ n35657 ;
  assign n45790 = n45789 ^ n40126 ;
  assign n45791 = n45790 ^ n33922 ;
  assign n45793 = n45792 ^ n45791 ;
  assign n46232 = n45890 ^ n45793 ;
  assign n45950 = n45887 ^ n45798 ;
  assign n46233 = n46232 ^ n45950 ;
  assign n45948 = n44490 ^ n44468 ;
  assign n45722 = n45248 ^ n45118 ;
  assign n45949 = n45948 ^ n45722 ;
  assign n45951 = n45950 ^ n45949 ;
  assign n45954 = n45884 ^ n45803 ;
  assign n45952 = n44496 ^ n44470 ;
  assign n45708 = n45245 ^ n45123 ;
  assign n45953 = n45952 ^ n45708 ;
  assign n45955 = n45954 ^ n45953 ;
  assign n45958 = n45881 ^ n45805 ;
  assign n45956 = n44502 ^ n44478 ;
  assign n45691 = n45242 ^ n45128 ;
  assign n45957 = n45956 ^ n45691 ;
  assign n45959 = n45958 ^ n45957 ;
  assign n45962 = n45879 ^ n45809 ;
  assign n45960 = n44506 ^ n44480 ;
  assign n45550 = n45239 ^ n45133 ;
  assign n45961 = n45960 ^ n45550 ;
  assign n45963 = n45962 ^ n45961 ;
  assign n45966 = n45875 ^ n45815 ;
  assign n45964 = n44512 ^ n44488 ;
  assign n45302 = n45236 ^ n45138 ;
  assign n45965 = n45964 ^ n45302 ;
  assign n45967 = n45966 ^ n45965 ;
  assign n45970 = n45873 ^ n45819 ;
  assign n45306 = n45233 ^ n45143 ;
  assign n45968 = n45306 ^ n44452 ;
  assign n45969 = n45968 ^ n44493 ;
  assign n45971 = n45970 ^ n45969 ;
  assign n45974 = n45869 ^ n45825 ;
  assign n45972 = n44495 ^ n44308 ;
  assign n45312 = n45230 ^ n45148 ;
  assign n45973 = n45972 ^ n45312 ;
  assign n45975 = n45974 ^ n45973 ;
  assign n45978 = n45867 ^ n45828 ;
  assign n45976 = n44500 ^ n44261 ;
  assign n45311 = n45227 ^ n45153 ;
  assign n45977 = n45976 ^ n45311 ;
  assign n45979 = n45978 ^ n45977 ;
  assign n45982 = n45863 ^ n45835 ;
  assign n46208 = n45982 ^ n45978 ;
  assign n45980 = n44509 ^ n44175 ;
  assign n45524 = n45225 ^ n45156 ;
  assign n45981 = n45980 ^ n45524 ;
  assign n45983 = n45982 ^ n45981 ;
  assign n45986 = n45860 ^ n45840 ;
  assign n45984 = n44511 ^ n44038 ;
  assign n45985 = n45984 ^ n45516 ;
  assign n45987 = n45986 ^ n45985 ;
  assign n45990 = n45857 ^ n45845 ;
  assign n45988 = n44518 ^ n44034 ;
  assign n45989 = n45988 ^ n45506 ;
  assign n45991 = n45990 ^ n45989 ;
  assign n46192 = n44520 ^ n44043 ;
  assign n46193 = n46192 ^ n45503 ;
  assign n45994 = n45853 ^ n45852 ;
  assign n45992 = n44524 ^ n44047 ;
  assign n45993 = n45992 ^ n45319 ;
  assign n45995 = n45994 ^ n45993 ;
  assign n46152 = n44086 ^ n35936 ;
  assign n46153 = n46152 ^ n40340 ;
  assign n46154 = n46153 ^ n2676 ;
  assign n46036 = n44113 ^ n43428 ;
  assign n46037 = n46036 ^ n44771 ;
  assign n46000 = n45257 ^ n45103 ;
  assign n45998 = n43961 ^ n43438 ;
  assign n45999 = n45998 ^ n45371 ;
  assign n46001 = n46000 ^ n45999 ;
  assign n45928 = n44819 ^ n44028 ;
  assign n45929 = n45928 ^ n45345 ;
  assign n45931 = n45930 ^ n45929 ;
  assign n45732 = n45251 ^ n45113 ;
  assign n45733 = n45732 ^ n45722 ;
  assign n45723 = n44027 ^ n43992 ;
  assign n45724 = n45723 ^ n45354 ;
  assign n45725 = n45724 ^ n45722 ;
  assign n45709 = n44471 ^ n43946 ;
  assign n45710 = n45709 ^ n45277 ;
  assign n45711 = n45710 ^ n45708 ;
  assign n45551 = n44481 ^ n43652 ;
  assign n45552 = n45551 ^ n44468 ;
  assign n45553 = n45552 ^ n45550 ;
  assign n45303 = n44485 ^ n43521 ;
  assign n45304 = n45303 ^ n44470 ;
  assign n45305 = n45304 ^ n45302 ;
  assign n45308 = n44490 ^ n43048 ;
  assign n45309 = n45308 ^ n44478 ;
  assign n45310 = n45309 ^ n45306 ;
  assign n45314 = n44502 ^ n43061 ;
  assign n45315 = n45314 ^ n44488 ;
  assign n45316 = n45315 ^ n45311 ;
  assign n45526 = n45524 ^ n45516 ;
  assign n45525 = n45524 ^ n45523 ;
  assign n45527 = n45526 ^ n45525 ;
  assign n45528 = n45521 & n45527 ;
  assign n45529 = n45528 ^ n45526 ;
  assign n45533 = n45524 ^ n45311 ;
  assign n45530 = n44506 ^ n43066 ;
  assign n45531 = n45530 ^ n44493 ;
  assign n45532 = n45531 ^ n45311 ;
  assign n45534 = n45533 ^ n45532 ;
  assign n45535 = n45529 & ~n45534 ;
  assign n45536 = n45535 ^ n45533 ;
  assign n45537 = n45316 & ~n45536 ;
  assign n45313 = n45312 ^ n45311 ;
  assign n45538 = n45537 ^ n45313 ;
  assign n45541 = n44496 ^ n43056 ;
  assign n45542 = n45541 ^ n44480 ;
  assign n45539 = n45312 ^ n45306 ;
  assign n45540 = n45539 ^ n45306 ;
  assign n45543 = n45542 ^ n45540 ;
  assign n45544 = n45538 & n45543 ;
  assign n45545 = n45544 ^ n45539 ;
  assign n45546 = n45310 & ~n45545 ;
  assign n45307 = n45306 ^ n45302 ;
  assign n45547 = n45546 ^ n45307 ;
  assign n45548 = ~n45305 & ~n45547 ;
  assign n45549 = n45548 ^ n45304 ;
  assign n45693 = n45550 ^ n45549 ;
  assign n45694 = ~n45553 & n45693 ;
  assign n45692 = n45691 ^ n45550 ;
  assign n45695 = n45694 ^ n45692 ;
  assign n45696 = n44475 ^ n43665 ;
  assign n45697 = n45696 ^ n44907 ;
  assign n45705 = n45697 ^ n45691 ;
  assign n45706 = n45695 & n45705 ;
  assign n45707 = n45706 ^ n45697 ;
  assign n45719 = n45708 ^ n45707 ;
  assign n45720 = n45711 & ~n45719 ;
  assign n45721 = n45720 ^ n45710 ;
  assign n45730 = n45722 ^ n45721 ;
  assign n45731 = ~n45725 & ~n45730 ;
  assign n45734 = n45733 ^ n45731 ;
  assign n45735 = n44784 ^ n44071 ;
  assign n45736 = n45735 ^ n45349 ;
  assign n45925 = n45736 ^ n45732 ;
  assign n45926 = ~n45734 & n45925 ;
  assign n45927 = n45926 ^ n45736 ;
  assign n46005 = n45929 ^ n45927 ;
  assign n46006 = n45931 & n46005 ;
  assign n46007 = n46006 ^ n45930 ;
  assign n46002 = n45260 ^ n45098 ;
  assign n46003 = n46002 ^ n46000 ;
  assign n46004 = n46003 ^ n46002 ;
  assign n46008 = n46007 ^ n46004 ;
  assign n46009 = ~n46001 & n46008 ;
  assign n46010 = n46009 ^ n46003 ;
  assign n46013 = n45263 ^ n45093 ;
  assign n46015 = n46013 ^ n46002 ;
  assign n46011 = n43960 ^ n43446 ;
  assign n46012 = n46011 ^ n45297 ;
  assign n46014 = n46013 ^ n46012 ;
  assign n46016 = n46015 ^ n46014 ;
  assign n46017 = ~n46010 & ~n46016 ;
  assign n46018 = n46017 ^ n46015 ;
  assign n46021 = n45266 ^ n45091 ;
  assign n46023 = n46021 ^ n46013 ;
  assign n46019 = n44011 ^ n43436 ;
  assign n46020 = n46019 ^ n44724 ;
  assign n46022 = n46021 ^ n46020 ;
  assign n46024 = n46023 ^ n46022 ;
  assign n46025 = n46018 & n46024 ;
  assign n46026 = n46025 ^ n46023 ;
  assign n46029 = n45269 ^ n45086 ;
  assign n46031 = n46029 ^ n46021 ;
  assign n46027 = n44117 ^ n43430 ;
  assign n46028 = n46027 ^ n44774 ;
  assign n46030 = n46029 ^ n46028 ;
  assign n46032 = n46031 ^ n46030 ;
  assign n46033 = ~n46026 & ~n46032 ;
  assign n46034 = n46033 ^ n46031 ;
  assign n46047 = n46037 ^ n46034 ;
  assign n46048 = n46047 ^ n42622 ;
  assign n46049 = n46028 ^ n46026 ;
  assign n46050 = n46049 ^ n42632 ;
  assign n46052 = n46012 ^ n46010 ;
  assign n46053 = n46052 ^ n42640 ;
  assign n46054 = n46007 ^ n46001 ;
  assign n46055 = n46054 ^ n42641 ;
  assign n45932 = n45931 ^ n45927 ;
  assign n45933 = n45932 ^ n43328 ;
  assign n45737 = n45736 ^ n45734 ;
  assign n45738 = n45737 ^ n43146 ;
  assign n45726 = n45725 ^ n45721 ;
  assign n45727 = n45726 ^ n43050 ;
  assign n45712 = n45711 ^ n45707 ;
  assign n45713 = n45712 ^ n43054 ;
  assign n45698 = n45697 ^ n45695 ;
  assign n45699 = n45698 ^ n43059 ;
  assign n45643 = n45547 ^ n45304 ;
  assign n45556 = n45545 ^ n45309 ;
  assign n45557 = n45556 ^ n43074 ;
  assign n45558 = n45542 ^ n45538 ;
  assign n45559 = n45558 ^ n43081 ;
  assign n45560 = n45531 ^ n45529 ;
  assign n45561 = n45560 ^ n43086 ;
  assign n45626 = n45625 ^ n45562 ;
  assign n45627 = ~n45563 & n45626 ;
  assign n45628 = n45627 ^ n43091 ;
  assign n45629 = n45628 ^ n45560 ;
  assign n45630 = ~n45561 & ~n45629 ;
  assign n45631 = n45630 ^ n43086 ;
  assign n45632 = n45631 ^ n43172 ;
  assign n45633 = n45536 ^ n45315 ;
  assign n45634 = n45633 ^ n45631 ;
  assign n45635 = ~n45632 & ~n45634 ;
  assign n45636 = n45635 ^ n43172 ;
  assign n45637 = n45636 ^ n45558 ;
  assign n45638 = ~n45559 & ~n45637 ;
  assign n45639 = n45638 ^ n43081 ;
  assign n45640 = n45639 ^ n45556 ;
  assign n45641 = ~n45557 & n45640 ;
  assign n45642 = n45641 ^ n43074 ;
  assign n45644 = n45643 ^ n45642 ;
  assign n45645 = n45643 ^ n43069 ;
  assign n45646 = n45644 & ~n45645 ;
  assign n45647 = n45646 ^ n43069 ;
  assign n45554 = n45553 ^ n45549 ;
  assign n45687 = n45647 ^ n45554 ;
  assign n45688 = n45647 ^ n43064 ;
  assign n45689 = ~n45687 & ~n45688 ;
  assign n45690 = n45689 ^ n43064 ;
  assign n45702 = n45698 ^ n45690 ;
  assign n45703 = n45699 & ~n45702 ;
  assign n45704 = n45703 ^ n43059 ;
  assign n45716 = n45712 ^ n45704 ;
  assign n45717 = ~n45713 & n45716 ;
  assign n45718 = n45717 ^ n43054 ;
  assign n45739 = n45726 ^ n45718 ;
  assign n45740 = ~n45727 & ~n45739 ;
  assign n45741 = n45740 ^ n43050 ;
  assign n45922 = n45741 ^ n45737 ;
  assign n45923 = n45738 & n45922 ;
  assign n45924 = n45923 ^ n43146 ;
  assign n46056 = n45932 ^ n45924 ;
  assign n46057 = ~n45933 & ~n46056 ;
  assign n46058 = n46057 ^ n43328 ;
  assign n46059 = n46058 ^ n46054 ;
  assign n46060 = n46055 & n46059 ;
  assign n46061 = n46060 ^ n42641 ;
  assign n46062 = n46061 ^ n46052 ;
  assign n46063 = n46053 & ~n46062 ;
  assign n46064 = n46063 ^ n42640 ;
  assign n46051 = n46020 ^ n46018 ;
  assign n46065 = n46064 ^ n46051 ;
  assign n46066 = n46064 ^ n42634 ;
  assign n46067 = ~n46065 & ~n46066 ;
  assign n46068 = n46067 ^ n42634 ;
  assign n46069 = n46068 ^ n46049 ;
  assign n46070 = n46050 & ~n46069 ;
  assign n46071 = n46070 ^ n42632 ;
  assign n46072 = n46071 ^ n46047 ;
  assign n46073 = n46048 & n46072 ;
  assign n46074 = n46073 ^ n42622 ;
  assign n46043 = n44063 ^ n43136 ;
  assign n46044 = n46043 ^ n44802 ;
  assign n46035 = n45273 ^ n1447 ;
  assign n46039 = n46035 ^ n46029 ;
  assign n46038 = n46037 ^ n46035 ;
  assign n46040 = n46039 ^ n46038 ;
  assign n46041 = n46034 & ~n46040 ;
  assign n46042 = n46041 ^ n46039 ;
  assign n46045 = n46044 ^ n46042 ;
  assign n46146 = n46074 ^ n46045 ;
  assign n46076 = n46071 ^ n46048 ;
  assign n46077 = n46051 ^ n42634 ;
  assign n46078 = n46077 ^ n46064 ;
  assign n45555 = n45554 ^ n43064 ;
  assign n45648 = n45647 ^ n45555 ;
  assign n45649 = n45645 ^ n45642 ;
  assign n45650 = n45639 ^ n45557 ;
  assign n45651 = n45636 ^ n45559 ;
  assign n45652 = n45633 ^ n45632 ;
  assign n45678 = ~n45653 & n45677 ;
  assign n45679 = n45628 ^ n43086 ;
  assign n45680 = n45679 ^ n45560 ;
  assign n45681 = ~n45678 & n45680 ;
  assign n45682 = ~n45652 & n45681 ;
  assign n45683 = ~n45651 & ~n45682 ;
  assign n45684 = ~n45650 & ~n45683 ;
  assign n45685 = n45649 & ~n45684 ;
  assign n45686 = n45648 & n45685 ;
  assign n45700 = n45699 ^ n45690 ;
  assign n45701 = n45686 & n45700 ;
  assign n45714 = n45713 ^ n45704 ;
  assign n45715 = ~n45701 & n45714 ;
  assign n45728 = n45727 ^ n45718 ;
  assign n45729 = n45715 & n45728 ;
  assign n45742 = n45741 ^ n45738 ;
  assign n45921 = ~n45729 & ~n45742 ;
  assign n45934 = n45933 ^ n45924 ;
  assign n46079 = n45921 & ~n45934 ;
  assign n46080 = n46058 ^ n46055 ;
  assign n46081 = ~n46079 & n46080 ;
  assign n46082 = n46061 ^ n46053 ;
  assign n46083 = ~n46081 & n46082 ;
  assign n46084 = n46078 & ~n46083 ;
  assign n46085 = n46068 ^ n46050 ;
  assign n46086 = ~n46084 & ~n46085 ;
  assign n46087 = ~n46076 & n46086 ;
  assign n46149 = n46146 ^ n46087 ;
  assign n46150 = n42665 & n46149 ;
  assign n46147 = n46087 ^ n46045 ;
  assign n46148 = ~n46146 & ~n46147 ;
  assign n46151 = n46150 ^ n46148 ;
  assign n46155 = n46154 ^ n46151 ;
  assign n46144 = n42665 ^ n42059 ;
  assign n46140 = n44056 ^ n43132 ;
  assign n46141 = n46140 ^ n46044 ;
  assign n46142 = n46141 ^ n44833 ;
  assign n45296 = n45295 ^ n45275 ;
  assign n46143 = n46142 ^ n45296 ;
  assign n46145 = n46144 ^ n46143 ;
  assign n46156 = n46155 ^ n46145 ;
  assign n46089 = n44009 ^ n2657 ;
  assign n46090 = n46089 ^ n40284 ;
  assign n46091 = n46090 ^ n34215 ;
  assign n46157 = n46156 ^ n46091 ;
  assign n46138 = n46044 ^ n46035 ;
  assign n46139 = n46042 & ~n46138 ;
  assign n46158 = n46157 ^ n46139 ;
  assign n46046 = n46045 ^ n42665 ;
  assign n46075 = n46074 ^ n46046 ;
  assign n46088 = n46087 ^ n46075 ;
  assign n46092 = n46091 ^ n46088 ;
  assign n46093 = n43942 ^ n35773 ;
  assign n46094 = n46093 ^ n38845 ;
  assign n46095 = n46094 ^ n34204 ;
  assign n46135 = n46095 ^ n46088 ;
  assign n46096 = n46086 ^ n46076 ;
  assign n46097 = n46096 ^ n46095 ;
  assign n46099 = n35731 ^ n2903 ;
  assign n46100 = n46099 ^ n40060 ;
  assign n46101 = n46100 ^ n34021 ;
  assign n46098 = n46085 ^ n46084 ;
  assign n46102 = n46101 ^ n46098 ;
  assign n46106 = n46083 ^ n46078 ;
  assign n46103 = n43738 ^ n34061 ;
  assign n46104 = n46103 ^ n40065 ;
  assign n46105 = n46104 ^ n33828 ;
  assign n46107 = n46106 ^ n46105 ;
  assign n46108 = n43743 ^ n2850 ;
  assign n46109 = n46108 ^ n40070 ;
  assign n46110 = n46109 ^ n33833 ;
  assign n46126 = n46110 ^ n46106 ;
  assign n46111 = n46082 ^ n46081 ;
  assign n46112 = n46111 ^ n46110 ;
  assign n46114 = n35529 ^ n1774 ;
  assign n46115 = n46114 ^ n40075 ;
  assign n46116 = n46115 ^ n33838 ;
  assign n46113 = n46080 ^ n46079 ;
  assign n46117 = n46116 ^ n46113 ;
  assign n45935 = n45934 ^ n45921 ;
  assign n45299 = n43751 ^ n1739 ;
  assign n45300 = n45299 ^ n1091 ;
  assign n45301 = n45300 ^ n33845 ;
  assign n45936 = n45935 ^ n45301 ;
  assign n45743 = n45742 ^ n45729 ;
  assign n45744 = n45743 ^ n45301 ;
  assign n45748 = n45728 ^ n45715 ;
  assign n45745 = n43757 ^ n1730 ;
  assign n45746 = n45745 ^ n40086 ;
  assign n45747 = n45746 ^ n1083 ;
  assign n45749 = n45748 ^ n45747 ;
  assign n45751 = n45714 ^ n45701 ;
  assign n930 = n929 ^ n893 ;
  assign n958 = n957 ^ n930 ;
  assign n965 = n964 ^ n958 ;
  assign n45752 = n45751 ^ n965 ;
  assign n45756 = n45700 ^ n45686 ;
  assign n45753 = n43763 ^ n35545 ;
  assign n45754 = n45753 ^ n40093 ;
  assign n45755 = n45754 ^ n949 ;
  assign n45757 = n45756 ^ n45755 ;
  assign n45761 = n45685 ^ n45648 ;
  assign n45762 = n45761 ^ n45760 ;
  assign n45907 = n45766 ^ n45761 ;
  assign n45763 = n45684 ^ n45649 ;
  assign n45767 = n45766 ^ n45763 ;
  assign n45769 = n43778 ^ n1574 ;
  assign n45770 = n45769 ^ n40106 ;
  assign n45771 = n45770 ^ n33880 ;
  assign n45904 = n45771 ^ n45763 ;
  assign n45768 = n45683 ^ n45650 ;
  assign n45772 = n45771 ^ n45768 ;
  assign n45776 = n45682 ^ n45651 ;
  assign n45901 = n45776 ^ n45768 ;
  assign n45773 = n43783 ^ n35563 ;
  assign n45774 = n45773 ^ n40111 ;
  assign n45775 = n45774 ^ n33909 ;
  assign n45777 = n45776 ^ n45775 ;
  assign n45782 = n45681 ^ n45652 ;
  assign n45778 = n43790 ^ n35558 ;
  assign n45779 = n45778 ^ n40117 ;
  assign n45780 = n45779 ^ n2957 ;
  assign n45783 = n45782 ^ n45780 ;
  assign n45785 = n43795 ^ n35568 ;
  assign n45786 = n45785 ^ n40122 ;
  assign n45787 = n45786 ^ n33917 ;
  assign n45784 = n45680 ^ n45678 ;
  assign n45788 = n45787 ^ n45784 ;
  assign n45891 = n45890 ^ n45791 ;
  assign n45892 = ~n45793 & n45891 ;
  assign n45893 = n45892 ^ n45792 ;
  assign n45894 = n45893 ^ n45787 ;
  assign n45895 = n45788 & ~n45894 ;
  assign n45896 = n45895 ^ n45787 ;
  assign n45897 = n45896 ^ n45780 ;
  assign n45898 = n45783 & n45897 ;
  assign n45781 = n45780 ^ n45775 ;
  assign n45899 = n45898 ^ n45781 ;
  assign n45900 = n45777 & ~n45899 ;
  assign n45902 = n45901 ^ n45900 ;
  assign n45903 = ~n45772 & n45902 ;
  assign n45905 = n45904 ^ n45903 ;
  assign n45906 = ~n45767 & n45905 ;
  assign n45908 = n45907 ^ n45906 ;
  assign n45909 = n45762 & n45908 ;
  assign n45910 = n45909 ^ n45761 ;
  assign n45911 = n45910 ^ n45755 ;
  assign n45912 = n45757 & ~n45911 ;
  assign n45913 = n45912 ^ n45756 ;
  assign n45914 = n45913 ^ n965 ;
  assign n45915 = n45752 & n45914 ;
  assign n45750 = n45748 ^ n965 ;
  assign n45916 = n45915 ^ n45750 ;
  assign n45917 = ~n45749 & ~n45916 ;
  assign n45918 = n45917 ^ n45748 ;
  assign n45919 = n45918 ^ n45301 ;
  assign n45920 = n45744 & ~n45919 ;
  assign n45937 = n45936 ^ n45920 ;
  assign n45938 = n35534 ^ n1759 ;
  assign n45939 = n45938 ^ n40079 ;
  assign n45940 = n45939 ^ n1262 ;
  assign n46118 = n45940 ^ n45935 ;
  assign n46119 = n45937 & ~n46118 ;
  assign n46120 = n46119 ^ n45940 ;
  assign n46121 = n46120 ^ n46113 ;
  assign n46122 = n46117 & ~n46121 ;
  assign n46123 = n46122 ^ n46116 ;
  assign n46124 = n46123 ^ n46110 ;
  assign n46125 = ~n46112 & n46124 ;
  assign n46127 = n46126 ^ n46125 ;
  assign n46128 = n46107 & n46127 ;
  assign n46129 = n46128 ^ n46106 ;
  assign n46130 = n46129 ^ n46098 ;
  assign n46131 = n46102 & ~n46130 ;
  assign n46132 = n46131 ^ n46101 ;
  assign n46133 = n46132 ^ n46095 ;
  assign n46134 = ~n46097 & n46133 ;
  assign n46136 = n46135 ^ n46134 ;
  assign n46137 = ~n46092 & n46136 ;
  assign n46159 = n46158 ^ n46137 ;
  assign n45996 = n44528 ^ n44049 ;
  assign n45997 = n45996 ^ n45321 ;
  assign n46160 = n46159 ^ n45997 ;
  assign n46163 = n46136 ^ n46091 ;
  assign n46185 = n46163 ^ n46159 ;
  assign n46161 = n44534 ^ n44152 ;
  assign n46162 = n46161 ^ n45327 ;
  assign n46164 = n46163 ^ n46162 ;
  assign n46167 = n46132 ^ n46097 ;
  assign n46165 = n44536 ^ n44144 ;
  assign n46166 = n46165 ^ n45331 ;
  assign n46168 = n46167 ^ n46166 ;
  assign n46174 = n44542 ^ n44134 ;
  assign n46175 = n46174 ^ n45333 ;
  assign n46169 = n44058 ^ n44023 ;
  assign n46170 = n46169 ^ n45339 ;
  assign n46171 = n46127 ^ n46105 ;
  assign n46172 = ~n46170 & n46171 ;
  assign n46176 = n46175 ^ n46172 ;
  assign n46177 = n46129 ^ n46102 ;
  assign n46178 = n46177 ^ n46172 ;
  assign n46179 = n46176 & n46178 ;
  assign n46173 = n46172 ^ n46167 ;
  assign n46180 = n46179 ^ n46173 ;
  assign n46181 = n46168 & ~n46180 ;
  assign n46182 = n46181 ^ n46167 ;
  assign n46183 = n46182 ^ n46163 ;
  assign n46184 = n46164 & n46183 ;
  assign n46186 = n46185 ^ n46184 ;
  assign n46187 = ~n46160 & ~n46186 ;
  assign n46188 = n46187 ^ n46159 ;
  assign n46189 = n46188 ^ n45993 ;
  assign n46190 = ~n45995 & n46189 ;
  assign n46191 = n46190 ^ n45994 ;
  assign n46194 = n46193 ^ n46191 ;
  assign n46195 = n45854 ^ n45849 ;
  assign n46198 = n46195 ^ n46191 ;
  assign n46199 = n46194 & n46198 ;
  assign n46196 = n46195 ^ n45990 ;
  assign n46200 = n46199 ^ n46196 ;
  assign n46201 = ~n45991 & ~n46200 ;
  assign n46202 = n46201 ^ n45990 ;
  assign n46203 = n46202 ^ n45986 ;
  assign n46204 = n45987 & n46203 ;
  assign n46205 = n46204 ^ n46202 ;
  assign n46206 = n46205 ^ n45981 ;
  assign n46207 = ~n45983 & ~n46206 ;
  assign n46209 = n46208 ^ n46207 ;
  assign n46210 = n45979 & n46209 ;
  assign n46211 = n46210 ^ n45978 ;
  assign n46212 = n46211 ^ n45973 ;
  assign n46213 = n45975 & ~n46212 ;
  assign n46214 = n46213 ^ n45974 ;
  assign n46215 = n46214 ^ n45969 ;
  assign n46216 = n45971 & ~n46215 ;
  assign n46217 = n46216 ^ n45970 ;
  assign n46218 = n46217 ^ n45965 ;
  assign n46219 = ~n45967 & n46218 ;
  assign n46220 = n46219 ^ n45966 ;
  assign n46221 = n46220 ^ n45961 ;
  assign n46222 = n45963 & ~n46221 ;
  assign n46223 = n46222 ^ n45962 ;
  assign n46224 = n46223 ^ n45957 ;
  assign n46225 = n45959 & ~n46224 ;
  assign n46226 = n46225 ^ n45958 ;
  assign n46227 = n46226 ^ n45953 ;
  assign n46228 = ~n45955 & ~n46227 ;
  assign n46229 = n46228 ^ n45954 ;
  assign n46230 = n46229 ^ n45950 ;
  assign n46231 = ~n45951 & ~n46230 ;
  assign n46234 = n46233 ^ n46231 ;
  assign n46521 = n45893 ^ n45788 ;
  assign n46522 = n46521 ^ n46232 ;
  assign n46523 = n46522 ^ n46521 ;
  assign n45946 = n44907 ^ n44485 ;
  assign n45947 = n45946 ^ n45732 ;
  assign n46524 = n46523 ^ n45947 ;
  assign n46525 = n46234 & ~n46524 ;
  assign n46526 = n46525 ^ n46522 ;
  assign n46529 = n46528 ^ n46526 ;
  assign n46530 = n46529 ^ n43652 ;
  assign n46236 = n46226 ^ n45955 ;
  assign n46237 = n46236 ^ n43056 ;
  assign n46239 = n46217 ^ n45967 ;
  assign n46240 = n46239 ^ n43071 ;
  assign n46241 = n46214 ^ n45971 ;
  assign n46242 = n46241 ^ n43076 ;
  assign n46244 = n46202 ^ n45987 ;
  assign n46245 = n46244 ^ n43093 ;
  assign n46280 = n46200 ^ n45989 ;
  assign n46246 = n46195 ^ n46193 ;
  assign n46247 = n46246 ^ n46191 ;
  assign n46248 = n46247 ^ n43102 ;
  assign n46249 = n46188 ^ n45995 ;
  assign n46250 = n46249 ^ n43106 ;
  assign n46251 = n46186 ^ n45997 ;
  assign n46252 = n46251 ^ n43110 ;
  assign n46253 = n46182 ^ n46164 ;
  assign n46254 = n46253 ^ n43114 ;
  assign n46255 = n46180 ^ n46166 ;
  assign n46256 = n46255 ^ n43118 ;
  assign n46259 = n46177 ^ n46176 ;
  assign n46257 = n46171 ^ n46170 ;
  assign n46258 = ~n43126 & ~n46257 ;
  assign n46260 = n46259 ^ n46258 ;
  assign n46261 = n46255 ^ n43120 ;
  assign n46262 = n46261 ^ n46255 ;
  assign n46263 = n46262 ^ n46258 ;
  assign n46264 = ~n46260 & n46263 ;
  assign n46265 = n46264 ^ n46261 ;
  assign n46266 = ~n46256 & ~n46265 ;
  assign n46267 = n46266 ^ n43118 ;
  assign n46268 = n46267 ^ n46253 ;
  assign n46269 = ~n46254 & ~n46268 ;
  assign n46270 = n46269 ^ n43114 ;
  assign n46271 = n46270 ^ n46251 ;
  assign n46272 = ~n46252 & ~n46271 ;
  assign n46273 = n46272 ^ n43110 ;
  assign n46274 = n46273 ^ n46249 ;
  assign n46275 = n46250 & ~n46274 ;
  assign n46276 = n46275 ^ n43106 ;
  assign n46277 = n46276 ^ n46247 ;
  assign n46278 = n46248 & ~n46277 ;
  assign n46279 = n46278 ^ n43102 ;
  assign n46281 = n46280 ^ n46279 ;
  assign n46282 = n46244 ^ n43095 ;
  assign n46283 = n46282 ^ n46279 ;
  assign n46284 = n46283 ^ n46244 ;
  assign n46285 = ~n46281 & n46284 ;
  assign n46286 = n46285 ^ n46282 ;
  assign n46287 = ~n46245 & n46286 ;
  assign n46288 = n46287 ^ n43093 ;
  assign n46243 = n46205 ^ n45983 ;
  assign n46289 = n46288 ^ n46243 ;
  assign n46290 = n46209 ^ n45977 ;
  assign n46291 = n46290 ^ n43088 ;
  assign n46292 = n46291 ^ n46288 ;
  assign n46293 = n46292 ^ n46290 ;
  assign n46294 = n46289 & n46293 ;
  assign n46295 = n46294 ^ n46291 ;
  assign n46296 = n46211 ^ n45975 ;
  assign n46298 = n46296 ^ n43495 ;
  assign n46297 = n46296 ^ n46290 ;
  assign n46299 = n46298 ^ n46297 ;
  assign n46300 = n46295 & ~n46299 ;
  assign n46301 = n46300 ^ n46298 ;
  assign n46303 = n46241 ^ n43083 ;
  assign n46302 = n46296 ^ n46241 ;
  assign n46304 = n46303 ^ n46302 ;
  assign n46305 = n46301 & n46304 ;
  assign n46306 = n46305 ^ n46303 ;
  assign n46307 = ~n46242 & ~n46306 ;
  assign n46308 = n46307 ^ n43076 ;
  assign n46309 = n46308 ^ n46239 ;
  assign n46310 = ~n46240 & ~n46309 ;
  assign n46311 = n46310 ^ n43071 ;
  assign n46312 = n46311 ^ n43066 ;
  assign n46313 = n46220 ^ n45963 ;
  assign n46314 = n46313 ^ n46311 ;
  assign n46315 = n46312 & ~n46314 ;
  assign n46316 = n46315 ^ n43066 ;
  assign n46238 = n46223 ^ n45959 ;
  assign n46317 = n46316 ^ n46238 ;
  assign n46318 = n46236 ^ n43061 ;
  assign n46319 = n46318 ^ n46236 ;
  assign n46320 = n46319 ^ n46238 ;
  assign n46321 = ~n46317 & ~n46320 ;
  assign n46322 = n46321 ^ n46318 ;
  assign n46323 = n46237 & ~n46322 ;
  assign n46324 = n46323 ^ n43056 ;
  assign n46325 = n46324 ^ n43048 ;
  assign n46326 = n46229 ^ n45951 ;
  assign n46327 = n46326 ^ n46324 ;
  assign n46328 = ~n46325 & n46327 ;
  assign n46329 = n46328 ^ n43048 ;
  assign n46330 = n46329 ^ n43521 ;
  assign n46235 = n46234 ^ n45947 ;
  assign n46518 = n46329 ^ n46235 ;
  assign n46519 = n46330 & n46518 ;
  assign n46520 = n46519 ^ n43521 ;
  assign n46531 = n46530 ^ n46520 ;
  assign n46331 = n46330 ^ n46235 ;
  assign n46332 = n46238 ^ n43061 ;
  assign n46333 = n46332 ^ n46316 ;
  assign n46334 = n46313 ^ n46312 ;
  assign n46335 = n46286 ^ n43093 ;
  assign n46336 = n46280 ^ n43095 ;
  assign n46337 = n46336 ^ n46279 ;
  assign n46338 = n46267 ^ n46254 ;
  assign n46339 = n46265 ^ n43118 ;
  assign n46340 = n46258 ^ n43120 ;
  assign n46341 = n46340 ^ n46259 ;
  assign n46342 = n46339 & ~n46341 ;
  assign n46343 = n46338 & ~n46342 ;
  assign n46344 = n46270 ^ n46252 ;
  assign n46345 = ~n46343 & n46344 ;
  assign n46346 = n46273 ^ n46250 ;
  assign n46347 = ~n46345 & ~n46346 ;
  assign n46348 = n46276 ^ n46248 ;
  assign n46349 = ~n46347 & n46348 ;
  assign n46350 = n46337 & n46349 ;
  assign n46351 = ~n46335 & n46350 ;
  assign n46352 = n46289 ^ n43088 ;
  assign n46353 = ~n46351 & n46352 ;
  assign n46354 = n46295 ^ n43495 ;
  assign n46355 = n46353 & n46354 ;
  assign n46356 = n46301 ^ n43083 ;
  assign n46357 = n46355 & ~n46356 ;
  assign n46358 = n46306 ^ n43076 ;
  assign n46359 = n46357 & ~n46358 ;
  assign n46360 = n46308 ^ n46240 ;
  assign n46361 = n46359 & n46360 ;
  assign n46362 = ~n46334 & ~n46361 ;
  assign n46363 = n46333 & n46362 ;
  assign n46364 = n46322 ^ n43056 ;
  assign n46365 = ~n46363 & ~n46364 ;
  assign n46366 = n46326 ^ n46325 ;
  assign n46367 = ~n46365 & n46366 ;
  assign n46517 = ~n46331 & ~n46367 ;
  assign n46532 = n46531 ^ n46517 ;
  assign n46514 = n44033 ^ n1632 ;
  assign n46515 = n46514 ^ n40862 ;
  assign n46516 = n46515 ^ n34517 ;
  assign n46533 = n46532 ^ n46516 ;
  assign n46754 = n46517 & n46531 ;
  assign n46648 = n45896 ^ n45783 ;
  assign n46654 = n46648 ^ n46521 ;
  assign n46652 = n46528 ^ n46521 ;
  assign n46653 = ~n46526 & ~n46652 ;
  assign n46655 = n46654 ^ n46653 ;
  assign n46649 = n46000 ^ n45354 ;
  assign n46650 = n46649 ^ n44475 ;
  assign n46690 = n46655 ^ n46650 ;
  assign n46752 = n46690 ^ n43665 ;
  assign n46691 = n46529 ^ n46520 ;
  assign n46692 = n46530 & n46691 ;
  assign n46693 = n46692 ^ n43652 ;
  assign n46753 = n46752 ^ n46693 ;
  assign n46816 = n46754 ^ n46753 ;
  assign n46817 = n46816 ^ n46516 ;
  assign n46818 = n46817 ^ n46816 ;
  assign n46368 = n46367 ^ n46331 ;
  assign n45943 = n44323 ^ n36322 ;
  assign n45944 = n45943 ^ n2984 ;
  assign n45945 = n45944 ^ n34522 ;
  assign n46369 = n46368 ^ n45945 ;
  assign n46510 = n46373 ^ n45945 ;
  assign n46370 = n46366 ^ n46365 ;
  assign n46374 = n46373 ^ n46370 ;
  assign n46378 = n46364 ^ n46363 ;
  assign n46375 = n44334 ^ n2966 ;
  assign n46376 = n46375 ^ n40874 ;
  assign n46377 = n46376 ^ n34553 ;
  assign n46379 = n46378 ^ n46377 ;
  assign n46381 = n44338 ^ n36335 ;
  assign n46382 = n46381 ^ n40879 ;
  assign n46383 = n46382 ^ n34558 ;
  assign n46504 = n46383 ^ n46377 ;
  assign n46380 = n46362 ^ n46333 ;
  assign n46384 = n46383 ^ n46380 ;
  assign n46386 = n44343 ^ n36342 ;
  assign n46387 = n46386 ^ n40884 ;
  assign n46388 = n46387 ^ n34563 ;
  assign n46501 = n46388 ^ n46383 ;
  assign n46385 = n46361 ^ n46334 ;
  assign n46389 = n46388 ^ n46385 ;
  assign n46393 = n46360 ^ n46359 ;
  assign n46390 = n44348 ^ n36347 ;
  assign n46391 = n46390 ^ n40889 ;
  assign n46392 = n46391 ^ n34569 ;
  assign n46394 = n46393 ^ n46392 ;
  assign n46398 = n46358 ^ n46357 ;
  assign n46395 = n44353 ^ n36351 ;
  assign n46396 = n46395 ^ n40895 ;
  assign n46397 = n46396 ^ n34574 ;
  assign n46399 = n46398 ^ n46397 ;
  assign n46403 = n46356 ^ n46355 ;
  assign n46400 = n44359 ^ n36357 ;
  assign n46401 = n46400 ^ n40902 ;
  assign n46402 = n46401 ^ n34580 ;
  assign n46404 = n46403 ^ n46402 ;
  assign n46482 = n46354 ^ n46353 ;
  assign n46408 = n46352 ^ n46351 ;
  assign n46405 = n44364 ^ n36367 ;
  assign n46406 = n46405 ^ n40911 ;
  assign n46407 = n46406 ^ n34586 ;
  assign n46409 = n46408 ^ n46407 ;
  assign n46470 = n46350 ^ n46335 ;
  assign n46413 = n46349 ^ n46337 ;
  assign n46410 = n44371 ^ n36402 ;
  assign n46411 = n46410 ^ n2072 ;
  assign n46412 = n46411 ^ n34613 ;
  assign n46414 = n46413 ^ n46412 ;
  assign n46418 = n46348 ^ n46347 ;
  assign n46415 = n44376 ^ n36377 ;
  assign n46416 = n46415 ^ n40448 ;
  assign n46417 = n46416 ^ n2064 ;
  assign n46419 = n46418 ^ n46417 ;
  assign n46423 = n46346 ^ n46345 ;
  assign n46420 = n44381 ^ n1970 ;
  assign n46421 = n46420 ^ n40424 ;
  assign n46422 = n46421 ^ n34621 ;
  assign n46424 = n46423 ^ n46422 ;
  assign n46426 = n44387 ^ n36384 ;
  assign n46427 = n46426 ^ n3089 ;
  assign n46428 = n46427 ^ n34625 ;
  assign n46460 = n46428 ^ n46423 ;
  assign n46425 = n46344 ^ n46343 ;
  assign n46429 = n46428 ^ n46425 ;
  assign n46431 = n43984 ^ n35785 ;
  assign n46432 = n46431 ^ n40363 ;
  assign n46433 = n46432 ^ n3081 ;
  assign n46430 = n46342 ^ n46338 ;
  assign n46434 = n46433 ^ n46430 ;
  assign n46436 = n3023 ^ n2783 ;
  assign n46437 = n46436 ^ n40372 ;
  assign n46438 = n46437 ^ n34632 ;
  assign n46435 = n46341 ^ n46339 ;
  assign n46439 = n46438 ^ n46435 ;
  assign n46440 = n43976 ^ n3230 ;
  assign n46441 = n46440 ^ n40367 ;
  assign n46442 = n46441 ^ n34054 ;
  assign n46443 = n46442 ^ n46341 ;
  assign n46444 = n44818 ^ n2724 ;
  assign n46445 = n46444 ^ n41244 ;
  assign n46446 = n46445 ^ n35198 ;
  assign n46447 = n46257 ^ n43126 ;
  assign n46448 = n46446 & n46447 ;
  assign n46449 = n46448 ^ n46442 ;
  assign n46450 = ~n46443 & ~n46449 ;
  assign n46451 = n46450 ^ n46341 ;
  assign n46452 = n46451 ^ n46435 ;
  assign n46453 = n46439 & n46452 ;
  assign n46454 = n46453 ^ n46438 ;
  assign n46455 = n46454 ^ n46430 ;
  assign n46456 = ~n46434 & n46455 ;
  assign n46457 = n46456 ^ n46433 ;
  assign n46458 = n46457 ^ n46428 ;
  assign n46459 = n46429 & n46458 ;
  assign n46461 = n46460 ^ n46459 ;
  assign n46462 = n46424 & n46461 ;
  assign n46463 = n46462 ^ n46423 ;
  assign n46464 = n46463 ^ n46417 ;
  assign n46465 = n46419 & ~n46464 ;
  assign n46466 = n46465 ^ n46418 ;
  assign n46467 = n46466 ^ n46412 ;
  assign n46468 = ~n46414 & ~n46467 ;
  assign n46469 = n46468 ^ n46413 ;
  assign n46471 = n46470 ^ n46469 ;
  assign n46472 = n44408 ^ n36372 ;
  assign n46473 = n46472 ^ n40916 ;
  assign n46474 = n46473 ^ n2165 ;
  assign n46477 = n46474 ^ n46469 ;
  assign n46478 = n46471 & ~n46477 ;
  assign n46475 = n46474 ^ n46407 ;
  assign n46479 = n46478 ^ n46475 ;
  assign n46480 = ~n46409 & ~n46479 ;
  assign n46481 = n46480 ^ n46408 ;
  assign n46483 = n46482 ^ n46481 ;
  assign n46484 = n44417 ^ n36362 ;
  assign n46485 = n46484 ^ n40906 ;
  assign n46486 = n46485 ^ n34591 ;
  assign n46487 = n46486 ^ n46481 ;
  assign n46488 = n46483 & ~n46487 ;
  assign n46489 = n46488 ^ n46486 ;
  assign n46490 = n46489 ^ n46402 ;
  assign n46491 = ~n46404 & ~n46490 ;
  assign n46492 = n46491 ^ n46403 ;
  assign n46493 = n46492 ^ n46397 ;
  assign n46494 = ~n46399 & n46493 ;
  assign n46495 = n46494 ^ n46398 ;
  assign n46496 = n46495 ^ n46392 ;
  assign n46497 = n46394 & n46496 ;
  assign n46498 = n46497 ^ n46393 ;
  assign n46499 = n46498 ^ n46388 ;
  assign n46500 = ~n46389 & n46499 ;
  assign n46502 = n46501 ^ n46500 ;
  assign n46503 = ~n46384 & n46502 ;
  assign n46505 = n46504 ^ n46503 ;
  assign n46506 = n46379 & ~n46505 ;
  assign n46507 = n46506 ^ n46378 ;
  assign n46508 = n46507 ^ n46370 ;
  assign n46509 = n46374 & ~n46508 ;
  assign n46511 = n46510 ^ n46509 ;
  assign n46512 = n46369 & ~n46511 ;
  assign n46513 = n46512 ^ n46368 ;
  assign n46819 = n46818 ^ n46513 ;
  assign n46820 = n46533 & n46819 ;
  assign n46821 = n46820 ^ n46817 ;
  assign n1659 = n1658 ^ n1030 ;
  assign n1675 = n1674 ^ n1659 ;
  assign n1679 = n1678 ^ n1675 ;
  assign n46826 = n46816 ^ n1679 ;
  assign n46822 = n44450 ^ n36317 ;
  assign n46823 = n46822 ^ n40857 ;
  assign n46824 = n46823 ^ n1669 ;
  assign n46825 = n46824 ^ n1679 ;
  assign n46827 = n46826 ^ n46825 ;
  assign n46828 = n46821 & n46827 ;
  assign n46829 = n46828 ^ n46826 ;
  assign n46694 = n46693 ^ n46690 ;
  assign n46651 = n46650 ^ n46648 ;
  assign n46656 = ~n46651 & n46655 ;
  assign n46657 = n46656 ^ n46650 ;
  assign n46645 = n45349 ^ n44471 ;
  assign n46646 = n46645 ^ n46002 ;
  assign n46568 = n45899 ^ n45776 ;
  assign n46647 = n46646 ^ n46568 ;
  assign n46695 = n46657 ^ n46647 ;
  assign n46696 = n46695 ^ n43665 ;
  assign n46697 = n46696 ^ n46690 ;
  assign n46698 = n46697 ^ n46695 ;
  assign n46699 = n46694 & ~n46698 ;
  assign n46700 = n46699 ^ n46696 ;
  assign n46756 = n46700 ^ n43946 ;
  assign n46755 = n46753 & n46754 ;
  assign n46814 = n46756 ^ n46755 ;
  assign n47113 = n46829 ^ n46814 ;
  assign n47111 = n45473 ^ n44774 ;
  assign n46862 = n46123 ^ n46112 ;
  assign n47112 = n47111 ^ n46862 ;
  assign n47114 = n47113 ^ n47112 ;
  assign n46974 = n46824 ^ n46821 ;
  assign n46972 = n45470 ^ n44724 ;
  assign n46745 = n46120 ^ n46117 ;
  assign n46973 = n46972 ^ n46745 ;
  assign n46975 = n46974 ^ n46973 ;
  assign n46534 = n46533 ^ n46513 ;
  assign n45941 = n45940 ^ n45937 ;
  assign n45298 = n45297 ^ n45296 ;
  assign n45942 = n45941 ^ n45298 ;
  assign n46535 = n46534 ^ n45942 ;
  assign n46539 = n46511 ^ n46368 ;
  assign n46537 = n45918 ^ n45744 ;
  assign n46536 = n46035 ^ n45371 ;
  assign n46538 = n46537 ^ n46536 ;
  assign n46540 = n46539 ^ n46538 ;
  assign n46544 = n46507 ^ n46374 ;
  assign n46542 = n45916 ^ n45747 ;
  assign n46541 = n46029 ^ n45345 ;
  assign n46543 = n46542 ^ n46541 ;
  assign n46545 = n46544 ^ n46543 ;
  assign n46549 = n46505 ^ n46378 ;
  assign n46547 = n45913 ^ n45752 ;
  assign n46546 = n46021 ^ n45349 ;
  assign n46548 = n46547 ^ n46546 ;
  assign n46550 = n46549 ^ n46548 ;
  assign n46554 = n46502 ^ n46380 ;
  assign n46552 = n45910 ^ n45757 ;
  assign n46551 = n46013 ^ n45354 ;
  assign n46553 = n46552 ^ n46551 ;
  assign n46555 = n46554 ^ n46553 ;
  assign n46559 = n46498 ^ n46389 ;
  assign n46557 = n45908 ^ n45760 ;
  assign n46556 = n46002 ^ n45277 ;
  assign n46558 = n46557 ^ n46556 ;
  assign n46560 = n46559 ^ n46558 ;
  assign n46564 = n46495 ^ n46394 ;
  assign n46562 = n45905 ^ n45766 ;
  assign n46561 = n46000 ^ n44907 ;
  assign n46563 = n46562 ^ n46561 ;
  assign n46565 = n46564 ^ n46563 ;
  assign n46567 = n45732 ^ n44470 ;
  assign n46569 = n46568 ^ n46567 ;
  assign n46566 = n46489 ^ n46404 ;
  assign n46570 = n46569 ^ n46566 ;
  assign n46933 = n45722 ^ n44478 ;
  assign n46934 = n46933 ^ n46648 ;
  assign n46574 = n46479 ^ n46408 ;
  assign n46935 = n46934 ^ n46574 ;
  assign n46575 = n45708 ^ n44480 ;
  assign n46576 = n46575 ^ n46521 ;
  assign n46577 = n46576 ^ n46574 ;
  assign n46580 = n46474 ^ n46470 ;
  assign n46581 = n46580 ^ n46469 ;
  assign n46578 = n45691 ^ n44488 ;
  assign n46579 = n46578 ^ n46232 ;
  assign n46582 = n46581 ^ n46579 ;
  assign n46585 = n46466 ^ n46414 ;
  assign n46583 = n45550 ^ n44493 ;
  assign n46584 = n46583 ^ n45950 ;
  assign n46586 = n46585 ^ n46584 ;
  assign n46588 = n45302 ^ n44495 ;
  assign n46589 = n46588 ^ n45954 ;
  assign n46587 = n46463 ^ n46419 ;
  assign n46590 = n46589 ^ n46587 ;
  assign n46594 = n46461 ^ n46422 ;
  assign n46591 = n45306 ^ n44500 ;
  assign n46592 = n46591 ^ n45958 ;
  assign n46595 = n46594 ^ n46592 ;
  assign n46597 = n45312 ^ n44509 ;
  assign n46598 = n46597 ^ n45962 ;
  assign n46596 = n46457 ^ n46429 ;
  assign n46599 = n46598 ^ n46596 ;
  assign n46604 = n46454 ^ n46434 ;
  assign n46602 = n45311 ^ n44511 ;
  assign n46603 = n46602 ^ n45966 ;
  assign n46605 = n46604 ^ n46603 ;
  assign n46608 = n46451 ^ n46439 ;
  assign n46606 = n45524 ^ n44518 ;
  assign n46607 = n46606 ^ n45970 ;
  assign n46609 = n46608 ^ n46607 ;
  assign n46612 = n46448 ^ n46443 ;
  assign n46610 = n45516 ^ n44520 ;
  assign n46611 = n46610 ^ n45974 ;
  assign n46613 = n46612 ^ n46611 ;
  assign n46616 = n46447 ^ n46446 ;
  assign n46614 = n45506 ^ n44524 ;
  assign n46615 = n46614 ^ n45978 ;
  assign n46617 = n46616 ^ n46615 ;
  assign n46743 = n44553 ^ n44063 ;
  assign n46744 = n46743 ^ n45460 ;
  assign n46746 = n46745 ^ n46744 ;
  assign n46620 = n44802 ^ n44117 ;
  assign n46621 = n46620 ^ n45473 ;
  assign n46622 = n46621 ^ n46537 ;
  assign n46627 = n44771 ^ n44011 ;
  assign n46628 = n46627 ^ n45470 ;
  assign n46629 = n46628 ^ n46542 ;
  assign n46630 = n44774 ^ n43960 ;
  assign n46631 = n46630 ^ n45296 ;
  assign n46632 = n46631 ^ n46547 ;
  assign n46633 = n46035 ^ n43961 ;
  assign n46634 = n46633 ^ n44724 ;
  assign n46635 = n46634 ^ n46552 ;
  assign n46636 = n46029 ^ n45297 ;
  assign n46637 = n46636 ^ n44819 ;
  assign n46638 = n46637 ^ n46557 ;
  assign n46639 = n45371 ^ n44784 ;
  assign n46640 = n46639 ^ n46021 ;
  assign n46641 = n46640 ^ n46562 ;
  assign n46642 = n46013 ^ n44027 ;
  assign n46643 = n46642 ^ n45345 ;
  assign n46572 = n45902 ^ n45771 ;
  assign n46644 = n46643 ^ n46572 ;
  assign n46658 = n46657 ^ n46568 ;
  assign n46659 = ~n46647 & n46658 ;
  assign n46660 = n46659 ^ n46646 ;
  assign n46661 = n46660 ^ n46572 ;
  assign n46662 = ~n46644 & ~n46661 ;
  assign n46663 = n46662 ^ n46643 ;
  assign n46664 = n46663 ^ n46562 ;
  assign n46665 = n46641 & n46664 ;
  assign n46666 = n46665 ^ n46640 ;
  assign n46667 = n46666 ^ n46557 ;
  assign n46668 = ~n46638 & n46667 ;
  assign n46669 = n46668 ^ n46637 ;
  assign n46670 = n46669 ^ n46552 ;
  assign n46671 = n46635 & n46670 ;
  assign n46672 = n46671 ^ n46634 ;
  assign n46673 = n46672 ^ n46631 ;
  assign n46674 = n46632 & ~n46673 ;
  assign n46675 = n46674 ^ n46547 ;
  assign n46676 = n46675 ^ n46542 ;
  assign n46677 = n46629 & n46676 ;
  assign n46678 = n46677 ^ n46628 ;
  assign n46623 = n44833 ^ n44113 ;
  assign n46624 = n46623 ^ n45464 ;
  assign n46625 = n46624 ^ n46537 ;
  assign n46626 = n46625 ^ n46624 ;
  assign n46679 = n46678 ^ n46626 ;
  assign n46680 = ~n46622 & n46679 ;
  assign n46681 = n46680 ^ n46625 ;
  assign n46740 = n46624 ^ n45941 ;
  assign n46741 = ~n46681 & ~n46740 ;
  assign n46742 = n46741 ^ n46624 ;
  assign n46747 = n46746 ^ n46742 ;
  assign n46748 = n46747 ^ n43136 ;
  assign n46683 = n46678 ^ n46622 ;
  assign n46684 = n46683 ^ n43430 ;
  assign n46686 = n46672 ^ n46632 ;
  assign n46687 = n46686 ^ n43446 ;
  assign n46688 = n46669 ^ n46635 ;
  assign n46689 = n46688 ^ n43438 ;
  assign n46701 = n46660 ^ n46644 ;
  assign n46703 = n46701 ^ n43946 ;
  assign n46702 = n46701 ^ n46695 ;
  assign n46704 = n46703 ^ n46702 ;
  assign n46705 = n46700 & ~n46704 ;
  assign n46706 = n46705 ^ n46703 ;
  assign n46707 = n46663 ^ n46641 ;
  assign n46709 = n46707 ^ n43992 ;
  assign n46708 = n46707 ^ n46701 ;
  assign n46710 = n46709 ^ n46708 ;
  assign n46711 = n46706 & ~n46710 ;
  assign n46712 = n46711 ^ n46709 ;
  assign n46713 = n46666 ^ n46638 ;
  assign n46715 = n46713 ^ n44071 ;
  assign n46714 = n46713 ^ n46707 ;
  assign n46716 = n46715 ^ n46714 ;
  assign n46717 = n46712 & ~n46716 ;
  assign n46718 = n46717 ^ n46715 ;
  assign n46720 = n46688 ^ n44028 ;
  assign n46719 = n46713 ^ n46688 ;
  assign n46721 = n46720 ^ n46719 ;
  assign n46722 = n46718 & ~n46721 ;
  assign n46723 = n46722 ^ n46720 ;
  assign n46724 = ~n46689 & ~n46723 ;
  assign n46725 = n46724 ^ n43438 ;
  assign n46726 = n46725 ^ n46686 ;
  assign n46727 = n46687 & ~n46726 ;
  assign n46728 = n46727 ^ n43446 ;
  assign n46685 = n46675 ^ n46629 ;
  assign n46729 = n46728 ^ n46685 ;
  assign n46730 = n46728 ^ n43436 ;
  assign n46731 = ~n46729 & ~n46730 ;
  assign n46732 = n46731 ^ n43436 ;
  assign n46733 = n46732 ^ n46683 ;
  assign n46734 = ~n46684 & n46733 ;
  assign n46735 = n46734 ^ n43430 ;
  assign n46682 = n46681 ^ n45941 ;
  assign n46736 = n46735 ^ n46682 ;
  assign n46737 = n46735 ^ n43428 ;
  assign n46738 = n46736 & n46737 ;
  assign n46739 = n46738 ^ n43428 ;
  assign n46749 = n46748 ^ n46739 ;
  assign n46750 = n46732 ^ n46684 ;
  assign n46751 = n46725 ^ n46687 ;
  assign n46757 = ~n46755 & ~n46756 ;
  assign n46758 = n46706 ^ n43992 ;
  assign n46759 = n46757 & ~n46758 ;
  assign n46760 = n46712 ^ n44071 ;
  assign n46761 = ~n46759 & n46760 ;
  assign n46762 = n46718 ^ n44028 ;
  assign n46763 = n46761 & n46762 ;
  assign n46764 = n46723 ^ n43438 ;
  assign n46765 = ~n46763 & ~n46764 ;
  assign n46766 = n46751 & ~n46765 ;
  assign n46767 = n46685 ^ n43436 ;
  assign n46768 = n46767 ^ n46728 ;
  assign n46769 = ~n46766 & n46768 ;
  assign n46770 = n46750 & ~n46769 ;
  assign n46771 = n46682 ^ n43428 ;
  assign n46772 = n46771 ^ n46735 ;
  assign n46773 = n46770 & n46772 ;
  assign n46874 = ~n46749 & ~n46773 ;
  assign n46867 = n44783 ^ n36683 ;
  assign n46868 = n46867 ^ n41153 ;
  assign n46869 = n46868 ^ n3158 ;
  assign n46863 = n46862 ^ n46140 ;
  assign n46864 = n46863 ^ n43136 ;
  assign n46865 = n46864 ^ n45456 ;
  assign n46861 = n46744 ^ n44549 ;
  assign n46866 = n46865 ^ n46861 ;
  assign n46870 = n46869 ^ n46866 ;
  assign n46775 = n44755 ^ n36545 ;
  assign n46776 = n46775 ^ n41206 ;
  assign n46777 = n46776 ^ n35042 ;
  assign n46871 = n46870 ^ n46777 ;
  assign n46859 = n46747 ^ n46739 ;
  assign n46860 = ~n46748 & n46859 ;
  assign n46872 = n46871 ^ n46860 ;
  assign n46857 = n46744 ^ n46742 ;
  assign n46858 = n46746 & n46857 ;
  assign n46873 = n46872 ^ n46858 ;
  assign n46875 = n46874 ^ n46873 ;
  assign n46774 = n46773 ^ n46749 ;
  assign n46778 = n46777 ^ n46774 ;
  assign n46782 = n46772 ^ n46770 ;
  assign n46779 = n44731 ^ n36502 ;
  assign n46780 = n46779 ^ n41212 ;
  assign n46781 = n46780 ^ n35115 ;
  assign n46783 = n46782 ^ n46781 ;
  assign n46787 = n46769 ^ n46750 ;
  assign n46784 = n44723 ^ n36292 ;
  assign n46785 = n46784 ^ n40988 ;
  assign n46786 = n46785 ^ n35047 ;
  assign n46788 = n46787 ^ n46786 ;
  assign n46790 = n44715 ^ n36288 ;
  assign n46791 = n46790 ^ n40815 ;
  assign n46792 = n46791 ^ n35051 ;
  assign n46789 = n46768 ^ n46766 ;
  assign n46793 = n46792 ^ n46789 ;
  assign n46795 = n44643 ^ n36298 ;
  assign n46796 = n46795 ^ n40839 ;
  assign n46797 = n46796 ^ n35057 ;
  assign n46794 = n46765 ^ n46751 ;
  assign n46798 = n46797 ^ n46794 ;
  assign n46799 = n46764 ^ n46763 ;
  assign n1389 = n1388 ^ n1370 ;
  assign n1390 = n1389 ^ n1286 ;
  assign n1400 = n1399 ^ n1390 ;
  assign n46800 = n46799 ^ n1400 ;
  assign n46804 = n46762 ^ n46761 ;
  assign n46801 = n44665 ^ n36304 ;
  assign n46802 = n46801 ^ n1231 ;
  assign n46803 = n46802 ^ n1362 ;
  assign n46805 = n46804 ^ n46803 ;
  assign n46806 = n46760 ^ n46759 ;
  assign n1186 = n1176 ^ n1125 ;
  assign n1214 = n1213 ^ n1186 ;
  assign n1221 = n1220 ^ n1214 ;
  assign n46807 = n46806 ^ n1221 ;
  assign n46809 = n44672 ^ n1048 ;
  assign n46810 = n46809 ^ n40851 ;
  assign n46811 = n46810 ^ n1205 ;
  assign n46833 = n46811 ^ n1221 ;
  assign n46808 = n46758 ^ n46757 ;
  assign n46812 = n46811 ^ n46808 ;
  assign n46815 = n46814 ^ n1679 ;
  assign n46830 = ~n46815 & n46829 ;
  assign n46813 = n46808 ^ n1679 ;
  assign n46831 = n46830 ^ n46813 ;
  assign n46832 = n46812 & ~n46831 ;
  assign n46834 = n46833 ^ n46832 ;
  assign n46835 = ~n46807 & ~n46834 ;
  assign n46836 = n46835 ^ n46806 ;
  assign n46837 = n46836 ^ n46803 ;
  assign n46838 = n46805 & n46837 ;
  assign n46839 = n46838 ^ n46804 ;
  assign n46840 = n46839 ^ n1400 ;
  assign n46841 = ~n46800 & ~n46840 ;
  assign n46842 = n46841 ^ n46799 ;
  assign n46843 = n46842 ^ n46794 ;
  assign n46844 = ~n46798 & ~n46843 ;
  assign n46845 = n46844 ^ n46797 ;
  assign n46846 = n46845 ^ n46792 ;
  assign n46847 = n46793 & n46846 ;
  assign n46848 = n46847 ^ n46792 ;
  assign n46849 = n46848 ^ n46786 ;
  assign n46850 = ~n46788 & ~n46849 ;
  assign n46851 = n46850 ^ n46787 ;
  assign n46852 = n46851 ^ n46781 ;
  assign n46853 = n46783 & n46852 ;
  assign n46854 = n46853 ^ n46782 ;
  assign n46855 = n46854 ^ n46777 ;
  assign n46856 = ~n46778 & n46855 ;
  assign n46876 = n46875 ^ n46856 ;
  assign n46905 = n46876 ^ n46616 ;
  assign n46618 = n45503 ^ n44528 ;
  assign n46619 = n46618 ^ n45982 ;
  assign n46877 = n46876 ^ n46619 ;
  assign n46880 = n46854 ^ n46778 ;
  assign n46878 = n45319 ^ n44534 ;
  assign n46879 = n46878 ^ n45986 ;
  assign n46881 = n46880 ^ n46879 ;
  assign n46884 = n45321 ^ n44536 ;
  assign n46885 = n46884 ^ n45990 ;
  assign n46882 = n46851 ^ n46783 ;
  assign n46886 = n46885 ^ n46882 ;
  assign n46889 = n45331 ^ n44023 ;
  assign n46890 = n46889 ^ n45994 ;
  assign n46891 = n46845 ^ n46793 ;
  assign n46892 = ~n46890 & n46891 ;
  assign n46887 = n45327 ^ n44542 ;
  assign n46888 = n46887 ^ n46195 ;
  assign n46893 = n46892 ^ n46888 ;
  assign n46894 = n46848 ^ n46788 ;
  assign n46895 = n46894 ^ n46892 ;
  assign n46896 = n46893 & ~n46895 ;
  assign n46897 = n46896 ^ n46892 ;
  assign n46898 = n46897 ^ n46882 ;
  assign n46899 = n46886 & ~n46898 ;
  assign n46883 = n46882 ^ n46880 ;
  assign n46900 = n46899 ^ n46883 ;
  assign n46901 = n46881 & n46900 ;
  assign n46902 = n46901 ^ n46880 ;
  assign n46903 = n46902 ^ n46876 ;
  assign n46904 = ~n46877 & ~n46903 ;
  assign n46906 = n46905 ^ n46904 ;
  assign n46907 = ~n46617 & n46906 ;
  assign n46908 = n46907 ^ n46616 ;
  assign n46909 = n46908 ^ n46611 ;
  assign n46910 = ~n46613 & ~n46909 ;
  assign n46911 = n46910 ^ n46612 ;
  assign n46912 = n46911 ^ n46607 ;
  assign n46913 = n46609 & ~n46912 ;
  assign n46914 = n46913 ^ n46608 ;
  assign n46915 = n46914 ^ n46603 ;
  assign n46916 = ~n46605 & n46915 ;
  assign n46917 = n46916 ^ n46604 ;
  assign n46918 = n46917 ^ n46596 ;
  assign n46919 = ~n46599 & ~n46918 ;
  assign n46600 = n46596 ^ n46592 ;
  assign n46920 = n46919 ^ n46600 ;
  assign n46921 = ~n46595 & ~n46920 ;
  assign n46593 = n46592 ^ n46589 ;
  assign n46922 = n46921 ^ n46593 ;
  assign n46923 = n46590 & ~n46922 ;
  assign n46924 = n46923 ^ n46589 ;
  assign n46925 = n46924 ^ n46585 ;
  assign n46926 = n46586 & ~n46925 ;
  assign n46927 = n46926 ^ n46585 ;
  assign n46928 = n46927 ^ n46579 ;
  assign n46929 = ~n46582 & n46928 ;
  assign n46930 = n46929 ^ n46581 ;
  assign n46931 = n46930 ^ n46574 ;
  assign n46932 = n46577 & n46931 ;
  assign n46936 = n46935 ^ n46932 ;
  assign n46937 = n46486 ^ n46483 ;
  assign n46938 = n46937 ^ n46934 ;
  assign n46939 = n46936 & n46938 ;
  assign n46940 = n46939 ^ n46934 ;
  assign n46571 = n45930 ^ n44468 ;
  assign n46573 = n46572 ^ n46571 ;
  assign n46941 = n46940 ^ n46573 ;
  assign n46942 = n46941 ^ n46566 ;
  assign n46943 = n46942 ^ n46573 ;
  assign n46944 = ~n46570 & n46943 ;
  assign n46945 = n46944 ^ n46941 ;
  assign n46947 = n46492 ^ n46399 ;
  assign n46948 = n46947 ^ n46564 ;
  assign n46946 = n46573 ^ n46564 ;
  assign n46949 = n46948 ^ n46946 ;
  assign n46950 = n46945 & ~n46949 ;
  assign n46951 = n46950 ^ n46946 ;
  assign n46952 = ~n46565 & n46951 ;
  assign n46953 = n46952 ^ n46564 ;
  assign n46954 = n46953 ^ n46558 ;
  assign n46955 = ~n46560 & n46954 ;
  assign n46956 = n46955 ^ n46559 ;
  assign n46957 = n46956 ^ n46553 ;
  assign n46958 = ~n46555 & n46957 ;
  assign n46959 = n46958 ^ n46554 ;
  assign n46960 = n46959 ^ n46548 ;
  assign n46961 = n46550 & n46960 ;
  assign n46962 = n46961 ^ n46549 ;
  assign n46963 = n46962 ^ n46543 ;
  assign n46964 = n46545 & ~n46963 ;
  assign n46965 = n46964 ^ n46544 ;
  assign n46966 = n46965 ^ n46538 ;
  assign n46967 = ~n46540 & n46966 ;
  assign n46968 = n46967 ^ n46539 ;
  assign n46969 = n46968 ^ n45942 ;
  assign n46970 = ~n46535 & n46969 ;
  assign n46971 = n46970 ^ n46534 ;
  assign n47108 = n46973 ^ n46971 ;
  assign n47109 = ~n46975 & n47108 ;
  assign n47110 = n47109 ^ n46974 ;
  assign n47115 = n47114 ^ n47110 ;
  assign n47389 = n47115 ^ n43960 ;
  assign n46976 = n46975 ^ n46971 ;
  assign n46977 = n46976 ^ n43961 ;
  assign n46978 = n46968 ^ n46535 ;
  assign n46979 = n46978 ^ n44819 ;
  assign n47092 = n46962 ^ n46545 ;
  assign n46981 = n46956 ^ n46555 ;
  assign n46982 = n46981 ^ n44475 ;
  assign n46983 = n46953 ^ n46560 ;
  assign n46984 = n46983 ^ n44481 ;
  assign n46985 = n46951 ^ n46563 ;
  assign n46986 = n46985 ^ n44485 ;
  assign n46987 = n46947 ^ n46945 ;
  assign n46988 = n46987 ^ n44490 ;
  assign n46990 = n46937 ^ n46936 ;
  assign n46991 = n46990 ^ n44502 ;
  assign n46992 = n46930 ^ n46577 ;
  assign n46993 = n46992 ^ n44506 ;
  assign n47058 = n46927 ^ n46582 ;
  assign n46995 = n46922 ^ n46587 ;
  assign n46996 = n46995 ^ n44308 ;
  assign n46998 = n46917 ^ n46599 ;
  assign n46999 = n46998 ^ n44175 ;
  assign n47038 = n46914 ^ n46605 ;
  assign n47000 = n46908 ^ n46613 ;
  assign n47001 = n47000 ^ n44043 ;
  assign n47021 = n46902 ^ n46877 ;
  assign n47003 = n46900 ^ n46879 ;
  assign n47004 = n47003 ^ n44152 ;
  assign n47012 = n46897 ^ n46886 ;
  assign n47005 = n46891 ^ n46890 ;
  assign n47006 = ~n44058 & ~n47005 ;
  assign n47007 = n47006 ^ n44134 ;
  assign n47008 = n46894 ^ n46893 ;
  assign n47009 = n47008 ^ n47006 ;
  assign n47010 = n47007 & n47009 ;
  assign n47011 = n47010 ^ n44134 ;
  assign n47013 = n47012 ^ n47011 ;
  assign n47014 = n47003 ^ n44144 ;
  assign n47015 = n47014 ^ n47003 ;
  assign n47016 = n47015 ^ n47011 ;
  assign n47017 = ~n47013 & ~n47016 ;
  assign n47018 = n47017 ^ n47014 ;
  assign n47019 = ~n47004 & ~n47018 ;
  assign n47020 = n47019 ^ n44152 ;
  assign n47022 = n47021 ^ n47020 ;
  assign n47023 = n47020 ^ n44049 ;
  assign n47024 = ~n47022 & ~n47023 ;
  assign n47025 = n47024 ^ n44049 ;
  assign n47002 = n46906 ^ n46615 ;
  assign n47026 = n47025 ^ n47002 ;
  assign n47027 = n47025 ^ n44047 ;
  assign n47028 = ~n47026 & ~n47027 ;
  assign n47029 = n47028 ^ n44047 ;
  assign n47030 = n47029 ^ n47000 ;
  assign n47031 = ~n47001 & n47030 ;
  assign n47032 = n47031 ^ n44043 ;
  assign n47033 = n47032 ^ n44034 ;
  assign n47034 = n46911 ^ n46609 ;
  assign n47035 = n47034 ^ n47032 ;
  assign n47036 = ~n47033 & n47035 ;
  assign n47037 = n47036 ^ n44034 ;
  assign n47039 = n47038 ^ n47037 ;
  assign n47040 = n46998 ^ n44038 ;
  assign n47041 = n47040 ^ n46998 ;
  assign n47042 = n47041 ^ n47037 ;
  assign n47043 = n47039 & n47042 ;
  assign n47044 = n47043 ^ n47040 ;
  assign n47045 = ~n46999 & n47044 ;
  assign n47046 = n47045 ^ n44175 ;
  assign n46997 = n46920 ^ n46594 ;
  assign n47047 = n47046 ^ n46997 ;
  assign n47048 = n47046 ^ n44261 ;
  assign n47049 = ~n47047 & ~n47048 ;
  assign n47050 = n47049 ^ n44261 ;
  assign n47051 = n47050 ^ n46995 ;
  assign n47052 = ~n46996 & n47051 ;
  assign n47053 = n47052 ^ n44308 ;
  assign n46994 = n46924 ^ n46586 ;
  assign n47054 = n47053 ^ n46994 ;
  assign n47055 = n47053 ^ n44452 ;
  assign n47056 = ~n47054 & n47055 ;
  assign n47057 = n47056 ^ n44452 ;
  assign n47059 = n47058 ^ n47057 ;
  assign n47060 = n46992 ^ n44512 ;
  assign n47061 = n47060 ^ n46992 ;
  assign n47062 = n47061 ^ n47057 ;
  assign n47063 = ~n47059 & ~n47062 ;
  assign n47064 = n47063 ^ n47060 ;
  assign n47065 = n46993 & ~n47064 ;
  assign n47066 = n47065 ^ n44506 ;
  assign n47067 = n47066 ^ n46990 ;
  assign n47068 = ~n46991 & ~n47067 ;
  assign n47069 = n47068 ^ n44502 ;
  assign n46989 = n46940 ^ n46570 ;
  assign n47070 = n47069 ^ n46989 ;
  assign n47071 = n46987 ^ n44496 ;
  assign n47072 = n47071 ^ n46989 ;
  assign n47073 = n47072 ^ n46987 ;
  assign n47074 = n47070 & ~n47073 ;
  assign n47075 = n47074 ^ n47071 ;
  assign n47076 = n46988 & ~n47075 ;
  assign n47077 = n47076 ^ n44490 ;
  assign n47078 = n47077 ^ n46985 ;
  assign n47079 = ~n46986 & ~n47078 ;
  assign n47080 = n47079 ^ n44485 ;
  assign n47081 = n47080 ^ n46983 ;
  assign n47082 = ~n46984 & n47081 ;
  assign n47083 = n47082 ^ n44481 ;
  assign n47084 = n47083 ^ n46981 ;
  assign n47085 = n46982 & n47084 ;
  assign n47086 = n47085 ^ n44475 ;
  assign n47087 = n47086 ^ n44471 ;
  assign n47088 = n46959 ^ n46550 ;
  assign n47089 = n47088 ^ n47086 ;
  assign n47090 = n47087 & n47089 ;
  assign n47091 = n47090 ^ n44471 ;
  assign n47093 = n47092 ^ n47091 ;
  assign n47094 = n47092 ^ n44027 ;
  assign n47095 = ~n47093 & n47094 ;
  assign n47096 = n47095 ^ n44027 ;
  assign n46980 = n46965 ^ n46540 ;
  assign n47097 = n47096 ^ n46980 ;
  assign n47098 = n47096 ^ n44784 ;
  assign n47099 = n47097 & n47098 ;
  assign n47100 = n47099 ^ n44784 ;
  assign n47101 = n47100 ^ n46978 ;
  assign n47102 = ~n46979 & n47101 ;
  assign n47103 = n47102 ^ n44819 ;
  assign n47104 = n47103 ^ n46976 ;
  assign n47105 = ~n46977 & n47104 ;
  assign n47106 = n47105 ^ n43961 ;
  assign n47390 = n47115 ^ n47106 ;
  assign n47391 = n47389 & n47390 ;
  assign n47392 = n47391 ^ n43960 ;
  assign n47386 = n46831 ^ n46811 ;
  assign n47379 = n45464 ^ n44771 ;
  assign n47380 = n47379 ^ n46171 ;
  assign n47381 = n47380 ^ n47113 ;
  assign n47382 = n47381 ^ n47380 ;
  assign n47383 = n47382 ^ n47110 ;
  assign n47384 = ~n47114 & ~n47383 ;
  assign n47385 = n47384 ^ n47381 ;
  assign n47387 = n47386 ^ n47385 ;
  assign n47388 = n47387 ^ n44011 ;
  assign n47393 = n47392 ^ n47388 ;
  assign n47107 = n47106 ^ n43960 ;
  assign n47116 = n47115 ^ n47107 ;
  assign n47117 = n47098 ^ n46980 ;
  assign n47118 = n47094 ^ n47091 ;
  assign n47119 = n47075 ^ n44490 ;
  assign n47120 = n47069 ^ n44496 ;
  assign n47121 = n47120 ^ n46989 ;
  assign n47122 = n47066 ^ n46991 ;
  assign n47123 = n47064 ^ n44506 ;
  assign n47124 = n47008 ^ n47007 ;
  assign n47125 = n47012 ^ n44144 ;
  assign n47126 = n47125 ^ n47011 ;
  assign n47127 = n47124 & n47126 ;
  assign n47128 = n47018 ^ n44152 ;
  assign n47129 = ~n47127 & n47128 ;
  assign n47130 = n47022 ^ n44049 ;
  assign n47131 = ~n47129 & n47130 ;
  assign n47132 = n47002 ^ n44047 ;
  assign n47133 = n47132 ^ n47025 ;
  assign n47134 = ~n47131 & n47133 ;
  assign n47135 = n47029 ^ n47001 ;
  assign n47136 = ~n47134 & n47135 ;
  assign n47137 = n47034 ^ n47033 ;
  assign n47138 = n47136 & ~n47137 ;
  assign n47139 = n47038 ^ n44038 ;
  assign n47140 = n47139 ^ n47037 ;
  assign n47141 = n47138 & ~n47140 ;
  assign n47142 = n47044 ^ n44175 ;
  assign n47143 = ~n47141 & n47142 ;
  assign n47144 = n46997 ^ n44261 ;
  assign n47145 = n47144 ^ n47046 ;
  assign n47146 = n47143 & n47145 ;
  assign n47147 = n47050 ^ n46996 ;
  assign n47148 = n47146 & ~n47147 ;
  assign n47149 = n46994 ^ n44452 ;
  assign n47150 = n47149 ^ n47053 ;
  assign n47151 = n47148 & n47150 ;
  assign n47152 = n47057 ^ n44512 ;
  assign n47153 = n47152 ^ n47058 ;
  assign n47154 = n47151 & ~n47153 ;
  assign n47155 = n47123 & ~n47154 ;
  assign n47156 = ~n47122 & n47155 ;
  assign n47157 = ~n47121 & ~n47156 ;
  assign n47158 = ~n47119 & ~n47157 ;
  assign n47159 = n47077 ^ n46986 ;
  assign n47160 = ~n47158 & ~n47159 ;
  assign n47161 = n47080 ^ n46984 ;
  assign n47162 = n47160 & n47161 ;
  assign n47163 = n47083 ^ n46982 ;
  assign n47164 = n47162 & ~n47163 ;
  assign n47165 = n47088 ^ n47087 ;
  assign n47166 = ~n47164 & n47165 ;
  assign n47167 = ~n47118 & n47166 ;
  assign n47168 = ~n47117 & ~n47167 ;
  assign n47169 = n47100 ^ n46979 ;
  assign n47170 = n47168 & ~n47169 ;
  assign n47171 = n47103 ^ n46977 ;
  assign n47172 = ~n47170 & n47171 ;
  assign n47378 = n47116 & ~n47172 ;
  assign n47394 = n47393 ^ n47378 ;
  assign n47398 = n47397 ^ n47394 ;
  assign n47173 = n47172 ^ n47116 ;
  assign n44024 = n37055 ^ n1447 ;
  assign n44025 = n44024 ^ n41625 ;
  assign n44026 = n44025 ^ n2850 ;
  assign n47174 = n47173 ^ n44026 ;
  assign n47178 = n47171 ^ n47170 ;
  assign n47175 = n2798 ^ n1429 ;
  assign n47176 = n47175 ^ n41630 ;
  assign n47177 = n47176 ^ n35529 ;
  assign n47179 = n47178 ^ n47177 ;
  assign n47184 = n47169 ^ n47168 ;
  assign n47180 = n45090 ^ n1322 ;
  assign n47181 = n47180 ^ n1747 ;
  assign n47182 = n47181 ^ n35534 ;
  assign n47185 = n47184 ^ n47182 ;
  assign n47186 = n47167 ^ n47117 ;
  assign n1723 = n1716 ^ n1307 ;
  assign n1733 = n1732 ^ n1723 ;
  assign n1740 = n1739 ^ n1733 ;
  assign n47187 = n47186 ^ n1740 ;
  assign n47191 = n47166 ^ n47118 ;
  assign n47188 = n45096 ^ n1699 ;
  assign n47189 = n47188 ^ n41640 ;
  assign n47190 = n47189 ^ n1730 ;
  assign n47192 = n47191 ^ n47190 ;
  assign n47196 = n47165 ^ n47164 ;
  assign n47193 = n45101 ^ n1690 ;
  assign n47194 = n47193 ^ n41645 ;
  assign n47195 = n47194 ^ n929 ;
  assign n47197 = n47196 ^ n47195 ;
  assign n47199 = n45106 ^ n37071 ;
  assign n47200 = n47199 ^ n827 ;
  assign n47201 = n47200 ^ n35545 ;
  assign n47360 = n47201 ^ n47195 ;
  assign n47198 = n47163 ^ n47162 ;
  assign n47202 = n47201 ^ n47198 ;
  assign n47203 = n45111 ^ n37067 ;
  assign n47204 = n47203 ^ n41652 ;
  assign n47205 = n47204 ^ n819 ;
  assign n47357 = n47205 ^ n47198 ;
  assign n47206 = n47161 ^ n47160 ;
  assign n47207 = n47206 ^ n47205 ;
  assign n47211 = n47159 ^ n47158 ;
  assign n47208 = n45116 ^ n722 ;
  assign n47209 = n47208 ^ n41657 ;
  assign n47210 = n47209 ^ n35551 ;
  assign n47212 = n47211 ^ n47210 ;
  assign n47214 = n45121 ^ n37078 ;
  assign n47215 = n47214 ^ n41662 ;
  assign n47216 = n47215 ^ n1574 ;
  assign n47213 = n47157 ^ n47119 ;
  assign n47217 = n47216 ^ n47213 ;
  assign n47223 = n47156 ^ n47121 ;
  assign n47220 = n45126 ^ n37083 ;
  assign n47221 = n47220 ^ n41667 ;
  assign n47222 = n47221 ^ n35563 ;
  assign n47224 = n47223 ^ n47222 ;
  assign n47226 = n45131 ^ n37089 ;
  assign n47227 = n47226 ^ n41674 ;
  assign n47228 = n47227 ^ n35558 ;
  assign n47346 = n47228 ^ n47223 ;
  assign n47225 = n47155 ^ n47122 ;
  assign n47229 = n47228 ^ n47225 ;
  assign n47231 = n45137 ^ n37094 ;
  assign n47232 = n47231 ^ n41679 ;
  assign n47233 = n47232 ^ n35568 ;
  assign n47230 = n47154 ^ n47123 ;
  assign n47234 = n47233 ^ n47230 ;
  assign n47236 = n45142 ^ n37098 ;
  assign n47237 = n47236 ^ n41684 ;
  assign n47238 = n47237 ^ n35657 ;
  assign n47235 = n47153 ^ n47151 ;
  assign n47239 = n47238 ^ n47235 ;
  assign n47241 = n45146 ^ n37105 ;
  assign n47242 = n47241 ^ n41689 ;
  assign n47243 = n47242 ^ n35573 ;
  assign n47337 = n47243 ^ n47238 ;
  assign n47240 = n47150 ^ n47148 ;
  assign n47244 = n47243 ^ n47240 ;
  assign n47248 = n47147 ^ n47146 ;
  assign n47245 = n45151 ^ n37109 ;
  assign n47246 = n47245 ^ n2396 ;
  assign n47247 = n47246 ^ n35578 ;
  assign n47249 = n47248 ^ n47247 ;
  assign n47251 = n45156 ^ n37115 ;
  assign n47252 = n47251 ^ n41695 ;
  assign n47253 = n47252 ^ n2391 ;
  assign n47331 = n47253 ^ n47247 ;
  assign n47250 = n47145 ^ n47143 ;
  assign n47254 = n47253 ^ n47250 ;
  assign n47256 = n47142 ^ n47141 ;
  assign n2235 = n2234 ^ n2201 ;
  assign n2269 = n2268 ^ n2235 ;
  assign n2279 = n2278 ^ n2269 ;
  assign n47257 = n47256 ^ n2279 ;
  assign n47259 = n45165 ^ n37122 ;
  assign n47260 = n47259 ^ n41752 ;
  assign n47261 = n47260 ^ n2260 ;
  assign n47258 = n47140 ^ n47138 ;
  assign n47262 = n47261 ^ n47258 ;
  assign n47266 = n47137 ^ n47136 ;
  assign n47263 = n45169 ^ n2124 ;
  assign n47264 = n47263 ^ n41702 ;
  assign n47265 = n47264 ^ n35590 ;
  assign n47267 = n47266 ^ n47265 ;
  assign n47269 = n45177 ^ n37128 ;
  assign n47270 = n47269 ^ n41708 ;
  assign n47271 = n47270 ^ n35594 ;
  assign n47268 = n47135 ^ n47134 ;
  assign n47272 = n47271 ^ n47268 ;
  assign n47274 = n45181 ^ n37132 ;
  assign n47275 = n47274 ^ n41738 ;
  assign n47276 = n47275 ^ n35624 ;
  assign n47317 = n47276 ^ n47271 ;
  assign n47273 = n47133 ^ n47131 ;
  assign n47277 = n47276 ^ n47273 ;
  assign n47279 = n45186 ^ n37137 ;
  assign n47280 = n47279 ^ n41712 ;
  assign n47281 = n47280 ^ n35616 ;
  assign n47314 = n47281 ^ n47276 ;
  assign n47278 = n47130 ^ n47129 ;
  assign n47282 = n47281 ^ n47278 ;
  assign n47286 = n47128 ^ n47127 ;
  assign n47311 = n47286 ^ n47278 ;
  assign n47283 = n45192 ^ n36535 ;
  assign n47284 = n47283 ^ n41717 ;
  assign n47285 = n47284 ^ n35612 ;
  assign n47287 = n47286 ^ n47285 ;
  assign n47291 = n47126 ^ n47124 ;
  assign n47308 = n47291 ^ n47286 ;
  assign n47288 = n45196 ^ n36491 ;
  assign n47289 = n47288 ^ n41721 ;
  assign n47290 = n47289 ^ n35599 ;
  assign n47292 = n47291 ^ n47290 ;
  assign n47298 = n40998 ^ n35828 ;
  assign n47299 = n47298 ^ n45200 ;
  assign n47300 = n47299 ^ n35604 ;
  assign n47293 = n47005 ^ n44058 ;
  assign n47294 = n45412 ^ n3173 ;
  assign n47295 = n47294 ^ n41838 ;
  assign n47296 = n47295 ^ n35958 ;
  assign n47297 = n47293 & n47296 ;
  assign n47301 = n47300 ^ n47297 ;
  assign n47304 = n47297 ^ n47124 ;
  assign n47305 = ~n47301 & n47304 ;
  assign n47302 = n47290 ^ n47124 ;
  assign n47306 = n47305 ^ n47302 ;
  assign n47307 = ~n47292 & ~n47306 ;
  assign n47309 = n47308 ^ n47307 ;
  assign n47310 = ~n47287 & n47309 ;
  assign n47312 = n47311 ^ n47310 ;
  assign n47313 = n47282 & n47312 ;
  assign n47315 = n47314 ^ n47313 ;
  assign n47316 = ~n47277 & n47315 ;
  assign n47318 = n47317 ^ n47316 ;
  assign n47319 = n47272 & n47318 ;
  assign n47320 = n47319 ^ n47271 ;
  assign n47321 = n47320 ^ n47265 ;
  assign n47322 = n47267 & ~n47321 ;
  assign n47323 = n47322 ^ n47266 ;
  assign n47324 = n47323 ^ n47258 ;
  assign n47325 = n47262 & ~n47324 ;
  assign n47326 = n47325 ^ n47261 ;
  assign n47327 = n47326 ^ n2279 ;
  assign n47328 = ~n47257 & n47327 ;
  assign n47255 = n47253 ^ n2279 ;
  assign n47329 = n47328 ^ n47255 ;
  assign n47330 = n47254 & n47329 ;
  assign n47332 = n47331 ^ n47330 ;
  assign n47333 = ~n47249 & ~n47332 ;
  assign n47334 = n47333 ^ n47248 ;
  assign n47335 = n47334 ^ n47240 ;
  assign n47336 = n47244 & n47335 ;
  assign n47338 = n47337 ^ n47336 ;
  assign n47339 = ~n47239 & n47338 ;
  assign n47340 = n47339 ^ n47238 ;
  assign n47341 = n47340 ^ n47230 ;
  assign n47342 = n47234 & ~n47341 ;
  assign n47343 = n47342 ^ n47233 ;
  assign n47344 = n47343 ^ n47228 ;
  assign n47345 = n47229 & n47344 ;
  assign n47347 = n47346 ^ n47345 ;
  assign n47348 = n47224 & n47347 ;
  assign n47349 = n47348 ^ n47223 ;
  assign n47350 = n47349 ^ n47216 ;
  assign n47351 = ~n47217 & n47350 ;
  assign n47218 = n47216 ^ n47211 ;
  assign n47352 = n47351 ^ n47218 ;
  assign n47353 = n47212 & n47352 ;
  assign n47354 = n47353 ^ n47211 ;
  assign n47355 = n47354 ^ n47205 ;
  assign n47356 = n47207 & n47355 ;
  assign n47358 = n47357 ^ n47356 ;
  assign n47359 = ~n47202 & n47358 ;
  assign n47361 = n47360 ^ n47359 ;
  assign n47362 = n47197 & ~n47361 ;
  assign n47363 = n47362 ^ n47196 ;
  assign n47364 = n47363 ^ n47190 ;
  assign n47365 = n47192 & ~n47364 ;
  assign n47366 = n47365 ^ n47191 ;
  assign n47367 = n47366 ^ n1740 ;
  assign n47368 = n47187 & ~n47367 ;
  assign n47369 = n47368 ^ n47186 ;
  assign n47370 = n47369 ^ n47182 ;
  assign n47371 = ~n47185 & n47370 ;
  assign n47183 = n47182 ^ n47177 ;
  assign n47372 = n47371 ^ n47183 ;
  assign n47373 = n47179 & ~n47372 ;
  assign n47374 = n47373 ^ n47178 ;
  assign n47375 = n47374 ^ n44026 ;
  assign n47376 = ~n47174 & ~n47375 ;
  assign n47377 = n47376 ^ n47173 ;
  assign n47399 = n47398 ^ n47377 ;
  assign n47400 = n45990 ^ n45331 ;
  assign n47401 = n47400 ^ n46616 ;
  assign n47431 = n47399 & n47401 ;
  assign n47429 = n45986 ^ n45327 ;
  assign n47430 = n47429 ^ n46612 ;
  assign n47432 = n47431 ^ n47430 ;
  assign n47425 = ~n47378 & ~n47393 ;
  assign n47420 = n46834 ^ n46806 ;
  assign n47418 = n45460 ^ n44802 ;
  assign n47419 = n47418 ^ n46177 ;
  assign n47421 = n47420 ^ n47419 ;
  assign n47415 = n47386 ^ n47380 ;
  assign n47416 = ~n47385 & ~n47415 ;
  assign n47417 = n47416 ^ n47386 ;
  assign n47422 = n47421 ^ n47417 ;
  assign n47423 = n47422 ^ n44117 ;
  assign n47411 = n47392 ^ n47387 ;
  assign n47412 = n47392 ^ n44011 ;
  assign n47413 = n47411 & n47412 ;
  assign n47414 = n47413 ^ n44011 ;
  assign n47424 = n47423 ^ n47414 ;
  assign n47426 = n47425 ^ n47424 ;
  assign n47408 = n45440 ^ n37050 ;
  assign n47409 = n47408 ^ n41618 ;
  assign n47410 = n47409 ^ n35731 ;
  assign n47427 = n47426 ^ n47410 ;
  assign n47405 = n47394 ^ n47377 ;
  assign n47406 = ~n47398 & ~n47405 ;
  assign n47407 = n47406 ^ n47397 ;
  assign n47428 = n47427 ^ n47407 ;
  assign n47433 = n47432 ^ n47428 ;
  assign n47402 = n47401 ^ n47399 ;
  assign n47403 = n44023 & n47402 ;
  assign n47435 = n47433 ^ n47403 ;
  assign n47463 = n45982 ^ n45321 ;
  assign n47464 = n47463 ^ n46608 ;
  assign n47460 = n47430 ^ n47428 ;
  assign n47461 = n47432 & ~n47460 ;
  assign n47454 = n45434 ^ n37392 ;
  assign n47455 = n47454 ^ n41614 ;
  assign n47456 = n47455 ^ n35773 ;
  assign n47452 = n47424 & ~n47425 ;
  assign n47448 = n47422 ^ n47414 ;
  assign n47449 = ~n47423 & ~n47448 ;
  assign n47450 = n47449 ^ n44117 ;
  assign n47443 = n45456 ^ n44833 ;
  assign n47444 = n47443 ^ n46167 ;
  assign n47442 = n46836 ^ n46805 ;
  assign n47445 = n47444 ^ n47442 ;
  assign n47439 = n47420 ^ n47417 ;
  assign n47440 = ~n47421 & ~n47439 ;
  assign n47441 = n47440 ^ n47420 ;
  assign n47446 = n47445 ^ n47441 ;
  assign n47447 = n47446 ^ n44113 ;
  assign n47451 = n47450 ^ n47447 ;
  assign n47453 = n47452 ^ n47451 ;
  assign n47457 = n47456 ^ n47453 ;
  assign n47436 = n47410 ^ n47407 ;
  assign n47437 = ~n47427 & ~n47436 ;
  assign n47438 = n47437 ^ n47426 ;
  assign n47458 = n47457 ^ n47438 ;
  assign n47459 = n47458 ^ n47430 ;
  assign n47462 = n47461 ^ n47459 ;
  assign n47465 = n47464 ^ n47462 ;
  assign n47466 = n47465 ^ n44542 ;
  assign n47467 = n47466 ^ n47465 ;
  assign n47468 = n47467 ^ n47403 ;
  assign n47469 = n47435 & n47468 ;
  assign n47470 = n47469 ^ n47466 ;
  assign n47471 = n47470 ^ n44536 ;
  assign n47404 = n47403 ^ n44542 ;
  assign n47434 = n47433 ^ n47404 ;
  assign n47651 = n47471 ^ n47434 ;
  assign n47638 = n45852 ^ n37247 ;
  assign n47639 = n47638 ^ n2732 ;
  assign n47640 = n47639 ^ n3230 ;
  assign n47641 = n47640 ^ n47434 ;
  assign n47642 = n46154 ^ n38201 ;
  assign n47643 = n47642 ^ n42610 ;
  assign n47644 = n47643 ^ n2724 ;
  assign n47645 = n47402 ^ n44023 ;
  assign n47646 = n47644 & n47645 ;
  assign n47647 = n47646 ^ n47640 ;
  assign n47648 = n47641 & ~n47647 ;
  assign n47649 = n47648 ^ n47434 ;
  assign n47652 = n47651 ^ n47649 ;
  assign n48341 = n47655 ^ n47652 ;
  assign n47771 = n47320 ^ n47267 ;
  assign n48339 = n47771 ^ n45962 ;
  assign n48340 = n48339 ^ n46574 ;
  assign n48342 = n48341 ^ n48340 ;
  assign n48274 = n47646 ^ n47641 ;
  assign n48272 = n46581 ^ n45966 ;
  assign n47773 = n47318 ^ n47268 ;
  assign n48273 = n48272 ^ n47773 ;
  assign n48275 = n48274 ^ n48273 ;
  assign n48259 = n47645 ^ n47644 ;
  assign n47777 = n47315 ^ n47273 ;
  assign n48257 = n47777 ^ n46585 ;
  assign n48258 = n48257 ^ n45970 ;
  assign n48260 = n48259 ^ n48258 ;
  assign n47937 = n46163 ^ n45460 ;
  assign n47938 = n47937 ^ n46894 ;
  assign n47831 = n46891 ^ n46167 ;
  assign n47832 = n47831 ^ n45464 ;
  assign n47830 = n47363 ^ n47192 ;
  assign n47833 = n47832 ^ n47830 ;
  assign n47931 = n47366 ^ n47187 ;
  assign n47932 = n47931 ^ n47830 ;
  assign n47933 = n47932 ^ n47931 ;
  assign n47707 = n46177 ^ n45473 ;
  assign n47528 = n46842 ^ n46798 ;
  assign n47708 = n47707 ^ n47528 ;
  assign n47706 = n47361 ^ n47196 ;
  assign n47709 = n47708 ^ n47706 ;
  assign n47486 = n46839 ^ n46800 ;
  assign n47711 = n47486 ^ n45470 ;
  assign n47712 = n47711 ^ n46171 ;
  assign n47710 = n47358 ^ n47201 ;
  assign n47713 = n47712 ^ n47710 ;
  assign n47716 = n47354 ^ n47207 ;
  assign n47714 = n47442 ^ n45296 ;
  assign n47715 = n47714 ^ n46862 ;
  assign n47717 = n47716 ^ n47715 ;
  assign n47719 = n47420 ^ n46745 ;
  assign n47720 = n47719 ^ n46035 ;
  assign n47718 = n47352 ^ n47210 ;
  assign n47721 = n47720 ^ n47718 ;
  assign n47724 = n47349 ^ n47217 ;
  assign n47722 = n46029 ^ n45941 ;
  assign n47723 = n47722 ^ n47386 ;
  assign n47725 = n47724 ^ n47723 ;
  assign n47730 = n47347 ^ n47222 ;
  assign n47728 = n47113 ^ n46537 ;
  assign n47729 = n47728 ^ n46021 ;
  assign n47731 = n47730 ^ n47729 ;
  assign n47734 = n47343 ^ n47229 ;
  assign n47732 = n46974 ^ n46542 ;
  assign n47733 = n47732 ^ n46013 ;
  assign n47735 = n47734 ^ n47733 ;
  assign n47739 = n47340 ^ n47234 ;
  assign n47736 = n46547 ^ n46002 ;
  assign n47737 = n47736 ^ n46534 ;
  assign n47740 = n47739 ^ n47737 ;
  assign n47743 = n47338 ^ n47235 ;
  assign n47741 = n46539 ^ n46000 ;
  assign n47742 = n47741 ^ n46552 ;
  assign n47744 = n47743 ^ n47742 ;
  assign n47749 = n47334 ^ n47244 ;
  assign n47747 = n46544 ^ n45930 ;
  assign n47748 = n47747 ^ n46557 ;
  assign n47750 = n47749 ^ n47748 ;
  assign n47753 = n47332 ^ n47248 ;
  assign n47751 = n46549 ^ n45732 ;
  assign n47752 = n47751 ^ n46562 ;
  assign n47754 = n47753 ^ n47752 ;
  assign n47757 = n47329 ^ n47250 ;
  assign n47755 = n46554 ^ n45722 ;
  assign n47756 = n47755 ^ n46572 ;
  assign n47758 = n47757 ^ n47756 ;
  assign n47760 = n46568 ^ n45708 ;
  assign n47761 = n47760 ^ n46559 ;
  assign n47696 = n47326 ^ n47257 ;
  assign n47762 = n47761 ^ n47696 ;
  assign n47765 = n47323 ^ n47262 ;
  assign n47763 = n46648 ^ n45691 ;
  assign n47764 = n47763 ^ n46564 ;
  assign n47766 = n47765 ^ n47764 ;
  assign n47769 = n46947 ^ n46521 ;
  assign n47770 = n47769 ^ n45550 ;
  assign n47772 = n47771 ^ n47770 ;
  assign n47774 = n46566 ^ n46232 ;
  assign n47775 = n47774 ^ n45302 ;
  assign n47776 = n47775 ^ n47773 ;
  assign n47786 = n47777 ^ n47775 ;
  assign n47778 = n46937 ^ n45306 ;
  assign n47779 = n47778 ^ n45950 ;
  assign n47780 = n47779 ^ n47777 ;
  assign n47685 = n47312 ^ n47281 ;
  assign n47596 = n47309 ^ n47285 ;
  assign n47686 = n47685 ^ n47596 ;
  assign n47578 = n47306 ^ n47291 ;
  assign n47597 = n47596 ^ n47578 ;
  assign n47567 = n47300 ^ n47124 ;
  assign n47568 = n47567 ^ n47297 ;
  assign n47565 = n46587 ^ n45516 ;
  assign n47566 = n47565 ^ n45966 ;
  assign n47569 = n47568 ^ n47566 ;
  assign n47579 = n47578 ^ n47568 ;
  assign n47580 = n47579 ^ n47578 ;
  assign n47549 = n47296 ^ n47293 ;
  assign n47478 = n47451 & n47452 ;
  assign n47487 = n45339 ^ n44553 ;
  assign n47488 = n47487 ^ n46163 ;
  assign n47489 = n47488 ^ n47486 ;
  assign n47483 = n47442 ^ n47441 ;
  assign n47484 = ~n47445 & n47483 ;
  assign n47485 = n47484 ^ n47442 ;
  assign n47490 = n47489 ^ n47485 ;
  assign n47491 = n47490 ^ n44063 ;
  assign n47479 = n47450 ^ n47446 ;
  assign n47480 = n47450 ^ n44113 ;
  assign n47481 = ~n47479 & n47480 ;
  assign n47482 = n47481 ^ n44113 ;
  assign n47492 = n47491 ^ n47482 ;
  assign n47540 = ~n47478 & n47492 ;
  assign n47533 = n45408 ^ n37373 ;
  assign n47534 = n47533 ^ n41604 ;
  assign n47535 = n47534 ^ n35936 ;
  assign n47531 = n44063 ^ n44056 ;
  assign n47526 = n45333 ^ n44549 ;
  assign n47527 = n47526 ^ n46159 ;
  assign n47529 = n47528 ^ n47527 ;
  assign n47530 = n47529 ^ n47488 ;
  assign n47532 = n47531 ^ n47530 ;
  assign n47536 = n47535 ^ n47532 ;
  assign n47499 = n45429 ^ n37387 ;
  assign n47500 = n47499 ^ n41608 ;
  assign n47501 = n47500 ^ n2657 ;
  assign n47537 = n47536 ^ n47501 ;
  assign n47524 = n47490 ^ n47482 ;
  assign n47525 = ~n47491 & n47524 ;
  assign n47538 = n47537 ^ n47525 ;
  assign n47522 = n47486 ^ n47485 ;
  assign n47523 = n47489 & ~n47522 ;
  assign n47539 = n47538 ^ n47523 ;
  assign n47541 = n47540 ^ n47539 ;
  assign n47493 = n47492 ^ n47478 ;
  assign n47494 = n47493 ^ n47456 ;
  assign n47495 = n47494 ^ n47493 ;
  assign n47496 = n47495 ^ n47438 ;
  assign n47497 = n47457 & ~n47496 ;
  assign n47498 = n47497 ^ n47494 ;
  assign n47520 = n47501 ^ n47493 ;
  assign n47521 = ~n47498 & n47520 ;
  assign n47542 = n47541 ^ n47521 ;
  assign n47550 = n47549 ^ n47542 ;
  assign n47518 = n45974 ^ n45503 ;
  assign n47519 = n47518 ^ n46596 ;
  assign n47543 = n47542 ^ n47519 ;
  assign n47502 = n47501 ^ n47498 ;
  assign n47476 = n45978 ^ n45319 ;
  assign n47477 = n47476 ^ n46604 ;
  assign n47503 = n47502 ^ n47477 ;
  assign n47473 = n47464 ^ n47458 ;
  assign n47474 = ~n47462 & ~n47473 ;
  assign n47475 = n47474 ^ n47458 ;
  assign n47515 = n47477 ^ n47475 ;
  assign n47516 = n47503 & n47515 ;
  assign n47517 = n47516 ^ n47502 ;
  assign n47547 = n47519 ^ n47517 ;
  assign n47548 = n47543 & ~n47547 ;
  assign n47551 = n47550 ^ n47548 ;
  assign n47552 = n46594 ^ n45970 ;
  assign n47553 = n47552 ^ n45506 ;
  assign n47562 = n47553 ^ n47549 ;
  assign n47563 = n47551 & ~n47562 ;
  assign n47564 = n47563 ^ n47549 ;
  assign n47581 = n47580 ^ n47564 ;
  assign n47582 = ~n47569 & n47581 ;
  assign n47583 = n47582 ^ n47579 ;
  assign n47584 = n46585 ^ n45962 ;
  assign n47585 = n47584 ^ n45524 ;
  assign n47594 = n47585 ^ n47578 ;
  assign n47595 = ~n47583 & ~n47594 ;
  assign n47598 = n47597 ^ n47595 ;
  assign n47599 = n45958 ^ n45311 ;
  assign n47600 = n47599 ^ n46581 ;
  assign n47683 = n47600 ^ n47596 ;
  assign n47684 = ~n47598 & ~n47683 ;
  assign n47687 = n47686 ^ n47684 ;
  assign n47688 = n46574 ^ n45312 ;
  assign n47689 = n47688 ^ n45954 ;
  assign n47781 = n47689 ^ n47685 ;
  assign n47782 = n47687 & ~n47781 ;
  assign n47783 = n47782 ^ n47689 ;
  assign n47784 = n47783 ^ n47777 ;
  assign n47785 = ~n47780 & ~n47784 ;
  assign n47787 = n47786 ^ n47785 ;
  assign n47788 = n47776 & ~n47787 ;
  assign n47789 = n47788 ^ n47775 ;
  assign n47790 = n47789 ^ n47771 ;
  assign n47791 = ~n47772 & n47790 ;
  assign n47792 = n47791 ^ n47771 ;
  assign n47793 = n47792 ^ n47765 ;
  assign n47794 = n47766 & n47793 ;
  assign n47767 = n47765 ^ n47696 ;
  assign n47795 = n47794 ^ n47767 ;
  assign n47796 = ~n47762 & ~n47795 ;
  assign n47759 = n47757 ^ n47696 ;
  assign n47797 = n47796 ^ n47759 ;
  assign n47798 = n47758 & ~n47797 ;
  assign n47799 = n47798 ^ n47757 ;
  assign n47800 = n47799 ^ n47752 ;
  assign n47801 = n47754 & n47800 ;
  assign n47802 = n47801 ^ n47753 ;
  assign n47803 = n47802 ^ n47748 ;
  assign n47804 = n47750 & ~n47803 ;
  assign n47805 = n47804 ^ n47749 ;
  assign n47806 = n47805 ^ n47743 ;
  assign n47807 = n47744 & n47806 ;
  assign n47745 = n47743 ^ n47737 ;
  assign n47808 = n47807 ^ n47745 ;
  assign n47809 = n47740 & ~n47808 ;
  assign n47738 = n47737 ^ n47733 ;
  assign n47810 = n47809 ^ n47738 ;
  assign n47811 = ~n47735 & n47810 ;
  assign n47812 = n47811 ^ n47734 ;
  assign n47813 = n47812 ^ n47729 ;
  assign n47814 = ~n47731 & n47813 ;
  assign n47815 = n47814 ^ n47730 ;
  assign n47816 = n47815 ^ n47724 ;
  assign n47817 = ~n47725 & ~n47816 ;
  assign n47726 = n47724 ^ n47720 ;
  assign n47818 = n47817 ^ n47726 ;
  assign n47819 = ~n47721 & n47818 ;
  assign n47820 = n47819 ^ n47720 ;
  assign n47821 = n47820 ^ n47716 ;
  assign n47822 = ~n47717 & ~n47821 ;
  assign n47823 = n47822 ^ n47820 ;
  assign n47824 = n47823 ^ n47710 ;
  assign n47825 = ~n47713 & ~n47824 ;
  assign n47826 = n47825 ^ n47712 ;
  assign n47827 = n47826 ^ n47706 ;
  assign n47828 = n47709 & ~n47827 ;
  assign n47829 = n47828 ^ n47708 ;
  assign n47934 = n47933 ^ n47829 ;
  assign n47935 = ~n47833 & n47934 ;
  assign n47936 = n47935 ^ n47932 ;
  assign n47939 = n47938 ^ n47936 ;
  assign n47940 = n47939 ^ n44802 ;
  assign n47835 = n47826 ^ n47709 ;
  assign n47836 = n47835 ^ n44774 ;
  assign n47919 = n47823 ^ n47713 ;
  assign n47838 = n47818 ^ n47718 ;
  assign n47839 = n47838 ^ n45371 ;
  assign n47840 = n47815 ^ n47725 ;
  assign n47841 = n47840 ^ n45345 ;
  assign n47843 = n47810 ^ n47734 ;
  assign n47844 = n47843 ^ n45354 ;
  assign n47846 = n47805 ^ n47744 ;
  assign n47847 = n47846 ^ n44907 ;
  assign n47888 = n47802 ^ n47750 ;
  assign n47848 = n47799 ^ n47754 ;
  assign n47849 = n47848 ^ n44470 ;
  assign n47880 = n47797 ^ n47756 ;
  assign n47850 = n47795 ^ n47761 ;
  assign n47851 = n47850 ^ n44480 ;
  assign n47861 = n47787 ^ n47773 ;
  assign n47690 = n47689 ^ n47687 ;
  assign n47691 = n47690 ^ n44509 ;
  assign n47504 = n47503 ^ n47475 ;
  assign n47505 = n47504 ^ n44534 ;
  assign n47506 = n47465 ^ n44536 ;
  assign n47507 = n47470 & n47506 ;
  assign n47508 = n47507 ^ n44536 ;
  assign n47511 = n47508 ^ n47504 ;
  assign n47512 = n47505 & ~n47511 ;
  assign n47513 = n47512 ^ n44534 ;
  assign n47514 = n47513 ^ n44528 ;
  assign n47544 = n47543 ^ n47517 ;
  assign n47556 = n47544 ^ n47513 ;
  assign n47557 = n47514 & n47556 ;
  assign n47558 = n47557 ^ n44528 ;
  assign n47554 = n47553 ^ n47551 ;
  assign n47561 = n47558 ^ n47554 ;
  assign n47570 = n47569 ^ n47564 ;
  assign n47571 = n47570 ^ n44524 ;
  assign n47572 = n47571 ^ n47570 ;
  assign n47573 = n47572 ^ n47554 ;
  assign n47574 = ~n47561 & ~n47573 ;
  assign n47575 = n47574 ^ n47571 ;
  assign n47588 = n47570 ^ n44520 ;
  assign n47589 = n47575 & n47588 ;
  assign n47590 = n47589 ^ n44520 ;
  assign n47586 = n47585 ^ n47583 ;
  assign n47593 = n47590 ^ n47586 ;
  assign n47601 = n47600 ^ n47598 ;
  assign n47602 = n47601 ^ n44518 ;
  assign n47603 = n47602 ^ n47601 ;
  assign n47604 = n47603 ^ n47586 ;
  assign n47605 = ~n47593 & ~n47604 ;
  assign n47606 = n47605 ^ n47602 ;
  assign n47680 = n47601 ^ n44511 ;
  assign n47681 = ~n47606 & n47680 ;
  assign n47682 = n47681 ^ n44511 ;
  assign n47853 = n47690 ^ n47682 ;
  assign n47854 = n47691 & n47853 ;
  assign n47855 = n47854 ^ n44509 ;
  assign n47856 = n47855 ^ n44500 ;
  assign n47857 = n47783 ^ n47780 ;
  assign n47858 = n47857 ^ n47855 ;
  assign n47859 = ~n47856 & ~n47858 ;
  assign n47860 = n47859 ^ n44500 ;
  assign n47862 = n47861 ^ n47860 ;
  assign n47863 = n47861 ^ n44495 ;
  assign n47864 = n47862 & ~n47863 ;
  assign n47865 = n47864 ^ n44495 ;
  assign n47852 = n47789 ^ n47772 ;
  assign n47866 = n47865 ^ n47852 ;
  assign n47867 = n47792 ^ n47766 ;
  assign n47868 = n47867 ^ n44493 ;
  assign n47869 = n47868 ^ n47852 ;
  assign n47870 = n47869 ^ n47867 ;
  assign n47871 = n47866 & n47870 ;
  assign n47872 = n47871 ^ n47868 ;
  assign n47874 = n47850 ^ n44488 ;
  assign n47873 = n47867 ^ n47850 ;
  assign n47875 = n47874 ^ n47873 ;
  assign n47876 = n47872 & ~n47875 ;
  assign n47877 = n47876 ^ n47874 ;
  assign n47878 = n47851 & ~n47877 ;
  assign n47879 = n47878 ^ n44480 ;
  assign n47881 = n47880 ^ n47879 ;
  assign n47882 = n47880 ^ n44478 ;
  assign n47883 = ~n47881 & n47882 ;
  assign n47884 = n47883 ^ n44478 ;
  assign n47885 = n47884 ^ n47848 ;
  assign n47886 = ~n47849 & n47885 ;
  assign n47887 = n47886 ^ n44470 ;
  assign n47889 = n47888 ^ n47887 ;
  assign n47890 = n47846 ^ n44468 ;
  assign n47891 = n47890 ^ n47846 ;
  assign n47892 = n47891 ^ n47887 ;
  assign n47893 = ~n47889 & n47892 ;
  assign n47894 = n47893 ^ n47890 ;
  assign n47895 = ~n47847 & ~n47894 ;
  assign n47896 = n47895 ^ n44907 ;
  assign n47845 = n47808 ^ n47739 ;
  assign n47897 = n47896 ^ n47845 ;
  assign n47898 = n47896 ^ n45277 ;
  assign n47899 = n47897 & n47898 ;
  assign n47900 = n47899 ^ n45277 ;
  assign n47901 = n47900 ^ n47843 ;
  assign n47902 = ~n47844 & n47901 ;
  assign n47903 = n47902 ^ n45354 ;
  assign n47842 = n47812 ^ n47731 ;
  assign n47904 = n47903 ^ n47842 ;
  assign n47905 = n47840 ^ n45349 ;
  assign n47906 = n47905 ^ n47840 ;
  assign n47907 = n47906 ^ n47842 ;
  assign n47908 = n47904 & n47907 ;
  assign n47909 = n47908 ^ n47905 ;
  assign n47910 = ~n47841 & ~n47909 ;
  assign n47911 = n47910 ^ n45345 ;
  assign n47912 = n47911 ^ n47838 ;
  assign n47913 = n47839 & ~n47912 ;
  assign n47914 = n47913 ^ n45371 ;
  assign n47837 = n47820 ^ n47717 ;
  assign n47915 = n47914 ^ n47837 ;
  assign n47916 = n47914 ^ n45297 ;
  assign n47917 = n47915 & n47916 ;
  assign n47918 = n47917 ^ n45297 ;
  assign n47920 = n47919 ^ n47918 ;
  assign n47921 = n47919 ^ n44724 ;
  assign n47922 = ~n47920 & n47921 ;
  assign n47923 = n47922 ^ n44724 ;
  assign n47924 = n47923 ^ n47835 ;
  assign n47925 = ~n47836 & ~n47924 ;
  assign n47926 = n47925 ^ n44774 ;
  assign n47834 = n47833 ^ n47829 ;
  assign n47927 = n47926 ^ n47834 ;
  assign n47928 = n47926 ^ n44771 ;
  assign n47929 = ~n47927 & n47928 ;
  assign n47930 = n47929 ^ n44771 ;
  assign n47941 = n47940 ^ n47930 ;
  assign n47942 = n47837 ^ n45297 ;
  assign n47943 = n47942 ^ n47914 ;
  assign n47944 = n47911 ^ n47839 ;
  assign n47945 = n47909 ^ n45345 ;
  assign n47946 = n47842 ^ n45349 ;
  assign n47947 = n47946 ^ n47903 ;
  assign n47948 = n47894 ^ n44907 ;
  assign n47949 = n47887 ^ n44468 ;
  assign n47950 = n47949 ^ n47888 ;
  assign n47951 = n47877 ^ n44480 ;
  assign n47952 = n47872 ^ n44488 ;
  assign n47472 = n47434 & ~n47471 ;
  assign n47509 = n47508 ^ n47505 ;
  assign n47510 = ~n47472 & ~n47509 ;
  assign n47545 = n47544 ^ n47514 ;
  assign n47546 = ~n47510 & ~n47545 ;
  assign n47555 = n47554 ^ n44524 ;
  assign n47559 = n47558 ^ n47555 ;
  assign n47560 = ~n47546 & n47559 ;
  assign n47576 = n47575 ^ n44520 ;
  assign n47577 = ~n47560 & ~n47576 ;
  assign n47587 = n47586 ^ n44518 ;
  assign n47591 = n47590 ^ n47587 ;
  assign n47592 = n47577 & ~n47591 ;
  assign n47607 = n47606 ^ n44511 ;
  assign n47679 = n47592 & ~n47607 ;
  assign n47692 = n47691 ^ n47682 ;
  assign n47953 = ~n47679 & n47692 ;
  assign n47954 = n47857 ^ n47856 ;
  assign n47955 = n47953 & n47954 ;
  assign n47956 = n47863 ^ n47860 ;
  assign n47957 = n47955 & ~n47956 ;
  assign n47958 = n47852 ^ n44493 ;
  assign n47959 = n47958 ^ n47865 ;
  assign n47960 = n47957 & n47959 ;
  assign n47961 = n47952 & n47960 ;
  assign n47962 = n47951 & ~n47961 ;
  assign n47963 = n47882 ^ n47879 ;
  assign n47964 = n47962 & n47963 ;
  assign n47965 = n47884 ^ n47849 ;
  assign n47966 = ~n47964 & n47965 ;
  assign n47967 = n47950 & ~n47966 ;
  assign n47968 = n47948 & ~n47967 ;
  assign n47969 = n47845 ^ n45277 ;
  assign n47970 = n47969 ^ n47896 ;
  assign n47971 = n47968 & ~n47970 ;
  assign n47972 = n47900 ^ n47844 ;
  assign n47973 = n47971 & ~n47972 ;
  assign n47974 = ~n47947 & ~n47973 ;
  assign n47975 = ~n47945 & n47974 ;
  assign n47976 = n47944 & ~n47975 ;
  assign n47977 = ~n47943 & n47976 ;
  assign n47978 = n47921 ^ n47918 ;
  assign n47979 = ~n47977 & ~n47978 ;
  assign n47980 = n47923 ^ n47836 ;
  assign n47981 = ~n47979 & ~n47980 ;
  assign n47982 = n47834 ^ n44771 ;
  assign n47983 = n47982 ^ n47926 ;
  assign n47984 = ~n47981 & n47983 ;
  assign n48139 = ~n47941 & ~n47984 ;
  assign n48149 = n46159 ^ n45456 ;
  assign n48150 = n48149 ^ n46882 ;
  assign n48143 = n47369 ^ n47185 ;
  assign n48145 = n48143 ^ n47931 ;
  assign n48144 = n48143 ^ n47938 ;
  assign n48146 = n48145 ^ n48144 ;
  assign n48147 = n47936 & n48146 ;
  assign n48148 = n48147 ^ n48145 ;
  assign n48151 = n48150 ^ n48148 ;
  assign n48152 = n48151 ^ n44833 ;
  assign n48140 = n47939 ^ n47930 ;
  assign n48141 = n47940 & n48140 ;
  assign n48142 = n48141 ^ n44802 ;
  assign n48153 = n48152 ^ n48142 ;
  assign n48177 = n48139 & ~n48153 ;
  assign n48187 = n48151 ^ n48142 ;
  assign n48188 = ~n48152 & n48187 ;
  assign n48189 = n48188 ^ n44833 ;
  assign n48190 = n48189 ^ n44553 ;
  assign n48184 = n46880 ^ n45339 ;
  assign n48185 = n48184 ^ n45994 ;
  assign n48178 = n47372 ^ n47178 ;
  assign n48180 = n48178 ^ n48143 ;
  assign n48179 = n48178 ^ n48150 ;
  assign n48181 = n48180 ^ n48179 ;
  assign n48182 = ~n48148 & ~n48181 ;
  assign n48183 = n48182 ^ n48180 ;
  assign n48186 = n48185 ^ n48183 ;
  assign n48191 = n48190 ^ n48186 ;
  assign n48236 = ~n48177 & ~n48191 ;
  assign n48231 = n48185 ^ n46876 ;
  assign n48228 = n47374 ^ n47174 ;
  assign n48223 = n46091 ^ n2660 ;
  assign n48224 = n48223 ^ n42433 ;
  assign n48225 = n48224 ^ n36683 ;
  assign n48226 = n48225 ^ n46195 ;
  assign n48227 = n48226 ^ n47526 ;
  assign n48229 = n48228 ^ n48227 ;
  assign n48230 = n48229 ^ n44553 ;
  assign n48232 = n48231 ^ n48230 ;
  assign n48193 = n46095 ^ n38064 ;
  assign n48194 = n48193 ^ n42437 ;
  assign n48195 = n48194 ^ n36545 ;
  assign n48233 = n48232 ^ n48195 ;
  assign n48221 = n48189 ^ n48186 ;
  assign n48222 = n48190 & ~n48221 ;
  assign n48234 = n48233 ^ n48222 ;
  assign n48219 = n48185 ^ n48178 ;
  assign n48220 = n48183 & ~n48219 ;
  assign n48235 = n48234 ^ n48220 ;
  assign n48237 = n48236 ^ n48235 ;
  assign n48192 = n48191 ^ n48177 ;
  assign n48196 = n48195 ^ n48192 ;
  assign n48134 = n46101 ^ n38069 ;
  assign n48135 = n48134 ^ n42442 ;
  assign n48136 = n48135 ^ n36502 ;
  assign n47985 = n47984 ^ n47941 ;
  assign n48137 = n48136 ^ n47985 ;
  assign n47703 = n46105 ^ n38073 ;
  assign n47704 = n47703 ^ n42447 ;
  assign n47705 = n47704 ^ n36292 ;
  assign n47986 = n47985 ^ n47705 ;
  assign n47990 = n47983 ^ n47981 ;
  assign n47987 = n46110 ^ n2895 ;
  assign n47988 = n47987 ^ n42453 ;
  assign n47989 = n47988 ^ n36288 ;
  assign n47991 = n47990 ^ n47989 ;
  assign n47993 = n46116 ^ n38083 ;
  assign n47994 = n47993 ^ n42458 ;
  assign n47995 = n47994 ^ n36298 ;
  assign n47992 = n47980 ^ n47979 ;
  assign n47996 = n47995 ^ n47992 ;
  assign n48000 = n47978 ^ n47977 ;
  assign n48125 = n48000 ^ n47995 ;
  assign n47997 = n45940 ^ n38088 ;
  assign n47998 = n47997 ^ n42463 ;
  assign n47999 = n47998 ^ n1388 ;
  assign n48001 = n48000 ^ n47999 ;
  assign n48003 = n45301 ^ n1766 ;
  assign n48004 = n48003 ^ n1184 ;
  assign n48005 = n48004 ^ n36304 ;
  assign n48002 = n47976 ^ n47943 ;
  assign n48006 = n48005 ^ n48002 ;
  assign n48012 = n47975 ^ n47944 ;
  assign n48009 = n45747 ^ n1757 ;
  assign n48010 = n48009 ^ n42469 ;
  assign n48011 = n48010 ^ n1176 ;
  assign n48013 = n48012 ^ n48011 ;
  assign n48014 = n47974 ^ n47945 ;
  assign n1005 = n1004 ^ n965 ;
  assign n1039 = n1038 ^ n1005 ;
  assign n1049 = n1048 ^ n1039 ;
  assign n48015 = n48014 ^ n1049 ;
  assign n48016 = n45755 ^ n38098 ;
  assign n48017 = n48016 ^ n42476 ;
  assign n48018 = n48017 ^ n1030 ;
  assign n48114 = n48018 ^ n1049 ;
  assign n48019 = n47973 ^ n47947 ;
  assign n48020 = n48019 ^ n48018 ;
  assign n48024 = n47972 ^ n47971 ;
  assign n48025 = n48024 ^ n48023 ;
  assign n48029 = n47970 ^ n47968 ;
  assign n48030 = n48029 ^ n48028 ;
  assign n48032 = n45771 ^ n1595 ;
  assign n48033 = n48032 ^ n42488 ;
  assign n48034 = n48033 ^ n36322 ;
  assign n48105 = n48034 ^ n48028 ;
  assign n48031 = n47967 ^ n47948 ;
  assign n48035 = n48034 ^ n48031 ;
  assign n48037 = n45775 ^ n37643 ;
  assign n48038 = n48037 ^ n42493 ;
  assign n48039 = n48038 ^ n36327 ;
  assign n48102 = n48039 ^ n48034 ;
  assign n48036 = n47966 ^ n47950 ;
  assign n48040 = n48039 ^ n48036 ;
  assign n48044 = n47965 ^ n47964 ;
  assign n48041 = n45780 ^ n37647 ;
  assign n48042 = n48041 ^ n42499 ;
  assign n48043 = n48042 ^ n2966 ;
  assign n48045 = n48044 ^ n48043 ;
  assign n48049 = n47963 ^ n47962 ;
  assign n48096 = n48049 ^ n48044 ;
  assign n48046 = n45787 ^ n37652 ;
  assign n48047 = n48046 ^ n42505 ;
  assign n48048 = n48047 ^ n36335 ;
  assign n48050 = n48049 ^ n48048 ;
  assign n48055 = n47961 ^ n47951 ;
  assign n48051 = n45791 ^ n37658 ;
  assign n48052 = n48051 ^ n42511 ;
  assign n48053 = n48052 ^ n36342 ;
  assign n48056 = n48055 ^ n48053 ;
  assign n48060 = n47960 ^ n47952 ;
  assign n48057 = n45796 ^ n37665 ;
  assign n48058 = n48057 ^ n42515 ;
  assign n48059 = n48058 ^ n36347 ;
  assign n48061 = n48060 ^ n48059 ;
  assign n48065 = n47959 ^ n47957 ;
  assign n48062 = n45801 ^ n37669 ;
  assign n48063 = n48062 ^ n42520 ;
  assign n48064 = n48063 ^ n36351 ;
  assign n48066 = n48065 ^ n48064 ;
  assign n48082 = n47956 ^ n47955 ;
  assign n48074 = n47954 ^ n47953 ;
  assign n48071 = n45809 ^ n2359 ;
  assign n48072 = n48071 ^ n42530 ;
  assign n48073 = n48072 ^ n36362 ;
  assign n48075 = n48074 ^ n48073 ;
  assign n47693 = n47692 ^ n47679 ;
  assign n47676 = n45813 ^ n2341 ;
  assign n47677 = n47676 ^ n42028 ;
  assign n47678 = n47677 ^ n36367 ;
  assign n47694 = n47693 ^ n47678 ;
  assign n47609 = n45819 ^ n37733 ;
  assign n47610 = n47609 ^ n41953 ;
  assign n47611 = n47610 ^ n36372 ;
  assign n47608 = n47607 ^ n47592 ;
  assign n47612 = n47611 ^ n47608 ;
  assign n47616 = n47591 ^ n47577 ;
  assign n47613 = n45824 ^ n37686 ;
  assign n47614 = n47613 ^ n41957 ;
  assign n47615 = n47614 ^ n36402 ;
  assign n47617 = n47616 ^ n47615 ;
  assign n47619 = n45828 ^ n37691 ;
  assign n47620 = n47619 ^ n41962 ;
  assign n47621 = n47620 ^ n36377 ;
  assign n47669 = n47621 ^ n47615 ;
  assign n47618 = n47576 ^ n47560 ;
  assign n47622 = n47621 ^ n47618 ;
  assign n47624 = n45833 ^ n37720 ;
  assign n47625 = n47624 ^ n41967 ;
  assign n47626 = n47625 ^ n1970 ;
  assign n47666 = n47626 ^ n47621 ;
  assign n47623 = n47559 ^ n47546 ;
  assign n47627 = n47626 ^ n47623 ;
  assign n47631 = n47545 ^ n47510 ;
  assign n47628 = n45838 ^ n37695 ;
  assign n47629 = n47628 ^ n41991 ;
  assign n47630 = n47629 ^ n36384 ;
  assign n47632 = n47631 ^ n47630 ;
  assign n47634 = n45844 ^ n37700 ;
  assign n47635 = n47634 ^ n41972 ;
  assign n47636 = n47635 ^ n35785 ;
  assign n47660 = n47636 ^ n47631 ;
  assign n47633 = n47509 ^ n47472 ;
  assign n47637 = n47636 ^ n47633 ;
  assign n47656 = n47655 ^ n47649 ;
  assign n47657 = n47652 & n47656 ;
  assign n47650 = n47649 ^ n47636 ;
  assign n47658 = n47657 ^ n47650 ;
  assign n47659 = n47637 & n47658 ;
  assign n47661 = n47660 ^ n47659 ;
  assign n47662 = ~n47632 & ~n47661 ;
  assign n47663 = n47662 ^ n47631 ;
  assign n47664 = n47663 ^ n47626 ;
  assign n47665 = ~n47627 & ~n47664 ;
  assign n47667 = n47666 ^ n47665 ;
  assign n47668 = ~n47622 & n47667 ;
  assign n47670 = n47669 ^ n47668 ;
  assign n47671 = n47617 & ~n47670 ;
  assign n47672 = n47671 ^ n47616 ;
  assign n47673 = n47672 ^ n47608 ;
  assign n47674 = n47612 & ~n47673 ;
  assign n47675 = n47674 ^ n47611 ;
  assign n48077 = n47678 ^ n47675 ;
  assign n48078 = ~n47694 & n48077 ;
  assign n48076 = n48074 ^ n47678 ;
  assign n48079 = n48078 ^ n48076 ;
  assign n48080 = n48075 & n48079 ;
  assign n48081 = n48080 ^ n48074 ;
  assign n48083 = n48082 ^ n48081 ;
  assign n48067 = n37675 ^ n2430 ;
  assign n48068 = n48067 ^ n42526 ;
  assign n48069 = n48068 ^ n36357 ;
  assign n48084 = n48081 ^ n48069 ;
  assign n48085 = n48083 & n48084 ;
  assign n48070 = n48069 ^ n48064 ;
  assign n48086 = n48085 ^ n48070 ;
  assign n48087 = n48066 & ~n48086 ;
  assign n48088 = n48087 ^ n48065 ;
  assign n48089 = n48088 ^ n48059 ;
  assign n48090 = n48061 & ~n48089 ;
  assign n48091 = n48090 ^ n48060 ;
  assign n48092 = n48091 ^ n48053 ;
  assign n48093 = n48056 & n48092 ;
  assign n48054 = n48053 ^ n48048 ;
  assign n48094 = n48093 ^ n48054 ;
  assign n48095 = ~n48050 & ~n48094 ;
  assign n48097 = n48096 ^ n48095 ;
  assign n48098 = ~n48045 & n48097 ;
  assign n48099 = n48098 ^ n48044 ;
  assign n48100 = n48099 ^ n48039 ;
  assign n48101 = n48040 & ~n48100 ;
  assign n48103 = n48102 ^ n48101 ;
  assign n48104 = ~n48035 & n48103 ;
  assign n48106 = n48105 ^ n48104 ;
  assign n48107 = ~n48030 & ~n48106 ;
  assign n48108 = n48107 ^ n48029 ;
  assign n48109 = n48108 ^ n48023 ;
  assign n48110 = ~n48025 & n48109 ;
  assign n48111 = n48110 ^ n48024 ;
  assign n48112 = n48111 ^ n48018 ;
  assign n48113 = ~n48020 & ~n48112 ;
  assign n48115 = n48114 ^ n48113 ;
  assign n48116 = n48015 & ~n48115 ;
  assign n48117 = n48116 ^ n48014 ;
  assign n48118 = n48117 ^ n48011 ;
  assign n48119 = ~n48013 & ~n48118 ;
  assign n48120 = n48119 ^ n48012 ;
  assign n48007 = n48005 ^ n47999 ;
  assign n48008 = n48007 ^ n47999 ;
  assign n48121 = n48120 ^ n48008 ;
  assign n48122 = ~n48006 & ~n48121 ;
  assign n48123 = n48122 ^ n48007 ;
  assign n48124 = ~n48001 & ~n48123 ;
  assign n48126 = n48125 ^ n48124 ;
  assign n48127 = n47996 & ~n48126 ;
  assign n48128 = n48127 ^ n47995 ;
  assign n48129 = n48128 ^ n47989 ;
  assign n48130 = n47991 & ~n48129 ;
  assign n48131 = n48130 ^ n47990 ;
  assign n48132 = n48131 ^ n47705 ;
  assign n48133 = n47986 & ~n48132 ;
  assign n48138 = n48137 ^ n48133 ;
  assign n48154 = n48153 ^ n48139 ;
  assign n48174 = n48154 ^ n48136 ;
  assign n48175 = n48138 & ~n48174 ;
  assign n48176 = n48175 ^ n48136 ;
  assign n48217 = n48195 ^ n48176 ;
  assign n48218 = ~n48196 & n48217 ;
  assign n48238 = n48237 ^ n48218 ;
  assign n48215 = n46587 ^ n45974 ;
  assign n48216 = n48215 ^ n47685 ;
  assign n48239 = n48238 ^ n48216 ;
  assign n48170 = n47596 ^ n45978 ;
  assign n48171 = n48170 ^ n46594 ;
  assign n48155 = n48154 ^ n48138 ;
  assign n48172 = n48171 ^ n48155 ;
  assign n47701 = n47578 ^ n45982 ;
  assign n47702 = n47701 ^ n46596 ;
  assign n48156 = n48155 ^ n47702 ;
  assign n48160 = n46608 ^ n45990 ;
  assign n48161 = n48160 ^ n47549 ;
  assign n48162 = n48128 ^ n47991 ;
  assign n48163 = n48161 & n48162 ;
  assign n48157 = n46604 ^ n45986 ;
  assign n48158 = n48157 ^ n47568 ;
  assign n48164 = n48163 ^ n48158 ;
  assign n48165 = n48131 ^ n47986 ;
  assign n48166 = n48165 ^ n48158 ;
  assign n48167 = n48164 & n48166 ;
  assign n48159 = n48158 ^ n47702 ;
  assign n48168 = n48167 ^ n48159 ;
  assign n48169 = n48156 & n48168 ;
  assign n48173 = n48172 ^ n48169 ;
  assign n48197 = n48196 ^ n48176 ;
  assign n48212 = n48197 ^ n48171 ;
  assign n48213 = ~n48173 & ~n48212 ;
  assign n48214 = n48213 ^ n48171 ;
  assign n48254 = n48238 ^ n48214 ;
  assign n48255 = ~n48239 & n48254 ;
  assign n48256 = n48255 ^ n48238 ;
  assign n48269 = n48259 ^ n48256 ;
  assign n48270 = n48260 & n48269 ;
  assign n48271 = n48270 ^ n48259 ;
  assign n48336 = n48273 ^ n48271 ;
  assign n48337 = ~n48275 & n48336 ;
  assign n48338 = n48337 ^ n48274 ;
  assign n48421 = n48340 ^ n48338 ;
  assign n48422 = ~n48342 & n48421 ;
  assign n48423 = n48422 ^ n48341 ;
  assign n48419 = n47658 ^ n47633 ;
  assign n48417 = n47765 ^ n45958 ;
  assign n48418 = n48417 ^ n46937 ;
  assign n48420 = n48419 ^ n48418 ;
  assign n48504 = n48423 ^ n48420 ;
  assign n48206 = n48168 ^ n48155 ;
  assign n48199 = n48162 ^ n48161 ;
  assign n48200 = ~n45331 & n48199 ;
  assign n48201 = n48200 ^ n45327 ;
  assign n48202 = n48165 ^ n48164 ;
  assign n48203 = n48202 ^ n48200 ;
  assign n48204 = n48201 & ~n48203 ;
  assign n48205 = n48204 ^ n45327 ;
  assign n48207 = n48206 ^ n48205 ;
  assign n48208 = n48206 ^ n45321 ;
  assign n48209 = ~n48207 & ~n48208 ;
  assign n48210 = n48209 ^ n45321 ;
  assign n48198 = n48197 ^ n48173 ;
  assign n48211 = n48210 ^ n48198 ;
  assign n48240 = n48239 ^ n48214 ;
  assign n48241 = n48240 ^ n45319 ;
  assign n48242 = n48241 ^ n48198 ;
  assign n48243 = n48242 ^ n48240 ;
  assign n48244 = n48211 & ~n48243 ;
  assign n48245 = n48244 ^ n48241 ;
  assign n48261 = n48260 ^ n48256 ;
  assign n48263 = n48261 ^ n45503 ;
  assign n48262 = n48261 ^ n48240 ;
  assign n48264 = n48263 ^ n48262 ;
  assign n48265 = ~n48245 & ~n48264 ;
  assign n48266 = n48265 ^ n48263 ;
  assign n48276 = n48275 ^ n48271 ;
  assign n48278 = n48276 ^ n45506 ;
  assign n48277 = n48276 ^ n48261 ;
  assign n48279 = n48278 ^ n48277 ;
  assign n48280 = ~n48266 & ~n48279 ;
  assign n48281 = n48280 ^ n48278 ;
  assign n48345 = n48276 ^ n45516 ;
  assign n48346 = ~n48281 & n48345 ;
  assign n48347 = n48346 ^ n45516 ;
  assign n48343 = n48342 ^ n48338 ;
  assign n48500 = n48347 ^ n48343 ;
  assign n48501 = n48347 ^ n45524 ;
  assign n48502 = ~n48500 & n48501 ;
  assign n48503 = n48502 ^ n45524 ;
  assign n48505 = n48504 ^ n48503 ;
  assign n48506 = n48504 ^ n45311 ;
  assign n48507 = ~n48505 & ~n48506 ;
  assign n48508 = n48507 ^ n45311 ;
  assign n48593 = n48508 ^ n45312 ;
  assign n48424 = n48423 ^ n48418 ;
  assign n48425 = ~n48420 & n48424 ;
  assign n48426 = n48425 ^ n48419 ;
  assign n48415 = n47661 ^ n47630 ;
  assign n48413 = n47696 ^ n46566 ;
  assign n48414 = n48413 ^ n45954 ;
  assign n48416 = n48415 ^ n48414 ;
  assign n48498 = n48426 ^ n48416 ;
  assign n48594 = n48593 ^ n48498 ;
  assign n48595 = n48506 ^ n48503 ;
  assign n48246 = n48245 ^ n45503 ;
  assign n48247 = n48210 ^ n45319 ;
  assign n48248 = n48247 ^ n48198 ;
  assign n48249 = n48202 ^ n48201 ;
  assign n48250 = n48208 ^ n48205 ;
  assign n48251 = ~n48249 & n48250 ;
  assign n48252 = n48248 & ~n48251 ;
  assign n48253 = ~n48246 & ~n48252 ;
  assign n48267 = n48266 ^ n45506 ;
  assign n48268 = ~n48253 & ~n48267 ;
  assign n48282 = n48281 ^ n45516 ;
  assign n48335 = ~n48268 & n48282 ;
  assign n48344 = n48343 ^ n45524 ;
  assign n48348 = n48347 ^ n48344 ;
  assign n48596 = n48335 & n48348 ;
  assign n48597 = ~n48595 & n48596 ;
  assign n48598 = n48594 & ~n48597 ;
  assign n48499 = n48498 ^ n45312 ;
  assign n48509 = n48508 ^ n48498 ;
  assign n48510 = n48499 & ~n48509 ;
  assign n48511 = n48510 ^ n45312 ;
  assign n48409 = n47663 ^ n47627 ;
  assign n48429 = n48415 ^ n48409 ;
  assign n48427 = n48426 ^ n48415 ;
  assign n48428 = n48416 & ~n48427 ;
  assign n48430 = n48429 ^ n48428 ;
  assign n48410 = n46947 ^ n45950 ;
  assign n48411 = n48410 ^ n47757 ;
  assign n48496 = n48430 ^ n48411 ;
  assign n48497 = n48496 ^ n45306 ;
  assign n48599 = n48511 ^ n48497 ;
  assign n48600 = n48598 & n48599 ;
  assign n48512 = n48511 ^ n48496 ;
  assign n48513 = n48497 & n48512 ;
  assign n48514 = n48513 ^ n45306 ;
  assign n48407 = n47667 ^ n47618 ;
  assign n48432 = n48411 ^ n48407 ;
  assign n48412 = n48411 ^ n48409 ;
  assign n48431 = n48412 & n48430 ;
  assign n48433 = n48432 ^ n48431 ;
  assign n48405 = n46564 ^ n46232 ;
  assign n48406 = n48405 ^ n47753 ;
  assign n48494 = n48433 ^ n48406 ;
  assign n48495 = n48494 ^ n45302 ;
  assign n48601 = n48514 ^ n48495 ;
  assign n48602 = n48600 & ~n48601 ;
  assign n48515 = n48514 ^ n48494 ;
  assign n48516 = n48495 & ~n48515 ;
  assign n48517 = n48516 ^ n45302 ;
  assign n48408 = n48407 ^ n48406 ;
  assign n48434 = ~n48408 & ~n48433 ;
  assign n48435 = n48434 ^ n48407 ;
  assign n48403 = n47670 ^ n47616 ;
  assign n48401 = n46559 ^ n46521 ;
  assign n48402 = n48401 ^ n47749 ;
  assign n48404 = n48403 ^ n48402 ;
  assign n48492 = n48435 ^ n48404 ;
  assign n48493 = n48492 ^ n45550 ;
  assign n48603 = n48517 ^ n48493 ;
  assign n48604 = n48602 & ~n48603 ;
  assign n48518 = n48517 ^ n48492 ;
  assign n48519 = n48493 & n48518 ;
  assign n48520 = n48519 ^ n45550 ;
  assign n48436 = n48435 ^ n48402 ;
  assign n48437 = ~n48404 & ~n48436 ;
  assign n48438 = n48437 ^ n48403 ;
  assign n48399 = n47672 ^ n47612 ;
  assign n48397 = n47743 ^ n46554 ;
  assign n48398 = n48397 ^ n46648 ;
  assign n48400 = n48399 ^ n48398 ;
  assign n48490 = n48438 ^ n48400 ;
  assign n48491 = n48490 ^ n45691 ;
  assign n48605 = n48520 ^ n48491 ;
  assign n48606 = n48604 & ~n48605 ;
  assign n48521 = n48520 ^ n48490 ;
  assign n48522 = ~n48491 & ~n48521 ;
  assign n48523 = n48522 ^ n45691 ;
  assign n48439 = n48438 ^ n48398 ;
  assign n48440 = n48400 & ~n48439 ;
  assign n48441 = n48440 ^ n48399 ;
  assign n48394 = n47739 ^ n46568 ;
  assign n48395 = n48394 ^ n46549 ;
  assign n47695 = n47694 ^ n47675 ;
  assign n48396 = n48395 ^ n47695 ;
  assign n48488 = n48441 ^ n48396 ;
  assign n48489 = n48488 ^ n45708 ;
  assign n48607 = n48523 ^ n48489 ;
  assign n48608 = ~n48606 & n48607 ;
  assign n48524 = n48523 ^ n48488 ;
  assign n48525 = n48489 & ~n48524 ;
  assign n48526 = n48525 ^ n45708 ;
  assign n48392 = n48079 ^ n48073 ;
  assign n48444 = n48392 ^ n47695 ;
  assign n48442 = n48441 ^ n47695 ;
  assign n48443 = ~n48396 & ~n48442 ;
  assign n48445 = n48444 ^ n48443 ;
  assign n48390 = n46572 ^ n46544 ;
  assign n48391 = n48390 ^ n47734 ;
  assign n48486 = n48445 ^ n48391 ;
  assign n48487 = n48486 ^ n45722 ;
  assign n48609 = n48526 ^ n48487 ;
  assign n48610 = n48608 & n48609 ;
  assign n48527 = n48526 ^ n48486 ;
  assign n48528 = n48487 & n48527 ;
  assign n48529 = n48528 ^ n45722 ;
  assign n48451 = n48083 ^ n48069 ;
  assign n48448 = n46562 ^ n46539 ;
  assign n48449 = n48448 ^ n47730 ;
  assign n48483 = n48451 ^ n48449 ;
  assign n48393 = n48392 ^ n48391 ;
  assign n48446 = ~n48393 & ~n48445 ;
  assign n48447 = n48446 ^ n48392 ;
  assign n48484 = n48483 ^ n48447 ;
  assign n48485 = n48484 ^ n45732 ;
  assign n48611 = n48529 ^ n48485 ;
  assign n48612 = ~n48610 & n48611 ;
  assign n48530 = n48529 ^ n48484 ;
  assign n48531 = n48485 & ~n48530 ;
  assign n48532 = n48531 ^ n45732 ;
  assign n48450 = n48449 ^ n48447 ;
  assign n48454 = n48451 ^ n48447 ;
  assign n48455 = n48450 & ~n48454 ;
  assign n48388 = n48086 ^ n48065 ;
  assign n48452 = n48451 ^ n48388 ;
  assign n48456 = n48455 ^ n48452 ;
  assign n48386 = n47724 ^ n46557 ;
  assign n48387 = n48386 ^ n46534 ;
  assign n48481 = n48456 ^ n48387 ;
  assign n48482 = n48481 ^ n45930 ;
  assign n48613 = n48532 ^ n48482 ;
  assign n48614 = ~n48612 & n48613 ;
  assign n48389 = n48388 ^ n48387 ;
  assign n48457 = ~n48389 & ~n48456 ;
  assign n48458 = n48457 ^ n48388 ;
  assign n48384 = n48088 ^ n48061 ;
  assign n48382 = n46974 ^ n46552 ;
  assign n48383 = n48382 ^ n47718 ;
  assign n48385 = n48384 ^ n48383 ;
  assign n48480 = n48458 ^ n48385 ;
  assign n48591 = n48480 ^ n46000 ;
  assign n48533 = n48532 ^ n48481 ;
  assign n48534 = ~n48482 & ~n48533 ;
  assign n48535 = n48534 ^ n45930 ;
  assign n48592 = n48591 ^ n48535 ;
  assign n48725 = n48614 ^ n48592 ;
  assign n48646 = n48613 ^ n48612 ;
  assign n48726 = n48725 ^ n48646 ;
  assign n48643 = n46377 ^ n2975 ;
  assign n48644 = n48643 ^ n42894 ;
  assign n48645 = n48644 ^ n37078 ;
  assign n48647 = n48646 ^ n48645 ;
  assign n48651 = n48611 ^ n48610 ;
  assign n48722 = n48651 ^ n48646 ;
  assign n48648 = n46383 ^ n38578 ;
  assign n48649 = n48648 ^ n42899 ;
  assign n48650 = n48649 ^ n37083 ;
  assign n48652 = n48651 ^ n48650 ;
  assign n48653 = n46388 ^ n38583 ;
  assign n48654 = n48653 ^ n42904 ;
  assign n48655 = n48654 ^ n37089 ;
  assign n48719 = n48655 ^ n48651 ;
  assign n48656 = n48609 ^ n48608 ;
  assign n48657 = n48656 ^ n48655 ;
  assign n48661 = n48607 ^ n48606 ;
  assign n48658 = n46392 ^ n38589 ;
  assign n48659 = n48658 ^ n42910 ;
  assign n48660 = n48659 ^ n37094 ;
  assign n48662 = n48661 ^ n48660 ;
  assign n48666 = n48605 ^ n48604 ;
  assign n48663 = n46397 ^ n38593 ;
  assign n48664 = n48663 ^ n42917 ;
  assign n48665 = n48664 ^ n37098 ;
  assign n48667 = n48666 ^ n48665 ;
  assign n48671 = n48603 ^ n48602 ;
  assign n48668 = n46402 ^ n38599 ;
  assign n48669 = n48668 ^ n42921 ;
  assign n48670 = n48669 ^ n37105 ;
  assign n48672 = n48671 ^ n48670 ;
  assign n48676 = n48601 ^ n48600 ;
  assign n48707 = n48676 ^ n48671 ;
  assign n48673 = n46486 ^ n38604 ;
  assign n48674 = n48673 ^ n42926 ;
  assign n48675 = n48674 ^ n37109 ;
  assign n48677 = n48676 ^ n48675 ;
  assign n48679 = n46407 ^ n38608 ;
  assign n48680 = n48679 ^ n42931 ;
  assign n48681 = n48680 ^ n37115 ;
  assign n48704 = n48681 ^ n48675 ;
  assign n48678 = n48599 ^ n48598 ;
  assign n48682 = n48681 ^ n48678 ;
  assign n48684 = n46474 ^ n38614 ;
  assign n48685 = n48684 ^ n42936 ;
  assign n48686 = n48685 ^ n2234 ;
  assign n48683 = n48597 ^ n48594 ;
  assign n48687 = n48686 ^ n48683 ;
  assign n48689 = n46412 ^ n38620 ;
  assign n48690 = n48689 ^ n2132 ;
  assign n48691 = n48690 ^ n37122 ;
  assign n48698 = n48691 ^ n48686 ;
  assign n48688 = n48596 ^ n48595 ;
  assign n48692 = n48691 ^ n48688 ;
  assign n48349 = n48348 ^ n48335 ;
  assign n48332 = n46417 ^ n38624 ;
  assign n48333 = n48332 ^ n42943 ;
  assign n48334 = n48333 ^ n2124 ;
  assign n48350 = n48349 ^ n48334 ;
  assign n48283 = n48282 ^ n48268 ;
  assign n47698 = n46422 ^ n2015 ;
  assign n47699 = n47698 ^ n42947 ;
  assign n47700 = n47699 ^ n37128 ;
  assign n48284 = n48283 ^ n47700 ;
  assign n48286 = n46428 ^ n38632 ;
  assign n48287 = n48286 ^ n42952 ;
  assign n48288 = n48287 ^ n37132 ;
  assign n48328 = n48288 ^ n47700 ;
  assign n48285 = n48267 ^ n48253 ;
  assign n48289 = n48288 ^ n48285 ;
  assign n48291 = n46433 ^ n38636 ;
  assign n48292 = n48291 ^ n42957 ;
  assign n48293 = n48292 ^ n37137 ;
  assign n48325 = n48293 ^ n48288 ;
  assign n48290 = n48252 ^ n48246 ;
  assign n48294 = n48293 ^ n48290 ;
  assign n48298 = n48251 ^ n48248 ;
  assign n48322 = n48298 ^ n48290 ;
  assign n48295 = n46438 ^ n3053 ;
  assign n48296 = n48295 ^ n42962 ;
  assign n48297 = n48296 ^ n36535 ;
  assign n48299 = n48298 ^ n48297 ;
  assign n48304 = n48250 ^ n48249 ;
  assign n48300 = n46442 ^ n38644 ;
  assign n48301 = n48300 ^ n42971 ;
  assign n48302 = n48301 ^ n36491 ;
  assign n48305 = n48304 ^ n48302 ;
  assign n48309 = n46869 ^ n38993 ;
  assign n48310 = n48309 ^ n43335 ;
  assign n48311 = n48310 ^ n3173 ;
  assign n48312 = n48199 ^ n45331 ;
  assign n48313 = n48311 & ~n48312 ;
  assign n48306 = n46446 ^ n2775 ;
  assign n48307 = n48306 ^ n42967 ;
  assign n48308 = n48307 ^ n35828 ;
  assign n48314 = n48313 ^ n48308 ;
  assign n48315 = n48313 ^ n48249 ;
  assign n48316 = ~n48314 & ~n48315 ;
  assign n48317 = n48316 ^ n48249 ;
  assign n48318 = n48317 ^ n48302 ;
  assign n48319 = n48305 & ~n48318 ;
  assign n48303 = n48302 ^ n48297 ;
  assign n48320 = n48319 ^ n48303 ;
  assign n48321 = ~n48299 & ~n48320 ;
  assign n48323 = n48322 ^ n48321 ;
  assign n48324 = ~n48294 & ~n48323 ;
  assign n48326 = n48325 ^ n48324 ;
  assign n48327 = n48289 & n48326 ;
  assign n48329 = n48328 ^ n48327 ;
  assign n48330 = n48284 & ~n48329 ;
  assign n48331 = n48330 ^ n48283 ;
  assign n48693 = n48334 ^ n48331 ;
  assign n48694 = ~n48350 & ~n48693 ;
  assign n48695 = n48694 ^ n48349 ;
  assign n48696 = n48695 ^ n48691 ;
  assign n48697 = n48692 & ~n48696 ;
  assign n48699 = n48698 ^ n48697 ;
  assign n48700 = ~n48687 & n48699 ;
  assign n48701 = n48700 ^ n48686 ;
  assign n48702 = n48701 ^ n48678 ;
  assign n48703 = n48682 & ~n48702 ;
  assign n48705 = n48704 ^ n48703 ;
  assign n48706 = ~n48677 & ~n48705 ;
  assign n48708 = n48707 ^ n48706 ;
  assign n48709 = ~n48672 & n48708 ;
  assign n48710 = n48709 ^ n48671 ;
  assign n48711 = n48710 ^ n48665 ;
  assign n48712 = ~n48667 & n48711 ;
  assign n48713 = n48712 ^ n48666 ;
  assign n48714 = n48713 ^ n48660 ;
  assign n48715 = n48662 & n48714 ;
  assign n48716 = n48715 ^ n48661 ;
  assign n48717 = n48716 ^ n48655 ;
  assign n48718 = ~n48657 & n48717 ;
  assign n48720 = n48719 ^ n48718 ;
  assign n48721 = ~n48652 & ~n48720 ;
  assign n48723 = n48722 ^ n48721 ;
  assign n48724 = n48647 & ~n48723 ;
  assign n48727 = n48726 ^ n48724 ;
  assign n48990 = n48732 ^ n48727 ;
  assign n49822 = n48990 ^ n47710 ;
  assign n48583 = n48108 ^ n48025 ;
  assign n49823 = n49822 ^ n48583 ;
  assign n48359 = n47578 ^ n46608 ;
  assign n48360 = n48359 ^ n48259 ;
  assign n48808 = n46797 ^ n38539 ;
  assign n48809 = n48808 ^ n43362 ;
  assign n48810 = n48809 ^ n37046 ;
  assign n48581 = n48178 ^ n46891 ;
  assign n48582 = n48581 ^ n46171 ;
  assign n48584 = n48583 ^ n48582 ;
  assign n48475 = n48103 ^ n48031 ;
  assign n48473 = n47931 ^ n47486 ;
  assign n48474 = n48473 ^ n46745 ;
  assign n48476 = n48475 ^ n48474 ;
  assign n48565 = n48106 ^ n48029 ;
  assign n48566 = n48565 ^ n48475 ;
  assign n48567 = n48566 ^ n48565 ;
  assign n48366 = n48099 ^ n48040 ;
  assign n48364 = n47442 ^ n45941 ;
  assign n48365 = n48364 ^ n47830 ;
  assign n48367 = n48366 ^ n48365 ;
  assign n48370 = n48097 ^ n48043 ;
  assign n48469 = n48370 ^ n48366 ;
  assign n48368 = n47706 ^ n46537 ;
  assign n48369 = n48368 ^ n47420 ;
  assign n48371 = n48370 ^ n48369 ;
  assign n48374 = n48094 ^ n48049 ;
  assign n48372 = n47710 ^ n47386 ;
  assign n48373 = n48372 ^ n46542 ;
  assign n48375 = n48374 ^ n48373 ;
  assign n48377 = n47716 ^ n47113 ;
  assign n48378 = n48377 ^ n46547 ;
  assign n48376 = n48091 ^ n48056 ;
  assign n48379 = n48378 ^ n48376 ;
  assign n48459 = n48458 ^ n48383 ;
  assign n48460 = n48385 & ~n48459 ;
  assign n48461 = n48460 ^ n48384 ;
  assign n48462 = n48461 ^ n48376 ;
  assign n48463 = ~n48379 & n48462 ;
  assign n48380 = n48376 ^ n48373 ;
  assign n48464 = n48463 ^ n48380 ;
  assign n48465 = ~n48375 & ~n48464 ;
  assign n48466 = n48465 ^ n48374 ;
  assign n48467 = n48466 ^ n48369 ;
  assign n48468 = n48371 & n48467 ;
  assign n48470 = n48469 ^ n48468 ;
  assign n48471 = ~n48367 & ~n48470 ;
  assign n48472 = n48471 ^ n48366 ;
  assign n48568 = n48567 ^ n48472 ;
  assign n48569 = n48476 & n48568 ;
  assign n48570 = n48569 ^ n48566 ;
  assign n48571 = n48143 ^ n46862 ;
  assign n48572 = n48571 ^ n47528 ;
  assign n48578 = n48572 ^ n48565 ;
  assign n48579 = ~n48570 & ~n48578 ;
  assign n48580 = n48579 ^ n48572 ;
  assign n48585 = n48584 ^ n48580 ;
  assign n48477 = n48476 ^ n48472 ;
  assign n48478 = n48477 ^ n46035 ;
  assign n48545 = n48464 ^ n48374 ;
  assign n48540 = n48461 ^ n48379 ;
  assign n48536 = n48535 ^ n48480 ;
  assign n48537 = n48535 ^ n46000 ;
  assign n48538 = n48536 & n48537 ;
  assign n48539 = n48538 ^ n46000 ;
  assign n48541 = n48540 ^ n48539 ;
  assign n48542 = n48540 ^ n46002 ;
  assign n48543 = ~n48541 & ~n48542 ;
  assign n48544 = n48543 ^ n46002 ;
  assign n48546 = n48545 ^ n48544 ;
  assign n48547 = n48545 ^ n46013 ;
  assign n48548 = n48546 & ~n48547 ;
  assign n48549 = n48548 ^ n46013 ;
  assign n48479 = n48466 ^ n48371 ;
  assign n48550 = n48549 ^ n48479 ;
  assign n48551 = n48470 ^ n48365 ;
  assign n48552 = n48551 ^ n46021 ;
  assign n48553 = n48552 ^ n48479 ;
  assign n48554 = n48553 ^ n48551 ;
  assign n48555 = n48550 & n48554 ;
  assign n48556 = n48555 ^ n48552 ;
  assign n48558 = n48477 ^ n46029 ;
  assign n48557 = n48551 ^ n48477 ;
  assign n48559 = n48558 ^ n48557 ;
  assign n48560 = ~n48556 & n48559 ;
  assign n48561 = n48560 ^ n48558 ;
  assign n48562 = ~n48478 & ~n48561 ;
  assign n48563 = n48562 ^ n46035 ;
  assign n48564 = n48563 ^ n45296 ;
  assign n48573 = n48572 ^ n48570 ;
  assign n48574 = n48573 ^ n48563 ;
  assign n48575 = n48564 & ~n48574 ;
  assign n48576 = n48575 ^ n45296 ;
  assign n48577 = n48576 ^ n45470 ;
  assign n48586 = n48585 ^ n48577 ;
  assign n48587 = n48573 ^ n48564 ;
  assign n48588 = n48561 ^ n46035 ;
  assign n48589 = n48556 ^ n46029 ;
  assign n48590 = n48547 ^ n48544 ;
  assign n48615 = n48592 & ~n48614 ;
  assign n48616 = n48539 ^ n46002 ;
  assign n48617 = n48616 ^ n48540 ;
  assign n48618 = n48615 & n48617 ;
  assign n48619 = ~n48590 & n48618 ;
  assign n48620 = n48479 ^ n46021 ;
  assign n48621 = n48620 ^ n48549 ;
  assign n48622 = ~n48619 & ~n48621 ;
  assign n48623 = n48589 & n48622 ;
  assign n48624 = n48588 & ~n48623 ;
  assign n48625 = n48587 & n48624 ;
  assign n48780 = n48586 & ~n48625 ;
  assign n48775 = n48111 ^ n48020 ;
  assign n48776 = n48775 ^ n48583 ;
  assign n48773 = n48583 ^ n48580 ;
  assign n48774 = n48584 & n48773 ;
  assign n48777 = n48776 ^ n48774 ;
  assign n48771 = n46894 ^ n46177 ;
  assign n48772 = n48771 ^ n48228 ;
  assign n48778 = n48777 ^ n48772 ;
  assign n48767 = n48585 ^ n48576 ;
  assign n48768 = ~n48577 & ~n48767 ;
  assign n48769 = n48768 ^ n45470 ;
  assign n48770 = n48769 ^ n45473 ;
  assign n48779 = n48778 ^ n48770 ;
  assign n48781 = n48780 ^ n48779 ;
  assign n48626 = n48625 ^ n48586 ;
  assign n48361 = n46803 ^ n38548 ;
  assign n48362 = n48361 ^ n1333 ;
  assign n48363 = n48362 ^ n2798 ;
  assign n48627 = n48626 ^ n48363 ;
  assign n48628 = n48624 ^ n48587 ;
  assign n1288 = n1278 ^ n1221 ;
  assign n1316 = n1315 ^ n1288 ;
  assign n1323 = n1322 ^ n1316 ;
  assign n48629 = n48628 ^ n1323 ;
  assign n48633 = n48623 ^ n48588 ;
  assign n48630 = n46811 ^ n1135 ;
  assign n48631 = n48630 ^ n43381 ;
  assign n48632 = n48631 ^ n1307 ;
  assign n48634 = n48633 ^ n48632 ;
  assign n48636 = n48622 ^ n48589 ;
  assign n1680 = n1679 ^ n1117 ;
  assign n1696 = n1695 ^ n1680 ;
  assign n1700 = n1699 ^ n1696 ;
  assign n48637 = n48636 ^ n1700 ;
  assign n48747 = n48621 ^ n48619 ;
  assign n48639 = n46516 ^ n1653 ;
  assign n48640 = n48639 ^ n43029 ;
  assign n48641 = n48640 ^ n37071 ;
  assign n48638 = n48618 ^ n48590 ;
  assign n48642 = n48641 ^ n48638 ;
  assign n48728 = n48617 ^ n48615 ;
  assign n48733 = n48732 ^ n48728 ;
  assign n48729 = n48728 ^ n48725 ;
  assign n48734 = n48733 ^ n48729 ;
  assign n48735 = ~n48727 & ~n48734 ;
  assign n48736 = n48735 ^ n48729 ;
  assign n48738 = n45945 ^ n38566 ;
  assign n48739 = n48738 ^ n2993 ;
  assign n48740 = n48739 ^ n37067 ;
  assign n48741 = n48740 ^ n48638 ;
  assign n48737 = n48728 ^ n48638 ;
  assign n48742 = n48741 ^ n48737 ;
  assign n48743 = ~n48736 & n48742 ;
  assign n48744 = n48743 ^ n48737 ;
  assign n48745 = ~n48642 & n48744 ;
  assign n48746 = n48745 ^ n48641 ;
  assign n48748 = n48747 ^ n48746 ;
  assign n48749 = n46824 ^ n38559 ;
  assign n48750 = n48749 ^ n43387 ;
  assign n48751 = n48750 ^ n1690 ;
  assign n48754 = n48751 ^ n48746 ;
  assign n48755 = n48748 & n48754 ;
  assign n48752 = n48751 ^ n1700 ;
  assign n48756 = n48755 ^ n48752 ;
  assign n48757 = ~n48637 & n48756 ;
  assign n48635 = n48633 ^ n1700 ;
  assign n48758 = n48757 ^ n48635 ;
  assign n48759 = ~n48634 & ~n48758 ;
  assign n48760 = n48759 ^ n48633 ;
  assign n48761 = n48760 ^ n1323 ;
  assign n48762 = n48629 & n48761 ;
  assign n48763 = n48762 ^ n48628 ;
  assign n48764 = n48763 ^ n48363 ;
  assign n48765 = n48627 & ~n48764 ;
  assign n48766 = n48765 ^ n48626 ;
  assign n48782 = n48781 ^ n48766 ;
  assign n48800 = n38544 ^ n1400 ;
  assign n48801 = n48800 ^ n43371 ;
  assign n48802 = n48801 ^ n37055 ;
  assign n49603 = n48802 ^ n48766 ;
  assign n48806 = ~n48782 & n49603 ;
  assign n48793 = n48778 ^ n45473 ;
  assign n48794 = n48778 ^ n48769 ;
  assign n48795 = n48793 & n48794 ;
  assign n48796 = n48795 ^ n45473 ;
  assign n48797 = n48796 ^ n45464 ;
  assign n48790 = n46882 ^ n46167 ;
  assign n48791 = n48790 ^ n47399 ;
  assign n48784 = n48115 ^ n48014 ;
  assign n48785 = n48784 ^ n48775 ;
  assign n48786 = n48785 ^ n48772 ;
  assign n48787 = n48786 ^ n48784 ;
  assign n48788 = n48777 & n48787 ;
  assign n48789 = n48788 ^ n48785 ;
  assign n48792 = n48791 ^ n48789 ;
  assign n48798 = n48797 ^ n48792 ;
  assign n48783 = ~n48779 & ~n48780 ;
  assign n48799 = n48798 ^ n48783 ;
  assign n48803 = n48802 ^ n48799 ;
  assign n48807 = n48806 ^ n48803 ;
  assign n48811 = n48810 ^ n48807 ;
  assign n48846 = n48360 & ~n48811 ;
  assign n48844 = n47596 ^ n46604 ;
  assign n48845 = n48844 ^ n48274 ;
  assign n48847 = n48846 ^ n48845 ;
  assign n48838 = n46880 ^ n46163 ;
  assign n48839 = n48838 ^ n47428 ;
  assign n48835 = n48117 ^ n48013 ;
  assign n48836 = n48835 ^ n48784 ;
  assign n48833 = n48791 ^ n48784 ;
  assign n48834 = n48789 & n48833 ;
  assign n48837 = n48836 ^ n48834 ;
  assign n48840 = n48839 ^ n48837 ;
  assign n48829 = n48796 ^ n48792 ;
  assign n48830 = n48797 & ~n48829 ;
  assign n48831 = n48830 ^ n45464 ;
  assign n48832 = n48831 ^ n45460 ;
  assign n48841 = n48840 ^ n48832 ;
  assign n48828 = ~n48783 & ~n48798 ;
  assign n48842 = n48841 ^ n48828 ;
  assign n48823 = n46792 ^ n38746 ;
  assign n48824 = n48823 ^ n43415 ;
  assign n48825 = n48824 ^ n37050 ;
  assign n48826 = n48825 ^ n48799 ;
  assign n48821 = n48810 ^ n48799 ;
  assign n48822 = ~n48807 & ~n48821 ;
  assign n48827 = n48826 ^ n48822 ;
  assign n48843 = n48842 ^ n48827 ;
  assign n48848 = n48847 ^ n48843 ;
  assign n48812 = n48811 ^ n48360 ;
  assign n48819 = ~n45990 & ~n48812 ;
  assign n48820 = n48819 ^ n45986 ;
  assign n48849 = n48848 ^ n48820 ;
  assign n48886 = n46786 ^ n38763 ;
  assign n48887 = n48886 ^ n43357 ;
  assign n48888 = n48887 ^ n37392 ;
  assign n48882 = ~n48828 & n48841 ;
  assign n48867 = n48840 ^ n48831 ;
  assign n48873 = n48120 ^ n48006 ;
  assign n48871 = n46876 ^ n46159 ;
  assign n48872 = n48871 ^ n47458 ;
  assign n48874 = n48873 ^ n48872 ;
  assign n48868 = n48839 ^ n48835 ;
  assign n48869 = ~n48837 & n48868 ;
  assign n48870 = n48869 ^ n48835 ;
  assign n48875 = n48874 ^ n48870 ;
  assign n48876 = n48875 ^ n45460 ;
  assign n48877 = n48876 ^ n48875 ;
  assign n48878 = n48877 ^ n48831 ;
  assign n48879 = ~n48867 & n48878 ;
  assign n48880 = n48879 ^ n48876 ;
  assign n48881 = n48880 ^ n45456 ;
  assign n48883 = n48882 ^ n48881 ;
  assign n48884 = n48883 ^ n48825 ;
  assign n48865 = n48842 ^ n48825 ;
  assign n48866 = ~n48827 & ~n48865 ;
  assign n48885 = n48884 ^ n48866 ;
  assign n48889 = n48888 ^ n48885 ;
  assign n48863 = n48341 ^ n46596 ;
  assign n48864 = n48863 ^ n47685 ;
  assign n48890 = n48889 ^ n48864 ;
  assign n48860 = n48845 ^ n48843 ;
  assign n48861 = ~n48847 & ~n48860 ;
  assign n48862 = n48861 ^ n48845 ;
  assign n48891 = n48890 ^ n48862 ;
  assign n48855 = n48848 ^ n48819 ;
  assign n48856 = n48848 ^ n45986 ;
  assign n48857 = n48855 & n48856 ;
  assign n48858 = n48857 ^ n45986 ;
  assign n48859 = n48858 ^ n45982 ;
  assign n48892 = n48891 ^ n48859 ;
  assign n48903 = ~n48849 & ~n48892 ;
  assign n48933 = n46781 ^ n38812 ;
  assign n48934 = n48933 ^ n43353 ;
  assign n48935 = n48934 ^ n37387 ;
  assign n48931 = ~n48881 & n48882 ;
  assign n48927 = n48875 ^ n45456 ;
  assign n48928 = ~n48880 & ~n48927 ;
  assign n48929 = n48928 ^ n45456 ;
  assign n48923 = n46616 ^ n45994 ;
  assign n48924 = n48923 ^ n47502 ;
  assign n48917 = n48123 ^ n48000 ;
  assign n48918 = n48917 ^ n48873 ;
  assign n48919 = n48918 ^ n48917 ;
  assign n48920 = n48919 ^ n48870 ;
  assign n48921 = ~n48874 & ~n48920 ;
  assign n48922 = n48921 ^ n48918 ;
  assign n48925 = n48924 ^ n48922 ;
  assign n48926 = n48925 ^ n45339 ;
  assign n48930 = n48929 ^ n48926 ;
  assign n48932 = n48931 ^ n48930 ;
  assign n48936 = n48935 ^ n48932 ;
  assign n48914 = n48888 ^ n48883 ;
  assign n48915 = n48885 & ~n48914 ;
  assign n48916 = n48915 ^ n48888 ;
  assign n48937 = n48936 ^ n48916 ;
  assign n48912 = n47777 ^ n46594 ;
  assign n48913 = n48912 ^ n48419 ;
  assign n48938 = n48937 ^ n48913 ;
  assign n48909 = n48864 ^ n48862 ;
  assign n48910 = n48890 & ~n48909 ;
  assign n48911 = n48910 ^ n48889 ;
  assign n48939 = n48938 ^ n48911 ;
  assign n48904 = n48891 ^ n48858 ;
  assign n48905 = n48891 ^ n45982 ;
  assign n48906 = ~n48904 & ~n48905 ;
  assign n48907 = n48906 ^ n45982 ;
  assign n48908 = n48907 ^ n45978 ;
  assign n48940 = n48939 ^ n48908 ;
  assign n49336 = ~n48903 & ~n48940 ;
  assign n49204 = n48939 ^ n48907 ;
  assign n49087 = n48913 ^ n48911 ;
  assign n49088 = n48938 & ~n49087 ;
  assign n49089 = n49088 ^ n48937 ;
  assign n49076 = n47542 ^ n46195 ;
  assign n49077 = n49076 ^ n46612 ;
  assign n49078 = n49077 ^ n48924 ;
  assign n48975 = n48126 ^ n47992 ;
  assign n49079 = n49078 ^ n48975 ;
  assign n49080 = n49079 ^ n45333 ;
  assign n49070 = n48929 ^ n48925 ;
  assign n49073 = n49070 ^ n48931 ;
  assign n49074 = n45339 & ~n49073 ;
  assign n49071 = n48931 ^ n48925 ;
  assign n49072 = ~n49070 & n49071 ;
  assign n49075 = n49074 ^ n49072 ;
  assign n49081 = n49080 ^ n49075 ;
  assign n49067 = n46777 ^ n38949 ;
  assign n49068 = n49067 ^ n43338 ;
  assign n49069 = n49068 ^ n37373 ;
  assign n49082 = n49081 ^ n49069 ;
  assign n49083 = n49082 ^ n48935 ;
  assign n49065 = n48924 ^ n48917 ;
  assign n49066 = n48922 & ~n49065 ;
  assign n49084 = n49083 ^ n49066 ;
  assign n49063 = n48935 ^ n48916 ;
  assign n49064 = ~n48936 & n49063 ;
  assign n49085 = n49084 ^ n49064 ;
  assign n49061 = n48415 ^ n46587 ;
  assign n49062 = n49061 ^ n47773 ;
  assign n49086 = n49085 ^ n49062 ;
  assign n49205 = n49089 ^ n49086 ;
  assign n49206 = n49205 ^ n45978 ;
  assign n49207 = n49206 ^ n49205 ;
  assign n49208 = n49207 ^ n48907 ;
  assign n49209 = n49204 & n49208 ;
  assign n49210 = n49209 ^ n49206 ;
  assign n49337 = n49210 ^ n45974 ;
  assign n49338 = ~n49336 & ~n49337 ;
  assign n49059 = n48312 ^ n48311 ;
  assign n49092 = n49085 ^ n49059 ;
  assign n49090 = n49089 ^ n49062 ;
  assign n49091 = ~n49086 & ~n49090 ;
  assign n49093 = n49092 ^ n49091 ;
  assign n49057 = n47771 ^ n46585 ;
  assign n49058 = n49057 ^ n48409 ;
  assign n49211 = n49093 ^ n49058 ;
  assign n49213 = n49211 ^ n45974 ;
  assign n49212 = n49211 ^ n49205 ;
  assign n49214 = n49213 ^ n49212 ;
  assign n49215 = ~n49210 & n49214 ;
  assign n49216 = n49215 ^ n49213 ;
  assign n49339 = n49216 ^ n45970 ;
  assign n49340 = ~n49338 & n49339 ;
  assign n49060 = n49059 ^ n49058 ;
  assign n49094 = n49060 & ~n49093 ;
  assign n49095 = n49094 ^ n49059 ;
  assign n49054 = n48308 ^ n48249 ;
  assign n49055 = n49054 ^ n48313 ;
  assign n49052 = n48407 ^ n46581 ;
  assign n49053 = n49052 ^ n47765 ;
  assign n49056 = n49055 ^ n49053 ;
  assign n49217 = n49095 ^ n49056 ;
  assign n49219 = n49217 ^ n45970 ;
  assign n49218 = n49217 ^ n49211 ;
  assign n49220 = n49219 ^ n49218 ;
  assign n49221 = ~n49216 & n49220 ;
  assign n49222 = n49221 ^ n49219 ;
  assign n49341 = n49222 ^ n45966 ;
  assign n49342 = ~n49340 & ~n49341 ;
  assign n49050 = n48317 ^ n48305 ;
  assign n49098 = n49055 ^ n49050 ;
  assign n49096 = n49095 ^ n49053 ;
  assign n49097 = ~n49056 & n49096 ;
  assign n49099 = n49098 ^ n49097 ;
  assign n49048 = n48403 ^ n47696 ;
  assign n49049 = n49048 ^ n46574 ;
  assign n49202 = n49099 ^ n49049 ;
  assign n49224 = n49202 ^ n45966 ;
  assign n49223 = n49217 ^ n49202 ;
  assign n49225 = n49224 ^ n49223 ;
  assign n49226 = ~n49222 & n49225 ;
  assign n49227 = n49226 ^ n49224 ;
  assign n49343 = n49227 ^ n45962 ;
  assign n49344 = n49342 & ~n49343 ;
  assign n49051 = n49050 ^ n49049 ;
  assign n49100 = ~n49051 & n49099 ;
  assign n49101 = n49100 ^ n49050 ;
  assign n49046 = n48320 ^ n48298 ;
  assign n49044 = n47757 ^ n46937 ;
  assign n49045 = n49044 ^ n48399 ;
  assign n49047 = n49046 ^ n49045 ;
  assign n49201 = n49101 ^ n49047 ;
  assign n49345 = n49201 ^ n45958 ;
  assign n49203 = n49202 ^ n45962 ;
  assign n49228 = n49203 & ~n49227 ;
  assign n49229 = n49228 ^ n45962 ;
  assign n49346 = n49345 ^ n49229 ;
  assign n49347 = n49344 & n49346 ;
  assign n49230 = n49229 ^ n49201 ;
  assign n49102 = n49101 ^ n49045 ;
  assign n49103 = n49047 & ~n49102 ;
  assign n49104 = n49103 ^ n49046 ;
  assign n49041 = n47753 ^ n46566 ;
  assign n49042 = n49041 ^ n47695 ;
  assign n48956 = n48323 ^ n48293 ;
  assign n49043 = n49042 ^ n48956 ;
  assign n49199 = n49104 ^ n49043 ;
  assign n49231 = n49199 ^ n45958 ;
  assign n49232 = n49231 ^ n49199 ;
  assign n49233 = n49232 ^ n49201 ;
  assign n49234 = n49230 & ~n49233 ;
  assign n49235 = n49234 ^ n49231 ;
  assign n49348 = n49235 ^ n45954 ;
  assign n49349 = ~n49347 & ~n49348 ;
  assign n49200 = n49199 ^ n45954 ;
  assign n49236 = ~n49200 & ~n49235 ;
  assign n49237 = n49236 ^ n45954 ;
  assign n49105 = n49104 ^ n49042 ;
  assign n49106 = ~n49043 & ~n49105 ;
  assign n49107 = n49106 ^ n48956 ;
  assign n49038 = n47749 ^ n46947 ;
  assign n49039 = n49038 ^ n48392 ;
  assign n48951 = n48326 ^ n48285 ;
  assign n49040 = n49039 ^ n48951 ;
  assign n49197 = n49107 ^ n49040 ;
  assign n49198 = n49197 ^ n45950 ;
  assign n49350 = n49237 ^ n49198 ;
  assign n49351 = n49349 & n49350 ;
  assign n48945 = n48329 ^ n48283 ;
  assign n49110 = n48951 ^ n48945 ;
  assign n49108 = n49107 ^ n48951 ;
  assign n49109 = ~n49040 & n49108 ;
  assign n49111 = n49110 ^ n49109 ;
  assign n49035 = n48451 ^ n47743 ;
  assign n49036 = n49035 ^ n46564 ;
  assign n49196 = n49111 ^ n49036 ;
  assign n49352 = n49196 ^ n46232 ;
  assign n49238 = n49237 ^ n49197 ;
  assign n49239 = ~n49198 & ~n49238 ;
  assign n49240 = n49239 ^ n45950 ;
  assign n49353 = n49352 ^ n49240 ;
  assign n49354 = n49351 & ~n49353 ;
  assign n49241 = n49240 ^ n49196 ;
  assign n49037 = n49036 ^ n48945 ;
  assign n49112 = ~n49037 & ~n49111 ;
  assign n49113 = n49112 ^ n49036 ;
  assign n49032 = n47739 ^ n46559 ;
  assign n49033 = n49032 ^ n48388 ;
  assign n48351 = n48350 ^ n48331 ;
  assign n49034 = n49033 ^ n48351 ;
  assign n49194 = n49113 ^ n49034 ;
  assign n49242 = n49194 ^ n46232 ;
  assign n49243 = n49242 ^ n49194 ;
  assign n49244 = n49243 ^ n49196 ;
  assign n49245 = n49241 & ~n49244 ;
  assign n49246 = n49245 ^ n49242 ;
  assign n49335 = n49246 ^ n46521 ;
  assign n49471 = n49354 ^ n49335 ;
  assign n49468 = n47247 ^ n39255 ;
  assign n49469 = n49468 ^ n43804 ;
  assign n49470 = n49469 ^ n37669 ;
  assign n49472 = n49471 ^ n49470 ;
  assign n49474 = n47253 ^ n39261 ;
  assign n49475 = n49474 ^ n43809 ;
  assign n49476 = n49475 ^ n37675 ;
  assign n49536 = n49476 ^ n49470 ;
  assign n49473 = n49353 ^ n49351 ;
  assign n49477 = n49476 ^ n49473 ;
  assign n49478 = n49350 ^ n49349 ;
  assign n2316 = n2315 ^ n2279 ;
  assign n2350 = n2349 ^ n2316 ;
  assign n2360 = n2359 ^ n2350 ;
  assign n49479 = n49478 ^ n2360 ;
  assign n49481 = n47261 ^ n39268 ;
  assign n49482 = n49481 ^ n43817 ;
  assign n49483 = n49482 ^ n2341 ;
  assign n49480 = n49348 ^ n49347 ;
  assign n49484 = n49483 ^ n49480 ;
  assign n49488 = n49346 ^ n49344 ;
  assign n49485 = n47265 ^ n2193 ;
  assign n49486 = n49485 ^ n43823 ;
  assign n49487 = n49486 ^ n37733 ;
  assign n49489 = n49488 ^ n49487 ;
  assign n49491 = n47271 ^ n39274 ;
  assign n49492 = n49491 ^ n43828 ;
  assign n49493 = n49492 ^ n37686 ;
  assign n49490 = n49343 ^ n49342 ;
  assign n49494 = n49493 ^ n49490 ;
  assign n49498 = n49341 ^ n49340 ;
  assign n49495 = n47276 ^ n39279 ;
  assign n49496 = n49495 ^ n43833 ;
  assign n49497 = n49496 ^ n37691 ;
  assign n49499 = n49498 ^ n49497 ;
  assign n49503 = n49339 ^ n49338 ;
  assign n49500 = n47281 ^ n39296 ;
  assign n49501 = n49500 ^ n43839 ;
  assign n49502 = n49501 ^ n37720 ;
  assign n49504 = n49503 ^ n49502 ;
  assign n49508 = n49337 ^ n49336 ;
  assign n49505 = n47285 ^ n39284 ;
  assign n49506 = n49505 ^ n43843 ;
  assign n49507 = n49506 ^ n37695 ;
  assign n49509 = n49508 ^ n49507 ;
  assign n48898 = n47290 ^ n38797 ;
  assign n48899 = n48898 ^ n43849 ;
  assign n48900 = n48899 ^ n37700 ;
  assign n48893 = n48892 ^ n48849 ;
  assign n48901 = n48900 ^ n48893 ;
  assign n48356 = n47535 ^ n39714 ;
  assign n48357 = n48356 ^ n44106 ;
  assign n48358 = n48357 ^ n38201 ;
  assign n48813 = n48812 ^ n45990 ;
  assign n48814 = n48358 & n48813 ;
  assign n48353 = n47296 ^ n3194 ;
  assign n48354 = n48353 ^ n43856 ;
  assign n48355 = n48354 ^ n37247 ;
  assign n48815 = n48814 ^ n48355 ;
  assign n48948 = n48849 ^ n48355 ;
  assign n48853 = ~n48815 & ~n48948 ;
  assign n48816 = n47300 ^ n38754 ;
  assign n48817 = n48816 ^ n43853 ;
  assign n48818 = n48817 ^ n37704 ;
  assign n48850 = n48849 ^ n48818 ;
  assign n48854 = n48853 ^ n48850 ;
  assign n48896 = n48893 ^ n48818 ;
  assign n48897 = n48854 & ~n48896 ;
  assign n48902 = n48901 ^ n48897 ;
  assign n48941 = n48940 ^ n48903 ;
  assign n49510 = n48941 ^ n48900 ;
  assign n49511 = ~n48902 & n49510 ;
  assign n49512 = n49511 ^ n48900 ;
  assign n49513 = n49512 ^ n49507 ;
  assign n49514 = ~n49509 & ~n49513 ;
  assign n49515 = n49514 ^ n49508 ;
  assign n49516 = n49515 ^ n49502 ;
  assign n49517 = ~n49504 & ~n49516 ;
  assign n49518 = n49517 ^ n49502 ;
  assign n49519 = n49518 ^ n49497 ;
  assign n49520 = ~n49499 & ~n49519 ;
  assign n49521 = n49520 ^ n49498 ;
  assign n49522 = n49521 ^ n49490 ;
  assign n49523 = n49494 & n49522 ;
  assign n49524 = n49523 ^ n49493 ;
  assign n49525 = n49524 ^ n49487 ;
  assign n49526 = ~n49489 & ~n49525 ;
  assign n49527 = n49526 ^ n49488 ;
  assign n49528 = n49527 ^ n49480 ;
  assign n49529 = n49484 & n49528 ;
  assign n49530 = n49529 ^ n49483 ;
  assign n49531 = n49530 ^ n2360 ;
  assign n49532 = n49479 & ~n49531 ;
  assign n49533 = n49532 ^ n49478 ;
  assign n49534 = n49533 ^ n49473 ;
  assign n49535 = ~n49477 & n49534 ;
  assign n49537 = n49536 ^ n49535 ;
  assign n49538 = n49472 & ~n49537 ;
  assign n49539 = n49538 ^ n49471 ;
  assign n49355 = n49335 & n49354 ;
  assign n49114 = n49113 ^ n49033 ;
  assign n49115 = n49034 & ~n49114 ;
  assign n49116 = n49115 ^ n48351 ;
  assign n49029 = n48384 ^ n46554 ;
  assign n49030 = n49029 ^ n47734 ;
  assign n49028 = n48695 ^ n48692 ;
  assign n49031 = n49030 ^ n49028 ;
  assign n49193 = n49116 ^ n49031 ;
  assign n49333 = n49193 ^ n46648 ;
  assign n49195 = n49194 ^ n46521 ;
  assign n49247 = n49195 & n49246 ;
  assign n49248 = n49247 ^ n46521 ;
  assign n49334 = n49333 ^ n49248 ;
  assign n49466 = n49355 ^ n49334 ;
  assign n49463 = n47243 ^ n39251 ;
  assign n49464 = n49463 ^ n43799 ;
  assign n49465 = n49464 ^ n37665 ;
  assign n49467 = n49466 ^ n49465 ;
  assign n49821 = n49539 ^ n49467 ;
  assign n49824 = n49823 ^ n49821 ;
  assign n48998 = n48720 ^ n48650 ;
  assign n49825 = n48998 ^ n48475 ;
  assign n49826 = n49825 ^ n47718 ;
  assign n49803 = n49533 ^ n49477 ;
  assign n49827 = n49826 ^ n49803 ;
  assign n49002 = n48716 ^ n48657 ;
  assign n49830 = n49002 ^ n47724 ;
  assign n49831 = n49830 ^ n48366 ;
  assign n49829 = n49530 ^ n49479 ;
  assign n49832 = n49831 ^ n49829 ;
  assign n49835 = n49524 ^ n49489 ;
  assign n49833 = n48374 ^ n47734 ;
  assign n49006 = n48710 ^ n48667 ;
  assign n49834 = n49833 ^ n49006 ;
  assign n49836 = n49835 ^ n49834 ;
  assign n49842 = n49521 ^ n49494 ;
  assign n49012 = n48708 ^ n48670 ;
  assign n49840 = n49012 ^ n48376 ;
  assign n49841 = n49840 ^ n47739 ;
  assign n49843 = n49842 ^ n49841 ;
  assign n49846 = n49518 ^ n49499 ;
  assign n49844 = n48384 ^ n47743 ;
  assign n49016 = n48705 ^ n48676 ;
  assign n49845 = n49844 ^ n49016 ;
  assign n49847 = n49846 ^ n49845 ;
  assign n49022 = n48701 ^ n48682 ;
  assign n49849 = n49022 ^ n48388 ;
  assign n49850 = n49849 ^ n47749 ;
  assign n49848 = n49515 ^ n49504 ;
  assign n49851 = n49850 ^ n49848 ;
  assign n48894 = n48893 ^ n48854 ;
  assign n47697 = n47696 ^ n47695 ;
  assign n48352 = n48351 ^ n47697 ;
  assign n48895 = n48894 ^ n48352 ;
  assign n48949 = n48948 ^ n48814 ;
  assign n48946 = n48945 ^ n47765 ;
  assign n48947 = n48946 ^ n48399 ;
  assign n48950 = n48949 ^ n48947 ;
  assign n48954 = n48813 ^ n48358 ;
  assign n48952 = n48951 ^ n48403 ;
  assign n48953 = n48952 ^ n47771 ;
  assign n48955 = n48954 ^ n48953 ;
  assign n48969 = n48756 ^ n48636 ;
  assign n48967 = n48162 ^ n46882 ;
  assign n48968 = n48967 ^ n47458 ;
  assign n48970 = n48969 ^ n48968 ;
  assign n48977 = n48751 ^ n48747 ;
  assign n48978 = n48977 ^ n48746 ;
  assign n48974 = n47428 ^ n46894 ;
  assign n48976 = n48975 ^ n48974 ;
  assign n48979 = n48978 ^ n48976 ;
  assign n48981 = n48917 ^ n46891 ;
  assign n48982 = n48981 ^ n47399 ;
  assign n48980 = n48744 ^ n48641 ;
  assign n48983 = n48982 ^ n48980 ;
  assign n48985 = n48873 ^ n48228 ;
  assign n48986 = n48985 ^ n47528 ;
  assign n48984 = n48740 ^ n48736 ;
  assign n48987 = n48986 ^ n48984 ;
  assign n48991 = n48835 ^ n48178 ;
  assign n48992 = n48991 ^ n47486 ;
  assign n48993 = n48992 ^ n48990 ;
  assign n48994 = n48723 ^ n48645 ;
  assign n49148 = n48994 ^ n48992 ;
  assign n48995 = n48784 ^ n47442 ;
  assign n48996 = n48995 ^ n48143 ;
  assign n48997 = n48996 ^ n48994 ;
  assign n48999 = n47931 ^ n47420 ;
  assign n49000 = n48999 ^ n48775 ;
  assign n49001 = n49000 ^ n48998 ;
  assign n49003 = n48583 ^ n47830 ;
  assign n49004 = n49003 ^ n47386 ;
  assign n49005 = n49004 ^ n49002 ;
  assign n49007 = n48713 ^ n48662 ;
  assign n49139 = n49007 ^ n49002 ;
  assign n49009 = n47710 ^ n46974 ;
  assign n49010 = n49009 ^ n48475 ;
  assign n49011 = n49010 ^ n49006 ;
  assign n49013 = n48366 ^ n47716 ;
  assign n49014 = n49013 ^ n46534 ;
  assign n49015 = n49014 ^ n49012 ;
  assign n49017 = n48370 ^ n46539 ;
  assign n49018 = n49017 ^ n47718 ;
  assign n49019 = n49018 ^ n49016 ;
  assign n49020 = n48374 ^ n46544 ;
  assign n49021 = n49020 ^ n47724 ;
  assign n49023 = n49022 ^ n49021 ;
  assign n49026 = n48699 ^ n48683 ;
  assign n49024 = n48376 ^ n47730 ;
  assign n49025 = n49024 ^ n46549 ;
  assign n49027 = n49026 ^ n49025 ;
  assign n49119 = n49028 ^ n49025 ;
  assign n49117 = n49116 ^ n49028 ;
  assign n49118 = n49031 & n49117 ;
  assign n49120 = n49119 ^ n49118 ;
  assign n49121 = ~n49027 & n49120 ;
  assign n49122 = n49121 ^ n49026 ;
  assign n49123 = n49122 ^ n49021 ;
  assign n49124 = n49023 & n49123 ;
  assign n49125 = n49124 ^ n49022 ;
  assign n49126 = n49125 ^ n49016 ;
  assign n49127 = ~n49019 & n49126 ;
  assign n49128 = n49127 ^ n49018 ;
  assign n49129 = n49128 ^ n49012 ;
  assign n49130 = ~n49015 & ~n49129 ;
  assign n49131 = n49130 ^ n49014 ;
  assign n49132 = n49131 ^ n49006 ;
  assign n49133 = n49011 & ~n49132 ;
  assign n49008 = n49007 ^ n49006 ;
  assign n49134 = n49133 ^ n49008 ;
  assign n49135 = n47706 ^ n47113 ;
  assign n49136 = n49135 ^ n48565 ;
  assign n49137 = n49136 ^ n49007 ;
  assign n49138 = ~n49134 & ~n49137 ;
  assign n49140 = n49139 ^ n49138 ;
  assign n49141 = ~n49005 & ~n49140 ;
  assign n49142 = n49141 ^ n49004 ;
  assign n49143 = n49142 ^ n48998 ;
  assign n49144 = n49001 & n49143 ;
  assign n49145 = n49144 ^ n49000 ;
  assign n49146 = n49145 ^ n48994 ;
  assign n49147 = ~n48997 & n49146 ;
  assign n49149 = n49148 ^ n49147 ;
  assign n49150 = ~n48993 & ~n49149 ;
  assign n49151 = n49150 ^ n48992 ;
  assign n49152 = n49151 ^ n48984 ;
  assign n49153 = n48987 & ~n49152 ;
  assign n48988 = n48984 ^ n48982 ;
  assign n49154 = n49153 ^ n48988 ;
  assign n49155 = n48983 & n49154 ;
  assign n49156 = n49155 ^ n48982 ;
  assign n49157 = n49156 ^ n48976 ;
  assign n49158 = n48979 & ~n49157 ;
  assign n49159 = n49158 ^ n48978 ;
  assign n48971 = n48758 ^ n48632 ;
  assign n48972 = n48971 ^ n48969 ;
  assign n48973 = n48972 ^ n48971 ;
  assign n49160 = n49159 ^ n48973 ;
  assign n49161 = ~n48970 & n49160 ;
  assign n49162 = n49161 ^ n48972 ;
  assign n49164 = n47502 ^ n46880 ;
  assign n49165 = n49164 ^ n48165 ;
  assign n48965 = n48760 ^ n48629 ;
  assign n49166 = n49165 ^ n48965 ;
  assign n49163 = n48971 ^ n48965 ;
  assign n49167 = n49166 ^ n49163 ;
  assign n49168 = n49162 & n49167 ;
  assign n49169 = n49168 ^ n49163 ;
  assign n48963 = n48155 ^ n46876 ;
  assign n48964 = n48963 ^ n47542 ;
  assign n49174 = n49169 ^ n48964 ;
  assign n49175 = n49174 ^ n46159 ;
  assign n49176 = n49165 ^ n49162 ;
  assign n49177 = n49176 ^ n46163 ;
  assign n49306 = n49159 ^ n48970 ;
  assign n49179 = n49154 ^ n48980 ;
  assign n49180 = n49179 ^ n46171 ;
  assign n49181 = n49151 ^ n48987 ;
  assign n49182 = n49181 ^ n46862 ;
  assign n49286 = n49145 ^ n48997 ;
  assign n49184 = n49142 ^ n49001 ;
  assign n49185 = n49184 ^ n46537 ;
  assign n49278 = n49140 ^ n49004 ;
  assign n49186 = n49136 ^ n49134 ;
  assign n49187 = n49186 ^ n46547 ;
  assign n49269 = n49131 ^ n49011 ;
  assign n49188 = n49128 ^ n49015 ;
  assign n49189 = n49188 ^ n46557 ;
  assign n49191 = n49122 ^ n49023 ;
  assign n49192 = n49191 ^ n46572 ;
  assign n49253 = n49120 ^ n49026 ;
  assign n49249 = n49248 ^ n49193 ;
  assign n49250 = n49248 ^ n46648 ;
  assign n49251 = ~n49249 & ~n49250 ;
  assign n49252 = n49251 ^ n46648 ;
  assign n49254 = n49253 ^ n49252 ;
  assign n49255 = n49191 ^ n46568 ;
  assign n49256 = n49255 ^ n49191 ;
  assign n49257 = n49256 ^ n49252 ;
  assign n49258 = ~n49254 & n49257 ;
  assign n49259 = n49258 ^ n49255 ;
  assign n49260 = n49192 & n49259 ;
  assign n49261 = n49260 ^ n46572 ;
  assign n49190 = n49125 ^ n49019 ;
  assign n49262 = n49261 ^ n49190 ;
  assign n49263 = n49261 ^ n46562 ;
  assign n49264 = ~n49262 & n49263 ;
  assign n49265 = n49264 ^ n46562 ;
  assign n49266 = n49265 ^ n49188 ;
  assign n49267 = ~n49189 & ~n49266 ;
  assign n49268 = n49267 ^ n46557 ;
  assign n49270 = n49269 ^ n49268 ;
  assign n49271 = n49186 ^ n46552 ;
  assign n49272 = n49271 ^ n49186 ;
  assign n49273 = n49272 ^ n49268 ;
  assign n49274 = n49270 & n49273 ;
  assign n49275 = n49274 ^ n49271 ;
  assign n49276 = ~n49187 & n49275 ;
  assign n49277 = n49276 ^ n46547 ;
  assign n49279 = n49278 ^ n49277 ;
  assign n49280 = n49278 ^ n46542 ;
  assign n49281 = ~n49279 & ~n49280 ;
  assign n49282 = n49281 ^ n46542 ;
  assign n49283 = n49282 ^ n49184 ;
  assign n49284 = ~n49185 & n49283 ;
  assign n49285 = n49284 ^ n46537 ;
  assign n49287 = n49286 ^ n49285 ;
  assign n49288 = n49286 ^ n45941 ;
  assign n49289 = n49287 & ~n49288 ;
  assign n49290 = n49289 ^ n45941 ;
  assign n49183 = n49149 ^ n48990 ;
  assign n49291 = n49290 ^ n49183 ;
  assign n49292 = n49181 ^ n46745 ;
  assign n49293 = n49292 ^ n49181 ;
  assign n49294 = n49293 ^ n49183 ;
  assign n49295 = n49291 & n49294 ;
  assign n49296 = n49295 ^ n49292 ;
  assign n49297 = ~n49182 & ~n49296 ;
  assign n49298 = n49297 ^ n46862 ;
  assign n49299 = n49298 ^ n49179 ;
  assign n49300 = ~n49180 & ~n49299 ;
  assign n49301 = n49300 ^ n46171 ;
  assign n49178 = n49156 ^ n48979 ;
  assign n49302 = n49301 ^ n49178 ;
  assign n49303 = n49301 ^ n46177 ;
  assign n49304 = n49302 & n49303 ;
  assign n49305 = n49304 ^ n46177 ;
  assign n49307 = n49306 ^ n49305 ;
  assign n49308 = n49176 ^ n46167 ;
  assign n49309 = n49308 ^ n49176 ;
  assign n49310 = n49309 ^ n49305 ;
  assign n49311 = ~n49307 & ~n49310 ;
  assign n49312 = n49311 ^ n49308 ;
  assign n49313 = n49177 & ~n49312 ;
  assign n49314 = n49313 ^ n46163 ;
  assign n49315 = n49314 ^ n49174 ;
  assign n49316 = ~n49175 & ~n49315 ;
  assign n49317 = n49316 ^ n46159 ;
  assign n48966 = n48965 ^ n48964 ;
  assign n49170 = n48966 & n49169 ;
  assign n49171 = n49170 ^ n48965 ;
  assign n48961 = n48763 ^ n48627 ;
  assign n48959 = n47549 ^ n46616 ;
  assign n48960 = n48959 ^ n48197 ;
  assign n48962 = n48961 ^ n48960 ;
  assign n49172 = n49171 ^ n48962 ;
  assign n49173 = n49172 ^ n45994 ;
  assign n49318 = n49317 ^ n49173 ;
  assign n49319 = n49314 ^ n49175 ;
  assign n49320 = n49306 ^ n46167 ;
  assign n49321 = n49320 ^ n49305 ;
  assign n49322 = n49178 ^ n46177 ;
  assign n49323 = n49322 ^ n49301 ;
  assign n49324 = n49183 ^ n46745 ;
  assign n49325 = n49324 ^ n49290 ;
  assign n49326 = n49288 ^ n49285 ;
  assign n49327 = n49265 ^ n49189 ;
  assign n49328 = n49190 ^ n46562 ;
  assign n49329 = n49328 ^ n49261 ;
  assign n49330 = n49259 ^ n46572 ;
  assign n49331 = n49253 ^ n46568 ;
  assign n49332 = n49331 ^ n49252 ;
  assign n49356 = n49334 & n49355 ;
  assign n49357 = ~n49332 & ~n49356 ;
  assign n49358 = ~n49330 & n49357 ;
  assign n49359 = ~n49329 & ~n49358 ;
  assign n49360 = ~n49327 & ~n49359 ;
  assign n49361 = n49268 ^ n46552 ;
  assign n49362 = n49361 ^ n49269 ;
  assign n49363 = ~n49360 & ~n49362 ;
  assign n49364 = n49275 ^ n46547 ;
  assign n49365 = n49363 & ~n49364 ;
  assign n49366 = n49280 ^ n49277 ;
  assign n49367 = n49365 & ~n49366 ;
  assign n49368 = n49282 ^ n49185 ;
  assign n49369 = ~n49367 & ~n49368 ;
  assign n49370 = ~n49326 & n49369 ;
  assign n49371 = ~n49325 & ~n49370 ;
  assign n49372 = n49296 ^ n46862 ;
  assign n49373 = n49371 & ~n49372 ;
  assign n49374 = n49298 ^ n49180 ;
  assign n49375 = ~n49373 & ~n49374 ;
  assign n49376 = ~n49323 & ~n49375 ;
  assign n49377 = n49321 & ~n49376 ;
  assign n49378 = n49312 ^ n46163 ;
  assign n49379 = ~n49377 & ~n49378 ;
  assign n49380 = n49319 & n49379 ;
  assign n49615 = ~n49318 & ~n49380 ;
  assign n49608 = n48960 ^ n46195 ;
  assign n49605 = n47568 ^ n46612 ;
  assign n49606 = n49605 ^ n48238 ;
  assign n49604 = n49603 ^ n48781 ;
  assign n49607 = n49606 ^ n49604 ;
  assign n49609 = n49608 ^ n49607 ;
  assign n49610 = n49609 ^ n45994 ;
  assign n49600 = n47501 ^ n39660 ;
  assign n49601 = n49600 ^ n44086 ;
  assign n49602 = n49601 ^ n2660 ;
  assign n49611 = n49610 ^ n49602 ;
  assign n49382 = n47456 ^ n39593 ;
  assign n49383 = n49382 ^ n44009 ;
  assign n49384 = n49383 ^ n38064 ;
  assign n49612 = n49611 ^ n49384 ;
  assign n49597 = n49171 ^ n48960 ;
  assign n49598 = n49171 ^ n48961 ;
  assign n49599 = n49597 & n49598 ;
  assign n49613 = n49612 ^ n49599 ;
  assign n49594 = n49317 ^ n49172 ;
  assign n49595 = n49317 ^ n45994 ;
  assign n49596 = ~n49594 & n49595 ;
  assign n49614 = n49613 ^ n49596 ;
  assign n49616 = n49615 ^ n49614 ;
  assign n49381 = n49380 ^ n49318 ;
  assign n49385 = n49384 ^ n49381 ;
  assign n49389 = n49379 ^ n49319 ;
  assign n49386 = n47410 ^ n39597 ;
  assign n49387 = n49386 ^ n43942 ;
  assign n49388 = n49387 ^ n38069 ;
  assign n49390 = n49389 ^ n49388 ;
  assign n49392 = n47397 ^ n39603 ;
  assign n49393 = n49392 ^ n2903 ;
  assign n49394 = n49393 ^ n38073 ;
  assign n49588 = n49394 ^ n49389 ;
  assign n49391 = n49378 ^ n49377 ;
  assign n49395 = n49394 ^ n49391 ;
  assign n49399 = n49376 ^ n49321 ;
  assign n49396 = n44026 ^ n39609 ;
  assign n49397 = n49396 ^ n43738 ;
  assign n49398 = n49397 ^ n2895 ;
  assign n49400 = n49399 ^ n49398 ;
  assign n49404 = n49375 ^ n49323 ;
  assign n49401 = n47177 ^ n2813 ;
  assign n49402 = n49401 ^ n43743 ;
  assign n49403 = n49402 ^ n38083 ;
  assign n49405 = n49404 ^ n49403 ;
  assign n49406 = n47182 ^ n1436 ;
  assign n49407 = n49406 ^ n1774 ;
  assign n49408 = n49407 ^ n38088 ;
  assign n49579 = n49408 ^ n49403 ;
  assign n49409 = n49374 ^ n49373 ;
  assign n49410 = n49409 ^ n49408 ;
  assign n49411 = n49372 ^ n49371 ;
  assign n1750 = n1740 ^ n1421 ;
  assign n1760 = n1759 ^ n1750 ;
  assign n1767 = n1766 ^ n1760 ;
  assign n49412 = n49411 ^ n1767 ;
  assign n49416 = n49370 ^ n49325 ;
  assign n49413 = n47190 ^ n1720 ;
  assign n49414 = n49413 ^ n43751 ;
  assign n49415 = n49414 ^ n1757 ;
  assign n49417 = n49416 ^ n49415 ;
  assign n49421 = n49369 ^ n49326 ;
  assign n49418 = n47195 ^ n1711 ;
  assign n49419 = n49418 ^ n43757 ;
  assign n49420 = n49419 ^ n1004 ;
  assign n49422 = n49421 ^ n49420 ;
  assign n49426 = n49368 ^ n49367 ;
  assign n49423 = n47201 ^ n39212 ;
  assign n49424 = n49423 ^ n893 ;
  assign n49425 = n49424 ^ n38098 ;
  assign n49427 = n49426 ^ n49425 ;
  assign n49429 = n47205 ^ n39217 ;
  assign n49430 = n49429 ^ n43763 ;
  assign n49431 = n49430 ^ n885 ;
  assign n49564 = n49431 ^ n49425 ;
  assign n49428 = n49366 ^ n49365 ;
  assign n49432 = n49431 ^ n49428 ;
  assign n49434 = n47210 ^ n770 ;
  assign n49435 = n49434 ^ n43768 ;
  assign n49436 = n49435 ^ n37767 ;
  assign n49561 = n49436 ^ n49431 ;
  assign n49433 = n49364 ^ n49363 ;
  assign n49437 = n49436 ^ n49433 ;
  assign n49441 = n49362 ^ n49360 ;
  assign n49438 = n47216 ^ n39224 ;
  assign n49439 = n49438 ^ n43773 ;
  assign n49440 = n49439 ^ n1595 ;
  assign n49442 = n49441 ^ n49440 ;
  assign n49444 = n47222 ^ n39229 ;
  assign n49445 = n49444 ^ n43778 ;
  assign n49446 = n49445 ^ n37643 ;
  assign n49555 = n49446 ^ n49441 ;
  assign n49443 = n49359 ^ n49327 ;
  assign n49447 = n49446 ^ n49443 ;
  assign n49451 = n49358 ^ n49329 ;
  assign n49448 = n47228 ^ n39234 ;
  assign n49449 = n49448 ^ n43783 ;
  assign n49450 = n49449 ^ n37647 ;
  assign n49452 = n49451 ^ n49450 ;
  assign n49458 = n47233 ^ n39241 ;
  assign n49459 = n49458 ^ n43790 ;
  assign n49460 = n49459 ^ n37652 ;
  assign n49549 = n49460 ^ n49450 ;
  assign n49454 = n47238 ^ n39246 ;
  assign n49455 = n49454 ^ n43795 ;
  assign n49456 = n49455 ^ n37658 ;
  assign n49453 = n49356 ^ n49332 ;
  assign n49457 = n49456 ^ n49453 ;
  assign n49540 = n49539 ^ n49465 ;
  assign n49541 = n49467 & ~n49540 ;
  assign n49542 = n49541 ^ n49466 ;
  assign n49543 = n49542 ^ n49456 ;
  assign n49544 = ~n49457 & n49543 ;
  assign n49461 = n49460 ^ n49456 ;
  assign n49545 = n49544 ^ n49461 ;
  assign n49546 = n49357 ^ n49330 ;
  assign n49547 = n49546 ^ n49460 ;
  assign n49548 = n49545 & n49547 ;
  assign n49550 = n49549 ^ n49548 ;
  assign n49551 = n49452 & ~n49550 ;
  assign n49552 = n49551 ^ n49451 ;
  assign n49553 = n49552 ^ n49446 ;
  assign n49554 = ~n49447 & n49553 ;
  assign n49556 = n49555 ^ n49554 ;
  assign n49557 = n49442 & n49556 ;
  assign n49558 = n49557 ^ n49441 ;
  assign n49559 = n49558 ^ n49433 ;
  assign n49560 = ~n49437 & n49559 ;
  assign n49562 = n49561 ^ n49560 ;
  assign n49563 = ~n49432 & n49562 ;
  assign n49565 = n49564 ^ n49563 ;
  assign n49566 = ~n49427 & ~n49565 ;
  assign n49567 = n49566 ^ n49426 ;
  assign n49568 = n49567 ^ n49420 ;
  assign n49569 = n49422 & n49568 ;
  assign n49570 = n49569 ^ n49421 ;
  assign n49571 = n49570 ^ n49415 ;
  assign n49572 = n49417 & ~n49571 ;
  assign n49573 = n49572 ^ n49416 ;
  assign n49574 = n49573 ^ n1767 ;
  assign n49575 = ~n49412 & ~n49574 ;
  assign n49576 = n49575 ^ n49411 ;
  assign n49577 = n49576 ^ n49408 ;
  assign n49578 = ~n49410 & ~n49577 ;
  assign n49580 = n49579 ^ n49578 ;
  assign n49581 = n49405 & ~n49580 ;
  assign n49582 = n49581 ^ n49404 ;
  assign n49583 = n49582 ^ n49398 ;
  assign n49584 = n49400 & ~n49583 ;
  assign n49585 = n49584 ^ n49399 ;
  assign n49586 = n49585 ^ n49394 ;
  assign n49587 = n49395 & n49586 ;
  assign n49589 = n49588 ^ n49587 ;
  assign n49590 = n49390 & n49589 ;
  assign n49591 = n49590 ^ n49389 ;
  assign n49592 = n49591 ^ n49384 ;
  assign n49593 = ~n49385 & n49592 ;
  assign n49617 = n49616 ^ n49593 ;
  assign n49646 = n49617 ^ n48954 ;
  assign n48957 = n48956 ^ n47773 ;
  assign n48958 = n48957 ^ n48407 ;
  assign n49618 = n49617 ^ n48958 ;
  assign n49621 = n49591 ^ n49385 ;
  assign n49619 = n49046 ^ n48409 ;
  assign n49620 = n49619 ^ n47777 ;
  assign n49622 = n49621 ^ n49620 ;
  assign n49625 = n49589 ^ n49388 ;
  assign n49623 = n48415 ^ n47685 ;
  assign n49624 = n49623 ^ n49050 ;
  assign n49626 = n49625 ^ n49624 ;
  assign n49631 = n49585 ^ n49395 ;
  assign n49637 = n49631 ^ n49625 ;
  assign n49627 = n49582 ^ n49400 ;
  assign n49628 = n49059 ^ n48341 ;
  assign n49629 = n49628 ^ n47578 ;
  assign n49630 = n49627 & n49629 ;
  assign n49632 = n49631 ^ n49630 ;
  assign n49633 = n49055 ^ n48419 ;
  assign n49634 = n49633 ^ n47596 ;
  assign n49635 = n49634 ^ n49630 ;
  assign n49636 = n49632 & n49635 ;
  assign n49638 = n49637 ^ n49636 ;
  assign n49639 = ~n49626 & n49638 ;
  assign n49640 = n49639 ^ n49625 ;
  assign n49641 = n49640 ^ n49620 ;
  assign n49642 = ~n49622 & ~n49641 ;
  assign n49643 = n49642 ^ n49621 ;
  assign n49644 = n49643 ^ n48958 ;
  assign n49645 = ~n49618 & ~n49644 ;
  assign n49647 = n49646 ^ n49645 ;
  assign n49648 = n48955 & n49647 ;
  assign n49649 = n49648 ^ n48954 ;
  assign n49650 = n49649 ^ n48947 ;
  assign n49651 = ~n48950 & ~n49650 ;
  assign n49652 = n49651 ^ n48949 ;
  assign n48942 = n48941 ^ n48902 ;
  assign n48943 = n48942 ^ n48894 ;
  assign n48944 = n48943 ^ n48942 ;
  assign n49653 = n49652 ^ n48944 ;
  assign n49654 = ~n48895 & ~n49653 ;
  assign n49655 = n49654 ^ n48943 ;
  assign n49779 = n49512 ^ n49509 ;
  assign n49781 = n49779 ^ n48942 ;
  assign n49656 = n49028 ^ n48392 ;
  assign n49657 = n49656 ^ n47757 ;
  assign n49780 = n49779 ^ n49657 ;
  assign n49782 = n49781 ^ n49780 ;
  assign n49783 = n49655 & n49782 ;
  assign n49784 = n49783 ^ n49780 ;
  assign n49785 = n48451 ^ n47753 ;
  assign n49786 = n49785 ^ n49026 ;
  assign n49852 = n49786 ^ n49779 ;
  assign n49853 = n49784 & n49852 ;
  assign n49854 = n49853 ^ n49779 ;
  assign n49855 = n49854 ^ n49846 ;
  assign n49856 = n49855 ^ n49848 ;
  assign n49857 = n49856 ^ n49846 ;
  assign n49858 = n49851 & ~n49857 ;
  assign n49859 = n49858 ^ n49855 ;
  assign n49860 = ~n49847 & n49859 ;
  assign n49861 = n49860 ^ n49846 ;
  assign n49862 = n49861 ^ n49841 ;
  assign n49863 = ~n49843 & n49862 ;
  assign n49864 = n49863 ^ n49842 ;
  assign n49837 = n49527 ^ n49484 ;
  assign n49838 = n49837 ^ n49835 ;
  assign n49839 = n49838 ^ n49837 ;
  assign n49865 = n49864 ^ n49839 ;
  assign n49866 = n49836 & n49865 ;
  assign n49867 = n49866 ^ n49838 ;
  assign n49871 = n49837 ^ n49831 ;
  assign n49868 = n49007 ^ n47730 ;
  assign n49869 = n49868 ^ n48370 ;
  assign n49870 = n49869 ^ n49831 ;
  assign n49872 = n49871 ^ n49870 ;
  assign n49873 = n49867 & n49872 ;
  assign n49874 = n49873 ^ n49871 ;
  assign n49875 = ~n49832 & n49874 ;
  assign n49876 = n49875 ^ n49831 ;
  assign n49828 = n49537 ^ n49471 ;
  assign n49877 = n49876 ^ n49828 ;
  assign n49878 = n49877 ^ n49803 ;
  assign n49879 = n49878 ^ n49828 ;
  assign n49880 = n49827 & n49879 ;
  assign n49881 = n49880 ^ n49877 ;
  assign n49885 = n49828 ^ n49823 ;
  assign n49882 = n48994 ^ n48565 ;
  assign n49883 = n49882 ^ n47716 ;
  assign n49884 = n49883 ^ n49823 ;
  assign n49886 = n49885 ^ n49884 ;
  assign n49887 = ~n49881 & n49886 ;
  assign n49888 = n49887 ^ n49885 ;
  assign n49889 = n49824 & n49888 ;
  assign n49890 = n49889 ^ n49823 ;
  assign n49819 = n49542 ^ n49457 ;
  assign n49817 = n48984 ^ n47706 ;
  assign n49818 = n49817 ^ n48775 ;
  assign n49820 = n49819 ^ n49818 ;
  assign n49905 = n49890 ^ n49820 ;
  assign n49906 = n49905 ^ n47113 ;
  assign n49907 = n49883 ^ n49881 ;
  assign n49908 = n49907 ^ n46534 ;
  assign n49909 = n49876 ^ n49827 ;
  assign n49910 = n49909 ^ n46539 ;
  assign n49912 = n49869 ^ n49867 ;
  assign n49913 = n49912 ^ n46549 ;
  assign n49932 = n49864 ^ n49836 ;
  assign n49915 = n49859 ^ n49845 ;
  assign n49916 = n49915 ^ n46564 ;
  assign n49660 = n49652 ^ n48895 ;
  assign n49661 = n49660 ^ n46574 ;
  assign n49662 = n49649 ^ n48950 ;
  assign n49663 = n49662 ^ n46581 ;
  assign n49686 = n49647 ^ n48953 ;
  assign n49665 = n49640 ^ n49622 ;
  assign n49666 = n49665 ^ n46594 ;
  assign n49674 = n49638 ^ n49624 ;
  assign n49667 = n49629 ^ n49627 ;
  assign n49668 = ~n46608 & n49667 ;
  assign n49669 = n49668 ^ n46604 ;
  assign n49670 = n49635 ^ n49631 ;
  assign n49671 = n49670 ^ n49668 ;
  assign n49672 = ~n49669 & n49671 ;
  assign n49673 = n49672 ^ n46604 ;
  assign n49675 = n49674 ^ n49673 ;
  assign n49676 = n49674 ^ n46596 ;
  assign n49677 = ~n49675 & ~n49676 ;
  assign n49678 = n49677 ^ n46596 ;
  assign n49679 = n49678 ^ n49665 ;
  assign n49680 = ~n49666 & n49679 ;
  assign n49681 = n49680 ^ n46594 ;
  assign n49664 = n49643 ^ n49618 ;
  assign n49682 = n49681 ^ n49664 ;
  assign n49683 = n49681 ^ n46587 ;
  assign n49684 = ~n49682 & n49683 ;
  assign n49685 = n49684 ^ n46587 ;
  assign n49687 = n49686 ^ n49685 ;
  assign n49688 = n49686 ^ n46585 ;
  assign n49689 = ~n49687 & ~n49688 ;
  assign n49690 = n49689 ^ n46585 ;
  assign n49691 = n49690 ^ n49662 ;
  assign n49692 = n49663 & ~n49691 ;
  assign n49693 = n49692 ^ n46581 ;
  assign n49694 = n49693 ^ n49660 ;
  assign n49695 = ~n49661 & n49694 ;
  assign n49696 = n49695 ^ n46574 ;
  assign n49658 = n49657 ^ n49655 ;
  assign n49778 = n49696 ^ n49658 ;
  assign n49787 = n49786 ^ n49784 ;
  assign n49788 = n49787 ^ n46937 ;
  assign n49789 = n49788 ^ n49787 ;
  assign n49790 = n49789 ^ n49658 ;
  assign n49791 = n49778 & ~n49790 ;
  assign n49792 = n49791 ^ n49788 ;
  assign n49918 = n49787 ^ n46566 ;
  assign n49919 = ~n49792 & n49918 ;
  assign n49920 = n49919 ^ n46566 ;
  assign n49917 = n49854 ^ n49851 ;
  assign n49921 = n49920 ^ n49917 ;
  assign n49922 = n49920 ^ n46947 ;
  assign n49923 = n49921 & ~n49922 ;
  assign n49924 = n49923 ^ n46947 ;
  assign n49925 = n49924 ^ n49915 ;
  assign n49926 = ~n49916 & ~n49925 ;
  assign n49927 = n49926 ^ n46564 ;
  assign n49914 = n49861 ^ n49843 ;
  assign n49928 = n49927 ^ n49914 ;
  assign n49929 = n49927 ^ n46559 ;
  assign n49930 = n49928 & n49929 ;
  assign n49931 = n49930 ^ n46559 ;
  assign n49933 = n49932 ^ n49931 ;
  assign n49934 = n49912 ^ n46554 ;
  assign n49935 = n49934 ^ n49912 ;
  assign n49936 = n49935 ^ n49931 ;
  assign n49937 = ~n49933 & n49936 ;
  assign n49938 = n49937 ^ n49934 ;
  assign n49939 = ~n49913 & ~n49938 ;
  assign n49940 = n49939 ^ n46549 ;
  assign n49911 = n49874 ^ n49829 ;
  assign n49941 = n49940 ^ n49911 ;
  assign n49942 = n49940 ^ n46544 ;
  assign n49943 = ~n49941 & n49942 ;
  assign n49944 = n49943 ^ n46544 ;
  assign n49945 = n49944 ^ n49909 ;
  assign n49946 = n49910 & ~n49945 ;
  assign n49947 = n49946 ^ n46539 ;
  assign n49948 = n49947 ^ n49907 ;
  assign n49949 = ~n49908 & n49948 ;
  assign n49950 = n49949 ^ n46534 ;
  assign n49951 = n49950 ^ n46974 ;
  assign n49952 = n49888 ^ n49821 ;
  assign n49953 = n49952 ^ n49950 ;
  assign n49954 = n49951 & ~n49953 ;
  assign n49955 = n49954 ^ n46974 ;
  assign n49956 = n49955 ^ n49905 ;
  assign n49957 = ~n49906 & ~n49956 ;
  assign n49958 = n49957 ^ n47113 ;
  assign n49891 = n49890 ^ n49818 ;
  assign n49892 = n49820 & n49891 ;
  assign n49893 = n49892 ^ n49819 ;
  assign n49815 = n49546 ^ n49545 ;
  assign n49813 = n48784 ^ n47830 ;
  assign n49814 = n49813 ^ n48980 ;
  assign n49816 = n49815 ^ n49814 ;
  assign n49903 = n49893 ^ n49816 ;
  assign n49904 = n49903 ^ n47386 ;
  assign n50014 = n49958 ^ n49904 ;
  assign n49988 = n49924 ^ n49916 ;
  assign n49989 = n49917 ^ n46947 ;
  assign n49990 = n49989 ^ n49920 ;
  assign n49793 = n49792 ^ n46566 ;
  assign n49659 = n49658 ^ n46937 ;
  assign n49697 = n49696 ^ n49659 ;
  assign n49698 = n49670 ^ n49669 ;
  assign n49699 = n49676 ^ n49673 ;
  assign n49700 = ~n49698 & ~n49699 ;
  assign n49701 = n49678 ^ n49666 ;
  assign n49702 = ~n49700 & ~n49701 ;
  assign n49703 = n49682 ^ n46587 ;
  assign n49704 = ~n49702 & ~n49703 ;
  assign n49705 = n49688 ^ n49685 ;
  assign n49706 = ~n49704 & ~n49705 ;
  assign n49707 = n49690 ^ n49663 ;
  assign n49708 = ~n49706 & n49707 ;
  assign n49709 = n49693 ^ n49661 ;
  assign n49710 = n49708 & ~n49709 ;
  assign n49794 = ~n49697 & n49710 ;
  assign n49991 = ~n49793 & ~n49794 ;
  assign n49992 = ~n49990 & n49991 ;
  assign n49993 = ~n49988 & n49992 ;
  assign n49994 = n49914 ^ n46559 ;
  assign n49995 = n49994 ^ n49927 ;
  assign n49996 = n49993 & n49995 ;
  assign n49997 = n49932 ^ n46554 ;
  assign n49998 = n49997 ^ n49931 ;
  assign n49999 = n49996 & ~n49998 ;
  assign n50000 = n49938 ^ n46549 ;
  assign n50001 = ~n49999 & ~n50000 ;
  assign n50002 = n49911 ^ n46544 ;
  assign n50003 = n50002 ^ n49940 ;
  assign n50004 = n50001 & ~n50003 ;
  assign n50005 = n49944 ^ n46539 ;
  assign n50006 = n50005 ^ n49909 ;
  assign n50007 = ~n50004 & n50006 ;
  assign n50008 = n49947 ^ n49908 ;
  assign n50009 = ~n50007 & n50008 ;
  assign n50010 = n49952 ^ n49951 ;
  assign n50011 = ~n50009 & n50010 ;
  assign n50012 = n49955 ^ n49906 ;
  assign n50013 = n50011 & ~n50012 ;
  assign n50095 = n50014 ^ n50013 ;
  assign n50099 = n50098 ^ n50095 ;
  assign n50103 = n50012 ^ n50011 ;
  assign n50100 = n48034 ^ n1616 ;
  assign n50101 = n50100 ^ n44033 ;
  assign n50102 = n50101 ^ n38566 ;
  assign n50104 = n50103 ^ n50102 ;
  assign n50108 = n50010 ^ n50009 ;
  assign n50105 = n48039 ^ n40100 ;
  assign n50106 = n50105 ^ n44323 ;
  assign n50107 = n50106 ^ n38571 ;
  assign n50109 = n50108 ^ n50107 ;
  assign n50115 = n50008 ^ n50007 ;
  assign n50112 = n48043 ^ n40106 ;
  assign n50113 = n50112 ^ n44328 ;
  assign n50114 = n50113 ^ n2975 ;
  assign n50116 = n50115 ^ n50114 ;
  assign n50120 = n50006 ^ n50004 ;
  assign n50117 = n48048 ^ n40111 ;
  assign n50118 = n50117 ^ n44334 ;
  assign n50119 = n50118 ^ n38578 ;
  assign n50121 = n50120 ^ n50119 ;
  assign n50125 = n50003 ^ n50001 ;
  assign n50122 = n48053 ^ n40117 ;
  assign n50123 = n50122 ^ n44338 ;
  assign n50124 = n50123 ^ n38583 ;
  assign n50126 = n50125 ^ n50124 ;
  assign n50130 = n50000 ^ n49999 ;
  assign n50127 = n48059 ^ n40122 ;
  assign n50128 = n50127 ^ n44343 ;
  assign n50129 = n50128 ^ n38589 ;
  assign n50131 = n50130 ^ n50129 ;
  assign n50133 = n48064 ^ n40126 ;
  assign n50134 = n50133 ^ n44348 ;
  assign n50135 = n50134 ^ n38593 ;
  assign n50166 = n50135 ^ n50129 ;
  assign n50132 = n49998 ^ n49996 ;
  assign n50136 = n50135 ^ n50132 ;
  assign n50140 = n49995 ^ n49993 ;
  assign n50163 = n50140 ^ n50135 ;
  assign n50137 = n48069 ^ n40131 ;
  assign n50138 = n50137 ^ n44353 ;
  assign n50139 = n50138 ^ n38599 ;
  assign n50141 = n50140 ^ n50139 ;
  assign n50146 = n49992 ^ n49988 ;
  assign n50142 = n48073 ^ n2440 ;
  assign n50143 = n50142 ^ n44359 ;
  assign n50144 = n50143 ^ n38604 ;
  assign n50147 = n50146 ^ n50144 ;
  assign n50151 = n49991 ^ n49990 ;
  assign n50148 = n47678 ^ n2422 ;
  assign n50149 = n50148 ^ n44417 ;
  assign n50150 = n50149 ^ n38608 ;
  assign n50152 = n50151 ^ n50150 ;
  assign n49795 = n49794 ^ n49793 ;
  assign n50155 = n50151 ^ n49795 ;
  assign n49712 = n47615 ^ n40146 ;
  assign n49713 = n49712 ^ n44408 ;
  assign n49714 = n49713 ^ n38620 ;
  assign n49796 = n49795 ^ n49714 ;
  assign n49711 = n49710 ^ n49697 ;
  assign n49715 = n49714 ^ n49711 ;
  assign n49719 = n49709 ^ n49708 ;
  assign n49716 = n47621 ^ n40151 ;
  assign n49717 = n49716 ^ n44371 ;
  assign n49718 = n49717 ^ n38624 ;
  assign n49720 = n49719 ^ n49718 ;
  assign n49722 = n47626 ^ n40155 ;
  assign n49723 = n49722 ^ n44376 ;
  assign n49724 = n49723 ^ n2015 ;
  assign n49772 = n49724 ^ n49718 ;
  assign n49721 = n49707 ^ n49706 ;
  assign n49725 = n49724 ^ n49721 ;
  assign n49729 = n49705 ^ n49704 ;
  assign n49726 = n47630 ^ n40161 ;
  assign n49727 = n49726 ^ n44381 ;
  assign n49728 = n49727 ^ n38632 ;
  assign n49730 = n49729 ^ n49728 ;
  assign n49731 = n47636 ^ n40185 ;
  assign n49732 = n49731 ^ n44387 ;
  assign n49733 = n49732 ^ n38636 ;
  assign n49766 = n49733 ^ n49728 ;
  assign n49734 = n49703 ^ n49702 ;
  assign n49735 = n49734 ^ n49733 ;
  assign n49739 = n49701 ^ n49700 ;
  assign n49736 = n47655 ^ n40165 ;
  assign n49737 = n49736 ^ n43984 ;
  assign n49738 = n49737 ^ n3053 ;
  assign n49740 = n49739 ^ n49738 ;
  assign n49742 = n47640 ^ n40169 ;
  assign n49743 = n49742 ^ n2783 ;
  assign n49744 = n49743 ^ n38644 ;
  assign n49760 = n49744 ^ n49739 ;
  assign n49741 = n49699 ^ n49698 ;
  assign n49745 = n49744 ^ n49741 ;
  assign n49749 = n49667 ^ n46608 ;
  assign n49750 = n48225 ^ n2684 ;
  assign n49751 = n49750 ^ n44818 ;
  assign n49752 = n49751 ^ n38993 ;
  assign n49753 = ~n49749 & n49752 ;
  assign n49746 = n47644 ^ n40172 ;
  assign n49747 = n49746 ^ n43976 ;
  assign n49748 = n49747 ^ n2775 ;
  assign n49754 = n49753 ^ n49748 ;
  assign n49755 = n49753 ^ n49698 ;
  assign n49756 = ~n49754 & ~n49755 ;
  assign n49757 = n49756 ^ n49698 ;
  assign n49758 = n49757 ^ n49744 ;
  assign n49759 = ~n49745 & ~n49758 ;
  assign n49761 = n49760 ^ n49759 ;
  assign n49762 = n49740 & n49761 ;
  assign n49763 = n49762 ^ n49739 ;
  assign n49764 = n49763 ^ n49733 ;
  assign n49765 = ~n49735 & n49764 ;
  assign n49767 = n49766 ^ n49765 ;
  assign n49768 = n49730 & ~n49767 ;
  assign n49769 = n49768 ^ n49729 ;
  assign n49770 = n49769 ^ n49721 ;
  assign n49771 = n49725 & ~n49770 ;
  assign n49773 = n49772 ^ n49771 ;
  assign n49774 = n49720 & ~n49773 ;
  assign n49775 = n49774 ^ n49719 ;
  assign n49776 = n49775 ^ n49714 ;
  assign n49777 = n49715 & n49776 ;
  assign n49797 = n49796 ^ n49777 ;
  assign n49798 = n47611 ^ n40141 ;
  assign n49799 = n49798 ^ n44364 ;
  assign n49800 = n49799 ^ n38614 ;
  assign n50153 = n49800 ^ n49795 ;
  assign n50154 = n49797 & n50153 ;
  assign n50156 = n50155 ^ n50154 ;
  assign n50157 = ~n50152 & ~n50156 ;
  assign n50158 = n50157 ^ n50151 ;
  assign n50159 = n50158 ^ n50144 ;
  assign n50160 = ~n50147 & ~n50159 ;
  assign n50145 = n50144 ^ n50139 ;
  assign n50161 = n50160 ^ n50145 ;
  assign n50162 = n50141 & ~n50161 ;
  assign n50164 = n50163 ^ n50162 ;
  assign n50165 = ~n50136 & n50164 ;
  assign n50167 = n50166 ^ n50165 ;
  assign n50168 = ~n50131 & ~n50167 ;
  assign n50169 = n50168 ^ n50130 ;
  assign n50170 = n50169 ^ n50124 ;
  assign n50171 = n50126 & n50170 ;
  assign n50172 = n50171 ^ n50125 ;
  assign n50173 = n50172 ^ n50119 ;
  assign n50174 = ~n50121 & ~n50173 ;
  assign n50175 = n50174 ^ n50120 ;
  assign n50176 = n50175 ^ n50114 ;
  assign n50177 = n50116 & n50176 ;
  assign n50178 = n50177 ^ n50115 ;
  assign n50179 = n50178 ^ n50107 ;
  assign n50180 = ~n50109 & n50179 ;
  assign n50110 = n50107 ^ n50102 ;
  assign n50181 = n50180 ^ n50110 ;
  assign n50182 = ~n50104 & ~n50181 ;
  assign n50183 = n50182 ^ n50103 ;
  assign n50184 = n50183 ^ n50095 ;
  assign n50185 = ~n50099 & ~n50184 ;
  assign n50187 = n50186 ^ n50185 ;
  assign n49959 = n49958 ^ n49903 ;
  assign n49960 = n49904 & n49959 ;
  assign n49961 = n49960 ^ n47386 ;
  assign n49899 = n49550 ^ n49451 ;
  assign n49897 = n48835 ^ n47931 ;
  assign n49898 = n49897 ^ n48978 ;
  assign n49900 = n49899 ^ n49898 ;
  assign n49894 = n49893 ^ n49814 ;
  assign n49895 = ~n49816 & ~n49894 ;
  assign n49896 = n49895 ^ n49815 ;
  assign n49901 = n49900 ^ n49896 ;
  assign n49902 = n49901 ^ n47420 ;
  assign n50016 = n49961 ^ n49902 ;
  assign n50015 = n50013 & ~n50014 ;
  assign n50093 = n50016 ^ n50015 ;
  assign n50428 = n50187 ^ n50093 ;
  assign n50232 = n49570 ^ n49417 ;
  assign n51360 = n50428 ^ n50232 ;
  assign n51361 = n51360 ^ n48971 ;
  assign n50858 = n48660 ^ n40879 ;
  assign n50859 = n50858 ^ n45131 ;
  assign n50860 = n50859 ^ n39241 ;
  assign n50852 = n48655 ^ n40874 ;
  assign n50853 = n50852 ^ n45126 ;
  assign n50854 = n50853 ^ n39234 ;
  assign n50947 = n50860 ^ n50854 ;
  assign n50479 = n49821 ^ n48374 ;
  assign n50480 = n50479 ^ n49002 ;
  assign n50398 = n49775 ^ n49715 ;
  assign n50481 = n50480 ^ n50398 ;
  assign n50401 = n49773 ^ n49719 ;
  assign n50538 = n50401 ^ n50398 ;
  assign n50482 = n49828 ^ n49007 ;
  assign n50483 = n50482 ^ n48376 ;
  assign n50484 = n50483 ^ n50401 ;
  assign n50485 = n49803 ^ n48384 ;
  assign n50486 = n50485 ^ n49006 ;
  assign n50407 = n49769 ^ n49725 ;
  assign n50487 = n50486 ^ n50407 ;
  assign n50488 = n49829 ^ n49012 ;
  assign n50489 = n50488 ^ n48388 ;
  assign n50412 = n49767 ^ n49729 ;
  assign n50490 = n50489 ^ n50412 ;
  assign n50493 = n49763 ^ n49735 ;
  assign n50491 = n49016 ^ n48451 ;
  assign n50492 = n50491 ^ n49837 ;
  assign n50494 = n50493 ^ n50492 ;
  assign n50496 = n49022 ^ n48392 ;
  assign n50497 = n50496 ^ n49835 ;
  assign n50495 = n49761 ^ n49738 ;
  assign n50498 = n50497 ^ n50495 ;
  assign n50501 = n49757 ^ n49745 ;
  assign n50523 = n50501 ^ n50495 ;
  assign n50499 = n49842 ^ n49026 ;
  assign n50500 = n50499 ^ n47695 ;
  assign n50502 = n50501 ^ n50500 ;
  assign n50512 = n49748 ^ n49698 ;
  assign n50513 = n50512 ^ n49753 ;
  assign n50505 = n49752 ^ n49749 ;
  assign n50514 = n50513 ^ n50505 ;
  assign n50503 = n48403 ^ n48351 ;
  assign n50504 = n50503 ^ n49848 ;
  assign n50506 = n50505 ^ n50504 ;
  assign n50283 = n49573 ^ n49412 ;
  assign n50281 = n48889 ^ n48238 ;
  assign n50282 = n50281 ^ n47542 ;
  assign n50284 = n50283 ^ n50282 ;
  assign n50230 = n48197 ^ n47502 ;
  assign n50231 = n50230 ^ n48843 ;
  assign n50233 = n50232 ^ n50231 ;
  assign n50207 = n49567 ^ n49422 ;
  assign n50057 = n49565 ^ n49426 ;
  assign n50208 = n50207 ^ n50057 ;
  assign n50043 = n49562 ^ n49428 ;
  assign n50058 = n50057 ^ n50043 ;
  assign n50044 = n48162 ^ n47399 ;
  assign n50045 = n50044 ^ n48961 ;
  assign n50046 = n50045 ^ n50043 ;
  assign n50026 = n49558 ^ n49437 ;
  assign n50024 = n48975 ^ n48228 ;
  assign n50025 = n50024 ^ n48965 ;
  assign n50027 = n50026 ^ n50025 ;
  assign n49983 = n49556 ^ n49440 ;
  assign n49981 = n48917 ^ n48178 ;
  assign n49982 = n49981 ^ n48971 ;
  assign n49984 = n49983 ^ n49982 ;
  assign n49971 = n49552 ^ n49447 ;
  assign n49969 = n48873 ^ n48143 ;
  assign n49970 = n49969 ^ n48969 ;
  assign n49972 = n49971 ^ n49970 ;
  assign n49966 = n49898 ^ n49896 ;
  assign n49967 = n49900 & ~n49966 ;
  assign n49968 = n49967 ^ n49899 ;
  assign n49978 = n49970 ^ n49968 ;
  assign n49979 = ~n49972 & ~n49978 ;
  assign n49980 = n49979 ^ n49971 ;
  assign n50021 = n49982 ^ n49980 ;
  assign n50022 = n49984 & n50021 ;
  assign n50023 = n50022 ^ n49983 ;
  assign n50040 = n50025 ^ n50023 ;
  assign n50041 = n50027 & n50040 ;
  assign n50042 = n50041 ^ n50026 ;
  assign n50055 = n50043 ^ n50042 ;
  assign n50056 = ~n50046 & n50055 ;
  assign n50059 = n50058 ^ n50056 ;
  assign n50053 = n48165 ^ n47428 ;
  assign n50054 = n50053 ^ n49604 ;
  assign n50205 = n50057 ^ n50054 ;
  assign n50206 = n50059 & n50205 ;
  assign n50209 = n50208 ^ n50206 ;
  assign n50210 = n48811 ^ n48155 ;
  assign n50211 = n50210 ^ n47458 ;
  assign n50227 = n50211 ^ n50207 ;
  assign n50228 = n50209 & n50227 ;
  assign n50229 = n50228 ^ n50207 ;
  assign n50278 = n50232 ^ n50229 ;
  assign n50279 = ~n50233 & ~n50278 ;
  assign n50280 = n50279 ^ n50232 ;
  assign n50324 = n50283 ^ n50280 ;
  assign n50325 = n50284 & ~n50324 ;
  assign n50326 = n50325 ^ n50283 ;
  assign n50321 = n48937 ^ n47549 ;
  assign n50322 = n50321 ^ n48259 ;
  assign n50377 = n50326 ^ n50322 ;
  assign n50320 = n49576 ^ n49410 ;
  assign n50378 = n50326 ^ n50320 ;
  assign n50379 = n50377 & n50378 ;
  assign n50372 = n46616 ^ n46612 ;
  assign n50370 = n49580 ^ n49404 ;
  assign n50367 = n48274 ^ n47568 ;
  assign n50368 = n50367 ^ n49085 ;
  assign n50369 = n50368 ^ n50322 ;
  assign n50371 = n50370 ^ n50369 ;
  assign n50373 = n50372 ^ n50371 ;
  assign n50364 = n48195 ^ n40340 ;
  assign n50365 = n50364 ^ n44783 ;
  assign n50366 = n50365 ^ n38949 ;
  assign n50374 = n50373 ^ n50366 ;
  assign n50335 = n48136 ^ n40284 ;
  assign n50336 = n50335 ^ n44755 ;
  assign n50337 = n50336 ^ n38812 ;
  assign n50375 = n50374 ^ n50337 ;
  assign n50323 = n50322 ^ n50320 ;
  assign n50327 = n50326 ^ n50323 ;
  assign n50328 = n50327 ^ n46616 ;
  assign n50212 = n50211 ^ n50209 ;
  assign n50213 = n50212 ^ n46882 ;
  assign n50060 = n50059 ^ n50054 ;
  assign n50061 = n50060 ^ n46894 ;
  assign n49985 = n49984 ^ n49980 ;
  assign n49962 = n49961 ^ n49901 ;
  assign n49963 = ~n49902 & ~n49962 ;
  assign n49964 = n49963 ^ n47420 ;
  assign n49965 = n49964 ^ n47442 ;
  assign n49973 = n49972 ^ n49968 ;
  assign n49974 = n49973 ^ n49964 ;
  assign n49975 = n49965 & ~n49974 ;
  assign n49976 = n49975 ^ n47442 ;
  assign n50020 = n49985 ^ n49976 ;
  assign n50028 = n50027 ^ n50023 ;
  assign n50029 = n50028 ^ n47486 ;
  assign n50030 = n50029 ^ n50028 ;
  assign n50031 = n50030 ^ n49976 ;
  assign n50032 = ~n50020 & n50031 ;
  assign n50033 = n50032 ^ n50029 ;
  assign n50036 = n50028 ^ n47528 ;
  assign n50037 = n50033 & n50036 ;
  assign n50038 = n50037 ^ n47528 ;
  assign n50039 = n50038 ^ n46891 ;
  assign n50047 = n50046 ^ n50042 ;
  assign n50050 = n50047 ^ n50038 ;
  assign n50051 = n50039 & ~n50050 ;
  assign n50052 = n50051 ^ n46891 ;
  assign n50214 = n50060 ^ n50052 ;
  assign n50215 = n50061 & n50214 ;
  assign n50216 = n50215 ^ n46894 ;
  assign n50236 = n50216 ^ n50212 ;
  assign n50237 = n50213 & ~n50236 ;
  assign n50238 = n50237 ^ n46882 ;
  assign n50234 = n50233 ^ n50229 ;
  assign n50277 = n50238 ^ n50234 ;
  assign n50285 = n50284 ^ n50280 ;
  assign n50286 = n50285 ^ n46880 ;
  assign n50287 = n50286 ^ n50285 ;
  assign n50288 = n50287 ^ n50234 ;
  assign n50289 = n50277 & ~n50288 ;
  assign n50290 = n50289 ^ n50286 ;
  assign n50329 = n50285 ^ n46876 ;
  assign n50330 = n50290 & n50329 ;
  assign n50331 = n50330 ^ n46876 ;
  assign n50362 = n50331 ^ n50327 ;
  assign n50363 = n50328 & ~n50362 ;
  assign n50376 = n50375 ^ n50363 ;
  assign n50380 = n50379 ^ n50376 ;
  assign n50332 = n50331 ^ n50328 ;
  assign n50291 = n50290 ^ n46876 ;
  assign n50235 = n50234 ^ n46880 ;
  assign n50239 = n50238 ^ n50235 ;
  assign n50217 = n50216 ^ n50213 ;
  assign n49977 = n49976 ^ n47486 ;
  assign n49986 = n49985 ^ n49977 ;
  assign n49987 = n49973 ^ n49965 ;
  assign n50017 = ~n50015 & n50016 ;
  assign n50018 = n49987 & n50017 ;
  assign n50019 = ~n49986 & ~n50018 ;
  assign n50034 = n50033 ^ n47528 ;
  assign n50035 = n50019 & ~n50034 ;
  assign n50048 = n50047 ^ n50039 ;
  assign n50049 = ~n50035 & ~n50048 ;
  assign n50062 = n50061 ^ n50052 ;
  assign n50218 = ~n50049 & n50062 ;
  assign n50240 = n50217 & ~n50218 ;
  assign n50292 = n50239 & ~n50240 ;
  assign n50333 = ~n50291 & n50292 ;
  assign n50361 = ~n50332 & ~n50333 ;
  assign n50381 = n50380 ^ n50361 ;
  assign n50334 = n50333 ^ n50332 ;
  assign n50338 = n50337 ^ n50334 ;
  assign n50293 = n50292 ^ n50291 ;
  assign n50274 = n47705 ^ n38845 ;
  assign n50275 = n50274 ^ n44731 ;
  assign n50276 = n50275 ^ n38763 ;
  assign n50294 = n50293 ^ n50276 ;
  assign n50064 = n47999 ^ n40070 ;
  assign n50065 = n50064 ^ n44643 ;
  assign n50066 = n50065 ^ n38544 ;
  assign n50063 = n50062 ^ n50049 ;
  assign n50067 = n50066 ^ n50063 ;
  assign n50076 = n50048 ^ n50035 ;
  assign n50073 = n48005 ^ n40075 ;
  assign n50074 = n50073 ^ n1286 ;
  assign n50075 = n50074 ^ n38548 ;
  assign n50077 = n50076 ^ n50075 ;
  assign n50081 = n50034 ^ n50019 ;
  assign n50078 = n48011 ^ n40079 ;
  assign n50079 = n50078 ^ n44665 ;
  assign n50080 = n50079 ^ n1278 ;
  assign n50082 = n50081 ^ n50080 ;
  assign n50083 = n50018 ^ n49986 ;
  assign n1092 = n1091 ^ n1049 ;
  assign n1126 = n1125 ^ n1092 ;
  assign n1136 = n1135 ^ n1126 ;
  assign n50084 = n50083 ^ n1136 ;
  assign n50088 = n50017 ^ n49987 ;
  assign n50085 = n48018 ^ n40086 ;
  assign n50086 = n50085 ^ n44672 ;
  assign n50087 = n50086 ^ n1117 ;
  assign n50089 = n50088 ^ n50087 ;
  assign n50094 = n50093 ^ n50092 ;
  assign n50188 = n50094 & ~n50187 ;
  assign n50189 = n50188 ^ n50093 ;
  assign n50190 = n50189 ^ n50087 ;
  assign n50191 = ~n50089 & ~n50190 ;
  assign n50192 = n50191 ^ n50088 ;
  assign n50193 = n50192 ^ n1136 ;
  assign n50194 = n50084 & n50193 ;
  assign n50195 = n50194 ^ n50083 ;
  assign n50196 = n50195 ^ n50080 ;
  assign n50197 = ~n50082 & ~n50196 ;
  assign n50198 = n50197 ^ n50081 ;
  assign n50199 = n50198 ^ n50075 ;
  assign n50200 = ~n50077 & n50199 ;
  assign n50201 = n50200 ^ n50076 ;
  assign n50202 = n50201 ^ n50066 ;
  assign n50203 = ~n50067 & ~n50202 ;
  assign n50068 = n47995 ^ n40065 ;
  assign n50069 = n50068 ^ n44715 ;
  assign n50070 = n50069 ^ n38539 ;
  assign n50071 = n50070 ^ n50066 ;
  assign n50204 = n50203 ^ n50071 ;
  assign n50219 = n50218 ^ n50217 ;
  assign n50243 = n50219 ^ n50070 ;
  assign n50244 = n50204 & n50243 ;
  assign n50241 = n50240 ^ n50239 ;
  assign n50242 = n50241 ^ n50070 ;
  assign n50245 = n50244 ^ n50242 ;
  assign n50246 = n47989 ^ n40060 ;
  assign n50247 = n50246 ^ n44723 ;
  assign n50248 = n50247 ^ n38746 ;
  assign n50271 = n50248 ^ n50241 ;
  assign n50272 = ~n50245 & ~n50271 ;
  assign n50273 = n50272 ^ n50241 ;
  assign n50317 = n50276 ^ n50273 ;
  assign n50318 = ~n50294 & n50317 ;
  assign n50319 = n50318 ^ n50293 ;
  assign n50359 = n50337 ^ n50319 ;
  assign n50360 = ~n50338 & ~n50359 ;
  assign n50382 = n50381 ^ n50360 ;
  assign n50509 = n50505 ^ n50382 ;
  assign n50357 = n49779 ^ n48945 ;
  assign n50358 = n50357 ^ n48407 ;
  assign n50383 = n50382 ^ n50358 ;
  assign n50251 = n49046 ^ n48949 ;
  assign n50252 = n50251 ^ n48419 ;
  assign n49811 = n49050 ^ n48341 ;
  assign n49812 = n49811 ^ n48954 ;
  assign n50220 = n50219 ^ n50204 ;
  assign n50250 = ~n49812 & n50220 ;
  assign n50253 = n50252 ^ n50250 ;
  assign n50264 = n48956 ^ n48894 ;
  assign n50265 = n50264 ^ n48415 ;
  assign n50266 = n50265 ^ n50250 ;
  assign n50267 = n50266 ^ n50265 ;
  assign n50249 = n50248 ^ n50245 ;
  assign n50268 = n50267 ^ n50249 ;
  assign n50269 = n50253 & ~n50268 ;
  assign n50270 = n50269 ^ n50266 ;
  assign n50295 = n50294 ^ n50273 ;
  assign n50314 = n50295 ^ n50265 ;
  assign n50315 = ~n50270 & ~n50314 ;
  assign n50311 = n48951 ^ n48409 ;
  assign n50312 = n50311 ^ n48942 ;
  assign n50313 = n50312 ^ n50265 ;
  assign n50316 = n50315 ^ n50313 ;
  assign n50339 = n50338 ^ n50319 ;
  assign n50354 = n50339 ^ n50312 ;
  assign n50355 = n50316 & ~n50354 ;
  assign n50356 = n50355 ^ n50312 ;
  assign n50507 = n50382 ^ n50356 ;
  assign n50508 = n50383 & ~n50507 ;
  assign n50510 = n50509 ^ n50508 ;
  assign n50511 = n50506 & ~n50510 ;
  assign n50515 = n50514 ^ n50511 ;
  assign n50516 = n49028 ^ n48399 ;
  assign n50517 = n50516 ^ n49846 ;
  assign n50518 = n50517 ^ n50513 ;
  assign n50519 = n50515 & ~n50518 ;
  assign n50520 = n50519 ^ n50513 ;
  assign n50521 = n50520 ^ n50500 ;
  assign n50522 = ~n50502 & ~n50521 ;
  assign n50524 = n50523 ^ n50522 ;
  assign n50525 = ~n50498 & ~n50524 ;
  assign n50526 = n50525 ^ n50497 ;
  assign n50527 = n50526 ^ n50492 ;
  assign n50528 = n50494 & ~n50527 ;
  assign n50529 = n50528 ^ n50493 ;
  assign n50530 = n50529 ^ n50489 ;
  assign n50531 = n50490 & n50530 ;
  assign n50532 = n50531 ^ n50412 ;
  assign n50533 = n50532 ^ n50486 ;
  assign n50534 = ~n50487 & n50533 ;
  assign n50535 = n50534 ^ n50407 ;
  assign n50536 = n50535 ^ n50483 ;
  assign n50537 = ~n50484 & n50536 ;
  assign n50539 = n50538 ^ n50537 ;
  assign n50540 = n50481 & n50539 ;
  assign n50541 = n50540 ^ n50398 ;
  assign n50476 = n48998 ^ n48370 ;
  assign n50477 = n50476 ^ n49819 ;
  assign n49801 = n49800 ^ n49797 ;
  assign n50478 = n50477 ^ n49801 ;
  assign n50623 = n50541 ^ n50478 ;
  assign n50624 = n50623 ^ n47730 ;
  assign n50625 = n50539 ^ n50480 ;
  assign n50626 = n50625 ^ n47734 ;
  assign n50627 = n50535 ^ n50484 ;
  assign n50628 = n50627 ^ n47739 ;
  assign n50629 = n50532 ^ n50487 ;
  assign n50630 = n50629 ^ n47743 ;
  assign n50631 = n50529 ^ n50490 ;
  assign n50632 = n50631 ^ n47749 ;
  assign n50633 = n50526 ^ n50494 ;
  assign n50634 = n50633 ^ n47753 ;
  assign n50635 = n50524 ^ n50497 ;
  assign n50636 = n50635 ^ n47757 ;
  assign n50645 = n50517 ^ n50515 ;
  assign n50384 = n50383 ^ n50356 ;
  assign n50385 = n50384 ^ n47773 ;
  assign n50340 = n50339 ^ n50316 ;
  assign n50341 = n50340 ^ n47777 ;
  assign n50296 = n50295 ^ n50270 ;
  assign n50254 = n50253 ^ n50249 ;
  assign n50221 = n50220 ^ n49812 ;
  assign n50225 = ~n47578 & ~n50221 ;
  assign n50259 = n50254 ^ n50225 ;
  assign n50260 = n50254 ^ n47596 ;
  assign n50261 = n50259 & ~n50260 ;
  assign n50262 = n50261 ^ n47596 ;
  assign n50307 = n50296 ^ n50262 ;
  assign n50308 = n50296 ^ n47685 ;
  assign n50309 = n50307 & n50308 ;
  assign n50310 = n50309 ^ n47685 ;
  assign n50351 = n50340 ^ n50310 ;
  assign n50352 = ~n50341 & n50351 ;
  assign n50353 = n50352 ^ n47777 ;
  assign n50638 = n50384 ^ n50353 ;
  assign n50639 = ~n50385 & ~n50638 ;
  assign n50640 = n50639 ^ n47773 ;
  assign n50637 = n50510 ^ n50504 ;
  assign n50641 = n50640 ^ n50637 ;
  assign n50642 = n50640 ^ n47771 ;
  assign n50643 = ~n50641 & n50642 ;
  assign n50644 = n50643 ^ n47771 ;
  assign n50646 = n50645 ^ n50644 ;
  assign n50647 = n50520 ^ n50502 ;
  assign n50648 = n50647 ^ n47765 ;
  assign n50649 = n50648 ^ n50647 ;
  assign n50650 = n50649 ^ n50644 ;
  assign n50651 = ~n50646 & n50650 ;
  assign n50652 = n50651 ^ n50648 ;
  assign n50654 = n50635 ^ n47696 ;
  assign n50653 = n50647 ^ n50635 ;
  assign n50655 = n50654 ^ n50653 ;
  assign n50656 = ~n50652 & ~n50655 ;
  assign n50657 = n50656 ^ n50654 ;
  assign n50658 = ~n50636 & ~n50657 ;
  assign n50659 = n50658 ^ n47757 ;
  assign n50660 = n50659 ^ n50633 ;
  assign n50661 = n50634 & n50660 ;
  assign n50662 = n50661 ^ n47753 ;
  assign n50663 = n50662 ^ n50631 ;
  assign n50664 = n50632 & ~n50663 ;
  assign n50665 = n50664 ^ n47749 ;
  assign n50666 = n50665 ^ n50629 ;
  assign n50667 = n50630 & ~n50666 ;
  assign n50668 = n50667 ^ n47743 ;
  assign n50669 = n50668 ^ n50627 ;
  assign n50670 = ~n50628 & ~n50669 ;
  assign n50671 = n50670 ^ n47739 ;
  assign n50672 = n50671 ^ n50625 ;
  assign n50673 = n50626 & ~n50672 ;
  assign n50674 = n50673 ^ n47734 ;
  assign n50675 = n50674 ^ n50623 ;
  assign n50676 = n50624 & ~n50675 ;
  assign n50677 = n50676 ^ n47730 ;
  assign n50472 = n49815 ^ n48366 ;
  assign n50473 = n50472 ^ n48994 ;
  assign n50544 = n50473 ^ n49801 ;
  assign n50542 = n50541 ^ n49801 ;
  assign n50543 = n50478 & n50542 ;
  assign n50545 = n50544 ^ n50543 ;
  assign n50474 = n50156 ^ n50150 ;
  assign n50621 = n50545 ^ n50474 ;
  assign n50622 = n50621 ^ n47724 ;
  assign n50771 = n50677 ^ n50622 ;
  assign n50746 = n50644 ^ n47765 ;
  assign n50747 = n50746 ^ n50645 ;
  assign n50748 = n50637 ^ n47771 ;
  assign n50749 = n50748 ^ n50640 ;
  assign n50386 = n50385 ^ n50353 ;
  assign n50226 = n50225 ^ n47596 ;
  assign n50255 = n50254 ^ n50226 ;
  assign n50263 = n50262 ^ n47685 ;
  assign n50297 = n50296 ^ n50263 ;
  assign n50306 = n50255 & ~n50297 ;
  assign n50342 = n50341 ^ n50310 ;
  assign n50387 = ~n50306 & n50342 ;
  assign n50750 = ~n50386 & ~n50387 ;
  assign n50751 = n50749 & ~n50750 ;
  assign n50752 = ~n50747 & ~n50751 ;
  assign n50753 = n50652 ^ n47696 ;
  assign n50754 = n50752 & n50753 ;
  assign n50755 = n50657 ^ n47757 ;
  assign n50756 = n50754 & ~n50755 ;
  assign n50757 = n50659 ^ n50634 ;
  assign n50758 = ~n50756 & n50757 ;
  assign n50759 = n50662 ^ n50632 ;
  assign n50760 = n50758 & ~n50759 ;
  assign n50761 = n50665 ^ n47743 ;
  assign n50762 = n50761 ^ n50629 ;
  assign n50763 = n50760 & ~n50762 ;
  assign n50764 = n50668 ^ n50628 ;
  assign n50765 = n50763 & n50764 ;
  assign n50766 = n50671 ^ n50626 ;
  assign n50767 = n50765 & n50766 ;
  assign n50768 = n50674 ^ n47730 ;
  assign n50769 = n50768 ^ n50623 ;
  assign n50770 = ~n50767 & ~n50769 ;
  assign n50857 = n50771 ^ n50770 ;
  assign n50861 = n50860 ^ n50857 ;
  assign n50865 = n50769 ^ n50767 ;
  assign n50862 = n48665 ^ n40884 ;
  assign n50863 = n50862 ^ n45137 ;
  assign n50864 = n50863 ^ n39246 ;
  assign n50866 = n50865 ^ n50864 ;
  assign n50867 = n48670 ^ n40889 ;
  assign n50868 = n50867 ^ n45142 ;
  assign n50869 = n50868 ^ n39251 ;
  assign n50941 = n50869 ^ n50865 ;
  assign n50870 = n50766 ^ n50765 ;
  assign n50871 = n50870 ^ n50869 ;
  assign n50875 = n50764 ^ n50763 ;
  assign n50872 = n48675 ^ n40895 ;
  assign n50873 = n50872 ^ n45146 ;
  assign n50874 = n50873 ^ n39255 ;
  assign n50876 = n50875 ^ n50874 ;
  assign n50878 = n48681 ^ n40902 ;
  assign n50879 = n50878 ^ n45151 ;
  assign n50880 = n50879 ^ n39261 ;
  assign n50935 = n50880 ^ n50874 ;
  assign n50877 = n50762 ^ n50760 ;
  assign n50881 = n50880 ^ n50877 ;
  assign n50885 = n50759 ^ n50758 ;
  assign n50882 = n48686 ^ n40906 ;
  assign n50883 = n50882 ^ n45156 ;
  assign n50884 = n50883 ^ n2315 ;
  assign n50886 = n50885 ^ n50884 ;
  assign n50888 = n48691 ^ n40911 ;
  assign n50889 = n50888 ^ n2201 ;
  assign n50890 = n50889 ^ n39268 ;
  assign n50929 = n50890 ^ n50884 ;
  assign n50887 = n50757 ^ n50756 ;
  assign n50891 = n50890 ^ n50887 ;
  assign n50895 = n50755 ^ n50754 ;
  assign n50892 = n48334 ^ n40916 ;
  assign n50893 = n50892 ^ n45165 ;
  assign n50894 = n50893 ^ n2193 ;
  assign n50896 = n50895 ^ n50894 ;
  assign n50900 = n50753 ^ n50752 ;
  assign n50897 = n47700 ^ n2072 ;
  assign n50898 = n50897 ^ n45169 ;
  assign n50899 = n50898 ^ n39274 ;
  assign n50901 = n50900 ^ n50899 ;
  assign n50905 = n50751 ^ n50747 ;
  assign n50902 = n48288 ^ n40448 ;
  assign n50903 = n50902 ^ n45177 ;
  assign n50904 = n50903 ^ n39279 ;
  assign n50906 = n50905 ^ n50904 ;
  assign n50910 = n50750 ^ n50749 ;
  assign n50907 = n48293 ^ n40424 ;
  assign n50908 = n50907 ^ n45181 ;
  assign n50909 = n50908 ^ n39296 ;
  assign n50911 = n50910 ^ n50909 ;
  assign n50389 = n48297 ^ n3089 ;
  assign n50390 = n50389 ^ n45186 ;
  assign n50391 = n50390 ^ n39284 ;
  assign n50914 = n50910 ^ n50391 ;
  assign n50388 = n50387 ^ n50386 ;
  assign n50392 = n50391 ^ n50388 ;
  assign n50343 = n50342 ^ n50306 ;
  assign n50298 = n50297 ^ n50255 ;
  assign n49808 = n49069 ^ n41244 ;
  assign n49809 = n49808 ^ n45412 ;
  assign n49810 = n49809 ^ n39714 ;
  assign n50222 = n50221 ^ n47578 ;
  assign n50223 = n49810 & n50222 ;
  assign n49805 = n48311 ^ n40367 ;
  assign n49806 = n49805 ^ n45200 ;
  assign n49807 = n49806 ^ n3194 ;
  assign n50224 = n50223 ^ n49807 ;
  assign n50256 = n50255 ^ n50223 ;
  assign n50257 = ~n50224 & n50256 ;
  assign n50258 = n50257 ^ n50255 ;
  assign n50299 = n50298 ^ n50258 ;
  assign n50300 = n48308 ^ n40372 ;
  assign n50301 = n50300 ^ n45196 ;
  assign n50302 = n50301 ^ n38754 ;
  assign n50303 = n50302 ^ n50258 ;
  assign n50304 = ~n50299 & n50303 ;
  assign n50305 = n50304 ^ n50302 ;
  assign n50344 = n50343 ^ n50305 ;
  assign n50345 = n48302 ^ n40363 ;
  assign n50346 = n50345 ^ n45192 ;
  assign n50347 = n50346 ^ n38797 ;
  assign n50348 = n50347 ^ n50305 ;
  assign n50349 = n50344 & n50348 ;
  assign n50350 = n50349 ^ n50347 ;
  assign n50912 = n50391 ^ n50350 ;
  assign n50913 = ~n50392 & n50912 ;
  assign n50915 = n50914 ^ n50913 ;
  assign n50916 = ~n50911 & ~n50915 ;
  assign n50917 = n50916 ^ n50910 ;
  assign n50918 = n50917 ^ n50904 ;
  assign n50919 = ~n50906 & ~n50918 ;
  assign n50920 = n50919 ^ n50904 ;
  assign n50921 = n50920 ^ n50899 ;
  assign n50922 = ~n50901 & ~n50921 ;
  assign n50923 = n50922 ^ n50900 ;
  assign n50924 = n50923 ^ n50894 ;
  assign n50925 = n50896 & n50924 ;
  assign n50926 = n50925 ^ n50895 ;
  assign n50927 = n50926 ^ n50890 ;
  assign n50928 = ~n50891 & n50927 ;
  assign n50930 = n50929 ^ n50928 ;
  assign n50931 = ~n50886 & ~n50930 ;
  assign n50932 = n50931 ^ n50885 ;
  assign n50933 = n50932 ^ n50877 ;
  assign n50934 = ~n50881 & ~n50933 ;
  assign n50936 = n50935 ^ n50934 ;
  assign n50937 = n50876 & ~n50936 ;
  assign n50938 = n50937 ^ n50875 ;
  assign n50939 = n50938 ^ n50869 ;
  assign n50940 = n50871 & n50939 ;
  assign n50942 = n50941 ^ n50940 ;
  assign n50943 = ~n50866 & ~n50942 ;
  assign n50944 = n50943 ^ n50865 ;
  assign n50945 = n50944 ^ n50857 ;
  assign n50946 = n50861 & n50945 ;
  assign n50948 = n50947 ^ n50946 ;
  assign n50678 = n50677 ^ n50621 ;
  assign n50679 = n50622 & n50678 ;
  assign n50680 = n50679 ^ n47724 ;
  assign n50475 = n50474 ^ n50473 ;
  assign n50546 = ~n50475 & ~n50545 ;
  assign n50547 = n50546 ^ n50474 ;
  assign n50470 = n50158 ^ n50147 ;
  assign n50468 = n49899 ^ n48475 ;
  assign n50469 = n50468 ^ n48990 ;
  assign n50471 = n50470 ^ n50469 ;
  assign n50619 = n50547 ^ n50471 ;
  assign n50620 = n50619 ^ n47718 ;
  assign n50773 = n50680 ^ n50620 ;
  assign n50772 = n50770 & ~n50771 ;
  assign n50855 = n50773 ^ n50772 ;
  assign n51306 = n50948 ^ n50855 ;
  assign n51362 = n51361 ^ n51306 ;
  assign n50434 = n50183 ^ n50099 ;
  assign n51363 = n50434 ^ n50207 ;
  assign n51364 = n51363 ^ n48969 ;
  assign n51311 = n50944 ^ n50861 ;
  assign n51365 = n51364 ^ n51311 ;
  assign n51318 = n50942 ^ n50864 ;
  assign n51409 = n51318 ^ n51311 ;
  assign n51366 = n50057 ^ n48978 ;
  assign n50430 = n50181 ^ n50103 ;
  assign n51367 = n51366 ^ n50430 ;
  assign n51368 = n51367 ^ n51318 ;
  assign n50437 = n50178 ^ n50109 ;
  assign n51369 = n50437 ^ n50043 ;
  assign n51370 = n51369 ^ n48980 ;
  assign n51323 = n50938 ^ n50871 ;
  assign n51371 = n51370 ^ n51323 ;
  assign n51328 = n50936 ^ n50875 ;
  assign n51403 = n51370 ^ n51328 ;
  assign n51372 = n50026 ^ n48984 ;
  assign n50441 = n50175 ^ n50116 ;
  assign n51373 = n51372 ^ n50441 ;
  assign n51374 = n51373 ^ n51328 ;
  assign n51377 = n50932 ^ n50881 ;
  assign n51400 = n51377 ^ n51328 ;
  assign n51375 = n49983 ^ n48990 ;
  assign n50445 = n50172 ^ n50121 ;
  assign n51376 = n51375 ^ n50445 ;
  assign n51378 = n51377 ^ n51376 ;
  assign n51386 = n50930 ^ n50885 ;
  assign n51397 = n51386 ^ n51377 ;
  assign n51071 = n50474 ^ n49012 ;
  assign n51072 = n51071 ^ n49828 ;
  assign n51070 = n50915 ^ n50909 ;
  assign n51073 = n51072 ^ n51070 ;
  assign n51151 = n50917 ^ n50906 ;
  assign n51152 = n51151 ^ n51070 ;
  assign n51153 = n51152 ^ n51151 ;
  assign n50393 = n50392 ^ n50350 ;
  assign n49802 = n49801 ^ n49016 ;
  assign n49804 = n49803 ^ n49802 ;
  assign n50394 = n50393 ^ n49804 ;
  assign n50397 = n49829 ^ n49022 ;
  assign n50399 = n50398 ^ n50397 ;
  assign n50395 = n50347 ^ n50344 ;
  assign n50400 = n50399 ^ n50395 ;
  assign n50404 = n50302 ^ n50299 ;
  assign n50402 = n50401 ^ n49026 ;
  assign n50403 = n50402 ^ n49837 ;
  assign n50405 = n50404 ^ n50403 ;
  assign n50409 = n50255 ^ n49807 ;
  assign n50410 = n50409 ^ n50223 ;
  assign n51061 = n50410 ^ n50404 ;
  assign n50406 = n49835 ^ n49028 ;
  assign n50408 = n50407 ^ n50406 ;
  assign n50411 = n50410 ^ n50408 ;
  assign n50415 = n50222 ^ n49810 ;
  assign n50413 = n50412 ^ n48351 ;
  assign n50414 = n50413 ^ n49842 ;
  assign n50416 = n50415 ^ n50414 ;
  assign n51023 = n50493 ^ n48945 ;
  assign n51024 = n51023 ^ n49846 ;
  assign n50422 = n49627 ^ n48155 ;
  assign n50423 = n50422 ^ n48889 ;
  assign n50421 = n50189 ^ n50089 ;
  assign n50424 = n50423 ^ n50421 ;
  assign n50426 = n50370 ^ n48165 ;
  assign n50427 = n50426 ^ n48843 ;
  assign n50429 = n50428 ^ n50427 ;
  assign n50431 = n49604 ^ n48975 ;
  assign n50432 = n50431 ^ n50283 ;
  assign n50433 = n50432 ^ n50430 ;
  assign n50438 = n48961 ^ n48917 ;
  assign n50439 = n50438 ^ n50232 ;
  assign n50440 = n50439 ^ n50437 ;
  assign n50442 = n50207 ^ n48965 ;
  assign n50443 = n50442 ^ n48873 ;
  assign n50444 = n50443 ^ n50441 ;
  assign n50446 = n50057 ^ n48971 ;
  assign n50447 = n50446 ^ n48835 ;
  assign n50563 = n50447 ^ n50443 ;
  assign n50448 = n50447 ^ n50445 ;
  assign n50452 = n50169 ^ n50126 ;
  assign n50449 = n50043 ^ n48784 ;
  assign n50450 = n50449 ^ n48969 ;
  assign n50453 = n50452 ^ n50450 ;
  assign n50455 = n48978 ^ n48775 ;
  assign n50456 = n50455 ^ n50026 ;
  assign n50454 = n50167 ^ n50130 ;
  assign n50457 = n50456 ^ n50454 ;
  assign n50462 = n50164 ^ n50132 ;
  assign n50460 = n49983 ^ n48583 ;
  assign n50461 = n50460 ^ n48980 ;
  assign n50463 = n50462 ^ n50461 ;
  assign n50466 = n50161 ^ n50140 ;
  assign n50464 = n48984 ^ n48565 ;
  assign n50465 = n50464 ^ n49971 ;
  assign n50467 = n50466 ^ n50465 ;
  assign n50548 = n50547 ^ n50469 ;
  assign n50549 = n50471 & n50548 ;
  assign n50550 = n50549 ^ n50470 ;
  assign n50551 = n50550 ^ n50465 ;
  assign n50552 = ~n50467 & n50551 ;
  assign n50553 = n50552 ^ n50466 ;
  assign n50554 = n50553 ^ n50461 ;
  assign n50555 = n50463 & n50554 ;
  assign n50556 = n50555 ^ n50462 ;
  assign n50458 = n50454 ^ n50450 ;
  assign n50459 = n50458 ^ n50450 ;
  assign n50557 = n50556 ^ n50459 ;
  assign n50558 = ~n50457 & n50557 ;
  assign n50559 = n50558 ^ n50458 ;
  assign n50560 = ~n50453 & ~n50559 ;
  assign n50451 = n50450 ^ n50447 ;
  assign n50561 = n50560 ^ n50451 ;
  assign n50562 = n50448 & ~n50561 ;
  assign n50564 = n50563 ^ n50562 ;
  assign n50565 = ~n50444 & ~n50564 ;
  assign n50566 = n50565 ^ n50443 ;
  assign n50567 = n50566 ^ n50437 ;
  assign n50568 = n50440 & n50567 ;
  assign n50569 = n50568 ^ n50439 ;
  assign n50435 = n50434 ^ n50430 ;
  assign n50436 = n50435 ^ n50434 ;
  assign n50570 = n50569 ^ n50436 ;
  assign n50571 = ~n50433 & n50570 ;
  assign n50572 = n50571 ^ n50435 ;
  assign n50576 = n50434 ^ n50428 ;
  assign n50573 = n48811 ^ n48162 ;
  assign n50574 = n50573 ^ n50320 ;
  assign n50575 = n50574 ^ n50428 ;
  assign n50577 = n50576 ^ n50575 ;
  assign n50578 = n50572 & ~n50577 ;
  assign n50579 = n50578 ^ n50575 ;
  assign n50580 = n50429 & ~n50579 ;
  assign n50581 = n50580 ^ n50428 ;
  assign n50425 = n50192 ^ n50084 ;
  assign n50582 = n50581 ^ n50425 ;
  assign n50583 = n50582 ^ n50421 ;
  assign n50584 = n50583 ^ n50425 ;
  assign n50585 = n50424 & ~n50584 ;
  assign n50586 = n50585 ^ n50582 ;
  assign n50418 = n49625 ^ n48238 ;
  assign n50419 = n50418 ^ n49085 ;
  assign n50590 = n50425 ^ n50419 ;
  assign n50587 = n48937 ^ n48197 ;
  assign n50588 = n50587 ^ n49631 ;
  assign n50589 = n50588 ^ n50419 ;
  assign n50591 = n50590 ^ n50589 ;
  assign n50592 = n50586 & ~n50591 ;
  assign n50593 = n50592 ^ n50589 ;
  assign n50417 = n50195 ^ n50082 ;
  assign n50602 = n50593 ^ n50417 ;
  assign n50603 = n50602 ^ n47542 ;
  assign n50721 = n50581 ^ n50424 ;
  assign n50607 = n50569 ^ n50433 ;
  assign n50608 = n50607 ^ n48228 ;
  assign n50610 = n50564 ^ n50441 ;
  assign n50611 = n50610 ^ n48143 ;
  assign n50612 = n50561 ^ n50445 ;
  assign n50613 = n50612 ^ n47931 ;
  assign n50614 = n50559 ^ n50452 ;
  assign n50615 = n50614 ^ n47830 ;
  assign n50617 = n50553 ^ n50463 ;
  assign n50618 = n50617 ^ n47710 ;
  assign n50684 = n50550 ^ n50467 ;
  assign n50681 = n50680 ^ n50619 ;
  assign n50682 = ~n50620 & ~n50681 ;
  assign n50683 = n50682 ^ n47718 ;
  assign n50685 = n50684 ^ n50683 ;
  assign n50686 = n50684 ^ n47716 ;
  assign n50687 = n50685 & ~n50686 ;
  assign n50688 = n50687 ^ n47716 ;
  assign n50689 = n50688 ^ n50617 ;
  assign n50690 = ~n50618 & ~n50689 ;
  assign n50691 = n50690 ^ n47710 ;
  assign n50616 = n50556 ^ n50457 ;
  assign n50692 = n50691 ^ n50616 ;
  assign n50693 = n50691 ^ n47706 ;
  assign n50694 = n50692 & ~n50693 ;
  assign n50695 = n50694 ^ n47706 ;
  assign n50696 = n50695 ^ n50614 ;
  assign n50697 = n50615 & ~n50696 ;
  assign n50698 = n50697 ^ n47830 ;
  assign n50699 = n50698 ^ n50612 ;
  assign n50700 = n50613 & ~n50699 ;
  assign n50701 = n50700 ^ n47931 ;
  assign n50702 = n50701 ^ n50610 ;
  assign n50703 = ~n50611 & ~n50702 ;
  assign n50704 = n50703 ^ n48143 ;
  assign n50609 = n50566 ^ n50440 ;
  assign n50705 = n50704 ^ n50609 ;
  assign n50706 = n50607 ^ n48178 ;
  assign n50707 = n50706 ^ n50607 ;
  assign n50708 = n50707 ^ n50609 ;
  assign n50709 = n50705 & n50708 ;
  assign n50710 = n50709 ^ n50706 ;
  assign n50711 = ~n50608 & ~n50710 ;
  assign n50712 = n50711 ^ n48228 ;
  assign n50606 = n50574 ^ n50572 ;
  assign n50713 = n50712 ^ n50606 ;
  assign n50714 = n50712 ^ n47399 ;
  assign n50715 = n50713 & ~n50714 ;
  assign n50716 = n50715 ^ n47399 ;
  assign n50605 = n50579 ^ n50427 ;
  assign n50717 = n50716 ^ n50605 ;
  assign n50718 = n50716 ^ n47428 ;
  assign n50719 = n50717 & ~n50718 ;
  assign n50720 = n50719 ^ n47428 ;
  assign n50722 = n50721 ^ n50720 ;
  assign n50723 = n50721 ^ n47458 ;
  assign n50724 = ~n50722 & n50723 ;
  assign n50725 = n50724 ^ n47458 ;
  assign n50604 = n50588 ^ n50586 ;
  assign n50726 = n50725 ^ n50604 ;
  assign n50727 = n50725 ^ n47502 ;
  assign n50728 = ~n50726 & ~n50727 ;
  assign n50729 = n50728 ^ n47502 ;
  assign n50730 = n50729 ^ n50602 ;
  assign n50731 = ~n50603 & n50730 ;
  assign n50732 = n50731 ^ n47542 ;
  assign n50598 = n50198 ^ n50077 ;
  assign n50596 = n49059 ^ n48259 ;
  assign n50597 = n50596 ^ n49621 ;
  assign n50599 = n50598 ^ n50597 ;
  assign n50420 = n50419 ^ n50417 ;
  assign n50594 = ~n50420 & n50593 ;
  assign n50595 = n50594 ^ n50419 ;
  assign n50600 = n50599 ^ n50595 ;
  assign n51004 = n50732 ^ n50600 ;
  assign n50734 = n50604 ^ n47502 ;
  assign n50735 = n50734 ^ n50725 ;
  assign n50736 = n50720 ^ n47458 ;
  assign n50737 = n50736 ^ n50721 ;
  assign n50738 = n50605 ^ n47428 ;
  assign n50739 = n50738 ^ n50716 ;
  assign n50740 = n50714 ^ n50606 ;
  assign n50741 = n50695 ^ n50615 ;
  assign n50742 = n50616 ^ n47706 ;
  assign n50743 = n50742 ^ n50691 ;
  assign n50744 = n50688 ^ n50618 ;
  assign n50745 = n50686 ^ n50683 ;
  assign n50774 = ~n50772 & n50773 ;
  assign n50775 = n50745 & ~n50774 ;
  assign n50776 = ~n50744 & ~n50775 ;
  assign n50777 = ~n50743 & n50776 ;
  assign n50778 = n50741 & n50777 ;
  assign n50779 = n50698 ^ n47931 ;
  assign n50780 = n50779 ^ n50612 ;
  assign n50781 = ~n50778 & ~n50780 ;
  assign n50782 = n50701 ^ n50611 ;
  assign n50783 = n50781 & n50782 ;
  assign n50784 = n50609 ^ n48178 ;
  assign n50785 = n50784 ^ n50704 ;
  assign n50786 = ~n50783 & ~n50785 ;
  assign n50787 = n50710 ^ n48228 ;
  assign n50788 = n50786 & ~n50787 ;
  assign n50789 = n50740 & ~n50788 ;
  assign n50790 = n50739 & ~n50789 ;
  assign n50791 = n50737 & ~n50790 ;
  assign n50792 = n50735 & ~n50791 ;
  assign n50793 = n50729 ^ n50603 ;
  assign n50794 = n50792 & ~n50793 ;
  assign n51018 = n51004 ^ n50794 ;
  assign n51019 = n47549 & ~n51018 ;
  assign n51011 = n50201 ^ n50067 ;
  assign n51010 = n50367 ^ n49055 ;
  assign n51012 = n51011 ^ n51010 ;
  assign n51007 = n48935 ^ n41153 ;
  assign n51008 = n51007 ^ n45408 ;
  assign n51009 = n51008 ^ n39660 ;
  assign n51013 = n51012 ^ n51009 ;
  assign n51014 = n51013 ^ n49617 ;
  assign n51015 = n51014 ^ n50597 ;
  assign n50796 = n48888 ^ n41206 ;
  assign n50797 = n50796 ^ n45429 ;
  assign n50798 = n50797 ^ n39593 ;
  assign n51016 = n51015 ^ n50798 ;
  assign n51005 = n50794 ^ n50732 ;
  assign n51006 = ~n51004 & ~n51005 ;
  assign n51017 = n51016 ^ n51006 ;
  assign n51020 = n51019 ^ n51017 ;
  assign n51002 = n50597 ^ n50595 ;
  assign n51003 = n50599 & n51002 ;
  assign n51021 = n51020 ^ n51003 ;
  assign n50601 = n50600 ^ n47549 ;
  assign n50733 = n50732 ^ n50601 ;
  assign n50795 = n50794 ^ n50733 ;
  assign n50799 = n50798 ^ n50795 ;
  assign n50801 = n48825 ^ n41212 ;
  assign n50802 = n50801 ^ n45434 ;
  assign n50803 = n50802 ^ n39597 ;
  assign n50800 = n50793 ^ n50792 ;
  assign n50804 = n50803 ^ n50800 ;
  assign n50808 = n50789 ^ n50739 ;
  assign n50805 = n48363 ^ n40839 ;
  assign n50806 = n50805 ^ n1447 ;
  assign n50807 = n50806 ^ n2813 ;
  assign n50809 = n50808 ^ n50807 ;
  assign n50813 = n50788 ^ n50740 ;
  assign n1402 = n1370 ^ n1323 ;
  assign n1430 = n1429 ^ n1402 ;
  assign n1437 = n1436 ^ n1430 ;
  assign n50814 = n50813 ^ n1437 ;
  assign n50816 = n48632 ^ n1231 ;
  assign n50817 = n50816 ^ n45090 ;
  assign n50818 = n50817 ^ n1421 ;
  assign n50815 = n50787 ^ n50786 ;
  assign n50819 = n50818 ^ n50815 ;
  assign n50820 = n50785 ^ n50783 ;
  assign n1701 = n1700 ^ n1213 ;
  assign n1717 = n1716 ^ n1701 ;
  assign n1721 = n1720 ^ n1717 ;
  assign n50821 = n50820 ^ n1721 ;
  assign n50825 = n50782 ^ n50781 ;
  assign n50822 = n48751 ^ n40851 ;
  assign n50823 = n50822 ^ n45096 ;
  assign n50824 = n50823 ^ n1711 ;
  assign n50826 = n50825 ^ n50824 ;
  assign n50828 = n48641 ^ n1674 ;
  assign n50829 = n50828 ^ n45101 ;
  assign n50830 = n50829 ^ n39212 ;
  assign n50965 = n50830 ^ n50824 ;
  assign n50827 = n50780 ^ n50778 ;
  assign n50831 = n50830 ^ n50827 ;
  assign n50835 = n50777 ^ n50741 ;
  assign n50832 = n48740 ^ n40857 ;
  assign n50833 = n50832 ^ n45106 ;
  assign n50834 = n50833 ^ n39217 ;
  assign n50836 = n50835 ^ n50834 ;
  assign n50840 = n50776 ^ n50743 ;
  assign n50837 = n48732 ^ n40862 ;
  assign n50838 = n50837 ^ n45111 ;
  assign n50839 = n50838 ^ n770 ;
  assign n50841 = n50840 ^ n50839 ;
  assign n50845 = n50775 ^ n50744 ;
  assign n50842 = n48645 ^ n2984 ;
  assign n50843 = n50842 ^ n45116 ;
  assign n50844 = n50843 ^ n39224 ;
  assign n50846 = n50845 ^ n50844 ;
  assign n50850 = n50774 ^ n50745 ;
  assign n50847 = n48650 ^ n40869 ;
  assign n50848 = n50847 ^ n45121 ;
  assign n50849 = n50848 ^ n39229 ;
  assign n50851 = n50850 ^ n50849 ;
  assign n50856 = n50855 ^ n50854 ;
  assign n50949 = ~n50856 & ~n50948 ;
  assign n50950 = n50949 ^ n50855 ;
  assign n50951 = n50950 ^ n50849 ;
  assign n50952 = n50851 & n50951 ;
  assign n50953 = n50952 ^ n50850 ;
  assign n50954 = n50953 ^ n50844 ;
  assign n50955 = n50846 & ~n50954 ;
  assign n50956 = n50955 ^ n50845 ;
  assign n50957 = n50956 ^ n50839 ;
  assign n50958 = ~n50841 & ~n50957 ;
  assign n50959 = n50958 ^ n50840 ;
  assign n50960 = n50959 ^ n50834 ;
  assign n50961 = n50836 & n50960 ;
  assign n50962 = n50961 ^ n50835 ;
  assign n50963 = n50962 ^ n50827 ;
  assign n50964 = ~n50831 & n50963 ;
  assign n50966 = n50965 ^ n50964 ;
  assign n50967 = ~n50826 & ~n50966 ;
  assign n50968 = n50967 ^ n50825 ;
  assign n50969 = n50968 ^ n1721 ;
  assign n50970 = n50821 & n50969 ;
  assign n50971 = n50970 ^ n50820 ;
  assign n50972 = n50971 ^ n50815 ;
  assign n50973 = ~n50819 & n50972 ;
  assign n50974 = n50973 ^ n50818 ;
  assign n50975 = n50974 ^ n1437 ;
  assign n50976 = n50814 & ~n50975 ;
  assign n50977 = n50976 ^ n50813 ;
  assign n50810 = n50790 ^ n50737 ;
  assign n50811 = n50810 ^ n50807 ;
  assign n50812 = n50811 ^ n50810 ;
  assign n50978 = n50977 ^ n50812 ;
  assign n50979 = ~n50809 & n50978 ;
  assign n50980 = n50979 ^ n50811 ;
  assign n50981 = n50791 ^ n50735 ;
  assign n50986 = n50981 ^ n50810 ;
  assign n50982 = n48802 ^ n40815 ;
  assign n50983 = n50982 ^ n45294 ;
  assign n50984 = n50983 ^ n39609 ;
  assign n50985 = n50984 ^ n50981 ;
  assign n50987 = n50986 ^ n50985 ;
  assign n50988 = n50980 & n50987 ;
  assign n50989 = n50988 ^ n50986 ;
  assign n50994 = n50981 ^ n50803 ;
  assign n50990 = n48810 ^ n40988 ;
  assign n50991 = n50990 ^ n45440 ;
  assign n50992 = n50991 ^ n39603 ;
  assign n50993 = n50992 ^ n50803 ;
  assign n50995 = n50994 ^ n50993 ;
  assign n50996 = ~n50989 & ~n50995 ;
  assign n50997 = n50996 ^ n50994 ;
  assign n50998 = ~n50804 & ~n50997 ;
  assign n50999 = n50998 ^ n50803 ;
  assign n51000 = n50999 ^ n50798 ;
  assign n51001 = ~n50799 & n51000 ;
  assign n51022 = n51021 ^ n51001 ;
  assign n51025 = n51024 ^ n51022 ;
  assign n51027 = n50495 ^ n49848 ;
  assign n51028 = n51027 ^ n48951 ;
  assign n51052 = n51028 ^ n51022 ;
  assign n51026 = n50999 ^ n50799 ;
  assign n51029 = n51028 ^ n51026 ;
  assign n51032 = n50505 ^ n49050 ;
  assign n51033 = n51032 ^ n48894 ;
  assign n51034 = n50984 ^ n50980 ;
  assign n51035 = n51033 & n51034 ;
  assign n51030 = n50513 ^ n48942 ;
  assign n51031 = n51030 ^ n49046 ;
  assign n51036 = n51035 ^ n51031 ;
  assign n51038 = n50992 ^ n50989 ;
  assign n51037 = n50997 ^ n50800 ;
  assign n51039 = n51038 ^ n51037 ;
  assign n51040 = n51039 ^ n51035 ;
  assign n51041 = n51040 ^ n51037 ;
  assign n51042 = n51036 & ~n51041 ;
  assign n51043 = n51042 ^ n51039 ;
  assign n51047 = n51037 ^ n51028 ;
  assign n51044 = n50501 ^ n49779 ;
  assign n51045 = n51044 ^ n48956 ;
  assign n51046 = n51045 ^ n51028 ;
  assign n51048 = n51047 ^ n51046 ;
  assign n51049 = ~n51043 & ~n51048 ;
  assign n51050 = n51049 ^ n51047 ;
  assign n51051 = ~n51029 & n51050 ;
  assign n51053 = n51052 ^ n51051 ;
  assign n51054 = ~n51025 & n51053 ;
  assign n51055 = n51054 ^ n51024 ;
  assign n51056 = n51055 ^ n50414 ;
  assign n51057 = n50416 & ~n51056 ;
  assign n51058 = n51057 ^ n50415 ;
  assign n51059 = n51058 ^ n50408 ;
  assign n51060 = n50411 & ~n51059 ;
  assign n51062 = n51061 ^ n51060 ;
  assign n51063 = n50405 & n51062 ;
  assign n51064 = n51063 ^ n50404 ;
  assign n51065 = n51064 ^ n50395 ;
  assign n51066 = ~n50400 & ~n51065 ;
  assign n50396 = n50395 ^ n50393 ;
  assign n51067 = n51066 ^ n50396 ;
  assign n51068 = ~n50394 & n51067 ;
  assign n51069 = n51068 ^ n50393 ;
  assign n51154 = n51153 ^ n51069 ;
  assign n51155 = n51073 & n51154 ;
  assign n51156 = n51155 ^ n51152 ;
  assign n51256 = n49819 ^ n49007 ;
  assign n51257 = n51256 ^ n50466 ;
  assign n51259 = n51257 ^ n51151 ;
  assign n51157 = n49821 ^ n49006 ;
  assign n51158 = n51157 ^ n50470 ;
  assign n51258 = n51257 ^ n51158 ;
  assign n51260 = n51259 ^ n51258 ;
  assign n51261 = ~n51156 & n51260 ;
  assign n51262 = n51261 ^ n51259 ;
  assign n51280 = n50923 ^ n50896 ;
  assign n51282 = n51280 ^ n51257 ;
  assign n51263 = n50920 ^ n50901 ;
  assign n51281 = n51280 ^ n51263 ;
  assign n51283 = n51282 ^ n51281 ;
  assign n51284 = n51262 & ~n51283 ;
  assign n51285 = n51284 ^ n51282 ;
  assign n51379 = n50454 ^ n49899 ;
  assign n51380 = n51379 ^ n48998 ;
  assign n51382 = n51380 ^ n51280 ;
  assign n51286 = n49815 ^ n49002 ;
  assign n51287 = n51286 ^ n50462 ;
  assign n51381 = n51380 ^ n51287 ;
  assign n51383 = n51382 ^ n51381 ;
  assign n51384 = ~n51285 & ~n51383 ;
  assign n51385 = n51384 ^ n51382 ;
  assign n51389 = n51386 ^ n51380 ;
  assign n51387 = n50926 ^ n50891 ;
  assign n51388 = n51387 ^ n51386 ;
  assign n51390 = n51389 ^ n51388 ;
  assign n51391 = ~n51385 & ~n51390 ;
  assign n51392 = n51391 ^ n51389 ;
  assign n51393 = n50452 ^ n48994 ;
  assign n51394 = n51393 ^ n49971 ;
  assign n51395 = n51394 ^ n51386 ;
  assign n51396 = ~n51392 & n51395 ;
  assign n51398 = n51397 ^ n51396 ;
  assign n51399 = n51378 & ~n51398 ;
  assign n51401 = n51400 ^ n51399 ;
  assign n51402 = ~n51374 & n51401 ;
  assign n51404 = n51403 ^ n51402 ;
  assign n51405 = ~n51371 & n51404 ;
  assign n51406 = n51405 ^ n51323 ;
  assign n51407 = n51406 ^ n51367 ;
  assign n51408 = n51368 & n51407 ;
  assign n51410 = n51409 ^ n51408 ;
  assign n51411 = ~n51365 & n51410 ;
  assign n51412 = n51411 ^ n51311 ;
  assign n51413 = n51412 ^ n51361 ;
  assign n51414 = n51362 & ~n51413 ;
  assign n51415 = n51414 ^ n51306 ;
  assign n51357 = n50283 ^ n48965 ;
  assign n51358 = n51357 ^ n50421 ;
  assign n51302 = n50950 ^ n50851 ;
  assign n51359 = n51358 ^ n51302 ;
  assign n51519 = n51415 ^ n51359 ;
  assign n51475 = n51412 ^ n51362 ;
  assign n51476 = n51475 ^ n48835 ;
  assign n51511 = n51410 ^ n51364 ;
  assign n51477 = n51406 ^ n51368 ;
  assign n51478 = n51477 ^ n48775 ;
  assign n51503 = n51404 ^ n51323 ;
  assign n51479 = n51398 ^ n51376 ;
  assign n51480 = n51479 ^ n48475 ;
  assign n51490 = n51394 ^ n51392 ;
  assign n51481 = n51387 ^ n51385 ;
  assign n51482 = n51481 ^ n48370 ;
  assign n51159 = n51158 ^ n51156 ;
  assign n51266 = n51159 ^ n48384 ;
  assign n51076 = n51067 ^ n49804 ;
  assign n51077 = n51076 ^ n48451 ;
  assign n51078 = n51064 ^ n50400 ;
  assign n51079 = n51078 ^ n48392 ;
  assign n51080 = n51058 ^ n50411 ;
  assign n51081 = n51080 ^ n48399 ;
  assign n51082 = n51055 ^ n50416 ;
  assign n51083 = n51082 ^ n48403 ;
  assign n51102 = n51053 ^ n51024 ;
  assign n51084 = n51050 ^ n51026 ;
  assign n51085 = n51084 ^ n48409 ;
  assign n51093 = n51045 ^ n51043 ;
  assign n51088 = n51038 ^ n51036 ;
  assign n51086 = n51034 ^ n51033 ;
  assign n51087 = n48341 & n51086 ;
  assign n51089 = n51088 ^ n51087 ;
  assign n51090 = n51088 ^ n48419 ;
  assign n51091 = ~n51089 & n51090 ;
  assign n51092 = n51091 ^ n48419 ;
  assign n51094 = n51093 ^ n51092 ;
  assign n51095 = n51084 ^ n48415 ;
  assign n51096 = n51095 ^ n51084 ;
  assign n51097 = n51096 ^ n51092 ;
  assign n51098 = ~n51094 & ~n51097 ;
  assign n51099 = n51098 ^ n51095 ;
  assign n51100 = ~n51085 & ~n51099 ;
  assign n51101 = n51100 ^ n48409 ;
  assign n51103 = n51102 ^ n51101 ;
  assign n51104 = n51102 ^ n48407 ;
  assign n51105 = n51103 & n51104 ;
  assign n51106 = n51105 ^ n48407 ;
  assign n51107 = n51106 ^ n51082 ;
  assign n51108 = n51083 & n51107 ;
  assign n51109 = n51108 ^ n48403 ;
  assign n51110 = n51109 ^ n51080 ;
  assign n51111 = n51081 & ~n51110 ;
  assign n51112 = n51111 ^ n48399 ;
  assign n51113 = n51112 ^ n47695 ;
  assign n51114 = n51062 ^ n50403 ;
  assign n51115 = n51114 ^ n51112 ;
  assign n51116 = ~n51113 & ~n51115 ;
  assign n51117 = n51116 ^ n47695 ;
  assign n51118 = n51117 ^ n51078 ;
  assign n51119 = ~n51079 & ~n51118 ;
  assign n51120 = n51119 ^ n48392 ;
  assign n51121 = n51120 ^ n51076 ;
  assign n51122 = ~n51077 & ~n51121 ;
  assign n51123 = n51122 ^ n48451 ;
  assign n51074 = n51073 ^ n51069 ;
  assign n51146 = n51123 ^ n51074 ;
  assign n51147 = n51123 ^ n48388 ;
  assign n51148 = ~n51146 & ~n51147 ;
  assign n51149 = n51148 ^ n48388 ;
  assign n51267 = n51159 ^ n51149 ;
  assign n51268 = ~n51266 & n51267 ;
  assign n51269 = n51268 ^ n48384 ;
  assign n51264 = n51263 ^ n51262 ;
  assign n51279 = n51269 ^ n51264 ;
  assign n51288 = n51287 ^ n51285 ;
  assign n51289 = n51288 ^ n48376 ;
  assign n51290 = n51289 ^ n51264 ;
  assign n51291 = n51290 ^ n51288 ;
  assign n51292 = n51279 & ~n51291 ;
  assign n51293 = n51292 ^ n51289 ;
  assign n51484 = n51481 ^ n48374 ;
  assign n51483 = n51481 ^ n51288 ;
  assign n51485 = n51484 ^ n51483 ;
  assign n51486 = n51293 & n51485 ;
  assign n51487 = n51486 ^ n51484 ;
  assign n51488 = n51482 & n51487 ;
  assign n51489 = n51488 ^ n48370 ;
  assign n51491 = n51490 ^ n51489 ;
  assign n51492 = n51490 ^ n48366 ;
  assign n51493 = ~n51491 & ~n51492 ;
  assign n51494 = n51493 ^ n48366 ;
  assign n51495 = n51494 ^ n51479 ;
  assign n51496 = n51480 & ~n51495 ;
  assign n51497 = n51496 ^ n48475 ;
  assign n51498 = n51497 ^ n48565 ;
  assign n51499 = n51401 ^ n51373 ;
  assign n51500 = n51499 ^ n51497 ;
  assign n51501 = n51498 & ~n51500 ;
  assign n51502 = n51501 ^ n48565 ;
  assign n51504 = n51503 ^ n51502 ;
  assign n51505 = n51503 ^ n48583 ;
  assign n51506 = ~n51504 & ~n51505 ;
  assign n51507 = n51506 ^ n48583 ;
  assign n51508 = n51507 ^ n51477 ;
  assign n51509 = n51478 & ~n51508 ;
  assign n51510 = n51509 ^ n48775 ;
  assign n51512 = n51511 ^ n51510 ;
  assign n51513 = n51511 ^ n48784 ;
  assign n51514 = ~n51512 & n51513 ;
  assign n51515 = n51514 ^ n48784 ;
  assign n51516 = n51515 ^ n51475 ;
  assign n51517 = n51476 & n51516 ;
  assign n51518 = n51517 ^ n48835 ;
  assign n51520 = n51519 ^ n51518 ;
  assign n51521 = n51519 ^ n48873 ;
  assign n51522 = ~n51520 & ~n51521 ;
  assign n51523 = n51522 ^ n48873 ;
  assign n51355 = n50953 ^ n50846 ;
  assign n51418 = n51355 ^ n51302 ;
  assign n51416 = n51415 ^ n51358 ;
  assign n51417 = n51359 & ~n51416 ;
  assign n51419 = n51418 ^ n51417 ;
  assign n51353 = n50425 ^ n50320 ;
  assign n51354 = n51353 ^ n48961 ;
  assign n51473 = n51419 ^ n51354 ;
  assign n51474 = n51473 ^ n48917 ;
  assign n51571 = n51523 ^ n51474 ;
  assign n51551 = n51494 ^ n51480 ;
  assign n51552 = n51487 ^ n48370 ;
  assign n51265 = n51264 ^ n48376 ;
  assign n51270 = n51269 ^ n51265 ;
  assign n51075 = n51074 ^ n48388 ;
  assign n51124 = n51123 ^ n51075 ;
  assign n51125 = n51106 ^ n51083 ;
  assign n51126 = n51104 ^ n51101 ;
  assign n51127 = n51087 ^ n48419 ;
  assign n51128 = n51127 ^ n51088 ;
  assign n51129 = n51093 ^ n48415 ;
  assign n51130 = n51129 ^ n51092 ;
  assign n51131 = ~n51128 & n51130 ;
  assign n51132 = n51099 ^ n48409 ;
  assign n51133 = ~n51131 & n51132 ;
  assign n51134 = ~n51126 & ~n51133 ;
  assign n51135 = ~n51125 & ~n51134 ;
  assign n51136 = n51109 ^ n51081 ;
  assign n51137 = ~n51135 & ~n51136 ;
  assign n51138 = n51114 ^ n51113 ;
  assign n51139 = n51137 & n51138 ;
  assign n51140 = n51117 ^ n51079 ;
  assign n51141 = n51139 & ~n51140 ;
  assign n51142 = n51120 ^ n48451 ;
  assign n51143 = n51142 ^ n51076 ;
  assign n51144 = ~n51141 & ~n51143 ;
  assign n51145 = n51124 & n51144 ;
  assign n51150 = n51149 ^ n48384 ;
  assign n51160 = n51159 ^ n51150 ;
  assign n51271 = n51145 & ~n51160 ;
  assign n51278 = ~n51270 & n51271 ;
  assign n51294 = n51293 ^ n48374 ;
  assign n51553 = n51278 & n51294 ;
  assign n51554 = n51552 & ~n51553 ;
  assign n51555 = n51489 ^ n48366 ;
  assign n51556 = n51555 ^ n51490 ;
  assign n51557 = n51554 & n51556 ;
  assign n51558 = ~n51551 & ~n51557 ;
  assign n51559 = n51499 ^ n51498 ;
  assign n51560 = ~n51558 & n51559 ;
  assign n51561 = n51505 ^ n51502 ;
  assign n51562 = ~n51560 & n51561 ;
  assign n51563 = n51507 ^ n51478 ;
  assign n51564 = n51562 & n51563 ;
  assign n51565 = n51513 ^ n51510 ;
  assign n51566 = n51564 & n51565 ;
  assign n51567 = n51515 ^ n51476 ;
  assign n51568 = ~n51566 & ~n51567 ;
  assign n51569 = n51521 ^ n51518 ;
  assign n51570 = n51568 & ~n51569 ;
  assign n51622 = n51571 ^ n51570 ;
  assign n51619 = n49420 ^ n1732 ;
  assign n51620 = n51619 ^ n45747 ;
  assign n51621 = n51620 ^ n1091 ;
  assign n51623 = n51622 ^ n51621 ;
  assign n51627 = n51569 ^ n51568 ;
  assign n51624 = n49425 ^ n41640 ;
  assign n51625 = n51624 ^ n965 ;
  assign n51626 = n51625 ^ n40086 ;
  assign n51628 = n51627 ^ n51626 ;
  assign n51630 = n49431 ^ n41645 ;
  assign n51631 = n51630 ^ n45755 ;
  assign n51632 = n51631 ^ n957 ;
  assign n51696 = n51632 ^ n51627 ;
  assign n51629 = n51567 ^ n51566 ;
  assign n51633 = n51632 ^ n51629 ;
  assign n51637 = n51565 ^ n51564 ;
  assign n51634 = n49436 ^ n827 ;
  assign n51635 = n51634 ^ n45760 ;
  assign n51636 = n51635 ^ n40093 ;
  assign n51638 = n51637 ^ n51636 ;
  assign n51642 = n51563 ^ n51562 ;
  assign n51639 = n49440 ^ n41652 ;
  assign n51640 = n51639 ^ n45766 ;
  assign n51641 = n51640 ^ n1616 ;
  assign n51643 = n51642 ^ n51641 ;
  assign n51644 = n49446 ^ n41657 ;
  assign n51645 = n51644 ^ n45771 ;
  assign n51646 = n51645 ^ n40100 ;
  assign n51687 = n51646 ^ n51642 ;
  assign n51647 = n51561 ^ n51560 ;
  assign n51648 = n51647 ^ n51646 ;
  assign n51652 = n51559 ^ n51558 ;
  assign n51649 = n49450 ^ n41662 ;
  assign n51650 = n51649 ^ n45775 ;
  assign n51651 = n51650 ^ n40106 ;
  assign n51653 = n51652 ^ n51651 ;
  assign n51657 = n51557 ^ n51551 ;
  assign n51681 = n51657 ^ n51652 ;
  assign n51654 = n49460 ^ n41667 ;
  assign n51655 = n51654 ^ n45780 ;
  assign n51656 = n51655 ^ n40111 ;
  assign n51658 = n51657 ^ n51656 ;
  assign n51662 = n51556 ^ n51554 ;
  assign n51678 = n51662 ^ n51656 ;
  assign n51659 = n49456 ^ n41674 ;
  assign n51660 = n51659 ^ n45787 ;
  assign n51661 = n51660 ^ n40117 ;
  assign n51663 = n51662 ^ n51661 ;
  assign n51668 = n51553 ^ n51552 ;
  assign n51664 = n49465 ^ n41679 ;
  assign n51665 = n51664 ^ n45791 ;
  assign n51666 = n51665 ^ n40122 ;
  assign n51669 = n51668 ^ n51666 ;
  assign n51296 = n49470 ^ n41684 ;
  assign n51297 = n51296 ^ n45796 ;
  assign n51298 = n51297 ^ n40126 ;
  assign n51295 = n51294 ^ n51278 ;
  assign n51299 = n51298 ^ n51295 ;
  assign n51670 = n51666 ^ n51298 ;
  assign n51671 = n51670 ^ n51666 ;
  assign n51272 = n51271 ^ n51270 ;
  assign n51253 = n49476 ^ n41689 ;
  assign n51254 = n51253 ^ n45801 ;
  assign n51255 = n51254 ^ n40131 ;
  assign n51273 = n51272 ^ n51255 ;
  assign n51161 = n51160 ^ n51145 ;
  assign n2397 = n2396 ^ n2360 ;
  assign n2431 = n2430 ^ n2397 ;
  assign n2441 = n2440 ^ n2431 ;
  assign n51162 = n51161 ^ n2441 ;
  assign n51167 = n51144 ^ n51124 ;
  assign n51163 = n49483 ^ n41695 ;
  assign n51164 = n51163 ^ n45809 ;
  assign n51165 = n51164 ^ n2422 ;
  assign n51168 = n51167 ^ n51165 ;
  assign n51172 = n51143 ^ n51141 ;
  assign n51169 = n49487 ^ n2268 ;
  assign n51170 = n51169 ^ n45813 ;
  assign n51171 = n51170 ^ n40141 ;
  assign n51173 = n51172 ^ n51171 ;
  assign n51177 = n51140 ^ n51139 ;
  assign n51244 = n51177 ^ n51172 ;
  assign n51174 = n49493 ^ n41752 ;
  assign n51175 = n51174 ^ n45819 ;
  assign n51176 = n51175 ^ n40146 ;
  assign n51178 = n51177 ^ n51176 ;
  assign n51183 = n51138 ^ n51137 ;
  assign n51179 = n49497 ^ n41702 ;
  assign n51180 = n51179 ^ n45824 ;
  assign n51181 = n51180 ^ n40151 ;
  assign n51184 = n51183 ^ n51181 ;
  assign n51188 = n51134 ^ n51125 ;
  assign n51185 = n49507 ^ n41738 ;
  assign n51186 = n51185 ^ n45833 ;
  assign n51187 = n51186 ^ n40161 ;
  assign n51189 = n51188 ^ n51187 ;
  assign n51198 = n51133 ^ n51126 ;
  assign n51195 = n48900 ^ n41712 ;
  assign n51196 = n51195 ^ n45838 ;
  assign n51197 = n51196 ^ n40185 ;
  assign n51199 = n51198 ^ n51197 ;
  assign n51201 = n48818 ^ n41717 ;
  assign n51202 = n51201 ^ n45844 ;
  assign n51203 = n51202 ^ n40165 ;
  assign n51228 = n51203 ^ n51197 ;
  assign n51200 = n51132 ^ n51131 ;
  assign n51204 = n51203 ^ n51200 ;
  assign n51208 = n51130 ^ n51128 ;
  assign n51205 = n48355 ^ n41721 ;
  assign n51206 = n51205 ^ n45848 ;
  assign n51207 = n51206 ^ n40169 ;
  assign n51209 = n51208 ^ n51207 ;
  assign n51215 = n51086 ^ n48341 ;
  assign n51216 = n49602 ^ n41838 ;
  assign n51217 = n51216 ^ n46154 ;
  assign n51218 = n51217 ^ n2684 ;
  assign n51219 = n51215 & n51218 ;
  assign n51212 = n48358 ^ n40998 ;
  assign n51213 = n51212 ^ n45852 ;
  assign n51214 = n51213 ^ n40172 ;
  assign n51220 = n51219 ^ n51214 ;
  assign n51221 = n51214 ^ n51128 ;
  assign n51222 = n51220 & n51221 ;
  assign n51223 = n51222 ^ n51219 ;
  assign n51210 = n51207 ^ n51203 ;
  assign n51211 = n51210 ^ n51203 ;
  assign n51224 = n51223 ^ n51211 ;
  assign n51225 = n51209 & n51224 ;
  assign n51226 = n51225 ^ n51210 ;
  assign n51227 = ~n51204 & n51226 ;
  assign n51229 = n51228 ^ n51227 ;
  assign n51230 = ~n51199 & ~n51229 ;
  assign n51231 = n51230 ^ n51198 ;
  assign n51232 = n51231 ^ n51187 ;
  assign n51233 = n51189 & ~n51232 ;
  assign n51190 = n49502 ^ n41708 ;
  assign n51191 = n51190 ^ n45828 ;
  assign n51192 = n51191 ^ n40155 ;
  assign n51193 = n51192 ^ n51187 ;
  assign n51234 = n51233 ^ n51193 ;
  assign n51237 = n51192 ^ n51181 ;
  assign n51235 = n51136 ^ n51135 ;
  assign n51236 = n51235 ^ n51181 ;
  assign n51238 = n51237 ^ n51236 ;
  assign n51239 = n51234 & ~n51238 ;
  assign n51240 = n51239 ^ n51237 ;
  assign n51241 = ~n51184 & n51240 ;
  assign n51182 = n51181 ^ n51176 ;
  assign n51242 = n51241 ^ n51182 ;
  assign n51243 = n51178 & ~n51242 ;
  assign n51245 = n51244 ^ n51243 ;
  assign n51246 = n51173 & n51245 ;
  assign n51247 = n51246 ^ n51172 ;
  assign n51248 = n51247 ^ n51165 ;
  assign n51249 = n51168 & n51248 ;
  assign n51166 = n51165 ^ n51161 ;
  assign n51250 = n51249 ^ n51166 ;
  assign n51251 = ~n51162 & ~n51250 ;
  assign n51252 = n51251 ^ n51161 ;
  assign n51275 = n51255 ^ n51252 ;
  assign n51276 = ~n51273 & n51275 ;
  assign n51277 = n51276 ^ n51272 ;
  assign n51672 = n51671 ^ n51277 ;
  assign n51673 = n51299 & ~n51672 ;
  assign n51674 = n51673 ^ n51670 ;
  assign n51675 = n51669 & n51674 ;
  assign n51667 = n51666 ^ n51661 ;
  assign n51676 = n51675 ^ n51667 ;
  assign n51677 = ~n51663 & ~n51676 ;
  assign n51679 = n51678 ^ n51677 ;
  assign n51680 = n51658 & n51679 ;
  assign n51682 = n51681 ^ n51680 ;
  assign n51683 = n51653 & n51682 ;
  assign n51684 = n51683 ^ n51652 ;
  assign n51685 = n51684 ^ n51646 ;
  assign n51686 = ~n51648 & n51685 ;
  assign n51688 = n51687 ^ n51686 ;
  assign n51689 = n51643 & n51688 ;
  assign n51690 = n51689 ^ n51642 ;
  assign n51691 = n51690 ^ n51636 ;
  assign n51692 = n51638 & ~n51691 ;
  assign n51693 = n51692 ^ n51637 ;
  assign n51694 = n51693 ^ n51632 ;
  assign n51695 = ~n51633 & n51694 ;
  assign n51697 = n51696 ^ n51695 ;
  assign n51698 = n51628 & n51697 ;
  assign n51699 = n51698 ^ n51627 ;
  assign n51700 = n51699 ^ n51621 ;
  assign n51701 = n51623 & ~n51700 ;
  assign n51702 = n51701 ^ n51622 ;
  assign n51572 = ~n51570 & ~n51571 ;
  assign n51524 = n51523 ^ n51473 ;
  assign n51525 = ~n51474 & ~n51524 ;
  assign n51526 = n51525 ^ n48917 ;
  assign n51356 = n51355 ^ n51354 ;
  assign n51420 = ~n51356 & ~n51419 ;
  assign n51421 = n51420 ^ n51355 ;
  assign n51351 = n50956 ^ n50841 ;
  assign n51349 = n50370 ^ n49604 ;
  assign n51350 = n51349 ^ n50417 ;
  assign n51352 = n51351 ^ n51350 ;
  assign n51471 = n51421 ^ n51352 ;
  assign n51472 = n51471 ^ n48975 ;
  assign n51550 = n51526 ^ n51472 ;
  assign n51617 = n51572 ^ n51550 ;
  assign n51614 = n49415 ^ n1747 ;
  assign n51615 = n51614 ^ n45301 ;
  assign n51616 = n51615 ^ n40079 ;
  assign n51618 = n51617 ^ n51616 ;
  assign n52219 = n51702 ^ n51618 ;
  assign n51728 = n50977 ^ n50809 ;
  assign n52218 = n51728 ^ n51011 ;
  assign n52220 = n52219 ^ n52218 ;
  assign n51319 = n51318 ^ n49899 ;
  assign n51320 = n51319 ^ n50445 ;
  assign n51316 = n51245 ^ n51171 ;
  assign n51321 = n51320 ^ n51316 ;
  assign n51325 = n51242 ^ n51177 ;
  assign n51322 = n50452 ^ n49815 ;
  assign n51324 = n51323 ^ n51322 ;
  assign n51326 = n51325 ^ n51324 ;
  assign n51330 = n51240 ^ n51183 ;
  assign n51823 = n51330 ^ n51325 ;
  assign n51327 = n50454 ^ n49819 ;
  assign n51329 = n51328 ^ n51327 ;
  assign n51331 = n51330 ^ n51329 ;
  assign n51780 = n51223 ^ n51209 ;
  assign n51334 = n51221 ^ n51219 ;
  assign n51781 = n51780 ^ n51334 ;
  assign n51332 = n51151 ^ n50398 ;
  assign n51333 = n51332 ^ n49835 ;
  assign n51335 = n51334 ^ n51333 ;
  assign n51338 = n51218 ^ n51215 ;
  assign n51336 = n51070 ^ n49842 ;
  assign n51337 = n51336 ^ n50401 ;
  assign n51339 = n51338 ^ n51337 ;
  assign n51453 = n49617 ^ n49085 ;
  assign n51454 = n51453 ^ n50295 ;
  assign n51344 = n50959 ^ n50836 ;
  assign n51342 = n50598 ^ n49627 ;
  assign n51343 = n51342 ^ n48811 ;
  assign n51345 = n51344 ^ n51343 ;
  assign n51422 = n51421 ^ n51350 ;
  assign n51423 = n51352 & n51422 ;
  assign n51424 = n51423 ^ n51351 ;
  assign n51346 = n50962 ^ n50831 ;
  assign n51347 = n51346 ^ n51344 ;
  assign n51348 = n51347 ^ n51346 ;
  assign n51425 = n51424 ^ n51348 ;
  assign n51426 = n51345 & n51425 ;
  assign n51427 = n51426 ^ n51347 ;
  assign n51428 = n50966 ^ n50825 ;
  assign n51432 = n51428 ^ n51346 ;
  assign n51429 = n49631 ^ n48843 ;
  assign n51430 = n51429 ^ n51011 ;
  assign n51431 = n51430 ^ n51428 ;
  assign n51433 = n51432 ^ n51431 ;
  assign n51434 = n51427 & ~n51433 ;
  assign n51435 = n51434 ^ n51432 ;
  assign n51436 = n50968 ^ n50821 ;
  assign n51440 = n51436 ^ n51428 ;
  assign n51437 = n49625 ^ n48889 ;
  assign n51438 = n51437 ^ n50220 ;
  assign n51439 = n51438 ^ n51436 ;
  assign n51441 = n51440 ^ n51439 ;
  assign n51442 = n51435 & n51441 ;
  assign n51443 = n51442 ^ n51440 ;
  assign n51446 = n50971 ^ n50819 ;
  assign n51448 = n51446 ^ n51436 ;
  assign n51444 = n49621 ^ n48937 ;
  assign n51445 = n51444 ^ n50249 ;
  assign n51447 = n51446 ^ n51445 ;
  assign n51449 = n51448 ^ n51447 ;
  assign n51450 = n51443 & n51449 ;
  assign n51451 = n51450 ^ n51448 ;
  assign n51464 = n51454 ^ n51451 ;
  assign n51465 = n51464 ^ n48238 ;
  assign n51540 = n51445 ^ n51443 ;
  assign n51466 = n51438 ^ n51435 ;
  assign n51467 = n51466 ^ n48155 ;
  assign n51469 = n51424 ^ n51345 ;
  assign n51470 = n51469 ^ n48162 ;
  assign n51527 = n51526 ^ n51471 ;
  assign n51528 = ~n51472 & n51527 ;
  assign n51529 = n51528 ^ n48975 ;
  assign n51530 = n51529 ^ n51469 ;
  assign n51531 = ~n51470 & ~n51530 ;
  assign n51532 = n51531 ^ n48162 ;
  assign n51468 = n51430 ^ n51427 ;
  assign n51533 = n51532 ^ n51468 ;
  assign n51534 = n51532 ^ n48165 ;
  assign n51535 = ~n51533 & n51534 ;
  assign n51536 = n51535 ^ n48165 ;
  assign n51537 = n51536 ^ n51466 ;
  assign n51538 = n51467 & n51537 ;
  assign n51539 = n51538 ^ n48155 ;
  assign n51541 = n51540 ^ n51539 ;
  assign n51542 = n51540 ^ n48197 ;
  assign n51543 = ~n51541 & n51542 ;
  assign n51544 = n51543 ^ n48197 ;
  assign n51545 = n51544 ^ n51464 ;
  assign n51546 = n51465 & n51545 ;
  assign n51547 = n51546 ^ n48238 ;
  assign n51460 = n49059 ^ n48954 ;
  assign n51461 = n51460 ^ n50339 ;
  assign n51452 = n50974 ^ n50814 ;
  assign n51456 = n51452 ^ n51446 ;
  assign n51455 = n51454 ^ n51452 ;
  assign n51457 = n51456 ^ n51455 ;
  assign n51458 = n51451 & ~n51457 ;
  assign n51459 = n51458 ^ n51456 ;
  assign n51462 = n51461 ^ n51459 ;
  assign n51725 = n51547 ^ n51462 ;
  assign n51549 = n51529 ^ n51470 ;
  assign n51573 = n51550 & n51572 ;
  assign n51574 = ~n51549 & ~n51573 ;
  assign n51575 = n51468 ^ n48165 ;
  assign n51576 = n51575 ^ n51532 ;
  assign n51577 = ~n51574 & n51576 ;
  assign n51578 = n51536 ^ n51467 ;
  assign n51579 = ~n51577 & ~n51578 ;
  assign n51580 = n51542 ^ n51539 ;
  assign n51581 = ~n51579 & ~n51580 ;
  assign n51582 = n51544 ^ n51465 ;
  assign n51583 = n51581 & ~n51582 ;
  assign n51741 = n51725 ^ n51583 ;
  assign n51742 = n48259 & n51741 ;
  assign n51735 = n49384 ^ n46091 ;
  assign n51736 = n51735 ^ n41604 ;
  assign n51737 = n51736 ^ n40340 ;
  assign n51733 = n48274 ^ n48259 ;
  assign n51729 = n49055 ^ n48949 ;
  assign n51730 = n51729 ^ n51461 ;
  assign n51731 = n51730 ^ n50382 ;
  assign n51732 = n51731 ^ n51728 ;
  assign n51734 = n51733 ^ n51732 ;
  assign n51738 = n51737 ^ n51734 ;
  assign n51585 = n49388 ^ n41608 ;
  assign n51586 = n51585 ^ n46095 ;
  assign n51587 = n51586 ^ n40284 ;
  assign n51739 = n51738 ^ n51587 ;
  assign n51726 = n51583 ^ n51462 ;
  assign n51727 = ~n51725 & ~n51726 ;
  assign n51740 = n51739 ^ n51727 ;
  assign n51743 = n51742 ^ n51740 ;
  assign n51723 = n51461 ^ n51452 ;
  assign n51724 = n51459 & ~n51723 ;
  assign n51744 = n51743 ^ n51724 ;
  assign n51463 = n51462 ^ n48259 ;
  assign n51548 = n51547 ^ n51463 ;
  assign n51584 = n51583 ^ n51548 ;
  assign n51588 = n51587 ^ n51584 ;
  assign n51590 = n49394 ^ n41614 ;
  assign n51591 = n51590 ^ n46101 ;
  assign n51592 = n51591 ^ n38845 ;
  assign n51720 = n51592 ^ n51584 ;
  assign n51589 = n51582 ^ n51581 ;
  assign n51593 = n51592 ^ n51589 ;
  assign n51597 = n51580 ^ n51579 ;
  assign n51594 = n49398 ^ n41618 ;
  assign n51595 = n51594 ^ n46105 ;
  assign n51596 = n51595 ^ n40060 ;
  assign n51598 = n51597 ^ n51596 ;
  assign n51602 = n51578 ^ n51577 ;
  assign n51599 = n49403 ^ n2858 ;
  assign n51600 = n51599 ^ n46110 ;
  assign n51601 = n51600 ^ n40065 ;
  assign n51603 = n51602 ^ n51601 ;
  assign n51607 = n51576 ^ n51574 ;
  assign n51604 = n49408 ^ n41625 ;
  assign n51605 = n51604 ^ n46116 ;
  assign n51606 = n51605 ^ n40070 ;
  assign n51608 = n51607 ^ n51606 ;
  assign n51609 = n41630 ^ n1767 ;
  assign n51610 = n51609 ^ n45940 ;
  assign n51611 = n51610 ^ n40075 ;
  assign n51708 = n51611 ^ n51607 ;
  assign n51612 = n51573 ^ n51549 ;
  assign n51613 = n51612 ^ n51611 ;
  assign n51703 = n51702 ^ n51616 ;
  assign n51704 = n51618 & ~n51703 ;
  assign n51705 = n51704 ^ n51617 ;
  assign n51706 = n51705 ^ n51611 ;
  assign n51707 = ~n51613 & n51706 ;
  assign n51709 = n51708 ^ n51707 ;
  assign n51710 = ~n51608 & ~n51709 ;
  assign n51711 = n51710 ^ n51607 ;
  assign n51712 = n51711 ^ n51601 ;
  assign n51713 = ~n51603 & n51712 ;
  assign n51714 = n51713 ^ n51602 ;
  assign n51715 = n51714 ^ n51596 ;
  assign n51716 = n51598 & n51715 ;
  assign n51717 = n51716 ^ n51597 ;
  assign n51718 = n51717 ^ n51592 ;
  assign n51719 = ~n51593 & n51718 ;
  assign n51721 = n51720 ^ n51719 ;
  assign n51722 = ~n51588 & n51721 ;
  assign n51745 = n51744 ^ n51722 ;
  assign n51340 = n50407 ^ n50393 ;
  assign n51341 = n51340 ^ n49846 ;
  assign n51746 = n51745 ^ n51341 ;
  assign n51749 = n51721 ^ n51587 ;
  assign n51771 = n51749 ^ n51745 ;
  assign n51747 = n50412 ^ n50395 ;
  assign n51748 = n51747 ^ n49848 ;
  assign n51750 = n51749 ^ n51748 ;
  assign n51752 = n50493 ^ n50404 ;
  assign n51753 = n51752 ^ n49779 ;
  assign n51751 = n51717 ^ n51593 ;
  assign n51754 = n51753 ^ n51751 ;
  assign n51757 = n50415 ^ n48894 ;
  assign n51758 = n51757 ^ n50501 ;
  assign n51759 = n51711 ^ n51603 ;
  assign n51760 = n51758 & n51759 ;
  assign n51765 = n51760 ^ n51751 ;
  assign n51755 = n50495 ^ n50410 ;
  assign n51756 = n51755 ^ n48942 ;
  assign n51761 = n51760 ^ n51756 ;
  assign n51762 = n51714 ^ n51598 ;
  assign n51763 = n51762 ^ n51760 ;
  assign n51764 = ~n51761 & ~n51763 ;
  assign n51766 = n51765 ^ n51764 ;
  assign n51767 = ~n51754 & n51766 ;
  assign n51768 = n51767 ^ n51753 ;
  assign n51769 = n51768 ^ n51748 ;
  assign n51770 = n51750 & n51769 ;
  assign n51772 = n51771 ^ n51770 ;
  assign n51773 = n51746 & ~n51772 ;
  assign n51774 = n51773 ^ n51745 ;
  assign n51775 = n51774 ^ n51337 ;
  assign n51776 = n51339 & ~n51775 ;
  assign n51777 = n51776 ^ n51338 ;
  assign n51778 = n51777 ^ n51334 ;
  assign n51779 = n51335 & ~n51778 ;
  assign n51782 = n51781 ^ n51779 ;
  assign n51786 = n49837 ^ n49801 ;
  assign n51787 = n51786 ^ n51263 ;
  assign n51783 = n51226 ^ n51200 ;
  assign n51784 = n51783 ^ n51780 ;
  assign n51785 = n51784 ^ n51783 ;
  assign n51788 = n51787 ^ n51785 ;
  assign n51789 = ~n51782 & n51788 ;
  assign n51790 = n51789 ^ n51784 ;
  assign n51791 = n51229 ^ n51198 ;
  assign n51795 = n51791 ^ n51783 ;
  assign n51792 = n50474 ^ n49829 ;
  assign n51793 = n51792 ^ n51280 ;
  assign n51794 = n51793 ^ n51791 ;
  assign n51796 = n51795 ^ n51794 ;
  assign n51797 = ~n51790 & ~n51796 ;
  assign n51798 = n51797 ^ n51795 ;
  assign n51799 = n51231 ^ n51189 ;
  assign n51803 = n51799 ^ n51791 ;
  assign n51800 = n50470 ^ n49803 ;
  assign n51801 = n51800 ^ n51387 ;
  assign n51802 = n51801 ^ n51799 ;
  assign n51804 = n51803 ^ n51802 ;
  assign n51805 = n51798 & ~n51804 ;
  assign n51806 = n51805 ^ n51803 ;
  assign n51807 = n51235 ^ n51234 ;
  assign n51811 = n51807 ^ n51799 ;
  assign n51808 = n51386 ^ n49828 ;
  assign n51809 = n51808 ^ n50466 ;
  assign n51810 = n51809 ^ n51807 ;
  assign n51812 = n51811 ^ n51810 ;
  assign n51813 = n51806 & n51812 ;
  assign n51814 = n51813 ^ n51811 ;
  assign n51818 = n51807 ^ n51330 ;
  assign n51815 = n51377 ^ n49821 ;
  assign n51816 = n51815 ^ n50462 ;
  assign n51817 = n51816 ^ n51330 ;
  assign n51819 = n51818 ^ n51817 ;
  assign n51820 = n51814 & n51819 ;
  assign n51821 = n51820 ^ n51818 ;
  assign n51822 = ~n51331 & n51821 ;
  assign n51824 = n51823 ^ n51822 ;
  assign n51825 = ~n51326 & ~n51824 ;
  assign n51826 = n51825 ^ n51325 ;
  assign n51827 = n51826 ^ n51316 ;
  assign n51828 = n51321 & n51827 ;
  assign n51314 = n51247 ^ n51168 ;
  assign n51317 = n51316 ^ n51314 ;
  assign n51829 = n51828 ^ n51317 ;
  assign n51312 = n51311 ^ n50441 ;
  assign n51313 = n51312 ^ n49971 ;
  assign n51845 = n51829 ^ n51313 ;
  assign n51945 = n51845 ^ n48994 ;
  assign n51846 = n51826 ^ n51321 ;
  assign n51847 = n51846 ^ n48998 ;
  assign n51849 = n51821 ^ n51329 ;
  assign n51850 = n51849 ^ n49007 ;
  assign n51851 = n51816 ^ n51814 ;
  assign n51852 = n51851 ^ n49006 ;
  assign n51854 = n51801 ^ n51798 ;
  assign n51855 = n51854 ^ n49016 ;
  assign n51856 = n51793 ^ n51790 ;
  assign n51857 = n51856 ^ n49022 ;
  assign n51858 = n51787 ^ n51782 ;
  assign n51859 = n51858 ^ n49026 ;
  assign n51860 = n51777 ^ n51335 ;
  assign n51861 = n51860 ^ n49028 ;
  assign n51862 = n51774 ^ n51339 ;
  assign n51863 = n51862 ^ n48351 ;
  assign n51864 = n51772 ^ n51341 ;
  assign n51865 = n51864 ^ n48945 ;
  assign n51879 = n51768 ^ n51750 ;
  assign n51866 = n51766 ^ n51753 ;
  assign n51867 = n51866 ^ n48956 ;
  assign n51870 = n51762 ^ n51761 ;
  assign n51868 = n51759 ^ n51758 ;
  assign n51869 = ~n49050 & n51868 ;
  assign n51871 = n51870 ^ n51869 ;
  assign n51872 = n51866 ^ n49046 ;
  assign n51873 = n51872 ^ n51866 ;
  assign n51874 = n51873 ^ n51869 ;
  assign n51875 = ~n51871 & ~n51874 ;
  assign n51876 = n51875 ^ n51872 ;
  assign n51877 = ~n51867 & ~n51876 ;
  assign n51878 = n51877 ^ n48956 ;
  assign n51880 = n51879 ^ n51878 ;
  assign n51881 = n51879 ^ n48951 ;
  assign n51882 = ~n51880 & n51881 ;
  assign n51883 = n51882 ^ n48951 ;
  assign n51884 = n51883 ^ n51864 ;
  assign n51885 = ~n51865 & n51884 ;
  assign n51886 = n51885 ^ n48945 ;
  assign n51887 = n51886 ^ n51862 ;
  assign n51888 = ~n51863 & ~n51887 ;
  assign n51889 = n51888 ^ n48351 ;
  assign n51890 = n51889 ^ n51860 ;
  assign n51891 = ~n51861 & n51890 ;
  assign n51892 = n51891 ^ n49028 ;
  assign n51893 = n51892 ^ n51858 ;
  assign n51894 = n51859 & ~n51893 ;
  assign n51895 = n51894 ^ n49026 ;
  assign n51896 = n51895 ^ n51856 ;
  assign n51897 = ~n51857 & ~n51896 ;
  assign n51898 = n51897 ^ n49022 ;
  assign n51899 = n51898 ^ n51854 ;
  assign n51900 = ~n51855 & ~n51899 ;
  assign n51901 = n51900 ^ n49016 ;
  assign n51853 = n51809 ^ n51806 ;
  assign n51902 = n51901 ^ n51853 ;
  assign n51903 = n51901 ^ n49012 ;
  assign n51904 = ~n51902 & ~n51903 ;
  assign n51905 = n51904 ^ n49012 ;
  assign n51906 = n51905 ^ n51851 ;
  assign n51907 = ~n51852 & n51906 ;
  assign n51908 = n51907 ^ n49006 ;
  assign n51909 = n51908 ^ n51849 ;
  assign n51910 = ~n51850 & ~n51909 ;
  assign n51911 = n51910 ^ n49007 ;
  assign n51848 = n51824 ^ n51324 ;
  assign n51912 = n51911 ^ n51848 ;
  assign n51913 = n51911 ^ n49002 ;
  assign n51914 = n51912 & n51913 ;
  assign n51915 = n51914 ^ n49002 ;
  assign n51916 = n51915 ^ n51846 ;
  assign n51917 = ~n51847 & n51916 ;
  assign n51918 = n51917 ^ n48998 ;
  assign n51946 = n51945 ^ n51918 ;
  assign n51947 = n51915 ^ n51847 ;
  assign n51948 = n51848 ^ n49002 ;
  assign n51949 = n51948 ^ n51911 ;
  assign n51950 = n51853 ^ n49012 ;
  assign n51951 = n51950 ^ n51901 ;
  assign n51952 = n51869 ^ n49046 ;
  assign n51953 = n51952 ^ n51870 ;
  assign n51954 = n51876 ^ n48956 ;
  assign n51955 = n51953 & ~n51954 ;
  assign n51956 = n51881 ^ n51878 ;
  assign n51957 = ~n51955 & n51956 ;
  assign n51958 = n51883 ^ n51865 ;
  assign n51959 = ~n51957 & n51958 ;
  assign n51960 = n51886 ^ n51863 ;
  assign n51961 = ~n51959 & ~n51960 ;
  assign n51962 = n51889 ^ n51861 ;
  assign n51963 = ~n51961 & ~n51962 ;
  assign n51964 = n51892 ^ n51859 ;
  assign n51965 = n51963 & n51964 ;
  assign n51966 = n51895 ^ n51857 ;
  assign n51967 = n51965 & ~n51966 ;
  assign n51968 = n51898 ^ n51855 ;
  assign n51969 = ~n51967 & ~n51968 ;
  assign n51970 = n51951 & n51969 ;
  assign n51971 = n51905 ^ n51852 ;
  assign n51972 = n51970 & ~n51971 ;
  assign n51973 = n51908 ^ n51850 ;
  assign n51974 = n51972 & ~n51973 ;
  assign n51975 = n51949 & n51974 ;
  assign n51976 = ~n51947 & ~n51975 ;
  assign n51977 = n51946 & n51976 ;
  assign n51919 = n51918 ^ n51845 ;
  assign n51920 = n51918 ^ n48994 ;
  assign n51921 = ~n51919 & n51920 ;
  assign n51922 = n51921 ^ n48994 ;
  assign n51315 = n51314 ^ n51313 ;
  assign n51830 = ~n51315 & n51829 ;
  assign n51831 = n51830 ^ n51314 ;
  assign n51309 = n51250 ^ n2441 ;
  assign n51307 = n51306 ^ n50437 ;
  assign n51308 = n51307 ^ n49983 ;
  assign n51310 = n51309 ^ n51308 ;
  assign n51843 = n51831 ^ n51310 ;
  assign n51844 = n51843 ^ n48990 ;
  assign n51978 = n51922 ^ n51844 ;
  assign n51979 = ~n51977 & ~n51978 ;
  assign n51923 = n51922 ^ n51843 ;
  assign n51924 = n51844 & ~n51923 ;
  assign n51925 = n51924 ^ n48990 ;
  assign n51832 = n51831 ^ n51308 ;
  assign n51833 = ~n51310 & ~n51832 ;
  assign n51834 = n51833 ^ n51309 ;
  assign n51303 = n51302 ^ n50430 ;
  assign n51304 = n51303 ^ n50026 ;
  assign n51274 = n51273 ^ n51252 ;
  assign n51305 = n51304 ^ n51274 ;
  assign n51841 = n51834 ^ n51305 ;
  assign n51842 = n51841 ^ n48984 ;
  assign n51980 = n51925 ^ n51842 ;
  assign n51981 = ~n51979 & ~n51980 ;
  assign n51838 = n50434 ^ n50043 ;
  assign n51839 = n51838 ^ n51355 ;
  assign n51835 = n51834 ^ n51274 ;
  assign n51836 = ~n51305 & ~n51835 ;
  assign n51300 = n51299 ^ n51277 ;
  assign n51301 = n51300 ^ n51274 ;
  assign n51837 = n51836 ^ n51301 ;
  assign n51840 = n51839 ^ n51837 ;
  assign n51943 = n51840 ^ n48980 ;
  assign n51926 = n51925 ^ n51841 ;
  assign n51927 = ~n51842 & n51926 ;
  assign n51928 = n51927 ^ n48984 ;
  assign n51944 = n51943 ^ n51928 ;
  assign n52030 = n51981 ^ n51944 ;
  assign n52026 = n50114 ^ n42488 ;
  assign n52027 = n52026 ^ n46373 ;
  assign n52028 = n52027 ^ n2984 ;
  assign n52031 = n52030 ^ n52028 ;
  assign n52035 = n51980 ^ n51979 ;
  assign n52032 = n50119 ^ n42493 ;
  assign n52033 = n52032 ^ n46377 ;
  assign n52034 = n52033 ^ n40869 ;
  assign n52036 = n52035 ^ n52034 ;
  assign n52040 = n51978 ^ n51977 ;
  assign n52169 = n52040 ^ n52035 ;
  assign n52037 = n50124 ^ n42499 ;
  assign n52038 = n52037 ^ n46383 ;
  assign n52039 = n52038 ^ n40874 ;
  assign n52041 = n52040 ^ n52039 ;
  assign n52045 = n51976 ^ n51946 ;
  assign n52166 = n52045 ^ n52039 ;
  assign n52042 = n50129 ^ n42505 ;
  assign n52043 = n52042 ^ n46388 ;
  assign n52044 = n52043 ^ n40879 ;
  assign n52046 = n52045 ^ n52044 ;
  assign n52050 = n51975 ^ n51947 ;
  assign n52047 = n50135 ^ n42511 ;
  assign n52048 = n52047 ^ n46392 ;
  assign n52049 = n52048 ^ n40884 ;
  assign n52051 = n52050 ^ n52049 ;
  assign n52055 = n51974 ^ n51949 ;
  assign n52052 = n50139 ^ n42515 ;
  assign n52053 = n52052 ^ n46397 ;
  assign n52054 = n52053 ^ n40889 ;
  assign n52056 = n52055 ^ n52054 ;
  assign n52060 = n51973 ^ n51972 ;
  assign n52057 = n50144 ^ n42520 ;
  assign n52058 = n52057 ^ n46402 ;
  assign n52059 = n52058 ^ n40895 ;
  assign n52061 = n52060 ^ n52059 ;
  assign n52063 = n50150 ^ n42526 ;
  assign n52064 = n52063 ^ n46486 ;
  assign n52065 = n52064 ^ n40902 ;
  assign n52062 = n51971 ^ n51970 ;
  assign n52066 = n52065 ^ n52062 ;
  assign n52072 = n51969 ^ n51951 ;
  assign n52069 = n49800 ^ n42530 ;
  assign n52070 = n52069 ^ n46407 ;
  assign n52071 = n52070 ^ n40906 ;
  assign n52073 = n52072 ^ n52071 ;
  assign n52077 = n51968 ^ n51967 ;
  assign n52074 = n49714 ^ n42028 ;
  assign n52075 = n52074 ^ n46474 ;
  assign n52076 = n52075 ^ n40911 ;
  assign n52078 = n52077 ^ n52076 ;
  assign n52079 = n49718 ^ n41953 ;
  assign n52080 = n52079 ^ n46412 ;
  assign n52081 = n52080 ^ n40916 ;
  assign n52146 = n52081 ^ n52077 ;
  assign n52082 = n51966 ^ n51965 ;
  assign n52083 = n52082 ^ n52081 ;
  assign n52087 = n51964 ^ n51963 ;
  assign n52084 = n49724 ^ n41957 ;
  assign n52085 = n52084 ^ n46417 ;
  assign n52086 = n52085 ^ n2072 ;
  assign n52088 = n52087 ^ n52086 ;
  assign n52093 = n51962 ^ n51961 ;
  assign n52089 = n49728 ^ n41962 ;
  assign n52090 = n52089 ^ n46422 ;
  assign n52091 = n52090 ^ n40448 ;
  assign n52094 = n52093 ^ n52091 ;
  assign n52098 = n51960 ^ n51959 ;
  assign n52095 = n49733 ^ n41967 ;
  assign n52096 = n52095 ^ n46428 ;
  assign n52097 = n52096 ^ n40424 ;
  assign n52099 = n52098 ^ n52097 ;
  assign n52104 = n51958 ^ n51957 ;
  assign n52100 = n49738 ^ n41991 ;
  assign n52101 = n52100 ^ n46433 ;
  assign n52102 = n52101 ^ n3089 ;
  assign n52105 = n52104 ^ n52102 ;
  assign n52107 = n49744 ^ n41972 ;
  assign n52108 = n52107 ^ n46438 ;
  assign n52109 = n52108 ^ n40363 ;
  assign n52106 = n51956 ^ n51955 ;
  assign n52110 = n52109 ^ n52106 ;
  assign n52114 = n51954 ^ n51953 ;
  assign n52111 = n49748 ^ n41976 ;
  assign n52112 = n52111 ^ n46442 ;
  assign n52113 = n52112 ^ n40372 ;
  assign n52115 = n52114 ^ n52113 ;
  assign n52119 = n51868 ^ n49050 ;
  assign n52120 = n50366 ^ n42610 ;
  assign n52121 = n52120 ^ n46869 ;
  assign n52122 = n52121 ^ n41244 ;
  assign n52123 = ~n52119 & n52122 ;
  assign n52116 = n49752 ^ n2732 ;
  assign n52117 = n52116 ^ n46446 ;
  assign n52118 = n52117 ^ n40367 ;
  assign n52124 = n52123 ^ n52118 ;
  assign n52125 = n52123 ^ n51953 ;
  assign n52126 = ~n52124 & n52125 ;
  assign n52127 = n52126 ^ n51953 ;
  assign n52128 = n52127 ^ n52113 ;
  assign n52129 = n52115 & ~n52128 ;
  assign n52130 = n52129 ^ n52114 ;
  assign n52131 = n52130 ^ n52106 ;
  assign n52132 = ~n52110 & n52131 ;
  assign n52133 = n52132 ^ n52109 ;
  assign n52134 = n52133 ^ n52102 ;
  assign n52135 = n52105 & n52134 ;
  assign n52103 = n52102 ^ n52098 ;
  assign n52136 = n52135 ^ n52103 ;
  assign n52137 = n52099 & n52136 ;
  assign n52138 = n52137 ^ n52098 ;
  assign n52139 = n52138 ^ n52091 ;
  assign n52140 = ~n52094 & n52139 ;
  assign n52092 = n52091 ^ n52087 ;
  assign n52141 = n52140 ^ n52092 ;
  assign n52142 = ~n52088 & ~n52141 ;
  assign n52143 = n52142 ^ n52087 ;
  assign n52144 = n52143 ^ n52081 ;
  assign n52145 = n52083 & ~n52144 ;
  assign n52147 = n52146 ^ n52145 ;
  assign n52148 = n52078 & n52147 ;
  assign n52149 = n52148 ^ n52077 ;
  assign n52150 = n52149 ^ n52071 ;
  assign n52151 = n52073 & ~n52150 ;
  assign n52152 = n52151 ^ n52072 ;
  assign n52153 = n52152 ^ n52065 ;
  assign n52154 = ~n52066 & n52153 ;
  assign n52067 = n52065 ^ n52060 ;
  assign n52155 = n52154 ^ n52067 ;
  assign n52156 = ~n52061 & ~n52155 ;
  assign n52157 = n52156 ^ n52060 ;
  assign n52158 = n52157 ^ n52054 ;
  assign n52159 = n52056 & n52158 ;
  assign n52160 = n52159 ^ n52055 ;
  assign n52161 = n52160 ^ n52049 ;
  assign n52162 = ~n52051 & ~n52161 ;
  assign n52163 = n52162 ^ n52050 ;
  assign n52164 = n52163 ^ n52044 ;
  assign n52165 = ~n52046 & n52164 ;
  assign n52167 = n52166 ^ n52165 ;
  assign n52168 = n52041 & n52167 ;
  assign n52170 = n52169 ^ n52168 ;
  assign n52171 = ~n52036 & ~n52170 ;
  assign n52172 = n52171 ^ n52035 ;
  assign n52173 = n52172 ^ n52028 ;
  assign n52174 = ~n52031 & ~n52173 ;
  assign n51982 = n51944 & ~n51981 ;
  assign n51938 = n51674 ^ n51668 ;
  assign n51936 = n50428 ^ n50057 ;
  assign n51937 = n51936 ^ n51351 ;
  assign n51939 = n51938 ^ n51937 ;
  assign n51933 = n51839 ^ n51300 ;
  assign n51934 = ~n51837 & n51933 ;
  assign n51935 = n51934 ^ n51300 ;
  assign n51940 = n51939 ^ n51935 ;
  assign n51941 = n51940 ^ n48978 ;
  assign n51929 = n51928 ^ n51840 ;
  assign n51930 = n51928 ^ n48980 ;
  assign n51931 = n51929 & n51930 ;
  assign n51932 = n51931 ^ n48980 ;
  assign n51942 = n51941 ^ n51932 ;
  assign n52024 = n51982 ^ n51942 ;
  assign n52029 = n52028 ^ n52024 ;
  assign n52175 = n52174 ^ n52029 ;
  assign n52021 = n50107 ^ n42483 ;
  assign n52022 = n52021 ^ n45945 ;
  assign n52023 = n52022 ^ n40862 ;
  assign n52217 = n52175 ^ n52023 ;
  assign n52221 = n52220 ^ n52217 ;
  assign n52226 = n52172 ^ n52031 ;
  assign n52224 = n51699 ^ n51623 ;
  assign n52223 = n51452 ^ n50598 ;
  assign n52225 = n52224 ^ n52223 ;
  assign n52227 = n52226 ^ n52225 ;
  assign n52230 = n51693 ^ n51633 ;
  assign n52229 = n51436 ^ n50425 ;
  assign n52231 = n52230 ^ n52229 ;
  assign n52228 = n52167 ^ n52040 ;
  assign n52232 = n52231 ^ n52228 ;
  assign n52237 = n52163 ^ n52046 ;
  assign n52235 = n51690 ^ n51638 ;
  assign n52234 = n51428 ^ n50421 ;
  assign n52236 = n52235 ^ n52234 ;
  assign n52238 = n52237 ^ n52236 ;
  assign n52240 = n51351 ^ n50430 ;
  assign n52191 = n51682 ^ n51651 ;
  assign n52241 = n52240 ^ n52191 ;
  assign n52239 = n52155 ^ n52059 ;
  assign n52242 = n52241 ^ n52239 ;
  assign n52247 = n51355 ^ n50437 ;
  assign n52006 = n51679 ^ n51657 ;
  assign n52248 = n52247 ^ n52006 ;
  assign n52246 = n52152 ^ n52066 ;
  assign n52249 = n52248 ^ n52246 ;
  assign n52251 = n51302 ^ n50441 ;
  assign n51987 = n51676 ^ n51662 ;
  assign n52252 = n52251 ^ n51987 ;
  assign n52250 = n52149 ^ n52073 ;
  assign n52253 = n52252 ^ n52250 ;
  assign n52256 = n52147 ^ n52076 ;
  assign n52553 = n52256 ^ n52250 ;
  assign n52254 = n51306 ^ n50445 ;
  assign n52255 = n52254 ^ n51938 ;
  assign n52257 = n52256 ^ n52255 ;
  assign n52259 = n51311 ^ n50452 ;
  assign n52260 = n52259 ^ n51300 ;
  assign n52258 = n52143 ^ n52083 ;
  assign n52261 = n52260 ^ n52258 ;
  assign n52262 = n52141 ^ n52086 ;
  assign n52547 = n52262 ^ n52258 ;
  assign n52263 = n51274 ^ n50454 ;
  assign n52264 = n52263 ^ n51318 ;
  assign n52265 = n52264 ^ n52262 ;
  assign n52268 = n52138 ^ n52094 ;
  assign n52266 = n51323 ^ n50462 ;
  assign n52267 = n52266 ^ n51309 ;
  assign n52269 = n52268 ^ n52267 ;
  assign n52272 = n52136 ^ n52097 ;
  assign n52541 = n52272 ^ n52268 ;
  assign n52270 = n51328 ^ n50466 ;
  assign n52271 = n52270 ^ n51314 ;
  assign n52273 = n52272 ^ n52271 ;
  assign n52275 = n51316 ^ n50470 ;
  assign n52276 = n52275 ^ n51377 ;
  assign n52274 = n52133 ^ n52105 ;
  assign n52277 = n52276 ^ n52274 ;
  assign n52280 = n51386 ^ n50474 ;
  assign n52281 = n52280 ^ n51325 ;
  assign n52278 = n52130 ^ n52110 ;
  assign n52282 = n52281 ^ n52278 ;
  assign n52285 = n52127 ^ n52115 ;
  assign n52283 = n51387 ^ n49801 ;
  assign n52284 = n52283 ^ n51330 ;
  assign n52286 = n52285 ^ n52284 ;
  assign n52287 = n52118 ^ n51953 ;
  assign n52288 = n52287 ^ n52123 ;
  assign n52530 = n52288 ^ n52285 ;
  assign n52289 = n51807 ^ n50398 ;
  assign n52290 = n52289 ^ n51280 ;
  assign n52291 = n52290 ^ n52288 ;
  assign n52294 = n52122 ^ n52119 ;
  assign n52292 = n51799 ^ n50401 ;
  assign n52293 = n52292 ^ n51263 ;
  assign n52295 = n52294 ^ n52293 ;
  assign n52485 = n50337 ^ n42433 ;
  assign n52486 = n52485 ^ n46777 ;
  assign n52487 = n52486 ^ n41153 ;
  assign n52488 = n52487 ^ n51729 ;
  assign n52209 = n51709 ^ n51606 ;
  assign n52489 = n52488 ^ n52209 ;
  assign n52484 = n51022 ^ n50513 ;
  assign n52490 = n52489 ^ n52484 ;
  assign n52390 = n51026 ^ n48954 ;
  assign n52391 = n52390 ^ n50505 ;
  assign n52491 = n52490 ^ n52391 ;
  assign n52414 = n50276 ^ n42437 ;
  assign n52415 = n52414 ^ n46781 ;
  assign n52416 = n52415 ^ n41206 ;
  assign n52492 = n52491 ^ n52416 ;
  assign n52345 = n50382 ^ n49617 ;
  assign n52346 = n52345 ^ n51037 ;
  assign n52298 = n51452 ^ n49627 ;
  assign n52299 = n52298 ^ n50220 ;
  assign n52300 = n52299 ^ n52235 ;
  assign n52305 = n51688 ^ n51641 ;
  assign n52303 = n51446 ^ n51011 ;
  assign n52304 = n52303 ^ n50370 ;
  assign n52306 = n52305 ^ n52304 ;
  assign n52308 = n50598 ^ n50320 ;
  assign n52309 = n52308 ^ n51436 ;
  assign n52307 = n51684 ^ n51648 ;
  assign n52310 = n52309 ^ n52307 ;
  assign n52313 = n52307 ^ n52191 ;
  assign n52189 = n51428 ^ n50283 ;
  assign n52190 = n52189 ^ n50417 ;
  assign n52192 = n52191 ^ n52190 ;
  assign n52004 = n51346 ^ n50232 ;
  assign n52005 = n52004 ^ n50425 ;
  assign n52007 = n52006 ^ n52005 ;
  assign n51989 = n51938 ^ n51935 ;
  assign n51990 = n51939 & ~n51989 ;
  assign n51988 = n51987 ^ n51938 ;
  assign n51991 = n51990 ^ n51988 ;
  assign n51992 = n51344 ^ n50207 ;
  assign n51993 = n51992 ^ n50421 ;
  assign n52001 = n51993 ^ n51987 ;
  assign n52002 = ~n51991 & n52001 ;
  assign n52003 = n52002 ^ n51987 ;
  assign n52186 = n52005 ^ n52003 ;
  assign n52187 = ~n52007 & n52186 ;
  assign n52188 = n52187 ^ n52006 ;
  assign n52311 = n52191 ^ n52188 ;
  assign n52312 = ~n52192 & ~n52311 ;
  assign n52314 = n52313 ^ n52312 ;
  assign n52315 = n52310 & n52314 ;
  assign n52316 = n52315 ^ n52309 ;
  assign n52317 = n52316 ^ n52304 ;
  assign n52318 = ~n52306 & ~n52317 ;
  assign n52319 = n52318 ^ n52305 ;
  assign n52301 = n52235 ^ n52230 ;
  assign n52302 = n52301 ^ n52230 ;
  assign n52320 = n52319 ^ n52302 ;
  assign n52321 = n52300 & n52320 ;
  assign n52322 = n52321 ^ n52301 ;
  assign n52325 = n51697 ^ n51626 ;
  assign n52327 = n52325 ^ n52230 ;
  assign n52323 = n51728 ^ n49631 ;
  assign n52324 = n52323 ^ n50249 ;
  assign n52326 = n52325 ^ n52324 ;
  assign n52328 = n52327 ^ n52326 ;
  assign n52329 = ~n52322 & ~n52328 ;
  assign n52330 = n52329 ^ n52327 ;
  assign n52334 = n52325 ^ n52224 ;
  assign n52331 = n51034 ^ n50295 ;
  assign n52332 = n52331 ^ n49625 ;
  assign n52333 = n52332 ^ n52224 ;
  assign n52335 = n52334 ^ n52333 ;
  assign n52336 = ~n52330 & n52335 ;
  assign n52337 = n52336 ^ n52334 ;
  assign n52341 = n52224 ^ n52219 ;
  assign n52338 = n51038 ^ n50339 ;
  assign n52339 = n52338 ^ n49621 ;
  assign n52340 = n52339 ^ n52219 ;
  assign n52342 = n52341 ^ n52340 ;
  assign n52343 = n52337 & n52342 ;
  assign n52344 = n52343 ^ n52341 ;
  assign n52347 = n52346 ^ n52344 ;
  assign n52395 = n52347 ^ n49085 ;
  assign n52348 = n52339 ^ n52337 ;
  assign n52349 = n52348 ^ n48937 ;
  assign n52350 = n52332 ^ n52330 ;
  assign n52351 = n52350 ^ n48889 ;
  assign n52353 = n52319 ^ n52300 ;
  assign n52354 = n52353 ^ n48811 ;
  assign n52359 = n52314 ^ n52309 ;
  assign n52193 = n52192 ^ n52188 ;
  assign n52194 = n52193 ^ n48965 ;
  assign n52008 = n52007 ^ n52003 ;
  assign n52009 = n52008 ^ n48971 ;
  assign n51994 = n51993 ^ n51991 ;
  assign n51995 = n51994 ^ n48969 ;
  assign n51984 = n51940 ^ n51932 ;
  assign n51985 = n51941 & ~n51984 ;
  assign n51986 = n51985 ^ n48978 ;
  assign n51998 = n51994 ^ n51986 ;
  assign n51999 = ~n51995 & n51998 ;
  assign n52000 = n51999 ^ n48969 ;
  assign n52183 = n52008 ^ n52000 ;
  assign n52184 = ~n52009 & n52183 ;
  assign n52185 = n52184 ^ n48971 ;
  assign n52356 = n52193 ^ n52185 ;
  assign n52357 = ~n52194 & n52356 ;
  assign n52358 = n52357 ^ n48965 ;
  assign n52360 = n52359 ^ n52358 ;
  assign n52361 = n52359 ^ n48961 ;
  assign n52362 = n52360 & n52361 ;
  assign n52363 = n52362 ^ n48961 ;
  assign n52355 = n52316 ^ n52306 ;
  assign n52364 = n52363 ^ n52355 ;
  assign n52365 = n52363 ^ n49604 ;
  assign n52366 = ~n52364 & n52365 ;
  assign n52367 = n52366 ^ n49604 ;
  assign n52368 = n52367 ^ n52353 ;
  assign n52369 = ~n52354 & ~n52368 ;
  assign n52370 = n52369 ^ n48811 ;
  assign n52352 = n52324 ^ n52322 ;
  assign n52371 = n52370 ^ n52352 ;
  assign n52372 = n52370 ^ n48843 ;
  assign n52373 = ~n52371 & ~n52372 ;
  assign n52374 = n52373 ^ n48843 ;
  assign n52375 = n52374 ^ n52350 ;
  assign n52376 = n52351 & n52375 ;
  assign n52377 = n52376 ^ n48889 ;
  assign n52378 = n52377 ^ n52348 ;
  assign n52379 = ~n52349 & n52378 ;
  assign n52380 = n52379 ^ n48937 ;
  assign n52396 = n52395 ^ n52380 ;
  assign n52397 = n52361 ^ n52358 ;
  assign n52195 = n52194 ^ n52185 ;
  assign n51983 = ~n51942 & n51982 ;
  assign n51996 = n51995 ^ n51986 ;
  assign n51997 = n51983 & n51996 ;
  assign n52010 = n52009 ^ n52000 ;
  assign n52196 = ~n51997 & ~n52010 ;
  assign n52398 = ~n52195 & n52196 ;
  assign n52399 = ~n52397 & ~n52398 ;
  assign n52400 = n52355 ^ n49604 ;
  assign n52401 = n52400 ^ n52363 ;
  assign n52402 = n52399 & n52401 ;
  assign n52403 = n52367 ^ n52354 ;
  assign n52404 = ~n52402 & n52403 ;
  assign n52405 = n52352 ^ n48843 ;
  assign n52406 = n52405 ^ n52370 ;
  assign n52407 = ~n52404 & n52406 ;
  assign n52408 = n52374 ^ n52351 ;
  assign n52409 = ~n52407 & ~n52408 ;
  assign n52410 = n52377 ^ n52349 ;
  assign n52411 = ~n52409 & n52410 ;
  assign n52412 = ~n52396 & n52411 ;
  assign n52213 = n51705 ^ n51613 ;
  assign n52386 = n52346 ^ n52213 ;
  assign n52385 = n52219 ^ n52213 ;
  assign n52387 = n52386 ^ n52385 ;
  assign n52388 = n52344 & n52387 ;
  assign n52389 = n52388 ^ n52385 ;
  assign n52392 = n52391 ^ n52389 ;
  assign n52478 = n52412 ^ n52392 ;
  assign n52381 = n52380 ^ n52347 ;
  assign n52382 = n52380 ^ n49085 ;
  assign n52383 = n52381 & ~n52382 ;
  assign n52384 = n52383 ^ n49085 ;
  assign n52481 = n52412 ^ n52384 ;
  assign n52482 = n52478 & ~n52481 ;
  assign n52479 = n52478 ^ n52384 ;
  assign n52480 = ~n49059 & n52479 ;
  assign n52483 = n52482 ^ n52480 ;
  assign n52493 = n52492 ^ n52483 ;
  assign n52476 = n52391 ^ n52213 ;
  assign n52477 = n52389 & ~n52476 ;
  assign n52494 = n52493 ^ n52477 ;
  assign n52393 = n52392 ^ n49059 ;
  assign n52394 = n52393 ^ n52384 ;
  assign n52413 = n52412 ^ n52394 ;
  assign n52417 = n52416 ^ n52413 ;
  assign n52418 = n50248 ^ n42442 ;
  assign n52419 = n52418 ^ n46786 ;
  assign n52420 = n52419 ^ n41212 ;
  assign n52473 = n52420 ^ n52413 ;
  assign n52421 = n52411 ^ n52396 ;
  assign n52422 = n52421 ^ n52420 ;
  assign n52426 = n52410 ^ n52409 ;
  assign n52423 = n50070 ^ n42447 ;
  assign n52424 = n52423 ^ n46792 ;
  assign n52425 = n52424 ^ n40988 ;
  assign n52427 = n52426 ^ n52425 ;
  assign n52429 = n50066 ^ n42453 ;
  assign n52430 = n52429 ^ n46797 ;
  assign n52431 = n52430 ^ n40815 ;
  assign n52467 = n52431 ^ n52426 ;
  assign n52428 = n52408 ^ n52407 ;
  assign n52432 = n52431 ^ n52428 ;
  assign n52436 = n52406 ^ n52404 ;
  assign n52433 = n50075 ^ n42458 ;
  assign n52434 = n52433 ^ n1400 ;
  assign n52435 = n52434 ^ n40839 ;
  assign n52437 = n52436 ^ n52435 ;
  assign n52441 = n52403 ^ n52402 ;
  assign n52438 = n50080 ^ n42463 ;
  assign n52439 = n52438 ^ n46803 ;
  assign n52440 = n52439 ^ n1370 ;
  assign n52442 = n52441 ^ n52440 ;
  assign n52443 = n52401 ^ n52399 ;
  assign n1185 = n1184 ^ n1136 ;
  assign n1222 = n1221 ^ n1185 ;
  assign n1232 = n1231 ^ n1222 ;
  assign n52444 = n52443 ^ n1232 ;
  assign n52446 = n50087 ^ n42469 ;
  assign n52447 = n52446 ^ n46811 ;
  assign n52448 = n52447 ^ n1213 ;
  assign n52455 = n52448 ^ n52443 ;
  assign n52445 = n52398 ^ n52397 ;
  assign n52449 = n52448 ^ n52445 ;
  assign n52197 = n52196 ^ n52195 ;
  assign n52012 = n50098 ^ n42476 ;
  assign n52013 = n52012 ^ n46824 ;
  assign n52014 = n52013 ^ n1674 ;
  assign n52198 = n52197 ^ n52014 ;
  assign n52011 = n52010 ^ n51997 ;
  assign n52015 = n52014 ^ n52011 ;
  assign n52019 = n51996 ^ n51983 ;
  assign n52016 = n50102 ^ n1637 ;
  assign n52017 = n52016 ^ n46516 ;
  assign n52018 = n52017 ^ n40857 ;
  assign n52020 = n52019 ^ n52018 ;
  assign n52025 = n52024 ^ n52023 ;
  assign n52176 = ~n52025 & ~n52175 ;
  assign n52177 = n52176 ^ n52024 ;
  assign n52178 = n52177 ^ n52018 ;
  assign n52179 = n52020 & n52178 ;
  assign n52180 = n52179 ^ n52019 ;
  assign n52181 = n52180 ^ n52014 ;
  assign n52182 = ~n52015 & n52181 ;
  assign n52199 = n52198 ^ n52182 ;
  assign n52200 = n50092 ^ n1038 ;
  assign n52201 = n52200 ^ n1679 ;
  assign n52202 = n52201 ^ n40851 ;
  assign n52450 = n52202 ^ n52197 ;
  assign n52451 = ~n52199 & n52450 ;
  assign n52452 = n52451 ^ n52202 ;
  assign n52453 = n52452 ^ n52448 ;
  assign n52454 = n52449 & n52453 ;
  assign n52456 = n52455 ^ n52454 ;
  assign n52457 = n52444 & n52456 ;
  assign n52458 = n52457 ^ n52443 ;
  assign n52459 = n52458 ^ n52440 ;
  assign n52460 = n52442 & ~n52459 ;
  assign n52461 = n52460 ^ n52441 ;
  assign n52462 = n52461 ^ n52435 ;
  assign n52463 = ~n52437 & ~n52462 ;
  assign n52464 = n52463 ^ n52436 ;
  assign n52465 = n52464 ^ n52431 ;
  assign n52466 = ~n52432 & ~n52465 ;
  assign n52468 = n52467 ^ n52466 ;
  assign n52469 = ~n52427 & ~n52468 ;
  assign n52470 = n52469 ^ n52426 ;
  assign n52471 = n52470 ^ n52420 ;
  assign n52472 = ~n52422 & ~n52471 ;
  assign n52474 = n52473 ^ n52472 ;
  assign n52475 = ~n52417 & n52474 ;
  assign n52495 = n52494 ^ n52475 ;
  assign n52296 = n51151 ^ n50407 ;
  assign n52297 = n52296 ^ n51791 ;
  assign n52496 = n52495 ^ n52297 ;
  assign n52499 = n52474 ^ n52416 ;
  assign n52521 = n52499 ^ n52495 ;
  assign n52497 = n51070 ^ n50412 ;
  assign n52498 = n52497 ^ n51783 ;
  assign n52500 = n52499 ^ n52498 ;
  assign n52503 = n52470 ^ n52422 ;
  assign n52501 = n50493 ^ n50393 ;
  assign n52502 = n52501 ^ n51780 ;
  assign n52504 = n52503 ^ n52502 ;
  assign n52510 = n51334 ^ n50395 ;
  assign n52511 = n52510 ^ n50495 ;
  assign n52505 = n50501 ^ n50404 ;
  assign n52506 = n52505 ^ n51338 ;
  assign n52507 = n52464 ^ n52432 ;
  assign n52508 = n52506 & n52507 ;
  assign n52512 = n52511 ^ n52508 ;
  assign n52513 = n52468 ^ n52425 ;
  assign n52514 = n52513 ^ n52508 ;
  assign n52515 = n52512 & ~n52514 ;
  assign n52509 = n52508 ^ n52503 ;
  assign n52516 = n52515 ^ n52509 ;
  assign n52517 = n52504 & n52516 ;
  assign n52518 = n52517 ^ n52503 ;
  assign n52519 = n52518 ^ n52498 ;
  assign n52520 = ~n52500 & ~n52519 ;
  assign n52522 = n52521 ^ n52520 ;
  assign n52523 = n52496 & n52522 ;
  assign n52524 = n52523 ^ n52495 ;
  assign n52525 = n52524 ^ n52293 ;
  assign n52526 = ~n52295 & n52525 ;
  assign n52527 = n52526 ^ n52294 ;
  assign n52528 = n52527 ^ n52288 ;
  assign n52529 = n52291 & ~n52528 ;
  assign n52531 = n52530 ^ n52529 ;
  assign n52532 = n52286 & n52531 ;
  assign n52533 = n52532 ^ n52285 ;
  assign n52534 = n52533 ^ n52278 ;
  assign n52535 = ~n52282 & ~n52534 ;
  assign n52279 = n52278 ^ n52274 ;
  assign n52536 = n52535 ^ n52279 ;
  assign n52537 = n52277 & n52536 ;
  assign n52538 = n52537 ^ n52276 ;
  assign n52539 = n52538 ^ n52272 ;
  assign n52540 = n52273 & n52539 ;
  assign n52542 = n52541 ^ n52540 ;
  assign n52543 = ~n52269 & ~n52542 ;
  assign n52544 = n52543 ^ n52268 ;
  assign n52545 = n52544 ^ n52262 ;
  assign n52546 = ~n52265 & n52545 ;
  assign n52548 = n52547 ^ n52546 ;
  assign n52549 = n52261 & ~n52548 ;
  assign n52550 = n52549 ^ n52260 ;
  assign n52551 = n52550 ^ n52256 ;
  assign n52552 = n52257 & ~n52551 ;
  assign n52554 = n52553 ^ n52552 ;
  assign n52555 = ~n52253 & ~n52554 ;
  assign n52556 = n52555 ^ n52252 ;
  assign n52557 = n52556 ^ n52246 ;
  assign n52558 = ~n52249 & ~n52557 ;
  assign n52559 = n52558 ^ n52248 ;
  assign n52243 = n52157 ^ n52056 ;
  assign n52244 = n52243 ^ n52239 ;
  assign n52245 = n52244 ^ n52243 ;
  assign n52560 = n52559 ^ n52245 ;
  assign n52561 = ~n52242 & ~n52560 ;
  assign n52562 = n52561 ^ n52244 ;
  assign n52563 = n52160 ^ n52051 ;
  assign n52567 = n52563 ^ n52243 ;
  assign n52564 = n51344 ^ n50434 ;
  assign n52565 = n52564 ^ n52307 ;
  assign n52566 = n52565 ^ n52563 ;
  assign n52568 = n52567 ^ n52566 ;
  assign n52569 = n52562 & ~n52568 ;
  assign n52570 = n52569 ^ n52567 ;
  assign n52574 = n52563 ^ n52237 ;
  assign n52571 = n51346 ^ n50428 ;
  assign n52572 = n52571 ^ n52305 ;
  assign n52573 = n52572 ^ n52237 ;
  assign n52575 = n52574 ^ n52573 ;
  assign n52576 = n52570 & n52575 ;
  assign n52577 = n52576 ^ n52574 ;
  assign n52578 = n52238 & ~n52577 ;
  assign n52579 = n52578 ^ n52237 ;
  assign n52233 = n52170 ^ n52034 ;
  assign n52580 = n52579 ^ n52233 ;
  assign n52581 = n52580 ^ n52228 ;
  assign n52582 = n52581 ^ n52233 ;
  assign n52583 = ~n52232 & ~n52582 ;
  assign n52584 = n52583 ^ n52580 ;
  assign n52588 = n52233 ^ n52226 ;
  assign n52585 = n51446 ^ n50417 ;
  assign n52586 = n52585 ^ n52325 ;
  assign n52587 = n52586 ^ n52226 ;
  assign n52589 = n52588 ^ n52587 ;
  assign n52590 = ~n52584 & ~n52589 ;
  assign n52591 = n52590 ^ n52588 ;
  assign n52592 = n52227 & ~n52591 ;
  assign n52593 = n52592 ^ n52226 ;
  assign n52215 = n52177 ^ n52020 ;
  assign n52222 = n52217 ^ n52215 ;
  assign n52594 = n52593 ^ n52222 ;
  assign n52595 = n52594 ^ n52215 ;
  assign n52596 = n52221 & ~n52595 ;
  assign n52597 = n52596 ^ n52222 ;
  assign n52212 = n51034 ^ n50220 ;
  assign n52214 = n52213 ^ n52212 ;
  assign n52611 = n52597 ^ n52214 ;
  assign n52612 = n52611 ^ n49627 ;
  assign n52732 = n52593 ^ n52221 ;
  assign n52614 = n52579 ^ n52232 ;
  assign n52615 = n52614 ^ n50232 ;
  assign n52708 = n52572 ^ n52570 ;
  assign n52617 = n52559 ^ n52242 ;
  assign n52618 = n52617 ^ n50026 ;
  assign n52619 = n52556 ^ n52249 ;
  assign n52620 = n52619 ^ n49983 ;
  assign n52621 = n52554 ^ n52252 ;
  assign n52622 = n52621 ^ n49971 ;
  assign n52623 = n52550 ^ n52257 ;
  assign n52624 = n52623 ^ n49899 ;
  assign n52625 = n52548 ^ n52260 ;
  assign n52626 = n52625 ^ n49815 ;
  assign n52627 = n52544 ^ n52265 ;
  assign n52628 = n52627 ^ n49819 ;
  assign n52629 = n52542 ^ n52267 ;
  assign n52630 = n52629 ^ n49821 ;
  assign n52674 = n52536 ^ n52276 ;
  assign n52632 = n52533 ^ n52282 ;
  assign n52633 = n52632 ^ n49829 ;
  assign n52634 = n52531 ^ n52284 ;
  assign n52635 = n52634 ^ n49837 ;
  assign n52636 = n52527 ^ n52291 ;
  assign n52637 = n52636 ^ n49835 ;
  assign n52638 = n52524 ^ n52295 ;
  assign n52639 = n52638 ^ n49842 ;
  assign n52640 = n52522 ^ n52297 ;
  assign n52641 = n52640 ^ n49846 ;
  assign n52642 = n52518 ^ n52500 ;
  assign n52643 = n52642 ^ n49848 ;
  assign n52644 = n52516 ^ n52502 ;
  assign n52645 = n52644 ^ n49779 ;
  assign n52646 = n52507 ^ n52506 ;
  assign n52647 = n48894 & n52646 ;
  assign n52648 = n52647 ^ n48942 ;
  assign n52649 = n52513 ^ n52512 ;
  assign n52650 = n52649 ^ n52647 ;
  assign n52651 = ~n52648 & n52650 ;
  assign n52652 = n52651 ^ n48942 ;
  assign n52653 = n52652 ^ n52644 ;
  assign n52654 = ~n52645 & n52653 ;
  assign n52655 = n52654 ^ n49779 ;
  assign n52656 = n52655 ^ n52642 ;
  assign n52657 = ~n52643 & ~n52656 ;
  assign n52658 = n52657 ^ n49848 ;
  assign n52659 = n52658 ^ n52640 ;
  assign n52660 = n52641 & n52659 ;
  assign n52661 = n52660 ^ n49846 ;
  assign n52662 = n52661 ^ n52638 ;
  assign n52663 = ~n52639 & n52662 ;
  assign n52664 = n52663 ^ n49842 ;
  assign n52665 = n52664 ^ n52636 ;
  assign n52666 = n52637 & ~n52665 ;
  assign n52667 = n52666 ^ n49835 ;
  assign n52668 = n52667 ^ n52634 ;
  assign n52669 = ~n52635 & n52668 ;
  assign n52670 = n52669 ^ n49837 ;
  assign n52671 = n52670 ^ n52632 ;
  assign n52672 = ~n52633 & ~n52671 ;
  assign n52673 = n52672 ^ n49829 ;
  assign n52675 = n52674 ^ n52673 ;
  assign n52676 = n52674 ^ n49803 ;
  assign n52677 = n52675 & n52676 ;
  assign n52678 = n52677 ^ n49803 ;
  assign n52631 = n52538 ^ n52273 ;
  assign n52679 = n52678 ^ n52631 ;
  assign n52680 = n52678 ^ n49828 ;
  assign n52681 = n52679 & ~n52680 ;
  assign n52682 = n52681 ^ n49828 ;
  assign n52683 = n52682 ^ n52629 ;
  assign n52684 = ~n52630 & n52683 ;
  assign n52685 = n52684 ^ n49821 ;
  assign n52686 = n52685 ^ n52627 ;
  assign n52687 = ~n52628 & ~n52686 ;
  assign n52688 = n52687 ^ n49819 ;
  assign n52689 = n52688 ^ n52625 ;
  assign n52690 = ~n52626 & ~n52689 ;
  assign n52691 = n52690 ^ n49815 ;
  assign n52692 = n52691 ^ n52623 ;
  assign n52693 = ~n52624 & n52692 ;
  assign n52694 = n52693 ^ n49899 ;
  assign n52695 = n52694 ^ n52621 ;
  assign n52696 = n52622 & n52695 ;
  assign n52697 = n52696 ^ n49971 ;
  assign n52698 = n52697 ^ n52619 ;
  assign n52699 = n52620 & n52698 ;
  assign n52700 = n52699 ^ n49983 ;
  assign n52701 = n52700 ^ n52617 ;
  assign n52702 = n52618 & n52701 ;
  assign n52703 = n52702 ^ n50026 ;
  assign n52616 = n52565 ^ n52562 ;
  assign n52704 = n52703 ^ n52616 ;
  assign n52705 = n52703 ^ n50043 ;
  assign n52706 = n52704 & n52705 ;
  assign n52707 = n52706 ^ n50043 ;
  assign n52709 = n52708 ^ n52707 ;
  assign n52710 = n52577 ^ n52236 ;
  assign n52711 = n52710 ^ n50057 ;
  assign n52712 = n52711 ^ n52710 ;
  assign n52713 = n52712 ^ n52707 ;
  assign n52714 = ~n52709 & n52713 ;
  assign n52715 = n52714 ^ n52711 ;
  assign n52717 = n52614 ^ n50207 ;
  assign n52716 = n52710 ^ n52614 ;
  assign n52718 = n52717 ^ n52716 ;
  assign n52719 = ~n52715 & n52718 ;
  assign n52720 = n52719 ^ n52717 ;
  assign n52721 = n52615 & n52720 ;
  assign n52722 = n52721 ^ n50232 ;
  assign n52723 = n52722 ^ n50283 ;
  assign n52724 = n52586 ^ n52584 ;
  assign n52725 = n52724 ^ n52722 ;
  assign n52726 = ~n52723 & n52725 ;
  assign n52727 = n52726 ^ n50283 ;
  assign n52613 = n52591 ^ n52225 ;
  assign n52728 = n52727 ^ n52613 ;
  assign n52729 = n52727 ^ n50320 ;
  assign n52730 = ~n52728 & ~n52729 ;
  assign n52731 = n52730 ^ n50320 ;
  assign n52733 = n52732 ^ n52731 ;
  assign n52734 = n52611 ^ n50370 ;
  assign n52735 = n52734 ^ n52611 ;
  assign n52736 = n52735 ^ n52731 ;
  assign n52737 = ~n52733 & n52736 ;
  assign n52738 = n52737 ^ n52734 ;
  assign n52739 = ~n52612 & n52738 ;
  assign n52740 = n52739 ^ n49627 ;
  assign n52820 = n52740 ^ n49631 ;
  assign n52216 = n52215 ^ n52214 ;
  assign n52598 = n52216 & n52597 ;
  assign n52599 = n52598 ^ n52215 ;
  assign n52208 = n51038 ^ n50249 ;
  assign n52210 = n52209 ^ n52208 ;
  assign n52207 = n52180 ^ n52015 ;
  assign n52211 = n52210 ^ n52207 ;
  assign n52741 = n52599 ^ n52211 ;
  assign n52821 = n52820 ^ n52741 ;
  assign n52766 = n52700 ^ n52618 ;
  assign n52767 = n52682 ^ n52630 ;
  assign n52768 = n52631 ^ n49828 ;
  assign n52769 = n52768 ^ n52678 ;
  assign n52770 = n52670 ^ n52633 ;
  assign n52771 = n52652 ^ n52645 ;
  assign n52772 = n52649 ^ n52648 ;
  assign n52773 = ~n52771 & ~n52772 ;
  assign n52774 = n52655 ^ n52643 ;
  assign n52775 = ~n52773 & n52774 ;
  assign n52776 = n52658 ^ n52641 ;
  assign n52777 = ~n52775 & ~n52776 ;
  assign n52778 = n52661 ^ n52639 ;
  assign n52779 = ~n52777 & n52778 ;
  assign n52780 = n52664 ^ n52637 ;
  assign n52781 = ~n52779 & n52780 ;
  assign n52782 = n52667 ^ n52635 ;
  assign n52783 = n52781 & ~n52782 ;
  assign n52784 = ~n52770 & n52783 ;
  assign n52785 = n52676 ^ n52673 ;
  assign n52786 = ~n52784 & n52785 ;
  assign n52787 = ~n52769 & n52786 ;
  assign n52788 = ~n52767 & n52787 ;
  assign n52789 = n52685 ^ n52628 ;
  assign n52790 = n52788 & ~n52789 ;
  assign n52791 = n52688 ^ n52626 ;
  assign n52792 = n52790 & n52791 ;
  assign n52793 = n52691 ^ n52624 ;
  assign n52794 = ~n52792 & n52793 ;
  assign n52795 = n52694 ^ n52622 ;
  assign n52796 = n52794 & ~n52795 ;
  assign n52797 = n52697 ^ n52620 ;
  assign n52798 = ~n52796 & ~n52797 ;
  assign n52799 = ~n52766 & ~n52798 ;
  assign n52800 = n52616 ^ n50043 ;
  assign n52801 = n52800 ^ n52703 ;
  assign n52802 = ~n52799 & n52801 ;
  assign n52803 = n52708 ^ n50057 ;
  assign n52804 = n52803 ^ n52707 ;
  assign n52805 = n52802 & ~n52804 ;
  assign n52806 = n52715 ^ n50207 ;
  assign n52807 = n52805 & ~n52806 ;
  assign n52808 = n52720 ^ n50232 ;
  assign n52809 = ~n52807 & n52808 ;
  assign n52810 = n52724 ^ n52723 ;
  assign n52811 = n52809 & ~n52810 ;
  assign n52812 = n52613 ^ n50320 ;
  assign n52813 = n52812 ^ n52727 ;
  assign n52814 = ~n52811 & n52813 ;
  assign n52815 = n52731 ^ n50370 ;
  assign n52816 = n52815 ^ n52732 ;
  assign n52817 = n52814 & n52816 ;
  assign n52818 = n52738 ^ n49627 ;
  assign n52819 = ~n52817 & n52818 ;
  assign n52846 = n52821 ^ n52819 ;
  assign n52843 = n43371 ^ n1437 ;
  assign n52844 = n52843 ^ n47177 ;
  assign n52845 = n52844 ^ n41625 ;
  assign n52847 = n52846 ^ n52845 ;
  assign n52849 = n50818 ^ n1333 ;
  assign n52850 = n52849 ^ n47182 ;
  assign n52851 = n52850 ^ n41630 ;
  assign n52848 = n52818 ^ n52817 ;
  assign n52852 = n52851 ^ n52848 ;
  assign n1722 = n1721 ^ n1315 ;
  assign n1741 = n1740 ^ n1722 ;
  assign n1748 = n1747 ^ n1741 ;
  assign n53045 = n52848 ^ n1748 ;
  assign n52853 = n52816 ^ n52814 ;
  assign n52854 = n52853 ^ n1748 ;
  assign n52858 = n52813 ^ n52811 ;
  assign n52855 = n50824 ^ n43381 ;
  assign n52856 = n52855 ^ n47190 ;
  assign n52857 = n52856 ^ n1732 ;
  assign n52859 = n52858 ^ n52857 ;
  assign n52863 = n52810 ^ n52809 ;
  assign n52860 = n50830 ^ n1695 ;
  assign n52861 = n52860 ^ n47195 ;
  assign n52862 = n52861 ^ n41640 ;
  assign n52864 = n52863 ^ n52862 ;
  assign n52868 = n52808 ^ n52807 ;
  assign n52865 = n50834 ^ n43387 ;
  assign n52866 = n52865 ^ n47201 ;
  assign n52867 = n52866 ^ n41645 ;
  assign n52869 = n52868 ^ n52867 ;
  assign n52871 = n50839 ^ n43029 ;
  assign n52872 = n52871 ^ n47205 ;
  assign n52873 = n52872 ^ n827 ;
  assign n52870 = n52806 ^ n52805 ;
  assign n52874 = n52873 ^ n52870 ;
  assign n52878 = n52804 ^ n52802 ;
  assign n52875 = n50844 ^ n2993 ;
  assign n52876 = n52875 ^ n47210 ;
  assign n52877 = n52876 ^ n41652 ;
  assign n52879 = n52878 ^ n52877 ;
  assign n52881 = n50849 ^ n42890 ;
  assign n52882 = n52881 ^ n47216 ;
  assign n52883 = n52882 ^ n41657 ;
  assign n53027 = n52883 ^ n52878 ;
  assign n52880 = n52801 ^ n52799 ;
  assign n52884 = n52883 ^ n52880 ;
  assign n52888 = n52798 ^ n52766 ;
  assign n52885 = n50854 ^ n42894 ;
  assign n52886 = n52885 ^ n47222 ;
  assign n52887 = n52886 ^ n41662 ;
  assign n52889 = n52888 ^ n52887 ;
  assign n52893 = n52797 ^ n52796 ;
  assign n52890 = n50860 ^ n42899 ;
  assign n52891 = n52890 ^ n47228 ;
  assign n52892 = n52891 ^ n41667 ;
  assign n52894 = n52893 ^ n52892 ;
  assign n52898 = n52795 ^ n52794 ;
  assign n52895 = n50864 ^ n42904 ;
  assign n52896 = n52895 ^ n47233 ;
  assign n52897 = n52896 ^ n41674 ;
  assign n52899 = n52898 ^ n52897 ;
  assign n52903 = n52793 ^ n52792 ;
  assign n52900 = n50869 ^ n42910 ;
  assign n52901 = n52900 ^ n47238 ;
  assign n52902 = n52901 ^ n41679 ;
  assign n52904 = n52903 ^ n52902 ;
  assign n52908 = n52791 ^ n52790 ;
  assign n52905 = n50874 ^ n42917 ;
  assign n52906 = n52905 ^ n47243 ;
  assign n52907 = n52906 ^ n41684 ;
  assign n52909 = n52908 ^ n52907 ;
  assign n52913 = n52789 ^ n52788 ;
  assign n52910 = n50880 ^ n42921 ;
  assign n52911 = n52910 ^ n47247 ;
  assign n52912 = n52911 ^ n41689 ;
  assign n52914 = n52913 ^ n52912 ;
  assign n52918 = n52787 ^ n52767 ;
  assign n52915 = n50884 ^ n47253 ;
  assign n52916 = n52915 ^ n42926 ;
  assign n52917 = n52916 ^ n2396 ;
  assign n52919 = n52918 ^ n52917 ;
  assign n52923 = n52786 ^ n52769 ;
  assign n52920 = n50890 ^ n42931 ;
  assign n52921 = n52920 ^ n2279 ;
  assign n52922 = n52921 ^ n41695 ;
  assign n52924 = n52923 ^ n52922 ;
  assign n52928 = n52785 ^ n52784 ;
  assign n52925 = n50894 ^ n42936 ;
  assign n52926 = n52925 ^ n47261 ;
  assign n52927 = n52926 ^ n2268 ;
  assign n52929 = n52928 ^ n52927 ;
  assign n52930 = n50899 ^ n2132 ;
  assign n52931 = n52930 ^ n47265 ;
  assign n52932 = n52931 ^ n41752 ;
  assign n52997 = n52932 ^ n52928 ;
  assign n52933 = n52783 ^ n52770 ;
  assign n52934 = n52933 ^ n52932 ;
  assign n52938 = n52782 ^ n52781 ;
  assign n52935 = n50904 ^ n42943 ;
  assign n52936 = n52935 ^ n47271 ;
  assign n52937 = n52936 ^ n41702 ;
  assign n52939 = n52938 ^ n52937 ;
  assign n52944 = n52780 ^ n52779 ;
  assign n52940 = n50909 ^ n42947 ;
  assign n52941 = n52940 ^ n47276 ;
  assign n52942 = n52941 ^ n41708 ;
  assign n52945 = n52944 ^ n52942 ;
  assign n52949 = n52778 ^ n52777 ;
  assign n52946 = n50391 ^ n42952 ;
  assign n52947 = n52946 ^ n47281 ;
  assign n52948 = n52947 ^ n41738 ;
  assign n52950 = n52949 ^ n52948 ;
  assign n52952 = n50347 ^ n42957 ;
  assign n52953 = n52952 ^ n47285 ;
  assign n52954 = n52953 ^ n41712 ;
  assign n52986 = n52954 ^ n52949 ;
  assign n52951 = n52776 ^ n52775 ;
  assign n52955 = n52954 ^ n52951 ;
  assign n52959 = n52774 ^ n52773 ;
  assign n52956 = n50302 ^ n42962 ;
  assign n52957 = n52956 ^ n47290 ;
  assign n52958 = n52957 ^ n41717 ;
  assign n52960 = n52959 ^ n52958 ;
  assign n52964 = n52772 ^ n52771 ;
  assign n52961 = n49807 ^ n42971 ;
  assign n52962 = n52961 ^ n47300 ;
  assign n52963 = n52962 ^ n41721 ;
  assign n52965 = n52964 ^ n52963 ;
  assign n52969 = n51009 ^ n43335 ;
  assign n52970 = n52969 ^ n47535 ;
  assign n52971 = n52970 ^ n41838 ;
  assign n52972 = n52646 ^ n48894 ;
  assign n52973 = n52971 & n52972 ;
  assign n52966 = n49810 ^ n42967 ;
  assign n52967 = n52966 ^ n47296 ;
  assign n52968 = n52967 ^ n40998 ;
  assign n52974 = n52973 ^ n52968 ;
  assign n52975 = n52973 ^ n52772 ;
  assign n52976 = ~n52974 & ~n52975 ;
  assign n52977 = n52976 ^ n52772 ;
  assign n52978 = n52977 ^ n52963 ;
  assign n52979 = ~n52965 & ~n52978 ;
  assign n52980 = n52979 ^ n52963 ;
  assign n52981 = n52980 ^ n52958 ;
  assign n52982 = ~n52960 & ~n52981 ;
  assign n52983 = n52982 ^ n52959 ;
  assign n52984 = n52983 ^ n52954 ;
  assign n52985 = ~n52955 & ~n52984 ;
  assign n52987 = n52986 ^ n52985 ;
  assign n52988 = ~n52950 & ~n52987 ;
  assign n52989 = n52988 ^ n52949 ;
  assign n52990 = n52989 ^ n52942 ;
  assign n52991 = n52945 & ~n52990 ;
  assign n52943 = n52942 ^ n52938 ;
  assign n52992 = n52991 ^ n52943 ;
  assign n52993 = n52939 & n52992 ;
  assign n52994 = n52993 ^ n52938 ;
  assign n52995 = n52994 ^ n52932 ;
  assign n52996 = n52934 & n52995 ;
  assign n52998 = n52997 ^ n52996 ;
  assign n52999 = ~n52929 & ~n52998 ;
  assign n53000 = n52999 ^ n52928 ;
  assign n53001 = n53000 ^ n52922 ;
  assign n53002 = ~n52924 & n53001 ;
  assign n53003 = n53002 ^ n52923 ;
  assign n53004 = n53003 ^ n52917 ;
  assign n53005 = ~n52919 & n53004 ;
  assign n53006 = n53005 ^ n52918 ;
  assign n53007 = n53006 ^ n52912 ;
  assign n53008 = ~n52914 & n53007 ;
  assign n53009 = n53008 ^ n52913 ;
  assign n53010 = n53009 ^ n52907 ;
  assign n53011 = n52909 & n53010 ;
  assign n53012 = n53011 ^ n52908 ;
  assign n53013 = n53012 ^ n52902 ;
  assign n53014 = n52904 & ~n53013 ;
  assign n53015 = n53014 ^ n52903 ;
  assign n53016 = n53015 ^ n52897 ;
  assign n53017 = n52899 & ~n53016 ;
  assign n53018 = n53017 ^ n52898 ;
  assign n53019 = n53018 ^ n52892 ;
  assign n53020 = n52894 & ~n53019 ;
  assign n53021 = n53020 ^ n52893 ;
  assign n53022 = n53021 ^ n52887 ;
  assign n53023 = ~n52889 & ~n53022 ;
  assign n53024 = n53023 ^ n52888 ;
  assign n53025 = n53024 ^ n52883 ;
  assign n53026 = ~n52884 & ~n53025 ;
  assign n53028 = n53027 ^ n53026 ;
  assign n53029 = ~n52879 & ~n53028 ;
  assign n53030 = n53029 ^ n52878 ;
  assign n53031 = n53030 ^ n52870 ;
  assign n53032 = ~n52874 & ~n53031 ;
  assign n53033 = n53032 ^ n52873 ;
  assign n53034 = n53033 ^ n52867 ;
  assign n53035 = n52869 & ~n53034 ;
  assign n53036 = n53035 ^ n52868 ;
  assign n53037 = n53036 ^ n52862 ;
  assign n53038 = n52864 & ~n53037 ;
  assign n53039 = n53038 ^ n52863 ;
  assign n53040 = n53039 ^ n52857 ;
  assign n53041 = ~n52859 & ~n53040 ;
  assign n53042 = n53041 ^ n52858 ;
  assign n53043 = n53042 ^ n1748 ;
  assign n53044 = n52854 & ~n53043 ;
  assign n53046 = n53045 ^ n53044 ;
  assign n53047 = n52852 & ~n53046 ;
  assign n53048 = n53047 ^ n52851 ;
  assign n53049 = n53048 ^ n52845 ;
  assign n53050 = n52847 & ~n53049 ;
  assign n53051 = n53050 ^ n52846 ;
  assign n52600 = n52599 ^ n52210 ;
  assign n52601 = ~n52211 & n52600 ;
  assign n52602 = n52601 ^ n52599 ;
  assign n52204 = n51037 ^ n50295 ;
  assign n52205 = n52204 ^ n51759 ;
  assign n52203 = n52202 ^ n52199 ;
  assign n52206 = n52205 ^ n52203 ;
  assign n52746 = n52602 ^ n52206 ;
  assign n52742 = n52741 ^ n52740 ;
  assign n52743 = n52741 ^ n49631 ;
  assign n52744 = n52742 & ~n52743 ;
  assign n52745 = n52744 ^ n49631 ;
  assign n52747 = n52746 ^ n52745 ;
  assign n52823 = n52747 ^ n49625 ;
  assign n52822 = ~n52819 & ~n52821 ;
  assign n52841 = n52823 ^ n52822 ;
  assign n52838 = n50807 ^ n43362 ;
  assign n52839 = n52838 ^ n44026 ;
  assign n52840 = n52839 ^ n2858 ;
  assign n52842 = n52841 ^ n52840 ;
  assign n53093 = n53051 ^ n52842 ;
  assign n53091 = n51780 ^ n50404 ;
  assign n53092 = n53091 ^ n52294 ;
  assign n53134 = n53093 ^ n53092 ;
  assign n53189 = n53134 ^ n50501 ;
  assign n53186 = n51737 ^ n44106 ;
  assign n53187 = n53186 ^ n48225 ;
  assign n53188 = n53187 ^ n42610 ;
  assign n53300 = n53189 ^ n53188 ;
  assign n54021 = n52065 ^ n44353 ;
  assign n54022 = n54021 ^ n48675 ;
  assign n54023 = n54022 ^ n42921 ;
  assign n53273 = n53000 ^ n52924 ;
  assign n53272 = n52239 ^ n51274 ;
  assign n53274 = n53273 ^ n53272 ;
  assign n53135 = n50501 & ~n53134 ;
  assign n53136 = n53135 ^ n50495 ;
  assign n53052 = n53051 ^ n52840 ;
  assign n53053 = n52842 & ~n53052 ;
  assign n53054 = n53053 ^ n52841 ;
  assign n52607 = n51026 ^ n50339 ;
  assign n52608 = n52607 ^ n51762 ;
  assign n52606 = n52452 ^ n52449 ;
  assign n52609 = n52608 ^ n52606 ;
  assign n52603 = n52602 ^ n52203 ;
  assign n52604 = n52206 & n52603 ;
  assign n52605 = n52604 ^ n52205 ;
  assign n52610 = n52609 ^ n52605 ;
  assign n52825 = n52610 ^ n49621 ;
  assign n52748 = n52745 ^ n49625 ;
  assign n52749 = n52747 & n52748 ;
  assign n52750 = n52749 ^ n49625 ;
  assign n52826 = n52825 ^ n52750 ;
  assign n52824 = ~n52822 & n52823 ;
  assign n52836 = n52826 ^ n52824 ;
  assign n52833 = n50984 ^ n43415 ;
  assign n52834 = n52833 ^ n47397 ;
  assign n52835 = n52834 ^ n41618 ;
  assign n52837 = n52836 ^ n52835 ;
  assign n53096 = n53054 ^ n52837 ;
  assign n53094 = ~n53092 & n53093 ;
  assign n53089 = n51783 ^ n50395 ;
  assign n53090 = n53089 ^ n52288 ;
  assign n53095 = n53094 ^ n53090 ;
  assign n53137 = n53096 ^ n53095 ;
  assign n53138 = n53137 ^ n53135 ;
  assign n53139 = n53136 & ~n53138 ;
  assign n53140 = n53139 ^ n50495 ;
  assign n53141 = n53140 ^ n50493 ;
  assign n53097 = n53096 ^ n53090 ;
  assign n53098 = n53095 & ~n53097 ;
  assign n53099 = n53098 ^ n53094 ;
  assign n53086 = n51791 ^ n50393 ;
  assign n53087 = n53086 ^ n52285 ;
  assign n52829 = n50992 ^ n43357 ;
  assign n52830 = n52829 ^ n47410 ;
  assign n52831 = n52830 ^ n41614 ;
  assign n53057 = n52836 ^ n52831 ;
  assign n53055 = n53054 ^ n52835 ;
  assign n53056 = n52837 & ~n53055 ;
  assign n53058 = n53057 ^ n53056 ;
  assign n52827 = ~n52824 & ~n52826 ;
  assign n52761 = n51022 ^ n50382 ;
  assign n52762 = n52761 ^ n51751 ;
  assign n52755 = n52456 ^ n1232 ;
  assign n52756 = n52755 ^ n52606 ;
  assign n52757 = n52756 ^ n52755 ;
  assign n52758 = n52757 ^ n52605 ;
  assign n52759 = n52609 & n52758 ;
  assign n52760 = n52759 ^ n52756 ;
  assign n52763 = n52762 ^ n52760 ;
  assign n52764 = n52763 ^ n49617 ;
  assign n52751 = n52750 ^ n52610 ;
  assign n52752 = n52750 ^ n49621 ;
  assign n52753 = ~n52751 & ~n52752 ;
  assign n52754 = n52753 ^ n49621 ;
  assign n52765 = n52764 ^ n52754 ;
  assign n52828 = n52827 ^ n52765 ;
  assign n53084 = n53058 ^ n52828 ;
  assign n53088 = n53087 ^ n53084 ;
  assign n53142 = n53099 ^ n53088 ;
  assign n53143 = n53142 ^ n53140 ;
  assign n53144 = ~n53141 & n53143 ;
  assign n53145 = n53144 ^ n50493 ;
  assign n53100 = n53099 ^ n53084 ;
  assign n53101 = ~n53088 & ~n53100 ;
  assign n53081 = n51799 ^ n51070 ;
  assign n53082 = n53081 ^ n52278 ;
  assign n53085 = n53084 ^ n53082 ;
  assign n53102 = n53101 ^ n53085 ;
  assign n53076 = n50803 ^ n43353 ;
  assign n53077 = n53076 ^ n47456 ;
  assign n53078 = n53077 ^ n41608 ;
  assign n53074 = ~n52765 & n52827 ;
  assign n53068 = n50505 ^ n50415 ;
  assign n53069 = n53068 ^ n51749 ;
  assign n53067 = n52458 ^ n52442 ;
  assign n53070 = n53069 ^ n53067 ;
  assign n53064 = n52762 ^ n52755 ;
  assign n53065 = n52760 & n53064 ;
  assign n53066 = n53065 ^ n52755 ;
  assign n53071 = n53070 ^ n53066 ;
  assign n53072 = n53071 ^ n48954 ;
  assign n53061 = n52763 ^ n52754 ;
  assign n53062 = n52764 & n53061 ;
  assign n53063 = n53062 ^ n49617 ;
  assign n53073 = n53072 ^ n53063 ;
  assign n53075 = n53074 ^ n53073 ;
  assign n53079 = n53078 ^ n53075 ;
  assign n52832 = n52831 ^ n52828 ;
  assign n53059 = ~n52832 & n53058 ;
  assign n53060 = n53059 ^ n52831 ;
  assign n53080 = n53079 ^ n53060 ;
  assign n53132 = n53102 ^ n53080 ;
  assign n53133 = n53132 ^ n50412 ;
  assign n53166 = n53145 ^ n53133 ;
  assign n53167 = n53137 ^ n53136 ;
  assign n53168 = n53142 ^ n53141 ;
  assign n53169 = ~n53167 & ~n53168 ;
  assign n53170 = n53166 & ~n53169 ;
  assign n53146 = n53145 ^ n53132 ;
  assign n53147 = ~n53133 & ~n53146 ;
  assign n53148 = n53147 ^ n50412 ;
  assign n53164 = n53148 ^ n50407 ;
  assign n53127 = n53078 ^ n53060 ;
  assign n53128 = ~n53079 & n53127 ;
  assign n53120 = n48954 ^ n48949 ;
  assign n53116 = n50513 ^ n50410 ;
  assign n53117 = n53116 ^ n51745 ;
  assign n53118 = n53117 ^ n53069 ;
  assign n53115 = n52461 ^ n52437 ;
  assign n53119 = n53118 ^ n53115 ;
  assign n53121 = n53120 ^ n53119 ;
  assign n53112 = n50798 ^ n43338 ;
  assign n53113 = n53112 ^ n47501 ;
  assign n53114 = n53113 ^ n41604 ;
  assign n53122 = n53121 ^ n53114 ;
  assign n53123 = n53122 ^ n53078 ;
  assign n53110 = n53067 ^ n53066 ;
  assign n53111 = n53070 & ~n53110 ;
  assign n53124 = n53123 ^ n53111 ;
  assign n53108 = n53071 ^ n53063 ;
  assign n53109 = n53072 & ~n53108 ;
  assign n53125 = n53124 ^ n53109 ;
  assign n53107 = ~n53073 & ~n53074 ;
  assign n53126 = n53125 ^ n53107 ;
  assign n53129 = n53128 ^ n53126 ;
  assign n53105 = n51807 ^ n51151 ;
  assign n53106 = n53105 ^ n52274 ;
  assign n53130 = n53129 ^ n53106 ;
  assign n53083 = n53082 ^ n53080 ;
  assign n53103 = n53083 & n53102 ;
  assign n53104 = n53103 ^ n53082 ;
  assign n53131 = n53130 ^ n53104 ;
  assign n53165 = n53164 ^ n53131 ;
  assign n53181 = n53170 ^ n53165 ;
  assign n53177 = n51203 ^ n43843 ;
  assign n53178 = n53177 ^ n47636 ;
  assign n53179 = n53178 ^ n41991 ;
  assign n53182 = n53181 ^ n53179 ;
  assign n53190 = n53188 & ~n53189 ;
  assign n53183 = n51218 ^ n43856 ;
  assign n53184 = n53183 ^ n47644 ;
  assign n53185 = n53184 ^ n2732 ;
  assign n53191 = n53190 ^ n53185 ;
  assign n53192 = n51214 ^ n43853 ;
  assign n53193 = n53192 ^ n47640 ;
  assign n53194 = n53193 ^ n41976 ;
  assign n53195 = n53194 ^ n53167 ;
  assign n53196 = n53195 ^ n53185 ;
  assign n53197 = n53196 ^ n53194 ;
  assign n53198 = ~n53191 & ~n53197 ;
  assign n53199 = n53198 ^ n53195 ;
  assign n53204 = n53168 ^ n53167 ;
  assign n53200 = n51207 ^ n43849 ;
  assign n53201 = n53200 ^ n47655 ;
  assign n53202 = n53201 ^ n41972 ;
  assign n53205 = n53204 ^ n53202 ;
  assign n53203 = n53202 ^ n53194 ;
  assign n53206 = n53205 ^ n53203 ;
  assign n53207 = ~n53199 & ~n53206 ;
  assign n53208 = n53207 ^ n53203 ;
  assign n53211 = n53202 ^ n53179 ;
  assign n53209 = n53169 ^ n53166 ;
  assign n53210 = n53209 ^ n53179 ;
  assign n53212 = n53211 ^ n53210 ;
  assign n53213 = n53208 & ~n53212 ;
  assign n53214 = n53213 ^ n53211 ;
  assign n53215 = n53182 & n53214 ;
  assign n53171 = n53165 & ~n53170 ;
  assign n53149 = n53148 ^ n53131 ;
  assign n53155 = n51330 ^ n51263 ;
  assign n53156 = n53155 ^ n52272 ;
  assign n53152 = n52972 ^ n52971 ;
  assign n53153 = n53152 ^ n53129 ;
  assign n53150 = n53129 ^ n53104 ;
  assign n53151 = n53130 & n53150 ;
  assign n53154 = n53153 ^ n53151 ;
  assign n53157 = n53156 ^ n53154 ;
  assign n53158 = n53157 ^ n50407 ;
  assign n53159 = n53158 ^ n53157 ;
  assign n53160 = n53159 ^ n53131 ;
  assign n53161 = n53149 & ~n53160 ;
  assign n53162 = n53161 ^ n53158 ;
  assign n53163 = n53162 ^ n50401 ;
  assign n53172 = n53171 ^ n53163 ;
  assign n53180 = n53179 ^ n53172 ;
  assign n53216 = n53215 ^ n53180 ;
  assign n53173 = n51197 ^ n43839 ;
  assign n53174 = n53173 ^ n47630 ;
  assign n53175 = n53174 ^ n41967 ;
  assign n53271 = n53216 ^ n53175 ;
  assign n53275 = n53274 ^ n53271 ;
  assign n53279 = n53214 ^ n53181 ;
  assign n53887 = n53279 ^ n53274 ;
  assign n53277 = n52998 ^ n52927 ;
  assign n53276 = n52246 ^ n51309 ;
  assign n53278 = n53277 ^ n53276 ;
  assign n53280 = n53279 ^ n53278 ;
  assign n53284 = n53209 ^ n53208 ;
  assign n53282 = n52994 ^ n52934 ;
  assign n53281 = n52250 ^ n51314 ;
  assign n53283 = n53282 ^ n53281 ;
  assign n53285 = n53284 ^ n53283 ;
  assign n53286 = n53204 ^ n53199 ;
  assign n53881 = n53286 ^ n53284 ;
  assign n53288 = n52992 ^ n52937 ;
  assign n53287 = n52256 ^ n51316 ;
  assign n53289 = n53288 ^ n53287 ;
  assign n53290 = n53289 ^ n53286 ;
  assign n53294 = n53185 ^ n53167 ;
  assign n53295 = n53294 ^ n53190 ;
  assign n53292 = n52989 ^ n52945 ;
  assign n53291 = n52258 ^ n51325 ;
  assign n53293 = n53292 ^ n53291 ;
  assign n53296 = n53295 ^ n53293 ;
  assign n53298 = n52987 ^ n52948 ;
  assign n53297 = n52262 ^ n51330 ;
  assign n53299 = n53298 ^ n53297 ;
  assign n53301 = n53300 ^ n53299 ;
  assign n53440 = n53036 ^ n52864 ;
  assign n53437 = n51751 ^ n51037 ;
  assign n53438 = n53437 ^ n52507 ;
  assign n53310 = n53033 ^ n52869 ;
  assign n53308 = n51762 ^ n51038 ;
  assign n53309 = n53308 ^ n53115 ;
  assign n53311 = n53310 ^ n53309 ;
  assign n53314 = n53030 ^ n52874 ;
  assign n53433 = n53314 ^ n53310 ;
  assign n53312 = n51759 ^ n51034 ;
  assign n53313 = n53312 ^ n53067 ;
  assign n53315 = n53314 ^ n53313 ;
  assign n53318 = n53028 ^ n52877 ;
  assign n53316 = n52209 ^ n51728 ;
  assign n53317 = n53316 ^ n52755 ;
  assign n53319 = n53318 ^ n53317 ;
  assign n53322 = n53024 ^ n52884 ;
  assign n53320 = n52213 ^ n51452 ;
  assign n53321 = n53320 ^ n52606 ;
  assign n53323 = n53322 ^ n53321 ;
  assign n53326 = n53021 ^ n52889 ;
  assign n53324 = n52219 ^ n51446 ;
  assign n53325 = n53324 ^ n52203 ;
  assign n53327 = n53326 ^ n53325 ;
  assign n53330 = n53018 ^ n52894 ;
  assign n53328 = n52224 ^ n51436 ;
  assign n53329 = n53328 ^ n52207 ;
  assign n53331 = n53330 ^ n53329 ;
  assign n53334 = n53015 ^ n52899 ;
  assign n53332 = n52325 ^ n51428 ;
  assign n53333 = n53332 ^ n52215 ;
  assign n53335 = n53334 ^ n53333 ;
  assign n53337 = n52230 ^ n51346 ;
  assign n53338 = n53337 ^ n52217 ;
  assign n53336 = n53012 ^ n52904 ;
  assign n53339 = n53338 ^ n53336 ;
  assign n53342 = n53009 ^ n52909 ;
  assign n53340 = n52235 ^ n51344 ;
  assign n53341 = n53340 ^ n52226 ;
  assign n53343 = n53342 ^ n53341 ;
  assign n53345 = n52305 ^ n51351 ;
  assign n53346 = n53345 ^ n52233 ;
  assign n53344 = n53006 ^ n52914 ;
  assign n53347 = n53346 ^ n53344 ;
  assign n53241 = n53003 ^ n52919 ;
  assign n53405 = n53346 ^ n53241 ;
  assign n53348 = n52307 ^ n51355 ;
  assign n53349 = n53348 ^ n52228 ;
  assign n53350 = n53349 ^ n53241 ;
  assign n53351 = n52191 ^ n51302 ;
  assign n53352 = n53351 ^ n52237 ;
  assign n53353 = n53352 ^ n53273 ;
  assign n53399 = n53352 ^ n53277 ;
  assign n53354 = n52006 ^ n51306 ;
  assign n53355 = n53354 ^ n52563 ;
  assign n53356 = n53355 ^ n53277 ;
  assign n53357 = n51987 ^ n51311 ;
  assign n53358 = n53357 ^ n52243 ;
  assign n53359 = n53358 ^ n53282 ;
  assign n53360 = n51938 ^ n51318 ;
  assign n53361 = n53360 ^ n52239 ;
  assign n53362 = n53361 ^ n53288 ;
  assign n53363 = n51323 ^ n51300 ;
  assign n53364 = n53363 ^ n52246 ;
  assign n53365 = n53364 ^ n53292 ;
  assign n53366 = n51328 ^ n51274 ;
  assign n53367 = n53366 ^ n52250 ;
  assign n53368 = n53367 ^ n53298 ;
  assign n53369 = n51377 ^ n51309 ;
  assign n53370 = n53369 ^ n52256 ;
  assign n53303 = n52983 ^ n52955 ;
  assign n53371 = n53370 ^ n53303 ;
  assign n53373 = n51386 ^ n51314 ;
  assign n53374 = n53373 ^ n52258 ;
  assign n53381 = n53374 ^ n53370 ;
  assign n53372 = n52980 ^ n52960 ;
  assign n53375 = n53374 ^ n53372 ;
  assign n53257 = n52977 ^ n52965 ;
  assign n53255 = n51387 ^ n51316 ;
  assign n53256 = n53255 ^ n52262 ;
  assign n53258 = n53257 ^ n53256 ;
  assign n53230 = n52968 ^ n52772 ;
  assign n53231 = n53230 ^ n52973 ;
  assign n53232 = n53231 ^ n53152 ;
  assign n53228 = n53156 ^ n53152 ;
  assign n53229 = ~n53154 & n53228 ;
  assign n53233 = n53232 ^ n53229 ;
  assign n53234 = n51325 ^ n51280 ;
  assign n53235 = n53234 ^ n52268 ;
  assign n53252 = n53235 ^ n53231 ;
  assign n53253 = n53233 & ~n53252 ;
  assign n53254 = n53253 ^ n53235 ;
  assign n53376 = n53256 ^ n53254 ;
  assign n53377 = n53258 & ~n53376 ;
  assign n53378 = n53377 ^ n53257 ;
  assign n53379 = n53378 ^ n53372 ;
  assign n53380 = ~n53375 & n53379 ;
  assign n53382 = n53381 ^ n53380 ;
  assign n53383 = ~n53371 & ~n53382 ;
  assign n53384 = n53383 ^ n53370 ;
  assign n53385 = n53384 ^ n53298 ;
  assign n53386 = ~n53368 & n53385 ;
  assign n53387 = n53386 ^ n53298 ;
  assign n53388 = n53387 ^ n53364 ;
  assign n53389 = ~n53365 & n53388 ;
  assign n53390 = n53389 ^ n53292 ;
  assign n53391 = n53390 ^ n53361 ;
  assign n53392 = n53362 & n53391 ;
  assign n53393 = n53392 ^ n53288 ;
  assign n53394 = n53393 ^ n53358 ;
  assign n53395 = ~n53359 & n53394 ;
  assign n53396 = n53395 ^ n53282 ;
  assign n53397 = n53396 ^ n53277 ;
  assign n53398 = n53356 & ~n53397 ;
  assign n53400 = n53399 ^ n53398 ;
  assign n53401 = ~n53353 & ~n53400 ;
  assign n53402 = n53401 ^ n53273 ;
  assign n53403 = n53402 ^ n53241 ;
  assign n53404 = n53350 & n53403 ;
  assign n53406 = n53405 ^ n53404 ;
  assign n53407 = n53347 & n53406 ;
  assign n53408 = n53407 ^ n53346 ;
  assign n53409 = n53408 ^ n53342 ;
  assign n53410 = n53343 & ~n53409 ;
  assign n53411 = n53410 ^ n53342 ;
  assign n53412 = n53411 ^ n53334 ;
  assign n53413 = n53412 ^ n53336 ;
  assign n53414 = n53413 ^ n53334 ;
  assign n53415 = n53339 & ~n53414 ;
  assign n53416 = n53415 ^ n53412 ;
  assign n53417 = n53335 & ~n53416 ;
  assign n53418 = n53417 ^ n53334 ;
  assign n53419 = n53418 ^ n53329 ;
  assign n53420 = n53331 & ~n53419 ;
  assign n53421 = n53420 ^ n53330 ;
  assign n53422 = n53421 ^ n53325 ;
  assign n53423 = n53327 & n53422 ;
  assign n53424 = n53423 ^ n53326 ;
  assign n53425 = n53424 ^ n53321 ;
  assign n53426 = ~n53323 & ~n53425 ;
  assign n53427 = n53426 ^ n53322 ;
  assign n53428 = n53427 ^ n53317 ;
  assign n53429 = ~n53319 & ~n53428 ;
  assign n53430 = n53429 ^ n53318 ;
  assign n53431 = n53430 ^ n53314 ;
  assign n53432 = n53315 & ~n53431 ;
  assign n53434 = n53433 ^ n53432 ;
  assign n53435 = ~n53311 & n53434 ;
  assign n53436 = n53435 ^ n53310 ;
  assign n53439 = n53438 ^ n53436 ;
  assign n53551 = n53440 ^ n53439 ;
  assign n53449 = n53434 ^ n53309 ;
  assign n53450 = n53449 ^ n50249 ;
  assign n53543 = n53430 ^ n53315 ;
  assign n53451 = n53427 ^ n53319 ;
  assign n53452 = n53451 ^ n51011 ;
  assign n53535 = n53424 ^ n53323 ;
  assign n53453 = n53421 ^ n53327 ;
  assign n53454 = n53453 ^ n50417 ;
  assign n53526 = n53418 ^ n53331 ;
  assign n53455 = n53416 ^ n53333 ;
  assign n53456 = n53455 ^ n50421 ;
  assign n53458 = n53408 ^ n53343 ;
  assign n53459 = n53458 ^ n50434 ;
  assign n53509 = n53406 ^ n53344 ;
  assign n53461 = n53400 ^ n53273 ;
  assign n53462 = n53461 ^ n50441 ;
  assign n53463 = n53396 ^ n53356 ;
  assign n53464 = n53463 ^ n50445 ;
  assign n53465 = n53393 ^ n53359 ;
  assign n53466 = n53465 ^ n50452 ;
  assign n53467 = n53390 ^ n53362 ;
  assign n53468 = n53467 ^ n50454 ;
  assign n53469 = n53387 ^ n53365 ;
  assign n53470 = n53469 ^ n50462 ;
  assign n53471 = n53384 ^ n53368 ;
  assign n53472 = n53471 ^ n50466 ;
  assign n53474 = n53378 ^ n53375 ;
  assign n53475 = n53474 ^ n50474 ;
  assign n53236 = n53235 ^ n53233 ;
  assign n53224 = n53157 ^ n50401 ;
  assign n53225 = n53162 & ~n53224 ;
  assign n53226 = n53225 ^ n50401 ;
  assign n53251 = n53236 ^ n53226 ;
  assign n53259 = n53258 ^ n53254 ;
  assign n53260 = n53259 ^ n50398 ;
  assign n53261 = n53260 ^ n53226 ;
  assign n53262 = n53261 ^ n53259 ;
  assign n53263 = n53251 & n53262 ;
  assign n53264 = n53263 ^ n53260 ;
  assign n53477 = n53474 ^ n49801 ;
  assign n53476 = n53474 ^ n53259 ;
  assign n53478 = n53477 ^ n53476 ;
  assign n53479 = ~n53264 & n53478 ;
  assign n53480 = n53479 ^ n53477 ;
  assign n53481 = n53475 & n53480 ;
  assign n53482 = n53481 ^ n50474 ;
  assign n53473 = n53382 ^ n53303 ;
  assign n53483 = n53482 ^ n53473 ;
  assign n53484 = n53482 ^ n50470 ;
  assign n53485 = ~n53483 & ~n53484 ;
  assign n53486 = n53485 ^ n50470 ;
  assign n53487 = n53486 ^ n53471 ;
  assign n53488 = n53472 & ~n53487 ;
  assign n53489 = n53488 ^ n50466 ;
  assign n53490 = n53489 ^ n53469 ;
  assign n53491 = ~n53470 & ~n53490 ;
  assign n53492 = n53491 ^ n50462 ;
  assign n53493 = n53492 ^ n53467 ;
  assign n53494 = n53468 & ~n53493 ;
  assign n53495 = n53494 ^ n50454 ;
  assign n53496 = n53495 ^ n53465 ;
  assign n53497 = n53466 & ~n53496 ;
  assign n53498 = n53497 ^ n50452 ;
  assign n53499 = n53498 ^ n53463 ;
  assign n53500 = ~n53464 & n53499 ;
  assign n53501 = n53500 ^ n50445 ;
  assign n53502 = n53501 ^ n53461 ;
  assign n53503 = ~n53462 & n53502 ;
  assign n53504 = n53503 ^ n50441 ;
  assign n53460 = n53402 ^ n53350 ;
  assign n53505 = n53504 ^ n53460 ;
  assign n53506 = n53504 ^ n50437 ;
  assign n53507 = n53505 & n53506 ;
  assign n53508 = n53507 ^ n50437 ;
  assign n53510 = n53509 ^ n53508 ;
  assign n53511 = n53458 ^ n50430 ;
  assign n53512 = n53511 ^ n53458 ;
  assign n53513 = n53512 ^ n53508 ;
  assign n53514 = n53510 & n53513 ;
  assign n53515 = n53514 ^ n53511 ;
  assign n53516 = n53459 & n53515 ;
  assign n53517 = n53516 ^ n50434 ;
  assign n53457 = n53411 ^ n53339 ;
  assign n53518 = n53517 ^ n53457 ;
  assign n53519 = n53455 ^ n50428 ;
  assign n53520 = n53519 ^ n53457 ;
  assign n53521 = n53520 ^ n53455 ;
  assign n53522 = ~n53518 & n53521 ;
  assign n53523 = n53522 ^ n53519 ;
  assign n53524 = n53456 & n53523 ;
  assign n53525 = n53524 ^ n50421 ;
  assign n53527 = n53526 ^ n53525 ;
  assign n53528 = n53453 ^ n50425 ;
  assign n53529 = n53528 ^ n53525 ;
  assign n53530 = n53529 ^ n53453 ;
  assign n53531 = n53527 & n53530 ;
  assign n53532 = n53531 ^ n53528 ;
  assign n53533 = ~n53454 & n53532 ;
  assign n53534 = n53533 ^ n50417 ;
  assign n53536 = n53535 ^ n53534 ;
  assign n53537 = n53535 ^ n50598 ;
  assign n53538 = n53536 & n53537 ;
  assign n53539 = n53538 ^ n50598 ;
  assign n53540 = n53539 ^ n53451 ;
  assign n53541 = ~n53452 & n53540 ;
  assign n53542 = n53541 ^ n51011 ;
  assign n53544 = n53543 ^ n53542 ;
  assign n53545 = n53543 ^ n50220 ;
  assign n53546 = n53544 & ~n53545 ;
  assign n53547 = n53546 ^ n50220 ;
  assign n53548 = n53547 ^ n53449 ;
  assign n53549 = n53450 & n53548 ;
  assign n53550 = n53549 ^ n50249 ;
  assign n53552 = n53551 ^ n53550 ;
  assign n53553 = n53551 ^ n50295 ;
  assign n53554 = ~n53552 & ~n53553 ;
  assign n53555 = n53554 ^ n50295 ;
  assign n53446 = n53039 ^ n52859 ;
  assign n53444 = n51749 ^ n51026 ;
  assign n53445 = n53444 ^ n52513 ;
  assign n53447 = n53446 ^ n53445 ;
  assign n53441 = n53440 ^ n53436 ;
  assign n53442 = n53439 & n53441 ;
  assign n53443 = n53442 ^ n53440 ;
  assign n53448 = n53447 ^ n53443 ;
  assign n53556 = n53555 ^ n53448 ;
  assign n53561 = n53446 ^ n53443 ;
  assign n53562 = n53447 & ~n53561 ;
  assign n53563 = n53562 ^ n53446 ;
  assign n53559 = n53042 ^ n52854 ;
  assign n53557 = n51745 ^ n51022 ;
  assign n53558 = n53557 ^ n52503 ;
  assign n53560 = n53559 ^ n53558 ;
  assign n53564 = n53563 ^ n53560 ;
  assign n53565 = n53564 ^ n50339 ;
  assign n53566 = n53565 ^ n53448 ;
  assign n53567 = n53566 ^ n53564 ;
  assign n53568 = ~n53556 & n53567 ;
  assign n53569 = n53568 ^ n53565 ;
  assign n53576 = n53046 ^ n52851 ;
  assign n53574 = n51338 ^ n50415 ;
  assign n53575 = n53574 ^ n52499 ;
  assign n53577 = n53576 ^ n53575 ;
  assign n53570 = n53563 ^ n53559 ;
  assign n53571 = n53563 ^ n53558 ;
  assign n53572 = n53570 & ~n53571 ;
  assign n53573 = n53572 ^ n53559 ;
  assign n53578 = n53577 ^ n53573 ;
  assign n53580 = n53578 ^ n50382 ;
  assign n53579 = n53578 ^ n53564 ;
  assign n53581 = n53580 ^ n53579 ;
  assign n53582 = n53569 & ~n53581 ;
  assign n53583 = n53582 ^ n53580 ;
  assign n53584 = n53583 ^ n50505 ;
  assign n53585 = n53448 ^ n50339 ;
  assign n53586 = n53585 ^ n53555 ;
  assign n53587 = n53553 ^ n53550 ;
  assign n53588 = n53545 ^ n53542 ;
  assign n53589 = n53526 ^ n50425 ;
  assign n53590 = n53589 ^ n53525 ;
  assign n53591 = n53523 ^ n50421 ;
  assign n53592 = n53515 ^ n50434 ;
  assign n53593 = n53509 ^ n50430 ;
  assign n53594 = n53593 ^ n53508 ;
  assign n53595 = n53460 ^ n50437 ;
  assign n53596 = n53595 ^ n53504 ;
  assign n53597 = n53486 ^ n53472 ;
  assign n53598 = n53473 ^ n50470 ;
  assign n53599 = n53598 ^ n53482 ;
  assign n53223 = ~n53163 & ~n53171 ;
  assign n53227 = n53226 ^ n50398 ;
  assign n53237 = n53236 ^ n53227 ;
  assign n53250 = ~n53223 & n53237 ;
  assign n53265 = n53264 ^ n49801 ;
  assign n53600 = n53250 & ~n53265 ;
  assign n53601 = n53480 ^ n50474 ;
  assign n53602 = n53600 & ~n53601 ;
  assign n53603 = n53599 & ~n53602 ;
  assign n53604 = n53597 & n53603 ;
  assign n53605 = n53489 ^ n50462 ;
  assign n53606 = n53605 ^ n53469 ;
  assign n53607 = n53604 & ~n53606 ;
  assign n53608 = n53492 ^ n53468 ;
  assign n53609 = n53607 & ~n53608 ;
  assign n53610 = n53495 ^ n50452 ;
  assign n53611 = n53610 ^ n53465 ;
  assign n53612 = n53609 & ~n53611 ;
  assign n53613 = n53498 ^ n50445 ;
  assign n53614 = n53613 ^ n53463 ;
  assign n53615 = ~n53612 & ~n53614 ;
  assign n53616 = n53501 ^ n53462 ;
  assign n53617 = n53615 & ~n53616 ;
  assign n53618 = n53596 & ~n53617 ;
  assign n53619 = ~n53594 & ~n53618 ;
  assign n53620 = ~n53592 & ~n53619 ;
  assign n53621 = n53517 ^ n50428 ;
  assign n53622 = n53621 ^ n53457 ;
  assign n53623 = n53620 & n53622 ;
  assign n53624 = n53591 & n53623 ;
  assign n53625 = ~n53590 & ~n53624 ;
  assign n53626 = n53532 ^ n50417 ;
  assign n53627 = n53625 & ~n53626 ;
  assign n53628 = n53534 ^ n50598 ;
  assign n53629 = n53628 ^ n53535 ;
  assign n53630 = ~n53627 & ~n53629 ;
  assign n53631 = n53539 ^ n53452 ;
  assign n53632 = n53630 & ~n53631 ;
  assign n53633 = n53588 & ~n53632 ;
  assign n53634 = n53547 ^ n53450 ;
  assign n53635 = ~n53633 & n53634 ;
  assign n53636 = ~n53587 & ~n53635 ;
  assign n53637 = n53586 & ~n53636 ;
  assign n53638 = n53569 ^ n50382 ;
  assign n53639 = n53637 & ~n53638 ;
  assign n53841 = n53584 & ~n53639 ;
  assign n53833 = n53048 ^ n52847 ;
  assign n53831 = n51334 ^ n50410 ;
  assign n53832 = n53831 ^ n52495 ;
  assign n53834 = n53833 ^ n53832 ;
  assign n53835 = n53834 ^ n53575 ;
  assign n53836 = n53835 ^ n50514 ;
  assign n53828 = n51587 ^ n44086 ;
  assign n53829 = n53828 ^ n48195 ;
  assign n53830 = n53829 ^ n42433 ;
  assign n53837 = n53836 ^ n53830 ;
  assign n53305 = n51592 ^ n44009 ;
  assign n53306 = n53305 ^ n48136 ;
  assign n53307 = n53306 ^ n42437 ;
  assign n53838 = n53837 ^ n53307 ;
  assign n53826 = n53578 ^ n50505 ;
  assign n53827 = ~n53583 & ~n53826 ;
  assign n53839 = n53838 ^ n53827 ;
  assign n53824 = n53575 ^ n53573 ;
  assign n53825 = ~n53577 & n53824 ;
  assign n53840 = n53839 ^ n53825 ;
  assign n53842 = n53841 ^ n53840 ;
  assign n53640 = n53639 ^ n53584 ;
  assign n53641 = n53640 ^ n53307 ;
  assign n53645 = n53638 ^ n53637 ;
  assign n53642 = n51596 ^ n43942 ;
  assign n53643 = n53642 ^ n47705 ;
  assign n53644 = n53643 ^ n42442 ;
  assign n53646 = n53645 ^ n53644 ;
  assign n53648 = n51601 ^ n2903 ;
  assign n53649 = n53648 ^ n47989 ;
  assign n53650 = n53649 ^ n42447 ;
  assign n53818 = n53650 ^ n53644 ;
  assign n53647 = n53636 ^ n53586 ;
  assign n53651 = n53650 ^ n53647 ;
  assign n53655 = n53635 ^ n53587 ;
  assign n53652 = n51606 ^ n43738 ;
  assign n53653 = n53652 ^ n47995 ;
  assign n53654 = n53653 ^ n42453 ;
  assign n53656 = n53655 ^ n53654 ;
  assign n53662 = n51611 ^ n43743 ;
  assign n53663 = n53662 ^ n47999 ;
  assign n53664 = n53663 ^ n42458 ;
  assign n53812 = n53664 ^ n53654 ;
  assign n53658 = n51616 ^ n1774 ;
  assign n53659 = n53658 ^ n48005 ;
  assign n53660 = n53659 ^ n42463 ;
  assign n53657 = n53632 ^ n53588 ;
  assign n53661 = n53660 ^ n53657 ;
  assign n53670 = n53631 ^ n53630 ;
  assign n53667 = n51621 ^ n1759 ;
  assign n53668 = n53667 ^ n48011 ;
  assign n53669 = n53668 ^ n1184 ;
  assign n53671 = n53670 ^ n53669 ;
  assign n53675 = n53629 ^ n53627 ;
  assign n53672 = n51626 ^ n43751 ;
  assign n53673 = n53672 ^ n1049 ;
  assign n53674 = n53673 ^ n42469 ;
  assign n53676 = n53675 ^ n53674 ;
  assign n53681 = n53626 ^ n53625 ;
  assign n53677 = n51632 ^ n43757 ;
  assign n53678 = n53677 ^ n48018 ;
  assign n53679 = n53678 ^ n1038 ;
  assign n53682 = n53681 ^ n53679 ;
  assign n53686 = n53624 ^ n53590 ;
  assign n53683 = n51636 ^ n893 ;
  assign n53684 = n53683 ^ n48023 ;
  assign n53685 = n53684 ^ n42476 ;
  assign n53687 = n53686 ^ n53685 ;
  assign n53691 = n53623 ^ n53591 ;
  assign n53688 = n51641 ^ n43763 ;
  assign n53689 = n53688 ^ n48028 ;
  assign n53690 = n53689 ^ n1637 ;
  assign n53692 = n53691 ^ n53690 ;
  assign n53697 = n53622 ^ n53620 ;
  assign n53693 = n51646 ^ n43768 ;
  assign n53694 = n53693 ^ n48034 ;
  assign n53695 = n53694 ^ n42483 ;
  assign n53698 = n53697 ^ n53695 ;
  assign n53702 = n53619 ^ n53592 ;
  assign n53699 = n51651 ^ n43773 ;
  assign n53700 = n53699 ^ n48039 ;
  assign n53701 = n53700 ^ n42488 ;
  assign n53703 = n53702 ^ n53701 ;
  assign n53707 = n53618 ^ n53594 ;
  assign n53704 = n51656 ^ n43778 ;
  assign n53705 = n53704 ^ n48043 ;
  assign n53706 = n53705 ^ n42493 ;
  assign n53708 = n53707 ^ n53706 ;
  assign n53712 = n53617 ^ n53596 ;
  assign n53709 = n51661 ^ n43783 ;
  assign n53710 = n53709 ^ n48048 ;
  assign n53711 = n53710 ^ n42499 ;
  assign n53713 = n53712 ^ n53711 ;
  assign n53715 = n51666 ^ n43790 ;
  assign n53716 = n53715 ^ n48053 ;
  assign n53717 = n53716 ^ n42505 ;
  assign n53780 = n53717 ^ n53711 ;
  assign n53714 = n53616 ^ n53615 ;
  assign n53718 = n53717 ^ n53714 ;
  assign n53722 = n53614 ^ n53612 ;
  assign n53719 = n51298 ^ n43795 ;
  assign n53720 = n53719 ^ n48059 ;
  assign n53721 = n53720 ^ n42511 ;
  assign n53723 = n53722 ^ n53721 ;
  assign n53725 = n51255 ^ n43799 ;
  assign n53726 = n53725 ^ n48064 ;
  assign n53727 = n53726 ^ n42515 ;
  assign n53774 = n53727 ^ n53721 ;
  assign n53724 = n53611 ^ n53609 ;
  assign n53728 = n53727 ^ n53724 ;
  assign n53732 = n53608 ^ n53607 ;
  assign n53729 = n43804 ^ n2441 ;
  assign n53730 = n53729 ^ n48069 ;
  assign n53731 = n53730 ^ n42520 ;
  assign n53733 = n53732 ^ n53731 ;
  assign n53737 = n53606 ^ n53604 ;
  assign n53734 = n51165 ^ n43809 ;
  assign n53735 = n53734 ^ n48073 ;
  assign n53736 = n53735 ^ n42526 ;
  assign n53738 = n53737 ^ n53736 ;
  assign n53740 = n51171 ^ n2349 ;
  assign n53741 = n53740 ^ n47678 ;
  assign n53742 = n53741 ^ n42530 ;
  assign n53739 = n53603 ^ n53597 ;
  assign n53743 = n53742 ^ n53739 ;
  assign n53745 = n51176 ^ n43817 ;
  assign n53746 = n53745 ^ n47611 ;
  assign n53747 = n53746 ^ n42028 ;
  assign n53762 = n53747 ^ n53742 ;
  assign n53744 = n53602 ^ n53599 ;
  assign n53748 = n53747 ^ n53744 ;
  assign n53752 = n53601 ^ n53600 ;
  assign n53749 = n51181 ^ n43823 ;
  assign n53750 = n53749 ^ n47615 ;
  assign n53751 = n53750 ^ n41953 ;
  assign n53753 = n53752 ^ n53751 ;
  assign n53266 = n53265 ^ n53250 ;
  assign n53247 = n51192 ^ n43828 ;
  assign n53248 = n53247 ^ n47621 ;
  assign n53249 = n53248 ^ n41957 ;
  assign n53267 = n53266 ^ n53249 ;
  assign n53218 = n51187 ^ n43833 ;
  assign n53219 = n53218 ^ n47626 ;
  assign n53220 = n53219 ^ n41962 ;
  assign n53221 = n53220 ^ n53175 ;
  assign n53176 = n53175 ^ n53172 ;
  assign n53217 = n53176 & ~n53216 ;
  assign n53222 = n53221 ^ n53217 ;
  assign n53238 = n53237 ^ n53223 ;
  assign n53244 = n53238 ^ n53220 ;
  assign n53245 = n53222 & n53244 ;
  assign n53246 = n53245 ^ n53220 ;
  assign n53754 = n53249 ^ n53246 ;
  assign n53755 = n53267 & ~n53754 ;
  assign n53756 = n53755 ^ n53266 ;
  assign n53757 = n53756 ^ n53751 ;
  assign n53758 = n53753 & ~n53757 ;
  assign n53759 = n53758 ^ n53752 ;
  assign n53760 = n53759 ^ n53747 ;
  assign n53761 = ~n53748 & n53760 ;
  assign n53763 = n53762 ^ n53761 ;
  assign n53764 = n53743 & n53763 ;
  assign n53765 = n53764 ^ n53742 ;
  assign n53766 = n53765 ^ n53736 ;
  assign n53767 = ~n53738 & ~n53766 ;
  assign n53768 = n53767 ^ n53737 ;
  assign n53769 = n53768 ^ n53731 ;
  assign n53770 = ~n53733 & n53769 ;
  assign n53771 = n53770 ^ n53732 ;
  assign n53772 = n53771 ^ n53724 ;
  assign n53773 = ~n53728 & ~n53772 ;
  assign n53775 = n53774 ^ n53773 ;
  assign n53776 = ~n53723 & ~n53775 ;
  assign n53777 = n53776 ^ n53722 ;
  assign n53778 = n53777 ^ n53714 ;
  assign n53779 = n53718 & n53778 ;
  assign n53781 = n53780 ^ n53779 ;
  assign n53782 = ~n53713 & ~n53781 ;
  assign n53783 = n53782 ^ n53712 ;
  assign n53784 = n53783 ^ n53706 ;
  assign n53785 = ~n53708 & n53784 ;
  assign n53786 = n53785 ^ n53707 ;
  assign n53787 = n53786 ^ n53701 ;
  assign n53788 = n53703 & n53787 ;
  assign n53789 = n53788 ^ n53702 ;
  assign n53790 = n53789 ^ n53695 ;
  assign n53791 = n53698 & n53790 ;
  assign n53696 = n53695 ^ n53691 ;
  assign n53792 = n53791 ^ n53696 ;
  assign n53793 = n53692 & n53792 ;
  assign n53794 = n53793 ^ n53691 ;
  assign n53795 = n53794 ^ n53685 ;
  assign n53796 = ~n53687 & ~n53795 ;
  assign n53797 = n53796 ^ n53686 ;
  assign n53798 = n53797 ^ n53679 ;
  assign n53799 = n53682 & ~n53798 ;
  assign n53680 = n53679 ^ n53675 ;
  assign n53800 = n53799 ^ n53680 ;
  assign n53801 = n53676 & n53800 ;
  assign n53802 = n53801 ^ n53675 ;
  assign n53803 = n53802 ^ n53669 ;
  assign n53804 = ~n53671 & ~n53803 ;
  assign n53805 = n53804 ^ n53670 ;
  assign n53665 = n53664 ^ n53660 ;
  assign n53666 = n53665 ^ n53664 ;
  assign n53806 = n53805 ^ n53666 ;
  assign n53807 = n53661 & ~n53806 ;
  assign n53808 = n53807 ^ n53665 ;
  assign n53809 = n53634 ^ n53633 ;
  assign n53810 = n53809 ^ n53664 ;
  assign n53811 = n53808 & ~n53810 ;
  assign n53813 = n53812 ^ n53811 ;
  assign n53814 = ~n53656 & ~n53813 ;
  assign n53815 = n53814 ^ n53655 ;
  assign n53816 = n53815 ^ n53650 ;
  assign n53817 = ~n53651 & ~n53816 ;
  assign n53819 = n53818 ^ n53817 ;
  assign n53820 = ~n53646 & ~n53819 ;
  assign n53821 = n53820 ^ n53645 ;
  assign n53822 = n53821 ^ n53307 ;
  assign n53823 = n53641 & ~n53822 ;
  assign n53843 = n53842 ^ n53823 ;
  assign n53302 = n52268 ^ n51807 ;
  assign n53304 = n53303 ^ n53302 ;
  assign n53844 = n53843 ^ n53304 ;
  assign n53847 = n53821 ^ n53641 ;
  assign n53869 = n53847 ^ n53843 ;
  assign n53845 = n52272 ^ n51799 ;
  assign n53846 = n53845 ^ n53372 ;
  assign n53848 = n53847 ^ n53846 ;
  assign n53851 = n53819 ^ n53645 ;
  assign n53849 = n52274 ^ n51791 ;
  assign n53850 = n53849 ^ n53257 ;
  assign n53852 = n53851 ^ n53850 ;
  assign n53855 = n53813 ^ n53655 ;
  assign n53856 = n52285 ^ n51780 ;
  assign n53857 = n53856 ^ n53152 ;
  assign n53858 = ~n53855 & n53857 ;
  assign n53863 = n53858 ^ n53850 ;
  assign n53853 = n52278 ^ n51783 ;
  assign n53854 = n53853 ^ n53231 ;
  assign n53859 = n53858 ^ n53854 ;
  assign n53860 = n53815 ^ n53651 ;
  assign n53861 = n53860 ^ n53858 ;
  assign n53862 = ~n53859 & n53861 ;
  assign n53864 = n53863 ^ n53862 ;
  assign n53865 = n53852 & n53864 ;
  assign n53866 = n53865 ^ n53851 ;
  assign n53867 = n53866 ^ n53846 ;
  assign n53868 = ~n53848 & n53867 ;
  assign n53870 = n53869 ^ n53868 ;
  assign n53871 = ~n53844 & n53870 ;
  assign n53872 = n53871 ^ n53843 ;
  assign n53873 = n53872 ^ n53299 ;
  assign n53874 = n53301 & ~n53873 ;
  assign n53875 = n53874 ^ n53300 ;
  assign n53876 = n53875 ^ n53293 ;
  assign n53877 = ~n53296 & n53876 ;
  assign n53878 = n53877 ^ n53295 ;
  assign n53879 = n53878 ^ n53286 ;
  assign n53880 = n53290 & ~n53879 ;
  assign n53882 = n53881 ^ n53880 ;
  assign n53883 = ~n53285 & ~n53882 ;
  assign n53884 = n53883 ^ n53284 ;
  assign n53885 = n53884 ^ n53279 ;
  assign n53886 = ~n53280 & ~n53885 ;
  assign n53888 = n53887 ^ n53886 ;
  assign n53889 = ~n53275 & ~n53888 ;
  assign n53890 = n53889 ^ n53274 ;
  assign n53240 = n52243 ^ n51300 ;
  assign n53242 = n53241 ^ n53240 ;
  assign n53239 = n53238 ^ n53222 ;
  assign n53243 = n53242 ^ n53239 ;
  assign n53898 = n53890 ^ n53243 ;
  assign n53972 = n53898 ^ n51323 ;
  assign n53899 = n53888 ^ n53271 ;
  assign n53900 = n53899 ^ n51328 ;
  assign n53902 = n53882 ^ n53283 ;
  assign n53903 = n53902 ^ n51386 ;
  assign n53905 = n53875 ^ n53296 ;
  assign n53906 = n53905 ^ n51280 ;
  assign n53908 = n53866 ^ n53848 ;
  assign n53909 = n53908 ^ n51070 ;
  assign n53912 = n53857 ^ n53855 ;
  assign n53913 = n50404 & ~n53912 ;
  assign n53911 = n53860 ^ n53859 ;
  assign n53914 = n53913 ^ n53911 ;
  assign n53915 = n53913 ^ n50395 ;
  assign n53916 = n53914 & ~n53915 ;
  assign n53917 = n53916 ^ n50395 ;
  assign n53910 = n53864 ^ n53851 ;
  assign n53918 = n53917 ^ n53910 ;
  assign n53919 = n53908 ^ n50393 ;
  assign n53920 = n53919 ^ n53908 ;
  assign n53921 = n53920 ^ n53910 ;
  assign n53922 = n53918 & ~n53921 ;
  assign n53923 = n53922 ^ n53919 ;
  assign n53924 = ~n53909 & n53923 ;
  assign n53925 = n53924 ^ n51070 ;
  assign n53926 = n53925 ^ n51151 ;
  assign n53927 = n53870 ^ n53304 ;
  assign n53928 = n53927 ^ n53925 ;
  assign n53929 = ~n53926 & n53928 ;
  assign n53930 = n53929 ^ n51151 ;
  assign n53907 = n53872 ^ n53301 ;
  assign n53931 = n53930 ^ n53907 ;
  assign n53932 = n53930 ^ n51263 ;
  assign n53933 = n53931 & ~n53932 ;
  assign n53934 = n53933 ^ n51263 ;
  assign n53935 = n53934 ^ n53905 ;
  assign n53936 = ~n53906 & n53935 ;
  assign n53937 = n53936 ^ n51280 ;
  assign n53904 = n53878 ^ n53290 ;
  assign n53938 = n53937 ^ n53904 ;
  assign n53939 = n53937 ^ n51387 ;
  assign n53940 = ~n53938 & n53939 ;
  assign n53941 = n53940 ^ n51387 ;
  assign n53942 = n53941 ^ n53902 ;
  assign n53943 = n53903 & ~n53942 ;
  assign n53944 = n53943 ^ n51386 ;
  assign n53901 = n53884 ^ n53280 ;
  assign n53945 = n53944 ^ n53901 ;
  assign n53946 = n53899 ^ n51377 ;
  assign n53947 = n53946 ^ n53899 ;
  assign n53948 = n53947 ^ n53901 ;
  assign n53949 = n53945 & n53948 ;
  assign n53950 = n53949 ^ n53946 ;
  assign n53951 = ~n53900 & n53950 ;
  assign n53952 = n53951 ^ n51328 ;
  assign n53973 = n53972 ^ n53952 ;
  assign n53974 = n53915 ^ n53911 ;
  assign n53975 = n53910 ^ n50393 ;
  assign n53976 = n53975 ^ n53917 ;
  assign n53977 = ~n53974 & ~n53976 ;
  assign n53978 = n53923 ^ n51070 ;
  assign n53979 = ~n53977 & n53978 ;
  assign n53980 = n53927 ^ n53926 ;
  assign n53981 = ~n53979 & n53980 ;
  assign n53982 = n53932 ^ n53907 ;
  assign n53983 = ~n53981 & n53982 ;
  assign n53984 = n53934 ^ n53906 ;
  assign n53985 = ~n53983 & ~n53984 ;
  assign n53986 = n53939 ^ n53904 ;
  assign n53987 = n53985 & n53986 ;
  assign n53988 = n53941 ^ n51386 ;
  assign n53989 = n53988 ^ n53902 ;
  assign n53990 = n53987 & n53989 ;
  assign n53991 = n53901 ^ n51377 ;
  assign n53992 = n53991 ^ n53944 ;
  assign n53993 = ~n53990 & ~n53992 ;
  assign n53994 = n53950 ^ n51328 ;
  assign n53995 = n53993 & ~n53994 ;
  assign n53996 = ~n53973 & n53995 ;
  assign n53953 = n53952 ^ n53898 ;
  assign n53954 = n53952 ^ n51323 ;
  assign n53955 = n53953 & n53954 ;
  assign n53956 = n53955 ^ n51323 ;
  assign n53894 = n52563 ^ n51938 ;
  assign n53895 = n53894 ^ n53344 ;
  assign n53268 = n53267 ^ n53246 ;
  assign n53269 = n53268 ^ n53239 ;
  assign n53270 = n53269 ^ n53268 ;
  assign n53891 = n53890 ^ n53270 ;
  assign n53892 = n53243 & ~n53891 ;
  assign n53893 = n53892 ^ n53269 ;
  assign n53896 = n53895 ^ n53893 ;
  assign n53897 = n53896 ^ n51318 ;
  assign n53971 = n53956 ^ n53897 ;
  assign n54020 = n53996 ^ n53971 ;
  assign n54024 = n54023 ^ n54020 ;
  assign n54028 = n53995 ^ n53973 ;
  assign n54117 = n54028 ^ n54023 ;
  assign n54025 = n52071 ^ n44359 ;
  assign n54026 = n54025 ^ n48681 ;
  assign n54027 = n54026 ^ n42926 ;
  assign n54029 = n54028 ^ n54027 ;
  assign n54033 = n53994 ^ n53993 ;
  assign n54114 = n54033 ^ n54027 ;
  assign n54030 = n52076 ^ n44417 ;
  assign n54031 = n54030 ^ n48686 ;
  assign n54032 = n54031 ^ n42931 ;
  assign n54034 = n54033 ^ n54032 ;
  assign n54039 = n53992 ^ n53990 ;
  assign n54035 = n52081 ^ n44364 ;
  assign n54036 = n54035 ^ n48691 ;
  assign n54037 = n54036 ^ n42936 ;
  assign n54040 = n54039 ^ n54037 ;
  assign n54044 = n53989 ^ n53987 ;
  assign n54041 = n52086 ^ n44408 ;
  assign n54042 = n54041 ^ n48334 ;
  assign n54043 = n54042 ^ n2132 ;
  assign n54045 = n54044 ^ n54043 ;
  assign n54049 = n53986 ^ n53985 ;
  assign n54046 = n52091 ^ n44371 ;
  assign n54047 = n54046 ^ n47700 ;
  assign n54048 = n54047 ^ n42943 ;
  assign n54050 = n54049 ^ n54048 ;
  assign n54054 = n53984 ^ n53983 ;
  assign n54051 = n52097 ^ n44376 ;
  assign n54052 = n54051 ^ n48288 ;
  assign n54053 = n54052 ^ n42947 ;
  assign n54055 = n54054 ^ n54053 ;
  assign n54057 = n52102 ^ n44381 ;
  assign n54058 = n54057 ^ n48293 ;
  assign n54059 = n54058 ^ n42952 ;
  assign n54056 = n53982 ^ n53981 ;
  assign n54060 = n54059 ^ n54056 ;
  assign n54064 = n53980 ^ n53979 ;
  assign n54097 = n54064 ^ n54059 ;
  assign n54061 = n52109 ^ n44387 ;
  assign n54062 = n54061 ^ n48297 ;
  assign n54063 = n54062 ^ n42957 ;
  assign n54065 = n54064 ^ n54063 ;
  assign n54069 = n53978 ^ n53977 ;
  assign n54094 = n54069 ^ n54063 ;
  assign n54066 = n52113 ^ n43984 ;
  assign n54067 = n54066 ^ n48302 ;
  assign n54068 = n54067 ^ n42962 ;
  assign n54070 = n54069 ^ n54068 ;
  assign n54072 = n52118 ^ n2783 ;
  assign n54073 = n54072 ^ n48308 ;
  assign n54074 = n54073 ^ n42971 ;
  assign n54091 = n54074 ^ n54068 ;
  assign n54071 = n53976 ^ n53974 ;
  assign n54075 = n54074 ^ n54071 ;
  assign n54079 = n53912 ^ n50404 ;
  assign n54080 = n52487 ^ n44818 ;
  assign n54081 = n54080 ^ n49069 ;
  assign n54082 = n54081 ^ n43335 ;
  assign n54083 = ~n54079 & n54082 ;
  assign n54076 = n52122 ^ n43976 ;
  assign n54077 = n54076 ^ n48311 ;
  assign n54078 = n54077 ^ n42967 ;
  assign n54084 = n54083 ^ n54078 ;
  assign n54085 = n54074 ^ n53974 ;
  assign n54086 = n54085 ^ n54074 ;
  assign n54087 = n54086 ^ n54078 ;
  assign n54088 = ~n54084 & ~n54087 ;
  assign n54089 = n54088 ^ n54085 ;
  assign n54090 = ~n54075 & ~n54089 ;
  assign n54092 = n54091 ^ n54090 ;
  assign n54093 = ~n54070 & ~n54092 ;
  assign n54095 = n54094 ^ n54093 ;
  assign n54096 = n54065 & n54095 ;
  assign n54098 = n54097 ^ n54096 ;
  assign n54099 = ~n54060 & n54098 ;
  assign n54100 = n54099 ^ n54059 ;
  assign n54101 = n54100 ^ n54053 ;
  assign n54102 = ~n54055 & ~n54101 ;
  assign n54103 = n54102 ^ n54054 ;
  assign n54104 = n54103 ^ n54048 ;
  assign n54105 = ~n54050 & ~n54104 ;
  assign n54106 = n54105 ^ n54048 ;
  assign n54107 = n54106 ^ n54043 ;
  assign n54108 = ~n54045 & ~n54107 ;
  assign n54109 = n54108 ^ n54044 ;
  assign n54110 = n54109 ^ n54037 ;
  assign n54111 = n54040 & ~n54110 ;
  assign n54038 = n54037 ^ n54032 ;
  assign n54112 = n54111 ^ n54038 ;
  assign n54113 = ~n54034 & ~n54112 ;
  assign n54115 = n54114 ^ n54113 ;
  assign n54116 = ~n54029 & n54115 ;
  assign n54118 = n54117 ^ n54116 ;
  assign n54119 = n54024 & ~n54118 ;
  assign n54120 = n54119 ^ n54023 ;
  assign n53999 = n52059 ^ n44348 ;
  assign n54000 = n53999 ^ n48670 ;
  assign n54001 = n54000 ^ n42917 ;
  assign n53997 = n53971 & n53996 ;
  assign n53967 = n53756 ^ n53753 ;
  assign n53960 = n53342 ^ n52237 ;
  assign n53961 = n53960 ^ n51987 ;
  assign n53963 = n53961 ^ n53268 ;
  assign n53962 = n53961 ^ n53895 ;
  assign n53964 = n53963 ^ n53962 ;
  assign n53965 = n53893 & ~n53964 ;
  assign n53966 = n53965 ^ n53963 ;
  assign n53968 = n53967 ^ n53966 ;
  assign n53969 = n53968 ^ n51311 ;
  assign n53957 = n53956 ^ n53896 ;
  assign n53958 = n53897 & n53957 ;
  assign n53959 = n53958 ^ n51318 ;
  assign n53970 = n53969 ^ n53959 ;
  assign n53998 = n53997 ^ n53970 ;
  assign n54002 = n54001 ^ n53998 ;
  assign n54190 = n54120 ^ n54002 ;
  assign n54187 = n53786 ^ n53703 ;
  assign n54188 = n54187 ^ n52215 ;
  assign n54189 = n54188 ^ n53314 ;
  assign n54191 = n54190 ^ n54189 ;
  assign n54195 = n54118 ^ n54020 ;
  assign n54652 = n54195 ^ n54189 ;
  assign n54192 = n53783 ^ n53708 ;
  assign n54193 = n54192 ^ n53318 ;
  assign n54194 = n54193 ^ n52217 ;
  assign n54196 = n54195 ^ n54194 ;
  assign n54200 = n54115 ^ n54028 ;
  assign n54197 = n53781 ^ n53712 ;
  assign n54198 = n54197 ^ n52226 ;
  assign n54199 = n54198 ^ n53322 ;
  assign n54201 = n54200 ^ n54199 ;
  assign n54638 = n54112 ^ n54033 ;
  assign n54631 = n54109 ^ n54040 ;
  assign n54639 = n54638 ^ n54631 ;
  assign n54205 = n54106 ^ n54045 ;
  assign n54632 = n54631 ^ n54205 ;
  assign n54202 = n53771 ^ n53728 ;
  assign n54203 = n54202 ^ n52237 ;
  assign n54204 = n54203 ^ n53334 ;
  assign n54206 = n54205 ^ n54204 ;
  assign n54210 = n54103 ^ n54050 ;
  assign n54208 = n53768 ^ n53733 ;
  assign n54207 = n53336 ^ n52563 ;
  assign n54209 = n54208 ^ n54207 ;
  assign n54211 = n54210 ^ n54209 ;
  assign n54214 = n54100 ^ n54055 ;
  assign n54212 = n53342 ^ n52243 ;
  assign n54164 = n53765 ^ n53738 ;
  assign n54213 = n54212 ^ n54164 ;
  assign n54215 = n54214 ^ n54213 ;
  assign n54218 = n54098 ^ n54056 ;
  assign n54216 = n53344 ^ n52239 ;
  assign n54141 = n53763 ^ n53739 ;
  assign n54217 = n54216 ^ n54141 ;
  assign n54219 = n54218 ^ n54217 ;
  assign n54221 = n53241 ^ n52246 ;
  assign n54006 = n53759 ^ n53748 ;
  assign n54222 = n54221 ^ n54006 ;
  assign n54619 = n54222 ^ n54218 ;
  assign n54224 = n53967 ^ n52250 ;
  assign n54225 = n54224 ^ n53273 ;
  assign n54220 = n54092 ^ n54069 ;
  assign n54226 = n54225 ^ n54220 ;
  assign n54229 = n54089 ^ n54071 ;
  assign n54227 = n53277 ^ n52256 ;
  assign n54228 = n54227 ^ n53268 ;
  assign n54230 = n54229 ^ n54228 ;
  assign n54233 = n54078 ^ n53974 ;
  assign n54234 = n54233 ^ n54083 ;
  assign n54231 = n53239 ^ n52258 ;
  assign n54232 = n54231 ^ n53282 ;
  assign n54235 = n54234 ^ n54232 ;
  assign n54237 = n53271 ^ n52262 ;
  assign n54238 = n54237 ^ n53288 ;
  assign n54236 = n54082 ^ n54079 ;
  assign n54239 = n54238 ^ n54236 ;
  assign n54534 = n53080 ^ n52294 ;
  assign n54535 = n54534 ^ n51338 ;
  assign n54533 = n53805 ^ n53661 ;
  assign n54536 = n54535 ^ n54533 ;
  assign n54484 = n53800 ^ n53674 ;
  assign n54482 = n52499 ^ n51749 ;
  assign n54483 = n54482 ^ n53096 ;
  assign n54485 = n54484 ^ n54483 ;
  assign n54517 = n53084 ^ n52495 ;
  assign n54518 = n54517 ^ n51745 ;
  assign n54245 = n53833 ^ n51762 ;
  assign n54246 = n54245 ^ n52513 ;
  assign n54174 = n53794 ^ n53687 ;
  assign n54247 = n54246 ^ n54174 ;
  assign n54252 = n52507 ^ n51759 ;
  assign n54253 = n54252 ^ n53576 ;
  assign n54179 = n53792 ^ n53690 ;
  assign n54254 = n54253 ^ n54179 ;
  assign n54183 = n53789 ^ n53698 ;
  assign n54308 = n54183 ^ n54179 ;
  assign n54255 = n53446 ^ n52213 ;
  assign n54256 = n54255 ^ n53067 ;
  assign n54257 = n54256 ^ n54187 ;
  assign n54299 = n54256 ^ n54192 ;
  assign n54258 = n53440 ^ n52219 ;
  assign n54259 = n54258 ^ n52755 ;
  assign n54260 = n54259 ^ n54192 ;
  assign n54261 = n53310 ^ n52606 ;
  assign n54262 = n54261 ^ n52224 ;
  assign n54263 = n54262 ^ n54197 ;
  assign n54264 = n53777 ^ n53718 ;
  assign n54293 = n54264 ^ n54262 ;
  assign n54265 = n52325 ^ n52203 ;
  assign n54266 = n54265 ^ n53314 ;
  assign n54267 = n54266 ^ n54264 ;
  assign n54269 = n53318 ^ n52230 ;
  assign n54270 = n54269 ^ n52207 ;
  assign n54268 = n53775 ^ n53722 ;
  assign n54271 = n54270 ^ n54268 ;
  assign n54272 = n52235 ^ n52215 ;
  assign n54273 = n54272 ^ n53322 ;
  assign n54274 = n54273 ^ n54202 ;
  assign n54284 = n54273 ^ n54208 ;
  assign n54165 = n53330 ^ n52226 ;
  assign n54166 = n54165 ^ n52307 ;
  assign n54167 = n54166 ^ n54164 ;
  assign n54275 = n54208 ^ n54164 ;
  assign n54276 = n54275 ^ n54208 ;
  assign n54139 = n52233 ^ n52191 ;
  assign n54140 = n54139 ^ n53334 ;
  assign n54142 = n54141 ^ n54140 ;
  assign n54007 = n54006 ^ n53961 ;
  assign n54004 = n53967 ^ n53961 ;
  assign n54005 = n53966 & n54004 ;
  assign n54008 = n54007 ^ n54005 ;
  assign n54009 = n53336 ^ n52228 ;
  assign n54010 = n54009 ^ n52006 ;
  assign n54136 = n54010 ^ n54006 ;
  assign n54137 = n54008 & ~n54136 ;
  assign n54138 = n54137 ^ n54010 ;
  assign n54161 = n54140 ^ n54138 ;
  assign n54162 = ~n54142 & n54161 ;
  assign n54163 = n54162 ^ n54141 ;
  assign n54277 = n54276 ^ n54163 ;
  assign n54278 = n54167 & ~n54277 ;
  assign n54279 = n54278 ^ n54275 ;
  assign n54280 = n53326 ^ n52305 ;
  assign n54281 = n54280 ^ n52217 ;
  assign n54282 = n54281 ^ n54208 ;
  assign n54283 = ~n54279 & n54282 ;
  assign n54285 = n54284 ^ n54283 ;
  assign n54286 = ~n54274 & ~n54285 ;
  assign n54287 = n54286 ^ n54273 ;
  assign n54288 = n54287 ^ n54268 ;
  assign n54289 = n54271 & n54288 ;
  assign n54290 = n54289 ^ n54268 ;
  assign n54291 = n54290 ^ n54264 ;
  assign n54292 = ~n54267 & n54291 ;
  assign n54294 = n54293 ^ n54292 ;
  assign n54295 = ~n54263 & ~n54294 ;
  assign n54296 = n54295 ^ n54262 ;
  assign n54297 = n54296 ^ n54192 ;
  assign n54298 = n54260 & n54297 ;
  assign n54300 = n54299 ^ n54298 ;
  assign n54301 = ~n54257 & n54300 ;
  assign n54302 = n54301 ^ n54256 ;
  assign n54303 = n54302 ^ n54183 ;
  assign n54304 = n53115 ^ n52209 ;
  assign n54305 = n54304 ^ n53559 ;
  assign n54306 = n54305 ^ n54183 ;
  assign n54307 = n54303 & ~n54306 ;
  assign n54309 = n54308 ^ n54307 ;
  assign n54310 = n54254 & ~n54309 ;
  assign n54311 = n54310 ^ n54253 ;
  assign n54248 = n53093 ^ n51751 ;
  assign n54249 = n54248 ^ n52503 ;
  assign n54250 = n54249 ^ n54174 ;
  assign n54251 = n54250 ^ n54249 ;
  assign n54312 = n54311 ^ n54251 ;
  assign n54313 = ~n54247 & ~n54312 ;
  assign n54314 = n54313 ^ n54250 ;
  assign n54315 = n53797 ^ n53682 ;
  assign n54486 = n54315 ^ n54249 ;
  assign n54487 = n54314 & n54486 ;
  assign n54488 = n54487 ^ n54249 ;
  assign n54519 = n54518 ^ n54488 ;
  assign n54520 = n54519 ^ n54484 ;
  assign n54521 = n54520 ^ n54518 ;
  assign n54522 = ~n54485 & ~n54521 ;
  assign n54523 = n54522 ^ n54519 ;
  assign n54524 = n53802 ^ n53671 ;
  assign n54537 = n54524 ^ n54518 ;
  assign n54538 = ~n54523 & ~n54537 ;
  assign n54539 = n54538 ^ n54518 ;
  assign n54593 = n54539 ^ n54535 ;
  assign n54594 = ~n54536 & n54593 ;
  assign n54589 = n53129 ^ n50415 ;
  assign n54586 = n53831 ^ n52288 ;
  assign n54585 = n53809 ^ n53808 ;
  assign n54587 = n54586 ^ n54585 ;
  assign n54588 = n54587 ^ n54535 ;
  assign n54590 = n54589 ^ n54588 ;
  assign n54581 = n52416 ^ n44783 ;
  assign n54582 = n54581 ^ n48935 ;
  assign n54583 = n54582 ^ n43338 ;
  assign n54318 = n54311 ^ n54247 ;
  assign n54319 = n54318 ^ n51038 ;
  assign n54365 = n54309 ^ n54253 ;
  assign n54320 = n54300 ^ n54187 ;
  assign n54321 = n54320 ^ n51452 ;
  assign n54352 = n54296 ^ n54260 ;
  assign n54322 = n54294 ^ n54197 ;
  assign n54323 = n54322 ^ n51436 ;
  assign n54324 = n54290 ^ n54267 ;
  assign n54325 = n54324 ^ n51428 ;
  assign n54326 = n54287 ^ n54271 ;
  assign n54327 = n54326 ^ n51346 ;
  assign n54329 = n54281 ^ n54279 ;
  assign n54330 = n54329 ^ n51351 ;
  assign n54168 = n54167 ^ n54163 ;
  assign n54012 = n53968 ^ n53959 ;
  assign n54013 = ~n53969 & n54012 ;
  assign n54014 = n54013 ^ n51311 ;
  assign n54015 = n54014 ^ n51306 ;
  assign n54011 = n54010 ^ n54008 ;
  assign n54144 = n54014 ^ n54011 ;
  assign n54145 = n54015 & ~n54144 ;
  assign n54146 = n54145 ^ n51306 ;
  assign n54147 = n54146 ^ n51302 ;
  assign n54143 = n54142 ^ n54138 ;
  assign n54157 = n54146 ^ n54143 ;
  assign n54158 = n54147 & ~n54157 ;
  assign n54159 = n54158 ^ n51302 ;
  assign n54331 = n54168 ^ n54159 ;
  assign n54332 = n54329 ^ n51355 ;
  assign n54333 = n54332 ^ n54329 ;
  assign n54334 = n54333 ^ n54168 ;
  assign n54335 = n54331 & n54334 ;
  assign n54336 = n54335 ^ n54332 ;
  assign n54337 = n54330 & n54336 ;
  assign n54338 = n54337 ^ n51351 ;
  assign n54328 = n54285 ^ n54202 ;
  assign n54339 = n54338 ^ n54328 ;
  assign n54340 = n54338 ^ n51344 ;
  assign n54341 = ~n54339 & n54340 ;
  assign n54342 = n54341 ^ n51344 ;
  assign n54343 = n54342 ^ n54326 ;
  assign n54344 = n54327 & ~n54343 ;
  assign n54345 = n54344 ^ n51346 ;
  assign n54346 = n54345 ^ n54324 ;
  assign n54347 = ~n54325 & n54346 ;
  assign n54348 = n54347 ^ n51428 ;
  assign n54349 = n54348 ^ n54322 ;
  assign n54350 = ~n54323 & n54349 ;
  assign n54351 = n54350 ^ n51436 ;
  assign n54353 = n54352 ^ n54351 ;
  assign n54354 = n54352 ^ n51446 ;
  assign n54355 = n54353 & ~n54354 ;
  assign n54356 = n54355 ^ n51446 ;
  assign n54357 = n54356 ^ n54320 ;
  assign n54358 = ~n54321 & ~n54357 ;
  assign n54359 = n54358 ^ n51452 ;
  assign n54360 = n54359 ^ n51728 ;
  assign n54361 = n54306 ^ n54302 ;
  assign n54362 = n54361 ^ n54359 ;
  assign n54363 = ~n54360 & n54362 ;
  assign n54364 = n54363 ^ n51728 ;
  assign n54366 = n54365 ^ n54364 ;
  assign n54367 = n54365 ^ n51034 ;
  assign n54368 = n54366 & n54367 ;
  assign n54369 = n54368 ^ n51034 ;
  assign n54370 = n54369 ^ n54318 ;
  assign n54371 = n54319 & n54370 ;
  assign n54372 = n54371 ^ n51038 ;
  assign n54316 = n54315 ^ n54314 ;
  assign n54317 = n54316 ^ n51037 ;
  assign n54373 = n54372 ^ n54317 ;
  assign n54374 = n54356 ^ n54321 ;
  assign n54375 = n54354 ^ n54351 ;
  assign n54376 = n54348 ^ n54323 ;
  assign n54377 = n54342 ^ n54327 ;
  assign n54378 = n54328 ^ n51344 ;
  assign n54379 = n54378 ^ n54338 ;
  assign n54160 = n54159 ^ n51355 ;
  assign n54169 = n54168 ^ n54160 ;
  assign n54003 = n53970 & n53997 ;
  assign n54016 = n54015 ^ n54011 ;
  assign n54135 = ~n54003 & n54016 ;
  assign n54148 = n54147 ^ n54143 ;
  assign n54170 = n54135 & n54148 ;
  assign n54380 = ~n54169 & ~n54170 ;
  assign n54381 = n54336 ^ n51351 ;
  assign n54382 = ~n54380 & ~n54381 ;
  assign n54383 = ~n54379 & ~n54382 ;
  assign n54384 = ~n54377 & n54383 ;
  assign n54385 = n54345 ^ n54325 ;
  assign n54386 = n54384 & n54385 ;
  assign n54387 = ~n54376 & ~n54386 ;
  assign n54388 = ~n54375 & n54387 ;
  assign n54389 = n54374 & ~n54388 ;
  assign n54390 = n54361 ^ n54360 ;
  assign n54391 = n54389 & n54390 ;
  assign n54392 = n54367 ^ n54364 ;
  assign n54393 = ~n54391 & n54392 ;
  assign n54394 = n54369 ^ n54319 ;
  assign n54395 = ~n54393 & n54394 ;
  assign n54481 = ~n54373 & ~n54395 ;
  assign n54491 = n54372 ^ n54316 ;
  assign n54492 = ~n54317 & ~n54491 ;
  assign n54493 = n54492 ^ n51037 ;
  assign n54489 = n54488 ^ n54485 ;
  assign n54490 = n54489 ^ n51026 ;
  assign n54494 = n54493 ^ n54490 ;
  assign n54512 = ~n54481 & n54494 ;
  assign n54525 = n54524 ^ n54523 ;
  assign n54526 = n54525 ^ n51022 ;
  assign n54513 = n54493 ^ n54489 ;
  assign n54514 = n54493 ^ n51026 ;
  assign n54515 = n54513 & ~n54514 ;
  assign n54516 = n54515 ^ n51026 ;
  assign n54527 = n54526 ^ n54516 ;
  assign n54546 = n54512 & n54527 ;
  assign n54542 = n54525 ^ n54516 ;
  assign n54543 = ~n54526 & n54542 ;
  assign n54544 = n54543 ^ n51022 ;
  assign n54574 = n54546 ^ n54544 ;
  assign n54540 = n54539 ^ n54536 ;
  assign n54576 = n54544 ^ n54540 ;
  assign n54579 = n54574 & ~n54576 ;
  assign n54577 = n54576 ^ n54546 ;
  assign n54578 = n50415 & n54577 ;
  assign n54580 = n54579 ^ n54578 ;
  assign n54584 = n54583 ^ n54580 ;
  assign n54591 = n54590 ^ n54584 ;
  assign n54508 = n52420 ^ n44755 ;
  assign n54509 = n54508 ^ n48888 ;
  assign n54510 = n54509 ^ n43353 ;
  assign n54592 = n54591 ^ n54510 ;
  assign n54595 = n54594 ^ n54592 ;
  assign n54495 = n54494 ^ n54481 ;
  assign n54396 = n54395 ^ n54373 ;
  assign n54242 = n52435 ^ n44715 ;
  assign n54243 = n54242 ^ n48802 ;
  assign n54244 = n54243 ^ n43362 ;
  assign n54397 = n54396 ^ n54244 ;
  assign n54401 = n54394 ^ n54393 ;
  assign n54398 = n52440 ^ n44643 ;
  assign n54399 = n54398 ^ n48363 ;
  assign n54400 = n54399 ^ n43371 ;
  assign n54402 = n54401 ^ n54400 ;
  assign n54403 = n54392 ^ n54391 ;
  assign n1287 = n1286 ^ n1232 ;
  assign n1324 = n1323 ^ n1287 ;
  assign n1334 = n1333 ^ n1324 ;
  assign n54404 = n54403 ^ n1334 ;
  assign n54406 = n52448 ^ n44665 ;
  assign n54407 = n54406 ^ n48632 ;
  assign n54408 = n54407 ^ n1315 ;
  assign n54471 = n54408 ^ n1334 ;
  assign n54405 = n54390 ^ n54389 ;
  assign n54409 = n54408 ^ n54405 ;
  assign n54413 = n54388 ^ n54374 ;
  assign n54410 = n52202 ^ n1125 ;
  assign n54411 = n54410 ^ n1700 ;
  assign n54412 = n54411 ^ n43381 ;
  assign n54414 = n54413 ^ n54412 ;
  assign n54418 = n54387 ^ n54375 ;
  assign n54415 = n48751 ^ n44672 ;
  assign n54416 = n54415 ^ n52014 ;
  assign n54417 = n54416 ^ n1695 ;
  assign n54419 = n54418 ^ n54417 ;
  assign n54423 = n54386 ^ n54376 ;
  assign n54420 = n52018 ^ n1658 ;
  assign n54421 = n54420 ^ n48641 ;
  assign n54422 = n54421 ^ n43387 ;
  assign n54424 = n54423 ^ n54422 ;
  assign n54428 = n54385 ^ n54384 ;
  assign n54459 = n54428 ^ n54422 ;
  assign n54425 = n52023 ^ n44450 ;
  assign n54426 = n54425 ^ n48740 ;
  assign n54427 = n54426 ^ n43029 ;
  assign n54429 = n54428 ^ n54427 ;
  assign n54431 = n52028 ^ n44033 ;
  assign n54432 = n54431 ^ n48732 ;
  assign n54433 = n54432 ^ n2993 ;
  assign n54456 = n54433 ^ n54427 ;
  assign n54430 = n54383 ^ n54377 ;
  assign n54434 = n54433 ^ n54430 ;
  assign n54438 = n54382 ^ n54379 ;
  assign n54435 = n52034 ^ n44323 ;
  assign n54436 = n54435 ^ n48645 ;
  assign n54437 = n54436 ^ n42890 ;
  assign n54439 = n54438 ^ n54437 ;
  assign n54443 = n54381 ^ n54380 ;
  assign n54440 = n52039 ^ n44328 ;
  assign n54441 = n54440 ^ n48650 ;
  assign n54442 = n54441 ^ n42894 ;
  assign n54444 = n54443 ^ n54442 ;
  assign n54152 = n52044 ^ n44334 ;
  assign n54153 = n54152 ^ n48655 ;
  assign n54154 = n54153 ^ n42899 ;
  assign n54127 = n52049 ^ n44338 ;
  assign n54128 = n54127 ^ n48660 ;
  assign n54129 = n54128 ^ n42904 ;
  assign n54155 = n54154 ^ n54129 ;
  assign n54017 = n54016 ^ n54003 ;
  assign n54018 = n54017 ^ n54001 ;
  assign n54019 = n54018 ^ n54017 ;
  assign n54121 = n54120 ^ n54019 ;
  assign n54122 = n54002 & n54121 ;
  assign n54123 = n54122 ^ n54018 ;
  assign n54131 = n54129 ^ n54017 ;
  assign n54124 = n52054 ^ n44343 ;
  assign n54125 = n54124 ^ n48665 ;
  assign n54126 = n54125 ^ n42910 ;
  assign n54130 = n54129 ^ n54126 ;
  assign n54132 = n54131 ^ n54130 ;
  assign n54133 = n54123 & n54132 ;
  assign n54134 = n54133 ^ n54131 ;
  assign n54149 = n54148 ^ n54135 ;
  assign n54150 = n54149 ^ n54129 ;
  assign n54151 = n54134 & ~n54150 ;
  assign n54156 = n54155 ^ n54151 ;
  assign n54171 = n54170 ^ n54169 ;
  assign n54445 = n54171 ^ n54154 ;
  assign n54446 = ~n54156 & n54445 ;
  assign n54447 = n54446 ^ n54171 ;
  assign n54448 = n54447 ^ n54442 ;
  assign n54449 = ~n54444 & ~n54448 ;
  assign n54450 = n54449 ^ n54443 ;
  assign n54451 = n54450 ^ n54437 ;
  assign n54452 = n54439 & n54451 ;
  assign n54453 = n54452 ^ n54438 ;
  assign n54454 = n54453 ^ n54433 ;
  assign n54455 = ~n54434 & n54454 ;
  assign n54457 = n54456 ^ n54455 ;
  assign n54458 = n54429 & ~n54457 ;
  assign n54460 = n54459 ^ n54458 ;
  assign n54461 = ~n54424 & ~n54460 ;
  assign n54462 = n54461 ^ n54423 ;
  assign n54463 = n54462 ^ n54417 ;
  assign n54464 = n54419 & n54463 ;
  assign n54465 = n54464 ^ n54418 ;
  assign n54466 = n54465 ^ n54412 ;
  assign n54467 = ~n54414 & ~n54466 ;
  assign n54468 = n54467 ^ n54413 ;
  assign n54469 = n54468 ^ n54405 ;
  assign n54470 = n54409 & n54469 ;
  assign n54472 = n54471 ^ n54470 ;
  assign n54473 = n54404 & ~n54472 ;
  assign n54474 = n54473 ^ n54403 ;
  assign n54475 = n54474 ^ n54400 ;
  assign n54476 = ~n54402 & ~n54475 ;
  assign n54477 = n54476 ^ n54401 ;
  assign n54478 = n54477 ^ n54244 ;
  assign n54479 = ~n54397 & n54478 ;
  assign n54480 = n54479 ^ n54396 ;
  assign n54496 = n54495 ^ n54480 ;
  assign n54500 = n52431 ^ n44723 ;
  assign n54501 = n54500 ^ n48810 ;
  assign n54502 = n54501 ^ n43415 ;
  assign n54505 = n54502 ^ n54480 ;
  assign n54506 = ~n54496 & ~n54505 ;
  assign n54497 = n52425 ^ n43357 ;
  assign n54498 = n54497 ^ n48825 ;
  assign n54499 = n54498 ^ n44731 ;
  assign n54503 = n54502 ^ n54499 ;
  assign n54507 = n54506 ^ n54503 ;
  assign n54528 = n54527 ^ n54512 ;
  assign n54529 = n54528 ^ n54510 ;
  assign n54511 = n54510 ^ n54499 ;
  assign n54530 = n54529 ^ n54511 ;
  assign n54531 = n54507 & n54530 ;
  assign n54532 = n54531 ^ n54511 ;
  assign n54541 = n54540 ^ n50415 ;
  assign n54545 = n54544 ^ n54541 ;
  assign n54547 = n54546 ^ n54545 ;
  assign n54572 = n54547 ^ n54510 ;
  assign n54573 = n54532 & ~n54572 ;
  assign n54596 = n54595 ^ n54573 ;
  assign n54548 = n54547 ^ n54532 ;
  assign n54240 = n53284 ^ n52272 ;
  assign n54241 = n54240 ^ n53298 ;
  assign n54549 = n54548 ^ n54241 ;
  assign n54552 = n54528 ^ n54507 ;
  assign n54550 = n53303 ^ n53286 ;
  assign n54551 = n54550 ^ n52274 ;
  assign n54553 = n54552 ^ n54551 ;
  assign n54558 = n53295 ^ n52278 ;
  assign n54559 = n54558 ^ n53372 ;
  assign n54565 = n54559 ^ n54551 ;
  assign n54554 = n53257 ^ n52285 ;
  assign n54555 = n54554 ^ n53300 ;
  assign n54556 = n54477 ^ n54397 ;
  assign n54557 = ~n54555 & n54556 ;
  assign n54560 = n54559 ^ n54557 ;
  assign n54561 = n54502 ^ n54495 ;
  assign n54562 = n54561 ^ n54480 ;
  assign n54563 = n54562 ^ n54557 ;
  assign n54564 = ~n54560 & ~n54563 ;
  assign n54566 = n54565 ^ n54564 ;
  assign n54567 = n54553 & n54566 ;
  assign n54568 = n54567 ^ n54552 ;
  assign n54569 = n54568 ^ n54241 ;
  assign n54570 = ~n54549 & ~n54569 ;
  assign n54571 = n54570 ^ n54548 ;
  assign n54597 = n54596 ^ n54571 ;
  assign n54598 = n53292 ^ n52268 ;
  assign n54599 = n54598 ^ n53279 ;
  assign n54602 = n54599 ^ n54571 ;
  assign n54603 = ~n54597 & ~n54602 ;
  assign n54600 = n54599 ^ n54238 ;
  assign n54604 = n54603 ^ n54600 ;
  assign n54605 = n54239 & ~n54604 ;
  assign n54606 = n54605 ^ n54238 ;
  assign n54607 = n54606 ^ n54234 ;
  assign n54608 = n54235 & n54607 ;
  assign n54609 = n54608 ^ n54234 ;
  assign n54610 = n54609 ^ n54228 ;
  assign n54611 = ~n54230 & ~n54610 ;
  assign n54612 = n54611 ^ n54229 ;
  assign n54613 = n54612 ^ n54220 ;
  assign n54614 = ~n54226 & ~n54613 ;
  assign n54223 = n54222 ^ n54220 ;
  assign n54615 = n54614 ^ n54223 ;
  assign n54616 = n54095 ^ n54064 ;
  assign n54617 = n54616 ^ n54222 ;
  assign n54618 = ~n54615 & ~n54617 ;
  assign n54620 = n54619 ^ n54618 ;
  assign n54621 = n54219 & ~n54620 ;
  assign n54622 = n54621 ^ n54218 ;
  assign n54623 = n54622 ^ n54213 ;
  assign n54624 = n54215 & ~n54623 ;
  assign n54625 = n54624 ^ n54214 ;
  assign n54626 = n54625 ^ n54209 ;
  assign n54627 = ~n54211 & ~n54626 ;
  assign n54628 = n54627 ^ n54210 ;
  assign n54629 = n54628 ^ n54205 ;
  assign n54630 = ~n54206 & ~n54629 ;
  assign n54633 = n54632 ^ n54630 ;
  assign n54634 = n54268 ^ n53330 ;
  assign n54635 = n54634 ^ n52228 ;
  assign n54636 = n54635 ^ n54631 ;
  assign n54637 = n54633 & ~n54636 ;
  assign n54640 = n54639 ^ n54637 ;
  assign n54643 = n54264 ^ n53326 ;
  assign n54644 = n54643 ^ n52233 ;
  assign n54641 = n54638 ^ n54199 ;
  assign n54642 = n54641 ^ n54199 ;
  assign n54645 = n54644 ^ n54642 ;
  assign n54646 = n54640 & n54645 ;
  assign n54647 = n54646 ^ n54641 ;
  assign n54648 = ~n54201 & ~n54647 ;
  assign n54649 = n54648 ^ n54200 ;
  assign n54650 = n54649 ^ n54195 ;
  assign n54651 = ~n54196 & ~n54650 ;
  assign n54653 = n54652 ^ n54651 ;
  assign n54654 = n54191 & n54653 ;
  assign n54655 = n54654 ^ n54190 ;
  assign n54184 = n54183 ^ n53310 ;
  assign n54185 = n54184 ^ n52207 ;
  assign n54182 = n54126 ^ n54123 ;
  assign n54186 = n54185 ^ n54182 ;
  assign n54674 = n54655 ^ n54186 ;
  assign n54827 = n54674 ^ n52230 ;
  assign n54675 = n54653 ^ n54190 ;
  assign n54676 = n54675 ^ n52235 ;
  assign n54677 = n54649 ^ n54196 ;
  assign n54678 = n54677 ^ n52305 ;
  assign n54679 = n54647 ^ n54200 ;
  assign n54680 = n54679 ^ n52307 ;
  assign n54681 = n54644 ^ n54640 ;
  assign n54682 = n54681 ^ n52191 ;
  assign n54683 = n54635 ^ n54633 ;
  assign n54684 = n54683 ^ n52006 ;
  assign n54685 = n54628 ^ n54206 ;
  assign n54686 = n54685 ^ n51987 ;
  assign n54687 = n54625 ^ n54211 ;
  assign n54688 = n54687 ^ n51938 ;
  assign n54690 = n54616 ^ n54615 ;
  assign n54691 = n54690 ^ n51309 ;
  assign n54731 = n54612 ^ n54226 ;
  assign n54692 = n54609 ^ n54230 ;
  assign n54693 = n54692 ^ n51316 ;
  assign n54695 = n54604 ^ n54236 ;
  assign n54696 = n54695 ^ n51330 ;
  assign n54699 = n54568 ^ n54549 ;
  assign n54700 = n54699 ^ n51799 ;
  assign n54708 = n54566 ^ n54552 ;
  assign n54701 = n54556 ^ n54555 ;
  assign n54702 = n51780 & ~n54701 ;
  assign n54703 = n54702 ^ n51783 ;
  assign n54704 = n54562 ^ n54560 ;
  assign n54705 = n54704 ^ n54702 ;
  assign n54706 = ~n54703 & n54705 ;
  assign n54707 = n54706 ^ n51783 ;
  assign n54709 = n54708 ^ n54707 ;
  assign n54710 = n54708 ^ n51791 ;
  assign n54711 = ~n54709 & n54710 ;
  assign n54712 = n54711 ^ n51791 ;
  assign n54713 = n54712 ^ n54699 ;
  assign n54714 = n54700 & ~n54713 ;
  assign n54715 = n54714 ^ n51799 ;
  assign n54697 = n54599 ^ n54596 ;
  assign n54698 = n54697 ^ n54571 ;
  assign n54716 = n54715 ^ n54698 ;
  assign n54717 = n54715 ^ n51807 ;
  assign n54718 = n54716 & n54717 ;
  assign n54719 = n54718 ^ n51807 ;
  assign n54720 = n54719 ^ n54695 ;
  assign n54721 = ~n54696 & n54720 ;
  assign n54722 = n54721 ^ n51330 ;
  assign n54694 = n54606 ^ n54235 ;
  assign n54723 = n54722 ^ n54694 ;
  assign n54724 = n54692 ^ n51325 ;
  assign n54725 = n54724 ^ n54692 ;
  assign n54726 = n54725 ^ n54694 ;
  assign n54727 = ~n54723 & ~n54726 ;
  assign n54728 = n54727 ^ n54724 ;
  assign n54729 = n54693 & ~n54728 ;
  assign n54730 = n54729 ^ n51316 ;
  assign n54732 = n54731 ^ n54730 ;
  assign n54733 = n54690 ^ n51314 ;
  assign n54734 = n54733 ^ n54690 ;
  assign n54735 = n54734 ^ n54730 ;
  assign n54736 = n54732 & n54735 ;
  assign n54737 = n54736 ^ n54733 ;
  assign n54738 = ~n54691 & ~n54737 ;
  assign n54739 = n54738 ^ n51309 ;
  assign n54689 = n54620 ^ n54217 ;
  assign n54740 = n54739 ^ n54689 ;
  assign n54741 = n54622 ^ n54215 ;
  assign n54742 = n54741 ^ n51274 ;
  assign n54743 = n54742 ^ n54689 ;
  assign n54744 = n54743 ^ n54741 ;
  assign n54745 = n54740 & n54744 ;
  assign n54746 = n54745 ^ n54742 ;
  assign n54748 = n54687 ^ n51300 ;
  assign n54747 = n54741 ^ n54687 ;
  assign n54749 = n54748 ^ n54747 ;
  assign n54750 = n54746 & n54749 ;
  assign n54751 = n54750 ^ n54748 ;
  assign n54752 = n54688 & n54751 ;
  assign n54753 = n54752 ^ n51938 ;
  assign n54754 = n54753 ^ n54685 ;
  assign n54755 = n54686 & n54754 ;
  assign n54756 = n54755 ^ n51987 ;
  assign n54757 = n54756 ^ n54683 ;
  assign n54758 = ~n54684 & n54757 ;
  assign n54759 = n54758 ^ n52006 ;
  assign n54760 = n54759 ^ n54681 ;
  assign n54761 = ~n54682 & ~n54760 ;
  assign n54762 = n54761 ^ n52191 ;
  assign n54763 = n54762 ^ n54679 ;
  assign n54764 = ~n54680 & ~n54763 ;
  assign n54765 = n54764 ^ n52307 ;
  assign n54766 = n54765 ^ n54677 ;
  assign n54767 = ~n54678 & ~n54766 ;
  assign n54768 = n54767 ^ n52305 ;
  assign n54769 = n54768 ^ n54675 ;
  assign n54770 = ~n54676 & n54769 ;
  assign n54771 = n54770 ^ n52235 ;
  assign n54828 = n54827 ^ n54771 ;
  assign n54829 = n54751 ^ n51938 ;
  assign n54830 = n54746 ^ n51300 ;
  assign n54831 = n54737 ^ n51309 ;
  assign n54832 = n54731 ^ n51314 ;
  assign n54833 = n54832 ^ n54730 ;
  assign n54834 = n54728 ^ n51316 ;
  assign n54835 = n54719 ^ n54696 ;
  assign n54836 = n54698 ^ n51807 ;
  assign n54837 = n54836 ^ n54715 ;
  assign n54838 = n54704 ^ n54703 ;
  assign n54839 = n54710 ^ n54707 ;
  assign n54840 = ~n54838 & n54839 ;
  assign n54841 = n54712 ^ n54700 ;
  assign n54842 = ~n54840 & ~n54841 ;
  assign n54843 = ~n54837 & ~n54842 ;
  assign n54844 = n54835 & ~n54843 ;
  assign n54845 = n54722 ^ n51325 ;
  assign n54846 = n54845 ^ n54694 ;
  assign n54847 = ~n54844 & ~n54846 ;
  assign n54848 = ~n54834 & n54847 ;
  assign n54849 = n54833 & n54848 ;
  assign n54850 = ~n54831 & ~n54849 ;
  assign n54851 = n54689 ^ n51274 ;
  assign n54852 = n54851 ^ n54739 ;
  assign n54853 = n54850 & ~n54852 ;
  assign n54854 = n54830 & n54853 ;
  assign n54855 = ~n54829 & n54854 ;
  assign n54856 = n54753 ^ n54686 ;
  assign n54857 = n54855 & n54856 ;
  assign n54858 = n54756 ^ n54684 ;
  assign n54859 = ~n54857 & ~n54858 ;
  assign n54860 = n54759 ^ n54682 ;
  assign n54861 = n54859 & ~n54860 ;
  assign n54862 = n54762 ^ n52307 ;
  assign n54863 = n54862 ^ n54679 ;
  assign n54864 = ~n54861 & ~n54863 ;
  assign n54865 = n54765 ^ n52305 ;
  assign n54866 = n54865 ^ n54677 ;
  assign n54867 = ~n54864 & ~n54866 ;
  assign n54868 = n54768 ^ n54676 ;
  assign n54869 = ~n54867 & ~n54868 ;
  assign n54870 = n54828 & n54869 ;
  assign n54772 = n54771 ^ n54674 ;
  assign n54773 = n54771 ^ n52230 ;
  assign n54774 = n54772 & ~n54773 ;
  assign n54775 = n54774 ^ n52230 ;
  assign n54825 = n54775 ^ n52325 ;
  assign n54656 = n54655 ^ n54182 ;
  assign n54657 = ~n54186 & n54656 ;
  assign n54658 = n54657 ^ n54182 ;
  assign n54178 = n53440 ^ n52203 ;
  assign n54180 = n54179 ^ n54178 ;
  assign n54177 = n54149 ^ n54134 ;
  assign n54181 = n54180 ^ n54177 ;
  assign n54672 = n54658 ^ n54181 ;
  assign n54826 = n54825 ^ n54672 ;
  assign n54906 = n54870 ^ n54826 ;
  assign n54902 = n52877 ^ n45106 ;
  assign n54903 = n54902 ^ n49436 ;
  assign n54904 = n54903 ^ n43763 ;
  assign n54907 = n54906 ^ n54904 ;
  assign n54911 = n54869 ^ n54828 ;
  assign n54908 = n52883 ^ n45111 ;
  assign n54909 = n54908 ^ n49440 ;
  assign n54910 = n54909 ^ n43768 ;
  assign n54912 = n54911 ^ n54910 ;
  assign n54918 = n54868 ^ n54867 ;
  assign n54915 = n52887 ^ n45116 ;
  assign n54916 = n54915 ^ n49446 ;
  assign n54917 = n54916 ^ n43773 ;
  assign n54919 = n54918 ^ n54917 ;
  assign n54921 = n52892 ^ n45121 ;
  assign n54922 = n54921 ^ n49450 ;
  assign n54923 = n54922 ^ n43778 ;
  assign n55060 = n54923 ^ n54917 ;
  assign n54920 = n54866 ^ n54864 ;
  assign n54924 = n54923 ^ n54920 ;
  assign n54928 = n54863 ^ n54861 ;
  assign n54925 = n52897 ^ n45126 ;
  assign n54926 = n54925 ^ n49460 ;
  assign n54927 = n54926 ^ n43783 ;
  assign n54929 = n54928 ^ n54927 ;
  assign n54934 = n54860 ^ n54859 ;
  assign n54930 = n52902 ^ n45131 ;
  assign n54931 = n54930 ^ n49456 ;
  assign n54932 = n54931 ^ n43790 ;
  assign n54935 = n54934 ^ n54932 ;
  assign n54939 = n54858 ^ n54857 ;
  assign n54936 = n52907 ^ n45137 ;
  assign n54937 = n54936 ^ n49465 ;
  assign n54938 = n54937 ^ n43795 ;
  assign n54940 = n54939 ^ n54938 ;
  assign n54944 = n54856 ^ n54855 ;
  assign n55049 = n54944 ^ n54939 ;
  assign n54941 = n52912 ^ n45142 ;
  assign n54942 = n54941 ^ n49470 ;
  assign n54943 = n54942 ^ n43799 ;
  assign n54945 = n54944 ^ n54943 ;
  assign n54949 = n54854 ^ n54829 ;
  assign n55046 = n54949 ^ n54943 ;
  assign n54946 = n52917 ^ n45146 ;
  assign n54947 = n54946 ^ n49476 ;
  assign n54948 = n54947 ^ n43804 ;
  assign n54950 = n54949 ^ n54948 ;
  assign n54951 = n52922 ^ n45151 ;
  assign n54952 = n54951 ^ n2360 ;
  assign n54953 = n54952 ^ n43809 ;
  assign n55043 = n54953 ^ n54949 ;
  assign n54954 = n54853 ^ n54830 ;
  assign n54955 = n54954 ^ n54953 ;
  assign n54959 = n54852 ^ n54850 ;
  assign n54956 = n52927 ^ n45156 ;
  assign n54957 = n54956 ^ n49483 ;
  assign n54958 = n54957 ^ n2349 ;
  assign n54960 = n54959 ^ n54958 ;
  assign n54964 = n54849 ^ n54831 ;
  assign n54961 = n52932 ^ n2201 ;
  assign n54962 = n54961 ^ n49487 ;
  assign n54963 = n54962 ^ n43817 ;
  assign n54965 = n54964 ^ n54963 ;
  assign n54967 = n52937 ^ n45165 ;
  assign n54968 = n54967 ^ n49493 ;
  assign n54969 = n54968 ^ n43823 ;
  assign n54966 = n54848 ^ n54833 ;
  assign n54970 = n54969 ^ n54966 ;
  assign n54975 = n54847 ^ n54834 ;
  assign n54971 = n52942 ^ n45169 ;
  assign n54972 = n54971 ^ n49497 ;
  assign n54973 = n54972 ^ n43828 ;
  assign n54976 = n54975 ^ n54973 ;
  assign n54978 = n52948 ^ n45177 ;
  assign n54979 = n54978 ^ n49502 ;
  assign n54980 = n54979 ^ n43833 ;
  assign n54977 = n54846 ^ n54844 ;
  assign n54981 = n54980 ^ n54977 ;
  assign n54985 = n54843 ^ n54835 ;
  assign n54982 = n52954 ^ n45181 ;
  assign n54983 = n54982 ^ n49507 ;
  assign n54984 = n54983 ^ n43839 ;
  assign n54986 = n54985 ^ n54984 ;
  assign n55014 = n52958 ^ n45186 ;
  assign n55015 = n55014 ^ n48900 ;
  assign n55016 = n55015 ^ n43843 ;
  assign n54988 = n52963 ^ n45192 ;
  assign n54989 = n54988 ^ n48818 ;
  assign n54990 = n54989 ^ n43849 ;
  assign n55017 = n55016 ^ n54990 ;
  assign n54987 = n54841 ^ n54840 ;
  assign n54991 = n54990 ^ n54987 ;
  assign n54993 = n52968 ^ n45196 ;
  assign n54994 = n54993 ^ n48355 ;
  assign n54995 = n54994 ^ n43853 ;
  assign n54992 = n54839 ^ n54838 ;
  assign n54996 = n54995 ^ n54992 ;
  assign n55000 = n53114 ^ n45412 ;
  assign n55001 = n55000 ^ n49602 ;
  assign n55002 = n55001 ^ n44106 ;
  assign n55003 = n54701 ^ n51780 ;
  assign n55004 = n55002 & ~n55003 ;
  assign n54997 = n52971 ^ n45200 ;
  assign n54998 = n54997 ^ n48358 ;
  assign n54999 = n54998 ^ n43856 ;
  assign n55005 = n55004 ^ n54999 ;
  assign n55006 = n55004 ^ n54838 ;
  assign n55007 = ~n55005 & ~n55006 ;
  assign n55008 = n55007 ^ n54838 ;
  assign n55009 = n55008 ^ n54992 ;
  assign n55010 = n54996 & n55009 ;
  assign n55011 = n55010 ^ n54995 ;
  assign n55012 = n55011 ^ n54990 ;
  assign n55013 = n54991 & n55012 ;
  assign n55018 = n55017 ^ n55013 ;
  assign n55019 = n54842 ^ n54837 ;
  assign n55020 = n55019 ^ n54985 ;
  assign n55021 = n55020 ^ n55016 ;
  assign n55022 = n55021 ^ n54985 ;
  assign n55023 = ~n55018 & ~n55022 ;
  assign n55024 = n55023 ^ n55020 ;
  assign n55025 = ~n54986 & n55024 ;
  assign n55026 = n55025 ^ n54985 ;
  assign n55027 = n55026 ^ n54977 ;
  assign n55028 = ~n54981 & ~n55027 ;
  assign n55029 = n55028 ^ n54980 ;
  assign n55030 = n55029 ^ n54973 ;
  assign n55031 = n54976 & n55030 ;
  assign n54974 = n54973 ^ n54969 ;
  assign n55032 = n55031 ^ n54974 ;
  assign n55033 = ~n54970 & n55032 ;
  assign n55034 = n55033 ^ n54969 ;
  assign n55035 = n55034 ^ n54963 ;
  assign n55036 = n54965 & n55035 ;
  assign n55037 = n55036 ^ n54963 ;
  assign n55038 = n55037 ^ n54958 ;
  assign n55039 = ~n54960 & ~n55038 ;
  assign n55040 = n55039 ^ n54959 ;
  assign n55041 = n55040 ^ n54953 ;
  assign n55042 = n54955 & ~n55041 ;
  assign n55044 = n55043 ^ n55042 ;
  assign n55045 = ~n54950 & ~n55044 ;
  assign n55047 = n55046 ^ n55045 ;
  assign n55048 = n54945 & n55047 ;
  assign n55050 = n55049 ^ n55048 ;
  assign n55051 = ~n54940 & ~n55050 ;
  assign n55052 = n55051 ^ n54939 ;
  assign n55053 = n55052 ^ n54932 ;
  assign n55054 = n54935 & ~n55053 ;
  assign n54933 = n54932 ^ n54928 ;
  assign n55055 = n55054 ^ n54933 ;
  assign n55056 = n54929 & n55055 ;
  assign n55057 = n55056 ^ n54928 ;
  assign n55058 = n55057 ^ n54920 ;
  assign n55059 = ~n54924 & n55058 ;
  assign n55061 = n55060 ^ n55059 ;
  assign n55062 = n54919 & ~n55061 ;
  assign n55063 = n55062 ^ n54918 ;
  assign n54913 = n54910 ^ n54904 ;
  assign n54914 = n54913 ^ n54904 ;
  assign n55064 = n55063 ^ n54914 ;
  assign n55065 = n54912 & n55064 ;
  assign n55066 = n55065 ^ n54913 ;
  assign n55067 = n54907 & n55066 ;
  assign n54871 = n54826 & n54870 ;
  assign n54673 = n54672 ^ n52325 ;
  assign n54776 = n54775 ^ n54672 ;
  assign n54777 = ~n54673 & ~n54776 ;
  assign n54778 = n54777 ^ n52325 ;
  assign n54780 = n54778 ^ n52224 ;
  assign n54659 = n54658 ^ n54177 ;
  assign n54660 = ~n54181 & n54659 ;
  assign n54661 = n54660 ^ n54180 ;
  assign n54173 = n53446 ^ n52606 ;
  assign n54175 = n54174 ^ n54173 ;
  assign n54172 = n54171 ^ n54156 ;
  assign n54176 = n54175 ^ n54172 ;
  assign n54671 = n54661 ^ n54176 ;
  assign n54824 = n54780 ^ n54671 ;
  assign n54897 = n54871 ^ n54824 ;
  assign n54905 = n54904 ^ n54897 ;
  assign n55068 = n55067 ^ n54905 ;
  assign n54898 = n52873 ^ n45101 ;
  assign n54899 = n54898 ^ n49431 ;
  assign n54900 = n54899 ^ n893 ;
  assign n55666 = n55068 ^ n54900 ;
  assign n55667 = n55666 ^ n54484 ;
  assign n55169 = n54465 ^ n54414 ;
  assign n55668 = n55667 ^ n55169 ;
  assign n55322 = n54202 ^ n54200 ;
  assign n55323 = n55322 ^ n53342 ;
  assign n55132 = n55024 ^ n54984 ;
  assign n55130 = n54638 ^ n54208 ;
  assign n55131 = n55130 ^ n53344 ;
  assign n55133 = n55132 ^ n55131 ;
  assign n55139 = n55019 ^ n55018 ;
  assign n55137 = n54631 ^ n54164 ;
  assign n55138 = n55137 ^ n53241 ;
  assign n55140 = n55139 ^ n55138 ;
  assign n55142 = n54141 ^ n53273 ;
  assign n55143 = n55142 ^ n54205 ;
  assign n55314 = n55143 ^ n55138 ;
  assign n55141 = n55011 ^ n54991 ;
  assign n55144 = n55143 ^ n55141 ;
  assign n55145 = n55008 ^ n54996 ;
  assign n55311 = n55145 ^ n55143 ;
  assign n55146 = n54006 ^ n53277 ;
  assign n55147 = n55146 ^ n54210 ;
  assign n55148 = n55147 ^ n55145 ;
  assign n55151 = n54999 ^ n54838 ;
  assign n55152 = n55151 ^ n55004 ;
  assign n55149 = n54214 ^ n53967 ;
  assign n55150 = n55149 ^ n53282 ;
  assign n55153 = n55152 ^ n55150 ;
  assign n55156 = n55003 ^ n55002 ;
  assign n55154 = n53288 ^ n53268 ;
  assign n55155 = n55154 ^ n54218 ;
  assign n55157 = n55156 ^ n55155 ;
  assign n55209 = n54472 ^ n54403 ;
  assign n55207 = n53847 ^ n52294 ;
  assign n55208 = n55207 ^ n53152 ;
  assign n55210 = n55209 ^ n55208 ;
  assign n55165 = n54468 ^ n54409 ;
  assign n55163 = n53851 ^ n53129 ;
  assign n55164 = n55163 ^ n52495 ;
  assign n55166 = n55165 ^ n55164 ;
  assign n55167 = n53080 ^ n52499 ;
  assign n55168 = n55167 ^ n53860 ;
  assign n55170 = n55169 ^ n55168 ;
  assign n55173 = n54462 ^ n54419 ;
  assign n55171 = n53084 ^ n52503 ;
  assign n55172 = n55171 ^ n53855 ;
  assign n55174 = n55173 ^ n55172 ;
  assign n55091 = n54585 ^ n52513 ;
  assign n55092 = n55091 ^ n53096 ;
  assign n54809 = n54457 ^ n54428 ;
  assign n55093 = n55092 ^ n54809 ;
  assign n54791 = n54450 ^ n54439 ;
  assign n54789 = n53576 ^ n53067 ;
  assign n54790 = n54789 ^ n54484 ;
  assign n54792 = n54791 ^ n54790 ;
  assign n54795 = n54453 ^ n54434 ;
  assign n54796 = n54795 ^ n54791 ;
  assign n54797 = n54796 ^ n54795 ;
  assign n54667 = n54447 ^ n54444 ;
  assign n54665 = n53559 ^ n52755 ;
  assign n54666 = n54665 ^ n54315 ;
  assign n54668 = n54667 ^ n54666 ;
  assign n54662 = n54661 ^ n54172 ;
  assign n54663 = n54176 & ~n54662 ;
  assign n54664 = n54663 ^ n54175 ;
  assign n54786 = n54666 ^ n54664 ;
  assign n54787 = ~n54668 & ~n54786 ;
  assign n54788 = n54787 ^ n54667 ;
  assign n54798 = n54797 ^ n54788 ;
  assign n54799 = ~n54792 & n54798 ;
  assign n54800 = n54799 ^ n54796 ;
  assign n54811 = n54809 ^ n54795 ;
  assign n54801 = n53833 ^ n53115 ;
  assign n54802 = n54801 ^ n54524 ;
  assign n54810 = n54809 ^ n54802 ;
  assign n54812 = n54811 ^ n54810 ;
  assign n54813 = n54800 & ~n54812 ;
  assign n54814 = n54813 ^ n54811 ;
  assign n54815 = n54533 ^ n52507 ;
  assign n54816 = n54815 ^ n53093 ;
  assign n55089 = n54816 ^ n54809 ;
  assign n55090 = ~n54814 & ~n55089 ;
  assign n55094 = n55093 ^ n55090 ;
  assign n55095 = n54460 ^ n54423 ;
  assign n55177 = n55095 ^ n55092 ;
  assign n55178 = ~n55094 & ~n55177 ;
  assign n55179 = n55178 ^ n55095 ;
  assign n55180 = n55179 ^ n55173 ;
  assign n55181 = ~n55174 & n55180 ;
  assign n55175 = n55173 ^ n55169 ;
  assign n55182 = n55181 ^ n55175 ;
  assign n55183 = ~n55170 & n55182 ;
  assign n55184 = n55183 ^ n55169 ;
  assign n55204 = n55184 ^ n55165 ;
  assign n55205 = ~n55166 & n55204 ;
  assign n55206 = n55205 ^ n55184 ;
  assign n55211 = n55210 ^ n55206 ;
  assign n55212 = n55211 ^ n51338 ;
  assign n55186 = n55182 ^ n55168 ;
  assign n55187 = n55186 ^ n51749 ;
  assign n55191 = n55179 ^ n55174 ;
  assign n55096 = n55095 ^ n55094 ;
  assign n55097 = n55096 ^ n51762 ;
  assign n54793 = n54792 ^ n54788 ;
  assign n54669 = n54668 ^ n54664 ;
  assign n54670 = n54669 ^ n52219 ;
  assign n54779 = n54778 ^ n54671 ;
  assign n54781 = ~n54779 & n54780 ;
  assign n54782 = n54781 ^ n52224 ;
  assign n54783 = n54782 ^ n54669 ;
  assign n54784 = ~n54670 & n54783 ;
  assign n54785 = n54784 ^ n52219 ;
  assign n54794 = n54793 ^ n54785 ;
  assign n54803 = n54802 ^ n54800 ;
  assign n54804 = n54803 ^ n52213 ;
  assign n54805 = n54804 ^ n54785 ;
  assign n54806 = n54805 ^ n54803 ;
  assign n54807 = ~n54794 & ~n54806 ;
  assign n54808 = n54807 ^ n54804 ;
  assign n54817 = n54816 ^ n54814 ;
  assign n54819 = n54817 ^ n52209 ;
  assign n54818 = n54817 ^ n54803 ;
  assign n54820 = n54819 ^ n54818 ;
  assign n54821 = n54808 & ~n54820 ;
  assign n54822 = n54821 ^ n54819 ;
  assign n55086 = n54817 ^ n51759 ;
  assign n55087 = n54822 & n55086 ;
  assign n55088 = n55087 ^ n51759 ;
  assign n55188 = n55096 ^ n55088 ;
  assign n55189 = n55097 & n55188 ;
  assign n55190 = n55189 ^ n51762 ;
  assign n55192 = n55191 ^ n55190 ;
  assign n55193 = n55186 ^ n51751 ;
  assign n55194 = n55193 ^ n55190 ;
  assign n55195 = n55194 ^ n55186 ;
  assign n55196 = n55192 & n55195 ;
  assign n55197 = n55196 ^ n55193 ;
  assign n55198 = ~n55187 & n55197 ;
  assign n55199 = n55198 ^ n51749 ;
  assign n55185 = n55184 ^ n55166 ;
  assign n55200 = n55199 ^ n55185 ;
  assign n55201 = n55199 ^ n51745 ;
  assign n55202 = ~n55200 & ~n55201 ;
  assign n55203 = n55202 ^ n51745 ;
  assign n55213 = n55212 ^ n55203 ;
  assign n55214 = n55197 ^ n51749 ;
  assign n55098 = n55097 ^ n55088 ;
  assign n54823 = n54822 ^ n51759 ;
  assign n54872 = ~n54824 & ~n54871 ;
  assign n54873 = n54782 ^ n54670 ;
  assign n54874 = n54872 & n54873 ;
  assign n54875 = n54785 ^ n52213 ;
  assign n54876 = n54875 ^ n54793 ;
  assign n54877 = ~n54874 & ~n54876 ;
  assign n54878 = n54808 ^ n52209 ;
  assign n54879 = n54877 & n54878 ;
  assign n55099 = n54823 & ~n54879 ;
  assign n55215 = n55098 & ~n55099 ;
  assign n55216 = n55191 ^ n51751 ;
  assign n55217 = n55216 ^ n55190 ;
  assign n55218 = ~n55215 & ~n55217 ;
  assign n55219 = n55214 & ~n55218 ;
  assign n55220 = n55185 ^ n51745 ;
  assign n55221 = n55220 ^ n55199 ;
  assign n55222 = n55219 & n55221 ;
  assign n55271 = n55213 & ~n55222 ;
  assign n55268 = n55211 ^ n55203 ;
  assign n55269 = ~n55212 & n55268 ;
  assign n55261 = n53078 ^ n45408 ;
  assign n55262 = n55261 ^ n49384 ;
  assign n55263 = n55262 ^ n44086 ;
  assign n55264 = n55263 ^ n51338 ;
  assign n55256 = n53231 ^ n52288 ;
  assign n55257 = n55256 ^ n53843 ;
  assign n55258 = n55257 ^ n55208 ;
  assign n55106 = n54474 ^ n54402 ;
  assign n55259 = n55258 ^ n55106 ;
  assign n55260 = n55259 ^ n51334 ;
  assign n55265 = n55264 ^ n55260 ;
  assign n55160 = n52831 ^ n45429 ;
  assign n55161 = n55160 ^ n49388 ;
  assign n55162 = n55161 ^ n44009 ;
  assign n55266 = n55265 ^ n55162 ;
  assign n55254 = n55208 ^ n55206 ;
  assign n55255 = n55210 & ~n55254 ;
  assign n55267 = n55266 ^ n55255 ;
  assign n55270 = n55269 ^ n55267 ;
  assign n55272 = n55271 ^ n55270 ;
  assign n55223 = n55222 ^ n55213 ;
  assign n55224 = n55223 ^ n55162 ;
  assign n55226 = n52835 ^ n45434 ;
  assign n55227 = n55226 ^ n49394 ;
  assign n55228 = n55227 ^ n43942 ;
  assign n55225 = n55221 ^ n55219 ;
  assign n55229 = n55228 ^ n55225 ;
  assign n55233 = n55218 ^ n55214 ;
  assign n55230 = n52840 ^ n45440 ;
  assign n55231 = n55230 ^ n49398 ;
  assign n55232 = n55231 ^ n2903 ;
  assign n55234 = n55233 ^ n55232 ;
  assign n55238 = n55217 ^ n55215 ;
  assign n55235 = n52845 ^ n45294 ;
  assign n55236 = n55235 ^ n49403 ;
  assign n55237 = n55236 ^ n43738 ;
  assign n55239 = n55238 ^ n55237 ;
  assign n55083 = n52851 ^ n1447 ;
  assign n55084 = n55083 ^ n49408 ;
  assign n55085 = n55084 ^ n43743 ;
  assign n55242 = n55237 ^ n55085 ;
  assign n55100 = n55099 ^ n55098 ;
  assign n55101 = n55100 ^ n55085 ;
  assign n54880 = n54879 ^ n54823 ;
  assign n1749 = n1748 ^ n1429 ;
  assign n1768 = n1767 ^ n1749 ;
  assign n1775 = n1774 ^ n1768 ;
  assign n54881 = n54880 ^ n1775 ;
  assign n54885 = n54878 ^ n54877 ;
  assign n55079 = n54885 ^ n54880 ;
  assign n54882 = n52857 ^ n45090 ;
  assign n54883 = n54882 ^ n49415 ;
  assign n54884 = n54883 ^ n1759 ;
  assign n54886 = n54885 ^ n54884 ;
  assign n54888 = n52862 ^ n1716 ;
  assign n54889 = n54888 ^ n49420 ;
  assign n54890 = n54889 ^ n43751 ;
  assign n55076 = n54890 ^ n54885 ;
  assign n54887 = n54876 ^ n54874 ;
  assign n54891 = n54890 ^ n54887 ;
  assign n54895 = n54873 ^ n54872 ;
  assign n55073 = n54895 ^ n54890 ;
  assign n54892 = n52867 ^ n45096 ;
  assign n54893 = n54892 ^ n49425 ;
  assign n54894 = n54893 ^ n43757 ;
  assign n54896 = n54895 ^ n54894 ;
  assign n55070 = n54900 ^ n54894 ;
  assign n54901 = n54900 ^ n54897 ;
  assign n55069 = ~n54901 & n55068 ;
  assign n55071 = n55070 ^ n55069 ;
  assign n55072 = ~n54896 & ~n55071 ;
  assign n55074 = n55073 ^ n55072 ;
  assign n55075 = n54891 & ~n55074 ;
  assign n55077 = n55076 ^ n55075 ;
  assign n55078 = n54886 & n55077 ;
  assign n55080 = n55079 ^ n55078 ;
  assign n55081 = n54881 & n55080 ;
  assign n55082 = n55081 ^ n54880 ;
  assign n55240 = n55085 ^ n55082 ;
  assign n55241 = ~n55101 & n55240 ;
  assign n55243 = n55242 ^ n55241 ;
  assign n55244 = ~n55239 & ~n55243 ;
  assign n55245 = n55244 ^ n55238 ;
  assign n55246 = n55245 ^ n55232 ;
  assign n55247 = ~n55234 & n55246 ;
  assign n55248 = n55247 ^ n55233 ;
  assign n55249 = n55248 ^ n55225 ;
  assign n55250 = n55229 & n55249 ;
  assign n55251 = n55250 ^ n55228 ;
  assign n55252 = n55251 ^ n55162 ;
  assign n55253 = n55224 & n55252 ;
  assign n55273 = n55272 ^ n55253 ;
  assign n55158 = n54616 ^ n53239 ;
  assign n55159 = n55158 ^ n53292 ;
  assign n55274 = n55273 ^ n55159 ;
  assign n55277 = n55251 ^ n55224 ;
  assign n55299 = n55277 ^ n55159 ;
  assign n55275 = n54220 ^ n53271 ;
  assign n55276 = n55275 ^ n53298 ;
  assign n55278 = n55277 ^ n55276 ;
  assign n55280 = n54229 ^ n53279 ;
  assign n55281 = n55280 ^ n53303 ;
  assign n55279 = n55248 ^ n55229 ;
  assign n55282 = n55281 ^ n55279 ;
  assign n55285 = n54236 ^ n53286 ;
  assign n55286 = n55285 ^ n53257 ;
  assign n55287 = n55243 ^ n55238 ;
  assign n55288 = ~n55286 & ~n55287 ;
  assign n55283 = n54234 ^ n53372 ;
  assign n55284 = n55283 ^ n53284 ;
  assign n55289 = n55288 ^ n55284 ;
  assign n55290 = n55245 ^ n55234 ;
  assign n55291 = n55290 ^ n55288 ;
  assign n55292 = ~n55289 & n55291 ;
  assign n55293 = n55292 ^ n55288 ;
  assign n55294 = n55293 ^ n55279 ;
  assign n55295 = ~n55282 & n55294 ;
  assign n55296 = n55295 ^ n55281 ;
  assign n55297 = n55296 ^ n55277 ;
  assign n55298 = n55278 & n55297 ;
  assign n55300 = n55299 ^ n55298 ;
  assign n55301 = n55274 & ~n55300 ;
  assign n55302 = n55301 ^ n55273 ;
  assign n55303 = n55302 ^ n55155 ;
  assign n55304 = n55157 & n55303 ;
  assign n55305 = n55304 ^ n55156 ;
  assign n55306 = n55305 ^ n55150 ;
  assign n55307 = n55153 & ~n55306 ;
  assign n55308 = n55307 ^ n55152 ;
  assign n55309 = n55308 ^ n55145 ;
  assign n55310 = ~n55148 & n55309 ;
  assign n55312 = n55311 ^ n55310 ;
  assign n55313 = ~n55144 & n55312 ;
  assign n55315 = n55314 ^ n55313 ;
  assign n55316 = ~n55140 & n55315 ;
  assign n55317 = n55316 ^ n55139 ;
  assign n55134 = n55026 ^ n54981 ;
  assign n55135 = n55134 ^ n55132 ;
  assign n55136 = n55135 ^ n55134 ;
  assign n55318 = n55317 ^ n55136 ;
  assign n55319 = ~n55133 & ~n55318 ;
  assign n55320 = n55319 ^ n55135 ;
  assign n55351 = n55323 ^ n55320 ;
  assign n55352 = n55351 ^ n52243 ;
  assign n55354 = n55315 ^ n55139 ;
  assign n55355 = n55354 ^ n52246 ;
  assign n55356 = n55312 ^ n55141 ;
  assign n55357 = n55356 ^ n52250 ;
  assign n55359 = n55305 ^ n55153 ;
  assign n55360 = n55359 ^ n52258 ;
  assign n55361 = n55302 ^ n55157 ;
  assign n55362 = n55361 ^ n52262 ;
  assign n55363 = n55300 ^ n55273 ;
  assign n55364 = n55363 ^ n52268 ;
  assign n55378 = n55296 ^ n55278 ;
  assign n55365 = n55293 ^ n55282 ;
  assign n55366 = n55365 ^ n52274 ;
  assign n55369 = n55290 ^ n55289 ;
  assign n55367 = n55287 ^ n55286 ;
  assign n55368 = n52285 & n55367 ;
  assign n55370 = n55369 ^ n55368 ;
  assign n55371 = n55365 ^ n52278 ;
  assign n55372 = n55371 ^ n55365 ;
  assign n55373 = n55372 ^ n55368 ;
  assign n55374 = n55370 & ~n55373 ;
  assign n55375 = n55374 ^ n55371 ;
  assign n55376 = ~n55366 & ~n55375 ;
  assign n55377 = n55376 ^ n52274 ;
  assign n55379 = n55378 ^ n55377 ;
  assign n55380 = n55363 ^ n52272 ;
  assign n55381 = n55380 ^ n55363 ;
  assign n55382 = n55381 ^ n55377 ;
  assign n55383 = ~n55379 & n55382 ;
  assign n55384 = n55383 ^ n55380 ;
  assign n55385 = ~n55364 & ~n55384 ;
  assign n55386 = n55385 ^ n52268 ;
  assign n55387 = n55386 ^ n55361 ;
  assign n55388 = ~n55362 & n55387 ;
  assign n55389 = n55388 ^ n52262 ;
  assign n55390 = n55389 ^ n55359 ;
  assign n55391 = n55360 & ~n55390 ;
  assign n55392 = n55391 ^ n52258 ;
  assign n55358 = n55308 ^ n55148 ;
  assign n55393 = n55392 ^ n55358 ;
  assign n55394 = n55356 ^ n52256 ;
  assign n55395 = n55394 ^ n55356 ;
  assign n55396 = n55395 ^ n55358 ;
  assign n55397 = n55393 & n55396 ;
  assign n55398 = n55397 ^ n55394 ;
  assign n55399 = n55357 & ~n55398 ;
  assign n55400 = n55399 ^ n52250 ;
  assign n55401 = n55400 ^ n55354 ;
  assign n55402 = ~n55355 & ~n55401 ;
  assign n55403 = n55402 ^ n52246 ;
  assign n55353 = n55317 ^ n55133 ;
  assign n55404 = n55403 ^ n55353 ;
  assign n55405 = n55403 ^ n52239 ;
  assign n55406 = n55404 & n55405 ;
  assign n55407 = n55406 ^ n52239 ;
  assign n55408 = n55407 ^ n55351 ;
  assign n55409 = n55352 & ~n55408 ;
  assign n55410 = n55409 ^ n52243 ;
  assign n55411 = n55410 ^ n52563 ;
  assign n55329 = n54268 ^ n53336 ;
  assign n55330 = n55329 ^ n54195 ;
  assign n55321 = n55029 ^ n54976 ;
  assign n55325 = n55321 ^ n55134 ;
  assign n55324 = n55323 ^ n55321 ;
  assign n55326 = n55325 ^ n55324 ;
  assign n55327 = n55320 & ~n55326 ;
  assign n55328 = n55327 ^ n55325 ;
  assign n55412 = n55330 ^ n55328 ;
  assign n55413 = n55412 ^ n55410 ;
  assign n55414 = n55411 & n55413 ;
  assign n55415 = n55414 ^ n52563 ;
  assign n55416 = n55415 ^ n52237 ;
  assign n55128 = n55032 ^ n54966 ;
  assign n55332 = n55321 ^ n55128 ;
  assign n55331 = n55330 ^ n55128 ;
  assign n55333 = n55332 ^ n55331 ;
  assign n55334 = n55328 & n55333 ;
  assign n55335 = n55334 ^ n55332 ;
  assign n55126 = n54264 ^ n53334 ;
  assign n55127 = n55126 ^ n54190 ;
  assign n55417 = n55335 ^ n55127 ;
  assign n55418 = n55417 ^ n55415 ;
  assign n55419 = ~n55416 & n55418 ;
  assign n55420 = n55419 ^ n52237 ;
  assign n55453 = n55420 ^ n52228 ;
  assign n55129 = n55128 ^ n55127 ;
  assign n55336 = n55129 & ~n55335 ;
  assign n55337 = n55336 ^ n55128 ;
  assign n55122 = n55034 ^ n54965 ;
  assign n55120 = n54197 ^ n53330 ;
  assign n55121 = n55120 ^ n54182 ;
  assign n55123 = n55122 ^ n55121 ;
  assign n55421 = n55337 ^ n55123 ;
  assign n55454 = n55453 ^ n55421 ;
  assign n55455 = n55417 ^ n55416 ;
  assign n55456 = n55412 ^ n55411 ;
  assign n55457 = n55368 ^ n52278 ;
  assign n55458 = n55457 ^ n55369 ;
  assign n55459 = n55375 ^ n52274 ;
  assign n55460 = ~n55458 & ~n55459 ;
  assign n55461 = n55378 ^ n52272 ;
  assign n55462 = n55461 ^ n55377 ;
  assign n55463 = ~n55460 & n55462 ;
  assign n55464 = n55384 ^ n52268 ;
  assign n55465 = ~n55463 & n55464 ;
  assign n55466 = n55386 ^ n55362 ;
  assign n55467 = ~n55465 & n55466 ;
  assign n55468 = n55389 ^ n55360 ;
  assign n55469 = ~n55467 & n55468 ;
  assign n55470 = n55358 ^ n52256 ;
  assign n55471 = n55470 ^ n55392 ;
  assign n55472 = n55469 & n55471 ;
  assign n55473 = n55398 ^ n52250 ;
  assign n55474 = n55472 & ~n55473 ;
  assign n55475 = n55400 ^ n55355 ;
  assign n55476 = ~n55474 & ~n55475 ;
  assign n55477 = n55404 ^ n52239 ;
  assign n55478 = n55476 & n55477 ;
  assign n55479 = n55407 ^ n52243 ;
  assign n55480 = n55479 ^ n55351 ;
  assign n55481 = n55478 & ~n55480 ;
  assign n55482 = n55456 & n55481 ;
  assign n55483 = ~n55455 & n55482 ;
  assign n55484 = n55454 & ~n55483 ;
  assign n55422 = n55421 ^ n55420 ;
  assign n55423 = n55421 ^ n52228 ;
  assign n55424 = ~n55422 & ~n55423 ;
  assign n55425 = n55424 ^ n52228 ;
  assign n55451 = n55425 ^ n52233 ;
  assign n55338 = n55337 ^ n55122 ;
  assign n55339 = ~n55123 & ~n55338 ;
  assign n55116 = n54177 ^ n53326 ;
  assign n55117 = n55116 ^ n54192 ;
  assign n55124 = n55122 ^ n55117 ;
  assign n55340 = n55339 ^ n55124 ;
  assign n55118 = n55037 ^ n54960 ;
  assign n55426 = n55340 ^ n55118 ;
  assign n55452 = n55451 ^ n55426 ;
  assign n55504 = n55484 ^ n55452 ;
  assign n55501 = n53721 ^ n45787 ;
  assign n55502 = n55501 ^ n50129 ;
  assign n55503 = n55502 ^ n44338 ;
  assign n55505 = n55504 ^ n55503 ;
  assign n55509 = n55483 ^ n55454 ;
  assign n55506 = n53727 ^ n45791 ;
  assign n55507 = n55506 ^ n50135 ;
  assign n55508 = n55507 ^ n44343 ;
  assign n55510 = n55509 ^ n55508 ;
  assign n55514 = n55482 ^ n55455 ;
  assign n55511 = n53731 ^ n45796 ;
  assign n55512 = n55511 ^ n50139 ;
  assign n55513 = n55512 ^ n44348 ;
  assign n55515 = n55514 ^ n55513 ;
  assign n55519 = n55481 ^ n55456 ;
  assign n55516 = n53736 ^ n45801 ;
  assign n55517 = n55516 ^ n50144 ;
  assign n55518 = n55517 ^ n44353 ;
  assign n55520 = n55519 ^ n55518 ;
  assign n55522 = n53742 ^ n2430 ;
  assign n55523 = n55522 ^ n50150 ;
  assign n55524 = n55523 ^ n44359 ;
  assign n55612 = n55524 ^ n55519 ;
  assign n55521 = n55480 ^ n55478 ;
  assign n55525 = n55524 ^ n55521 ;
  assign n55595 = n55475 ^ n55474 ;
  assign n55530 = n55473 ^ n55472 ;
  assign n55527 = n53249 ^ n45819 ;
  assign n55528 = n55527 ^ n49718 ;
  assign n55529 = n55528 ^ n44408 ;
  assign n55531 = n55530 ^ n55529 ;
  assign n55535 = n55471 ^ n55469 ;
  assign n55591 = n55535 ^ n55530 ;
  assign n55532 = n53220 ^ n45824 ;
  assign n55533 = n55532 ^ n49724 ;
  assign n55534 = n55533 ^ n44371 ;
  assign n55536 = n55535 ^ n55534 ;
  assign n55538 = n53175 ^ n45828 ;
  assign n55539 = n55538 ^ n49728 ;
  assign n55540 = n55539 ^ n44376 ;
  assign n55588 = n55540 ^ n55534 ;
  assign n55537 = n55468 ^ n55467 ;
  assign n55541 = n55540 ^ n55537 ;
  assign n55545 = n55466 ^ n55465 ;
  assign n55542 = n53179 ^ n45833 ;
  assign n55543 = n55542 ^ n49733 ;
  assign n55544 = n55543 ^ n44381 ;
  assign n55546 = n55545 ^ n55544 ;
  assign n55550 = n55464 ^ n55463 ;
  assign n55582 = n55550 ^ n55545 ;
  assign n55547 = n53202 ^ n45838 ;
  assign n55548 = n55547 ^ n49738 ;
  assign n55549 = n55548 ^ n44387 ;
  assign n55551 = n55550 ^ n55549 ;
  assign n55553 = n53194 ^ n45844 ;
  assign n55554 = n55553 ^ n49744 ;
  assign n55555 = n55554 ^ n43984 ;
  assign n55579 = n55555 ^ n55550 ;
  assign n55552 = n55462 ^ n55460 ;
  assign n55556 = n55555 ^ n55552 ;
  assign n55559 = n53185 ^ n45848 ;
  assign n55560 = n55559 ^ n49748 ;
  assign n55561 = n55560 ^ n2783 ;
  assign n55557 = n55459 ^ n55458 ;
  assign n55562 = n55561 ^ n55557 ;
  assign n55566 = n53830 ^ n46154 ;
  assign n55567 = n55566 ^ n50366 ;
  assign n55568 = n55567 ^ n44818 ;
  assign n55569 = n55367 ^ n52285 ;
  assign n55570 = n55568 & n55569 ;
  assign n55563 = n53188 ^ n45852 ;
  assign n55564 = n55563 ^ n49752 ;
  assign n55565 = n55564 ^ n43976 ;
  assign n55571 = n55570 ^ n55565 ;
  assign n55572 = n55570 ^ n55458 ;
  assign n55573 = ~n55571 & ~n55572 ;
  assign n55574 = n55573 ^ n55458 ;
  assign n55575 = n55574 ^ n55557 ;
  assign n55576 = ~n55562 & n55575 ;
  assign n55558 = n55557 ^ n55555 ;
  assign n55577 = n55576 ^ n55558 ;
  assign n55578 = ~n55556 & ~n55577 ;
  assign n55580 = n55579 ^ n55578 ;
  assign n55581 = n55551 & n55580 ;
  assign n55583 = n55582 ^ n55581 ;
  assign n55584 = ~n55546 & ~n55583 ;
  assign n55585 = n55584 ^ n55545 ;
  assign n55586 = n55585 ^ n55537 ;
  assign n55587 = n55541 & n55586 ;
  assign n55589 = n55588 ^ n55587 ;
  assign n55590 = ~n55536 & ~n55589 ;
  assign n55592 = n55591 ^ n55590 ;
  assign n55593 = n55531 & ~n55592 ;
  assign n55594 = n55593 ^ n55530 ;
  assign n55596 = n55595 ^ n55594 ;
  assign n55597 = n53751 ^ n45813 ;
  assign n55598 = n55597 ^ n49714 ;
  assign n55599 = n55598 ^ n44364 ;
  assign n55600 = n55599 ^ n55594 ;
  assign n55601 = ~n55596 & n55600 ;
  assign n55602 = n55601 ^ n55599 ;
  assign n55609 = n55602 ^ n55524 ;
  assign n55526 = n55477 ^ n55476 ;
  assign n55603 = n55602 ^ n55526 ;
  assign n55604 = n53747 ^ n45809 ;
  assign n55605 = n55604 ^ n49800 ;
  assign n55606 = n55605 ^ n44417 ;
  assign n55607 = n55606 ^ n55602 ;
  assign n55608 = n55603 & n55607 ;
  assign n55610 = n55609 ^ n55608 ;
  assign n55611 = ~n55525 & n55610 ;
  assign n55613 = n55612 ^ n55611 ;
  assign n55614 = n55520 & n55613 ;
  assign n55615 = n55614 ^ n55519 ;
  assign n55616 = n55615 ^ n55513 ;
  assign n55617 = ~n55515 & ~n55616 ;
  assign n55618 = n55617 ^ n55514 ;
  assign n55619 = n55618 ^ n55508 ;
  assign n55620 = n55510 & n55619 ;
  assign n55621 = n55620 ^ n55509 ;
  assign n55622 = n55621 ^ n55503 ;
  assign n55623 = ~n55505 & ~n55622 ;
  assign n55624 = n55623 ^ n55504 ;
  assign n55119 = n55118 ^ n55117 ;
  assign n55341 = ~n55119 & ~n55340 ;
  assign n55342 = n55341 ^ n55118 ;
  assign n55114 = n55040 ^ n54955 ;
  assign n55112 = n54187 ^ n53322 ;
  assign n55113 = n55112 ^ n54172 ;
  assign n55115 = n55114 ^ n55113 ;
  assign n55431 = n55342 ^ n55115 ;
  assign n55433 = n55431 ^ n52226 ;
  assign n55427 = n55426 ^ n55425 ;
  assign n55428 = n55426 ^ n52233 ;
  assign n55429 = ~n55427 & n55428 ;
  assign n55430 = n55429 ^ n52233 ;
  assign n55486 = n55433 ^ n55430 ;
  assign n55485 = n55452 & n55484 ;
  assign n55499 = n55486 ^ n55485 ;
  assign n55496 = n53717 ^ n45780 ;
  assign n55497 = n55496 ^ n50124 ;
  assign n55498 = n55497 ^ n44334 ;
  assign n55500 = n55499 ^ n55498 ;
  assign n55665 = n55624 ^ n55500 ;
  assign n55669 = n55668 ^ n55665 ;
  assign n55671 = n55063 ^ n54912 ;
  assign n55672 = n55671 ^ n55095 ;
  assign n55673 = n55672 ^ n54174 ;
  assign n55670 = n55618 ^ n55510 ;
  assign n55674 = n55673 ^ n55670 ;
  assign n55681 = n55615 ^ n55515 ;
  assign n55678 = n55061 ^ n54918 ;
  assign n55679 = n55678 ^ n54179 ;
  assign n55680 = n55679 ^ n54809 ;
  assign n55682 = n55681 ^ n55680 ;
  assign n55686 = n55613 ^ n55518 ;
  assign n56073 = n55686 ^ n55681 ;
  assign n55684 = n54795 ^ n54183 ;
  assign n55683 = n55057 ^ n54924 ;
  assign n55685 = n55684 ^ n55683 ;
  assign n55687 = n55686 ^ n55685 ;
  assign n55690 = n54791 ^ n54187 ;
  assign n55689 = n55055 ^ n54927 ;
  assign n55691 = n55690 ^ n55689 ;
  assign n56070 = n55691 ^ n55685 ;
  assign n55688 = n55610 ^ n55521 ;
  assign n55692 = n55691 ^ n55688 ;
  assign n55696 = n55607 ^ n55526 ;
  assign n55693 = n55052 ^ n54935 ;
  assign n55694 = n55693 ^ n54192 ;
  assign n55695 = n55694 ^ n54667 ;
  assign n55697 = n55696 ^ n55695 ;
  assign n55700 = n55599 ^ n55596 ;
  assign n55646 = n55050 ^ n54938 ;
  assign n55698 = n55646 ^ n54172 ;
  assign n55699 = n55698 ^ n54197 ;
  assign n55701 = n55700 ^ n55699 ;
  assign n55704 = n55592 ^ n55529 ;
  assign n55702 = n54264 ^ n54177 ;
  assign n55445 = n55047 ^ n54944 ;
  assign n55703 = n55702 ^ n55445 ;
  assign n55705 = n55704 ^ n55703 ;
  assign n55708 = n55589 ^ n55535 ;
  assign n55345 = n55044 ^ n54948 ;
  assign n55706 = n55345 ^ n54182 ;
  assign n55707 = n55706 ^ n54268 ;
  assign n55709 = n55708 ^ n55707 ;
  assign n55712 = n55585 ^ n55541 ;
  assign n55710 = n55114 ^ n54202 ;
  assign n55711 = n55710 ^ n54190 ;
  assign n55713 = n55712 ^ n55711 ;
  assign n55716 = n55583 ^ n55544 ;
  assign n55714 = n54208 ^ n54195 ;
  assign n55715 = n55714 ^ n55118 ;
  assign n55717 = n55716 ^ n55715 ;
  assign n55720 = n55580 ^ n55549 ;
  assign n55718 = n55122 ^ n54164 ;
  assign n55719 = n55718 ^ n54200 ;
  assign n55721 = n55720 ^ n55719 ;
  assign n55723 = n55128 ^ n54638 ;
  assign n55724 = n55723 ^ n54141 ;
  assign n56046 = n55724 ^ n55719 ;
  assign n55722 = n55577 ^ n55552 ;
  assign n55725 = n55724 ^ n55722 ;
  assign n55728 = n55574 ^ n55562 ;
  assign n55726 = n54631 ^ n54006 ;
  assign n55727 = n55726 ^ n55321 ;
  assign n55729 = n55728 ^ n55727 ;
  assign n55732 = n55134 ^ n53967 ;
  assign n55733 = n55732 ^ n54205 ;
  assign n56040 = n55733 ^ n55727 ;
  assign n55730 = n55565 ^ n55458 ;
  assign n55731 = n55730 ^ n55570 ;
  assign n55734 = n55733 ^ n55731 ;
  assign n55735 = n55569 ^ n55568 ;
  assign n56037 = n55735 ^ n55733 ;
  assign n55736 = n55132 ^ n54210 ;
  assign n55737 = n55736 ^ n53268 ;
  assign n55738 = n55737 ^ n55735 ;
  assign n56004 = n55139 ^ n53239 ;
  assign n56005 = n56004 ^ n54214 ;
  assign n55853 = n53843 ^ n53129 ;
  assign n55854 = n55853 ^ n54552 ;
  assign n55105 = n55077 ^ n54884 ;
  assign n55855 = n55854 ^ n55105 ;
  assign n55795 = n54562 ^ n53080 ;
  assign n55796 = n55795 ^ n53847 ;
  assign n55657 = n55074 ^ n54887 ;
  assign n55797 = n55796 ^ n55657 ;
  assign n55742 = n53851 ^ n53084 ;
  assign n55743 = n55742 ^ n54556 ;
  assign n55661 = n55071 ^ n54895 ;
  assign n55744 = n55743 ^ n55661 ;
  assign n55745 = n55106 ^ n53096 ;
  assign n55746 = n55745 ^ n53860 ;
  assign n55747 = n55746 ^ n55666 ;
  assign n55750 = n55066 ^ n54906 ;
  assign n55748 = n55209 ^ n53093 ;
  assign n55749 = n55748 ^ n53855 ;
  assign n55751 = n55750 ^ n55749 ;
  assign n55752 = n55165 ^ n54585 ;
  assign n55753 = n55752 ^ n53833 ;
  assign n55754 = n55753 ^ n55671 ;
  assign n55755 = n54533 ^ n53576 ;
  assign n55756 = n55755 ^ n55169 ;
  assign n55757 = n55756 ^ n55678 ;
  assign n55758 = n55173 ^ n54524 ;
  assign n55759 = n55758 ^ n53559 ;
  assign n55760 = n55759 ^ n55683 ;
  assign n55761 = n55095 ^ n54484 ;
  assign n55762 = n55761 ^ n53446 ;
  assign n55763 = n55762 ^ n55689 ;
  assign n55764 = n54809 ^ n53440 ;
  assign n55765 = n55764 ^ n54315 ;
  assign n55766 = n55765 ^ n55693 ;
  assign n55647 = n55646 ^ n55445 ;
  assign n55446 = n55445 ^ n55345 ;
  assign n55346 = n55345 ^ n55114 ;
  assign n55343 = n55342 ^ n55114 ;
  assign n55344 = n55115 & n55343 ;
  assign n55347 = n55346 ^ n55344 ;
  assign n55348 = n54667 ^ n53318 ;
  assign n55349 = n55348 ^ n54183 ;
  assign n55443 = n55349 ^ n55345 ;
  assign n55444 = n55347 & ~n55443 ;
  assign n55447 = n55446 ^ n55444 ;
  assign n55441 = n54179 ^ n53314 ;
  assign n55442 = n55441 ^ n54791 ;
  assign n55644 = n55445 ^ n55442 ;
  assign n55645 = n55447 & n55644 ;
  assign n55648 = n55647 ^ n55645 ;
  assign n55767 = n55765 ^ n55646 ;
  assign n55768 = n55767 ^ n55765 ;
  assign n55642 = n54795 ^ n54174 ;
  assign n55643 = n55642 ^ n53310 ;
  assign n55769 = n55768 ^ n55643 ;
  assign n55770 = n55648 & ~n55769 ;
  assign n55771 = n55770 ^ n55767 ;
  assign n55772 = n55766 & ~n55771 ;
  assign n55773 = n55772 ^ n55693 ;
  assign n55774 = n55773 ^ n55762 ;
  assign n55775 = n55763 & n55774 ;
  assign n55776 = n55775 ^ n55689 ;
  assign n55777 = n55776 ^ n55759 ;
  assign n55778 = n55760 & n55777 ;
  assign n55779 = n55778 ^ n55683 ;
  assign n55780 = n55779 ^ n55756 ;
  assign n55781 = n55757 & n55780 ;
  assign n55782 = n55781 ^ n55678 ;
  assign n55783 = n55782 ^ n55671 ;
  assign n55784 = n55754 & ~n55783 ;
  assign n55785 = n55784 ^ n55753 ;
  assign n55786 = n55785 ^ n55749 ;
  assign n55787 = ~n55751 & n55786 ;
  assign n55788 = n55787 ^ n55750 ;
  assign n55789 = n55788 ^ n55666 ;
  assign n55790 = n55747 & n55789 ;
  assign n55791 = n55790 ^ n55746 ;
  assign n55792 = n55791 ^ n55661 ;
  assign n55793 = ~n55744 & ~n55792 ;
  assign n55794 = n55793 ^ n55743 ;
  assign n55850 = n55794 ^ n55657 ;
  assign n55851 = ~n55797 & n55850 ;
  assign n55852 = n55851 ^ n55796 ;
  assign n55856 = n55855 ^ n55852 ;
  assign n55798 = n55797 ^ n55794 ;
  assign n55799 = n55798 ^ n52499 ;
  assign n55800 = n55791 ^ n55744 ;
  assign n55801 = n55800 ^ n52503 ;
  assign n55802 = n55788 ^ n55747 ;
  assign n55803 = n55802 ^ n52513 ;
  assign n55805 = n55782 ^ n55754 ;
  assign n55806 = n55805 ^ n53115 ;
  assign n55807 = n55779 ^ n55757 ;
  assign n55808 = n55807 ^ n53067 ;
  assign n55810 = n55773 ^ n55763 ;
  assign n55811 = n55810 ^ n52606 ;
  assign n55432 = n55431 ^ n55430 ;
  assign n55434 = ~n55432 & ~n55433 ;
  assign n55435 = n55434 ^ n52226 ;
  assign n55350 = n55349 ^ n55347 ;
  assign n55436 = n55435 ^ n55350 ;
  assign n55437 = n55435 ^ n52217 ;
  assign n55438 = ~n55436 & ~n55437 ;
  assign n55439 = n55438 ^ n52217 ;
  assign n55440 = n55439 ^ n52215 ;
  assign n55448 = n55447 ^ n55442 ;
  assign n55638 = n55448 ^ n55439 ;
  assign n55639 = n55440 & ~n55638 ;
  assign n55640 = n55639 ^ n52215 ;
  assign n55641 = n55640 ^ n52207 ;
  assign n55649 = n55648 ^ n55643 ;
  assign n55813 = n55649 ^ n55640 ;
  assign n55814 = n55641 & n55813 ;
  assign n55815 = n55814 ^ n52207 ;
  assign n55812 = n55771 ^ n55693 ;
  assign n55816 = n55815 ^ n55812 ;
  assign n55817 = n55810 ^ n52203 ;
  assign n55818 = n55817 ^ n55810 ;
  assign n55819 = n55818 ^ n55812 ;
  assign n55820 = ~n55816 & ~n55819 ;
  assign n55821 = n55820 ^ n55817 ;
  assign n55822 = ~n55811 & n55821 ;
  assign n55823 = n55822 ^ n52606 ;
  assign n55809 = n55776 ^ n55760 ;
  assign n55824 = n55823 ^ n55809 ;
  assign n55825 = n55807 ^ n52755 ;
  assign n55826 = n55825 ^ n55807 ;
  assign n55827 = n55826 ^ n55809 ;
  assign n55828 = ~n55824 & n55827 ;
  assign n55829 = n55828 ^ n55825 ;
  assign n55830 = ~n55808 & n55829 ;
  assign n55831 = n55830 ^ n53067 ;
  assign n55832 = n55831 ^ n55805 ;
  assign n55833 = ~n55806 & ~n55832 ;
  assign n55834 = n55833 ^ n53115 ;
  assign n55804 = n55785 ^ n55751 ;
  assign n55835 = n55834 ^ n55804 ;
  assign n55836 = n55802 ^ n52507 ;
  assign n55837 = n55836 ^ n55802 ;
  assign n55838 = n55837 ^ n55804 ;
  assign n55839 = ~n55835 & ~n55838 ;
  assign n55840 = n55839 ^ n55836 ;
  assign n55841 = ~n55803 & ~n55840 ;
  assign n55842 = n55841 ^ n52513 ;
  assign n55843 = n55842 ^ n55800 ;
  assign n55844 = n55801 & n55843 ;
  assign n55845 = n55844 ^ n52503 ;
  assign n55846 = n55845 ^ n55798 ;
  assign n55847 = n55799 & n55846 ;
  assign n55848 = n55847 ^ n52499 ;
  assign n55882 = n55856 ^ n55848 ;
  assign n55890 = n55080 ^ n1775 ;
  assign n55883 = n53300 ^ n53152 ;
  assign n55884 = n55883 ^ n54548 ;
  assign n55885 = n55884 ^ n55105 ;
  assign n55886 = n55885 ^ n55884 ;
  assign n55887 = n55886 ^ n55852 ;
  assign n55888 = n55855 & n55887 ;
  assign n55889 = n55888 ^ n55885 ;
  assign n55891 = n55890 ^ n55889 ;
  assign n55892 = n55891 ^ n52495 ;
  assign n55893 = n55892 ^ n55848 ;
  assign n55894 = n55893 ^ n55891 ;
  assign n55895 = n55882 & n55894 ;
  assign n55896 = n55895 ^ n55892 ;
  assign n56000 = n55891 ^ n52294 ;
  assign n56001 = n55896 & ~n56000 ;
  assign n55995 = n54596 ^ n52294 ;
  assign n55990 = n53307 ^ n44783 ;
  assign n55102 = n55101 ^ n55082 ;
  assign n55988 = n55102 ^ n53295 ;
  assign n55989 = n55988 ^ n46091 ;
  assign n55991 = n55990 ^ n55989 ;
  assign n55992 = n55991 ^ n50337 ;
  assign n55993 = n55992 ^ n55256 ;
  assign n55994 = n55993 ^ n55884 ;
  assign n55996 = n55995 ^ n55994 ;
  assign n55739 = n53644 ^ n46095 ;
  assign n55740 = n55739 ^ n50276 ;
  assign n55741 = n55740 ^ n44755 ;
  assign n55997 = n55996 ^ n55741 ;
  assign n55849 = n55848 ^ n52495 ;
  assign n55857 = n55856 ^ n55849 ;
  assign n55858 = n55845 ^ n55799 ;
  assign n55859 = n55840 ^ n52513 ;
  assign n55860 = n55812 ^ n52203 ;
  assign n55861 = n55860 ^ n55815 ;
  assign n55650 = n55649 ^ n55641 ;
  assign n55449 = n55448 ^ n55440 ;
  assign n55450 = n55437 ^ n55350 ;
  assign n55487 = ~n55485 & n55486 ;
  assign n55488 = n55450 & ~n55487 ;
  assign n55651 = ~n55449 & ~n55488 ;
  assign n55862 = n55650 & n55651 ;
  assign n55863 = n55861 & n55862 ;
  assign n55864 = n55821 ^ n52606 ;
  assign n55865 = ~n55863 & n55864 ;
  assign n55866 = n55809 ^ n52755 ;
  assign n55867 = n55866 ^ n55823 ;
  assign n55868 = n55865 & ~n55867 ;
  assign n55869 = n55829 ^ n53067 ;
  assign n55870 = ~n55868 & ~n55869 ;
  assign n55871 = n55831 ^ n53115 ;
  assign n55872 = n55871 ^ n55805 ;
  assign n55873 = n55870 & ~n55872 ;
  assign n55874 = n55834 ^ n52507 ;
  assign n55875 = n55874 ^ n55804 ;
  assign n55876 = ~n55873 & ~n55875 ;
  assign n55877 = ~n55859 & ~n55876 ;
  assign n55878 = n55842 ^ n55801 ;
  assign n55879 = ~n55877 & n55878 ;
  assign n55880 = n55858 & ~n55879 ;
  assign n55881 = n55857 & n55880 ;
  assign n55897 = n55896 ^ n52294 ;
  assign n55987 = ~n55881 & ~n55897 ;
  assign n55998 = n55997 ^ n55987 ;
  assign n55985 = n55890 ^ n55884 ;
  assign n55986 = n55889 & n55985 ;
  assign n55999 = n55998 ^ n55986 ;
  assign n56002 = n56001 ^ n55999 ;
  assign n55898 = n55897 ^ n55881 ;
  assign n55899 = n55898 ^ n55741 ;
  assign n55903 = n55880 ^ n55857 ;
  assign n55900 = n53650 ^ n46101 ;
  assign n55901 = n55900 ^ n50248 ;
  assign n55902 = n55901 ^ n44731 ;
  assign n55904 = n55903 ^ n55902 ;
  assign n55909 = n55879 ^ n55858 ;
  assign n55905 = n53654 ^ n46105 ;
  assign n55906 = n55905 ^ n50070 ;
  assign n55907 = n55906 ^ n44723 ;
  assign n55910 = n55909 ^ n55907 ;
  assign n55914 = n55878 ^ n55877 ;
  assign n55911 = n53664 ^ n46110 ;
  assign n55912 = n55911 ^ n50066 ;
  assign n55913 = n55912 ^ n44715 ;
  assign n55915 = n55914 ^ n55913 ;
  assign n55919 = n55876 ^ n55859 ;
  assign n55974 = n55919 ^ n55913 ;
  assign n55916 = n53660 ^ n46116 ;
  assign n55917 = n55916 ^ n50075 ;
  assign n55918 = n55917 ^ n44643 ;
  assign n55920 = n55919 ^ n55918 ;
  assign n55924 = n55875 ^ n55873 ;
  assign n55921 = n53669 ^ n45940 ;
  assign n55922 = n55921 ^ n50080 ;
  assign n55923 = n55922 ^ n1286 ;
  assign n55925 = n55924 ^ n55923 ;
  assign n55929 = n55872 ^ n55870 ;
  assign n55926 = n53674 ^ n45301 ;
  assign n55927 = n55926 ^ n1136 ;
  assign n55928 = n55927 ^ n44665 ;
  assign n55930 = n55929 ^ n55928 ;
  assign n55932 = n53679 ^ n45747 ;
  assign n55933 = n55932 ^ n50087 ;
  assign n55934 = n55933 ^ n1125 ;
  assign n55965 = n55934 ^ n55929 ;
  assign n55931 = n55869 ^ n55868 ;
  assign n55935 = n55934 ^ n55931 ;
  assign n55939 = n55867 ^ n55865 ;
  assign n55936 = n53685 ^ n965 ;
  assign n55937 = n55936 ^ n50092 ;
  assign n55938 = n55937 ^ n44672 ;
  assign n55940 = n55939 ^ n55938 ;
  assign n55942 = n53690 ^ n45755 ;
  assign n55943 = n55942 ^ n50098 ;
  assign n55944 = n55943 ^ n1658 ;
  assign n55959 = n55944 ^ n55939 ;
  assign n55941 = n55864 ^ n55863 ;
  assign n55945 = n55944 ^ n55941 ;
  assign n55949 = n55862 ^ n55861 ;
  assign n55946 = n53695 ^ n45760 ;
  assign n55947 = n55946 ^ n50102 ;
  assign n55948 = n55947 ^ n44450 ;
  assign n55950 = n55949 ^ n55948 ;
  assign n55633 = n53701 ^ n45766 ;
  assign n55634 = n55633 ^ n50107 ;
  assign n55635 = n55634 ^ n44033 ;
  assign n55953 = n55948 ^ n55635 ;
  assign n55109 = n53706 ^ n45771 ;
  assign n55110 = n55109 ^ n50114 ;
  assign n55111 = n55110 ^ n44323 ;
  assign n55636 = n55635 ^ n55111 ;
  assign n55489 = n55488 ^ n55449 ;
  assign n55490 = n55489 ^ n55111 ;
  assign n55494 = n55487 ^ n55450 ;
  assign n55491 = n53711 ^ n45775 ;
  assign n55492 = n55491 ^ n50119 ;
  assign n55493 = n55492 ^ n44328 ;
  assign n55495 = n55494 ^ n55493 ;
  assign n55625 = n55624 ^ n55498 ;
  assign n55626 = ~n55500 & n55625 ;
  assign n55627 = n55626 ^ n55499 ;
  assign n55628 = n55627 ^ n55493 ;
  assign n55629 = n55495 & n55628 ;
  assign n55630 = n55629 ^ n55494 ;
  assign n55631 = n55630 ^ n55111 ;
  assign n55632 = n55490 & n55631 ;
  assign n55637 = n55636 ^ n55632 ;
  assign n55652 = n55651 ^ n55650 ;
  assign n55951 = n55652 ^ n55635 ;
  assign n55952 = n55637 & n55951 ;
  assign n55954 = n55953 ^ n55952 ;
  assign n55955 = n55950 & ~n55954 ;
  assign n55956 = n55955 ^ n55949 ;
  assign n55957 = n55956 ^ n55944 ;
  assign n55958 = n55945 & n55957 ;
  assign n55960 = n55959 ^ n55958 ;
  assign n55961 = n55940 & n55960 ;
  assign n55962 = n55961 ^ n55939 ;
  assign n55963 = n55962 ^ n55934 ;
  assign n55964 = n55935 & n55963 ;
  assign n55966 = n55965 ^ n55964 ;
  assign n55967 = ~n55930 & ~n55966 ;
  assign n55968 = n55967 ^ n55929 ;
  assign n55969 = n55968 ^ n55923 ;
  assign n55970 = ~n55925 & n55969 ;
  assign n55971 = n55970 ^ n55924 ;
  assign n55972 = n55971 ^ n55919 ;
  assign n55973 = n55920 & ~n55972 ;
  assign n55975 = n55974 ^ n55973 ;
  assign n55976 = n55915 & ~n55975 ;
  assign n55977 = n55976 ^ n55914 ;
  assign n55978 = n55977 ^ n55907 ;
  assign n55979 = ~n55910 & n55978 ;
  assign n55908 = n55907 ^ n55903 ;
  assign n55980 = n55979 ^ n55908 ;
  assign n55981 = n55904 & n55980 ;
  assign n55982 = n55981 ^ n55903 ;
  assign n55983 = n55982 ^ n55741 ;
  assign n55984 = ~n55899 & n55983 ;
  assign n56003 = n56002 ^ n55984 ;
  assign n56006 = n56005 ^ n56003 ;
  assign n56009 = n55982 ^ n55899 ;
  assign n56031 = n56009 ^ n56005 ;
  assign n56007 = n54218 ^ n53271 ;
  assign n56008 = n56007 ^ n55141 ;
  assign n56010 = n56009 ^ n56008 ;
  assign n56013 = n55980 ^ n55902 ;
  assign n56011 = n55145 ^ n53279 ;
  assign n56012 = n56011 ^ n54616 ;
  assign n56014 = n56013 ^ n56012 ;
  assign n56017 = n55975 ^ n55914 ;
  assign n56018 = n55156 ^ n53286 ;
  assign n56019 = n56018 ^ n54229 ;
  assign n56020 = n56017 & ~n56019 ;
  assign n56025 = n56020 ^ n56013 ;
  assign n56015 = n54220 ^ n53284 ;
  assign n56016 = n56015 ^ n55152 ;
  assign n56021 = n56020 ^ n56016 ;
  assign n56022 = n55977 ^ n55910 ;
  assign n56023 = n56022 ^ n56020 ;
  assign n56024 = ~n56021 & ~n56023 ;
  assign n56026 = n56025 ^ n56024 ;
  assign n56027 = n56014 & n56026 ;
  assign n56028 = n56027 ^ n56013 ;
  assign n56029 = n56028 ^ n56008 ;
  assign n56030 = n56010 & n56029 ;
  assign n56032 = n56031 ^ n56030 ;
  assign n56033 = ~n56006 & ~n56032 ;
  assign n56034 = n56033 ^ n56005 ;
  assign n56035 = n56034 ^ n55735 ;
  assign n56036 = n55738 & n56035 ;
  assign n56038 = n56037 ^ n56036 ;
  assign n56039 = n55734 & ~n56038 ;
  assign n56041 = n56040 ^ n56039 ;
  assign n56042 = n55729 & n56041 ;
  assign n56043 = n56042 ^ n55728 ;
  assign n56044 = n56043 ^ n55722 ;
  assign n56045 = n55725 & ~n56044 ;
  assign n56047 = n56046 ^ n56045 ;
  assign n56048 = ~n55721 & n56047 ;
  assign n56049 = n56048 ^ n55720 ;
  assign n56050 = n56049 ^ n55715 ;
  assign n56051 = ~n55717 & ~n56050 ;
  assign n56052 = n56051 ^ n55716 ;
  assign n56053 = n56052 ^ n55711 ;
  assign n56054 = n55713 & ~n56053 ;
  assign n56055 = n56054 ^ n55712 ;
  assign n56056 = n56055 ^ n55707 ;
  assign n56057 = ~n55709 & n56056 ;
  assign n56058 = n56057 ^ n55708 ;
  assign n56059 = n56058 ^ n55703 ;
  assign n56060 = n55705 & ~n56059 ;
  assign n56061 = n56060 ^ n55704 ;
  assign n56062 = n56061 ^ n55699 ;
  assign n56063 = n55701 & n56062 ;
  assign n56064 = n56063 ^ n55700 ;
  assign n56065 = n56064 ^ n55695 ;
  assign n56066 = n55697 & ~n56065 ;
  assign n56067 = n56066 ^ n55696 ;
  assign n56068 = n56067 ^ n55688 ;
  assign n56069 = ~n55692 & n56068 ;
  assign n56071 = n56070 ^ n56069 ;
  assign n56072 = n55687 & ~n56071 ;
  assign n56074 = n56073 ^ n56072 ;
  assign n56075 = ~n55682 & ~n56074 ;
  assign n56076 = n56075 ^ n55681 ;
  assign n55675 = n55621 ^ n55505 ;
  assign n55676 = n55675 ^ n55670 ;
  assign n55677 = n55676 ^ n55675 ;
  assign n56077 = n56076 ^ n55677 ;
  assign n56078 = ~n55674 & n56077 ;
  assign n56079 = n56078 ^ n55676 ;
  assign n56083 = n55675 ^ n55668 ;
  assign n56080 = n55750 ^ n54315 ;
  assign n56081 = n56080 ^ n55173 ;
  assign n56082 = n56081 ^ n55668 ;
  assign n56084 = n56083 ^ n56082 ;
  assign n56085 = n56079 & ~n56084 ;
  assign n56086 = n56085 ^ n56083 ;
  assign n56087 = n55669 & ~n56086 ;
  assign n56088 = n56087 ^ n55668 ;
  assign n55663 = n55627 ^ n55495 ;
  assign n55660 = n55165 ^ n54524 ;
  assign n55662 = n55661 ^ n55660 ;
  assign n55664 = n55663 ^ n55662 ;
  assign n56225 = n56088 ^ n55664 ;
  assign n56114 = n56086 ^ n55665 ;
  assign n56115 = n56114 ^ n53446 ;
  assign n56117 = n56076 ^ n55674 ;
  assign n56118 = n56117 ^ n53310 ;
  assign n56119 = n56074 ^ n55680 ;
  assign n56120 = n56119 ^ n53314 ;
  assign n56121 = n56071 ^ n55686 ;
  assign n56122 = n56121 ^ n53318 ;
  assign n56123 = n56067 ^ n55692 ;
  assign n56124 = n56123 ^ n53322 ;
  assign n56125 = n56064 ^ n55697 ;
  assign n56126 = n56125 ^ n53326 ;
  assign n56127 = n56061 ^ n55701 ;
  assign n56128 = n56127 ^ n53330 ;
  assign n56129 = n56058 ^ n55705 ;
  assign n56130 = n56129 ^ n53334 ;
  assign n56131 = n56055 ^ n55709 ;
  assign n56132 = n56131 ^ n53336 ;
  assign n56133 = n56052 ^ n55713 ;
  assign n56134 = n56133 ^ n53342 ;
  assign n56135 = n56049 ^ n55717 ;
  assign n56136 = n56135 ^ n53344 ;
  assign n56138 = n56043 ^ n55725 ;
  assign n56139 = n56138 ^ n53273 ;
  assign n56140 = n56041 ^ n55728 ;
  assign n56141 = n56140 ^ n53277 ;
  assign n56170 = n56038 ^ n55731 ;
  assign n56142 = n56034 ^ n55738 ;
  assign n56143 = n56142 ^ n53288 ;
  assign n56161 = n56032 ^ n56003 ;
  assign n56144 = n56028 ^ n56010 ;
  assign n56145 = n56144 ^ n53298 ;
  assign n56153 = n56026 ^ n56012 ;
  assign n56146 = n56019 ^ n56017 ;
  assign n56147 = n53257 & ~n56146 ;
  assign n56148 = n56147 ^ n53372 ;
  assign n56149 = n56022 ^ n56021 ;
  assign n56150 = n56149 ^ n56147 ;
  assign n56151 = ~n56148 & ~n56150 ;
  assign n56152 = n56151 ^ n53372 ;
  assign n56154 = n56153 ^ n56152 ;
  assign n56155 = n56153 ^ n53303 ;
  assign n56156 = n56154 & n56155 ;
  assign n56157 = n56156 ^ n53303 ;
  assign n56158 = n56157 ^ n56144 ;
  assign n56159 = ~n56145 & ~n56158 ;
  assign n56160 = n56159 ^ n53298 ;
  assign n56162 = n56161 ^ n56160 ;
  assign n56163 = n56142 ^ n53292 ;
  assign n56164 = n56163 ^ n56142 ;
  assign n56165 = n56164 ^ n56160 ;
  assign n56166 = n56162 & n56165 ;
  assign n56167 = n56166 ^ n56163 ;
  assign n56168 = n56143 & n56167 ;
  assign n56169 = n56168 ^ n53288 ;
  assign n56171 = n56170 ^ n56169 ;
  assign n56172 = n56140 ^ n53282 ;
  assign n56173 = n56172 ^ n56140 ;
  assign n56174 = n56173 ^ n56169 ;
  assign n56175 = ~n56171 & n56174 ;
  assign n56176 = n56175 ^ n56172 ;
  assign n56177 = n56141 & n56176 ;
  assign n56178 = n56177 ^ n53277 ;
  assign n56179 = n56178 ^ n56138 ;
  assign n56180 = n56139 & n56179 ;
  assign n56181 = n56180 ^ n53273 ;
  assign n56137 = n56047 ^ n55720 ;
  assign n56182 = n56181 ^ n56137 ;
  assign n56183 = n56135 ^ n53241 ;
  assign n56184 = n56183 ^ n56135 ;
  assign n56185 = n56184 ^ n56137 ;
  assign n56186 = n56182 & ~n56185 ;
  assign n56187 = n56186 ^ n56183 ;
  assign n56188 = ~n56136 & n56187 ;
  assign n56189 = n56188 ^ n53344 ;
  assign n56190 = n56189 ^ n56133 ;
  assign n56191 = n56134 & n56190 ;
  assign n56192 = n56191 ^ n53342 ;
  assign n56193 = n56192 ^ n56131 ;
  assign n56194 = n56132 & n56193 ;
  assign n56195 = n56194 ^ n53336 ;
  assign n56196 = n56195 ^ n56129 ;
  assign n56197 = ~n56130 & n56196 ;
  assign n56198 = n56197 ^ n53334 ;
  assign n56199 = n56198 ^ n56127 ;
  assign n56200 = ~n56128 & n56199 ;
  assign n56201 = n56200 ^ n53330 ;
  assign n56202 = n56201 ^ n56125 ;
  assign n56203 = ~n56126 & ~n56202 ;
  assign n56204 = n56203 ^ n53326 ;
  assign n56205 = n56204 ^ n56123 ;
  assign n56206 = ~n56124 & ~n56205 ;
  assign n56207 = n56206 ^ n53322 ;
  assign n56208 = n56207 ^ n56121 ;
  assign n56209 = ~n56122 & ~n56208 ;
  assign n56210 = n56209 ^ n53318 ;
  assign n56211 = n56210 ^ n56119 ;
  assign n56212 = ~n56120 & ~n56211 ;
  assign n56213 = n56212 ^ n53314 ;
  assign n56214 = n56213 ^ n56117 ;
  assign n56215 = n56118 & ~n56214 ;
  assign n56216 = n56215 ^ n53310 ;
  assign n56116 = n56081 ^ n56079 ;
  assign n56217 = n56216 ^ n56116 ;
  assign n56218 = n56114 ^ n53440 ;
  assign n56219 = n56218 ^ n56116 ;
  assign n56220 = n56219 ^ n56114 ;
  assign n56221 = ~n56217 & n56220 ;
  assign n56222 = n56221 ^ n56218 ;
  assign n56223 = n56115 & n56222 ;
  assign n56224 = n56223 ^ n53446 ;
  assign n56226 = n56225 ^ n56224 ;
  assign n55655 = n55630 ^ n55490 ;
  assign n56089 = n56088 ^ n55655 ;
  assign n56090 = n56089 ^ n55663 ;
  assign n56091 = n56090 ^ n55655 ;
  assign n56092 = ~n55664 & ~n56091 ;
  assign n56093 = n56092 ^ n56089 ;
  assign n55656 = n55209 ^ n54533 ;
  assign n55658 = n55657 ^ n55656 ;
  assign n56112 = n56093 ^ n55658 ;
  assign n56227 = n56112 ^ n53559 ;
  assign n56228 = n56227 ^ n56224 ;
  assign n56229 = n56228 ^ n56112 ;
  assign n56230 = n56226 & n56229 ;
  assign n56231 = n56230 ^ n56227 ;
  assign n56292 = n56231 ^ n53576 ;
  assign n56244 = n56222 ^ n53446 ;
  assign n56245 = n56149 ^ n56148 ;
  assign n56246 = n56155 ^ n56152 ;
  assign n56247 = n56245 & n56246 ;
  assign n56248 = n56157 ^ n56145 ;
  assign n56249 = ~n56247 & ~n56248 ;
  assign n56250 = n56161 ^ n53292 ;
  assign n56251 = n56250 ^ n56160 ;
  assign n56252 = ~n56249 & ~n56251 ;
  assign n56253 = n56167 ^ n53288 ;
  assign n56254 = ~n56252 & ~n56253 ;
  assign n56255 = n56170 ^ n53282 ;
  assign n56256 = n56255 ^ n56169 ;
  assign n56257 = ~n56254 & ~n56256 ;
  assign n56258 = n56176 ^ n53277 ;
  assign n56259 = n56257 & ~n56258 ;
  assign n56260 = n56178 ^ n56139 ;
  assign n56261 = n56259 & n56260 ;
  assign n56262 = n56137 ^ n53241 ;
  assign n56263 = n56262 ^ n56181 ;
  assign n56264 = ~n56261 & ~n56263 ;
  assign n56265 = n56187 ^ n53344 ;
  assign n56266 = n56264 & ~n56265 ;
  assign n56267 = n56189 ^ n56134 ;
  assign n56268 = n56266 & n56267 ;
  assign n56269 = n56192 ^ n56132 ;
  assign n56270 = n56268 & ~n56269 ;
  assign n56271 = n56195 ^ n56130 ;
  assign n56272 = n56270 & ~n56271 ;
  assign n56273 = n56198 ^ n56128 ;
  assign n56274 = ~n56272 & n56273 ;
  assign n56275 = n56201 ^ n56126 ;
  assign n56276 = n56274 & n56275 ;
  assign n56277 = n56204 ^ n56124 ;
  assign n56278 = ~n56276 & n56277 ;
  assign n56279 = n56207 ^ n56122 ;
  assign n56280 = ~n56278 & n56279 ;
  assign n56281 = n56210 ^ n56120 ;
  assign n56282 = ~n56280 & n56281 ;
  assign n56283 = n56213 ^ n56118 ;
  assign n56284 = n56282 & n56283 ;
  assign n56285 = n56216 ^ n53440 ;
  assign n56286 = n56285 ^ n56116 ;
  assign n56287 = n56284 & n56286 ;
  assign n56288 = ~n56244 & ~n56287 ;
  assign n56289 = n56225 ^ n53559 ;
  assign n56290 = n56289 ^ n56224 ;
  assign n56291 = n56288 & ~n56290 ;
  assign n56313 = n56292 ^ n56291 ;
  assign n56310 = n54417 ^ n46811 ;
  assign n56311 = n56310 ^ n50824 ;
  assign n56312 = n56311 ^ n1716 ;
  assign n56314 = n56313 ^ n56312 ;
  assign n56318 = n56290 ^ n56288 ;
  assign n56315 = n54422 ^ n1679 ;
  assign n56316 = n56315 ^ n50830 ;
  assign n56317 = n56316 ^ n45096 ;
  assign n56319 = n56318 ^ n56317 ;
  assign n56323 = n56287 ^ n56244 ;
  assign n56320 = n54427 ^ n46824 ;
  assign n56321 = n56320 ^ n50834 ;
  assign n56322 = n56321 ^ n45101 ;
  assign n56324 = n56323 ^ n56322 ;
  assign n56326 = n54433 ^ n46516 ;
  assign n56327 = n56326 ^ n50839 ;
  assign n56328 = n56327 ^ n45106 ;
  assign n56488 = n56328 ^ n56322 ;
  assign n56325 = n56286 ^ n56284 ;
  assign n56329 = n56328 ^ n56325 ;
  assign n56331 = n54437 ^ n45945 ;
  assign n56332 = n56331 ^ n50844 ;
  assign n56333 = n56332 ^ n45111 ;
  assign n56485 = n56333 ^ n56328 ;
  assign n56330 = n56283 ^ n56282 ;
  assign n56334 = n56333 ^ n56330 ;
  assign n56338 = n56281 ^ n56280 ;
  assign n56335 = n54442 ^ n46373 ;
  assign n56336 = n56335 ^ n50849 ;
  assign n56337 = n56336 ^ n45116 ;
  assign n56339 = n56338 ^ n56337 ;
  assign n56341 = n54154 ^ n46377 ;
  assign n56342 = n56341 ^ n50854 ;
  assign n56343 = n56342 ^ n45121 ;
  assign n56479 = n56343 ^ n56337 ;
  assign n56340 = n56279 ^ n56278 ;
  assign n56344 = n56343 ^ n56340 ;
  assign n56346 = n54129 ^ n46383 ;
  assign n56347 = n56346 ^ n50860 ;
  assign n56348 = n56347 ^ n45126 ;
  assign n56476 = n56348 ^ n56343 ;
  assign n56345 = n56277 ^ n56276 ;
  assign n56349 = n56348 ^ n56345 ;
  assign n56353 = n56275 ^ n56274 ;
  assign n56350 = n54126 ^ n46388 ;
  assign n56351 = n56350 ^ n50864 ;
  assign n56352 = n56351 ^ n45131 ;
  assign n56354 = n56353 ^ n56352 ;
  assign n56358 = n56273 ^ n56272 ;
  assign n56355 = n54001 ^ n46392 ;
  assign n56356 = n56355 ^ n50869 ;
  assign n56357 = n56356 ^ n45137 ;
  assign n56359 = n56358 ^ n56357 ;
  assign n56361 = n54023 ^ n46397 ;
  assign n56362 = n56361 ^ n50874 ;
  assign n56363 = n56362 ^ n45142 ;
  assign n56467 = n56363 ^ n56357 ;
  assign n56360 = n56271 ^ n56270 ;
  assign n56364 = n56363 ^ n56360 ;
  assign n56368 = n56269 ^ n56268 ;
  assign n56365 = n54027 ^ n50880 ;
  assign n56366 = n56365 ^ n46402 ;
  assign n56367 = n56366 ^ n45146 ;
  assign n56369 = n56368 ^ n56367 ;
  assign n56373 = n56267 ^ n56266 ;
  assign n56370 = n54032 ^ n46486 ;
  assign n56371 = n56370 ^ n50884 ;
  assign n56372 = n56371 ^ n45151 ;
  assign n56374 = n56373 ^ n56372 ;
  assign n56378 = n56265 ^ n56264 ;
  assign n56375 = n54037 ^ n46407 ;
  assign n56376 = n56375 ^ n50890 ;
  assign n56377 = n56376 ^ n45156 ;
  assign n56379 = n56378 ^ n56377 ;
  assign n56383 = n56263 ^ n56261 ;
  assign n56380 = n54043 ^ n46474 ;
  assign n56381 = n56380 ^ n50894 ;
  assign n56382 = n56381 ^ n2201 ;
  assign n56384 = n56383 ^ n56382 ;
  assign n56386 = n54048 ^ n46412 ;
  assign n56387 = n56386 ^ n50899 ;
  assign n56388 = n56387 ^ n45165 ;
  assign n56452 = n56388 ^ n56382 ;
  assign n56385 = n56260 ^ n56259 ;
  assign n56389 = n56388 ^ n56385 ;
  assign n56393 = n56258 ^ n56257 ;
  assign n56390 = n54053 ^ n46417 ;
  assign n56391 = n56390 ^ n50904 ;
  assign n56392 = n56391 ^ n45169 ;
  assign n56394 = n56393 ^ n56392 ;
  assign n56399 = n56253 ^ n56252 ;
  assign n56396 = n54063 ^ n46428 ;
  assign n56397 = n56396 ^ n50391 ;
  assign n56398 = n56397 ^ n45181 ;
  assign n56400 = n56399 ^ n56398 ;
  assign n56404 = n56251 ^ n56249 ;
  assign n56401 = n54068 ^ n46433 ;
  assign n56402 = n56401 ^ n50347 ;
  assign n56403 = n56402 ^ n45186 ;
  assign n56405 = n56404 ^ n56403 ;
  assign n56407 = n54074 ^ n46438 ;
  assign n56408 = n56407 ^ n50302 ;
  assign n56409 = n56408 ^ n45192 ;
  assign n56406 = n56248 ^ n56247 ;
  assign n56410 = n56409 ^ n56406 ;
  assign n56425 = n54078 ^ n46442 ;
  assign n56426 = n56425 ^ n49807 ;
  assign n56427 = n56426 ^ n45196 ;
  assign n56430 = n56427 ^ n56409 ;
  assign n56423 = n56246 ^ n56245 ;
  assign n56414 = n54583 ^ n46869 ;
  assign n56415 = n56414 ^ n51009 ;
  assign n56416 = n56415 ^ n45412 ;
  assign n56417 = n56146 ^ n53257 ;
  assign n56418 = n56416 & ~n56417 ;
  assign n56411 = n54082 ^ n46446 ;
  assign n56412 = n56411 ^ n49810 ;
  assign n56413 = n56412 ^ n45200 ;
  assign n56419 = n56418 ^ n56413 ;
  assign n56420 = n56418 ^ n56245 ;
  assign n56421 = ~n56419 & n56420 ;
  assign n56422 = n56421 ^ n56245 ;
  assign n56424 = n56423 ^ n56422 ;
  assign n56428 = n56427 ^ n56422 ;
  assign n56429 = n56424 & n56428 ;
  assign n56431 = n56430 ^ n56429 ;
  assign n56432 = n56410 & n56431 ;
  assign n56433 = n56432 ^ n56409 ;
  assign n56434 = n56433 ^ n56403 ;
  assign n56435 = ~n56405 & ~n56434 ;
  assign n56436 = n56435 ^ n56404 ;
  assign n56437 = n56436 ^ n56398 ;
  assign n56438 = n56400 & ~n56437 ;
  assign n56439 = n56438 ^ n56398 ;
  assign n56446 = n56439 ^ n56393 ;
  assign n56395 = n56256 ^ n56254 ;
  assign n56440 = n56439 ^ n56395 ;
  assign n56441 = n54059 ^ n46422 ;
  assign n56442 = n56441 ^ n50909 ;
  assign n56443 = n56442 ^ n45177 ;
  assign n56444 = n56443 ^ n56395 ;
  assign n56445 = ~n56440 & n56444 ;
  assign n56447 = n56446 ^ n56445 ;
  assign n56448 = n56394 & n56447 ;
  assign n56449 = n56448 ^ n56393 ;
  assign n56450 = n56449 ^ n56385 ;
  assign n56451 = ~n56389 & n56450 ;
  assign n56453 = n56452 ^ n56451 ;
  assign n56454 = n56384 & ~n56453 ;
  assign n56455 = n56454 ^ n56383 ;
  assign n56456 = n56455 ^ n56377 ;
  assign n56457 = ~n56379 & ~n56456 ;
  assign n56458 = n56457 ^ n56378 ;
  assign n56459 = n56458 ^ n56372 ;
  assign n56460 = n56374 & n56459 ;
  assign n56461 = n56460 ^ n56373 ;
  assign n56462 = n56461 ^ n56367 ;
  assign n56463 = ~n56369 & ~n56462 ;
  assign n56464 = n56463 ^ n56368 ;
  assign n56465 = n56464 ^ n56360 ;
  assign n56466 = ~n56364 & ~n56465 ;
  assign n56468 = n56467 ^ n56466 ;
  assign n56469 = n56359 & ~n56468 ;
  assign n56470 = n56469 ^ n56358 ;
  assign n56471 = n56470 ^ n56352 ;
  assign n56472 = ~n56354 & ~n56471 ;
  assign n56473 = n56472 ^ n56353 ;
  assign n56474 = n56473 ^ n56345 ;
  assign n56475 = ~n56349 & ~n56474 ;
  assign n56477 = n56476 ^ n56475 ;
  assign n56478 = n56344 & n56477 ;
  assign n56480 = n56479 ^ n56478 ;
  assign n56481 = ~n56339 & ~n56480 ;
  assign n56482 = n56481 ^ n56338 ;
  assign n56483 = n56482 ^ n56330 ;
  assign n56484 = n56334 & n56483 ;
  assign n56486 = n56485 ^ n56484 ;
  assign n56487 = n56329 & n56486 ;
  assign n56489 = n56488 ^ n56487 ;
  assign n56490 = ~n56324 & ~n56489 ;
  assign n56491 = n56490 ^ n56323 ;
  assign n56492 = n56491 ^ n56317 ;
  assign n56493 = n56319 & n56492 ;
  assign n56494 = n56493 ^ n56318 ;
  assign n56495 = n56494 ^ n56312 ;
  assign n56496 = n56314 & ~n56495 ;
  assign n56497 = n56496 ^ n56313 ;
  assign n56293 = ~n56291 & ~n56292 ;
  assign n55659 = n55658 ^ n55655 ;
  assign n56094 = n55659 & ~n56093 ;
  assign n56095 = n56094 ^ n55658 ;
  assign n55653 = n55652 ^ n55637 ;
  assign n55107 = n55106 ^ n55105 ;
  assign n55108 = n55107 ^ n54585 ;
  assign n55654 = n55653 ^ n55108 ;
  assign n56234 = n56095 ^ n55654 ;
  assign n56236 = n56234 ^ n53833 ;
  assign n56113 = n56112 ^ n53576 ;
  assign n56232 = n56113 & n56231 ;
  assign n56233 = n56232 ^ n53576 ;
  assign n56243 = n56236 ^ n56233 ;
  assign n56308 = n56293 ^ n56243 ;
  assign n56304 = n54412 ^ n1221 ;
  assign n56305 = n56304 ^ n1721 ;
  assign n56306 = n56305 ^ n45090 ;
  assign n56309 = n56308 ^ n56306 ;
  assign n57320 = n56497 ^ n56309 ;
  assign n57318 = n56013 ^ n55273 ;
  assign n57319 = n57318 ^ n54596 ;
  assign n57321 = n57320 ^ n57319 ;
  assign n57299 = n56494 ^ n56314 ;
  assign n57297 = n55277 ^ n54548 ;
  assign n57298 = n57297 ^ n56022 ;
  assign n57300 = n57299 ^ n57298 ;
  assign n57278 = n56491 ^ n56319 ;
  assign n57276 = n55279 ^ n54552 ;
  assign n57277 = n57276 ^ n56017 ;
  assign n57279 = n57278 ^ n57277 ;
  assign n57249 = n56489 ^ n56323 ;
  assign n57217 = n56486 ^ n56325 ;
  assign n57250 = n57249 ^ n57217 ;
  assign n57218 = n55287 ^ n54556 ;
  assign n56635 = n55968 ^ n55925 ;
  assign n57219 = n57218 ^ n56635 ;
  assign n57220 = n57219 ^ n57217 ;
  assign n57194 = n56482 ^ n56334 ;
  assign n57166 = n56480 ^ n56338 ;
  assign n57195 = n57194 ^ n57166 ;
  assign n56541 = n55962 ^ n55935 ;
  assign n57167 = n56541 ^ n55209 ;
  assign n57168 = n57167 ^ n55890 ;
  assign n57169 = n57168 ^ n57166 ;
  assign n57142 = n56477 ^ n56340 ;
  assign n56515 = n55960 ^ n55938 ;
  assign n57140 = n56515 ^ n55165 ;
  assign n57141 = n57140 ^ n55105 ;
  assign n57143 = n57142 ^ n57141 ;
  assign n57125 = n56473 ^ n56349 ;
  assign n56105 = n55956 ^ n55945 ;
  assign n57123 = n56105 ^ n55169 ;
  assign n57124 = n57123 ^ n55657 ;
  assign n57126 = n57125 ^ n57124 ;
  assign n57099 = n56470 ^ n56354 ;
  assign n57072 = n56468 ^ n56358 ;
  assign n57100 = n57099 ^ n57072 ;
  assign n57070 = n55666 ^ n55653 ;
  assign n57071 = n57070 ^ n55095 ;
  assign n57073 = n57072 ^ n57071 ;
  assign n57047 = n56464 ^ n56364 ;
  assign n57045 = n55750 ^ n54809 ;
  assign n57046 = n57045 ^ n55655 ;
  assign n57048 = n57047 ^ n57046 ;
  assign n57026 = n56461 ^ n56369 ;
  assign n57024 = n55663 ^ n54795 ;
  assign n57025 = n57024 ^ n55671 ;
  assign n57027 = n57026 ^ n57025 ;
  assign n57005 = n56458 ^ n56374 ;
  assign n57003 = n55678 ^ n55665 ;
  assign n57004 = n57003 ^ n54791 ;
  assign n57006 = n57005 ^ n57004 ;
  assign n56978 = n56455 ^ n56379 ;
  assign n56951 = n56453 ^ n56383 ;
  assign n56979 = n56978 ^ n56951 ;
  assign n56949 = n55689 ^ n55670 ;
  assign n56950 = n56949 ^ n54172 ;
  assign n56952 = n56951 ^ n56950 ;
  assign n56923 = n55681 ^ n54177 ;
  assign n56924 = n56923 ^ n55693 ;
  assign n56903 = n56447 ^ n56392 ;
  assign n56925 = n56924 ^ n56903 ;
  assign n56854 = n56436 ^ n56400 ;
  assign n56852 = n55345 ^ n54195 ;
  assign n56853 = n56852 ^ n55696 ;
  assign n56855 = n56854 ^ n56853 ;
  assign n56874 = n56444 ^ n56439 ;
  assign n56875 = n56874 ^ n56854 ;
  assign n56876 = n56875 ^ n56874 ;
  assign n56829 = n56433 ^ n56405 ;
  assign n56827 = n55700 ^ n55114 ;
  assign n56828 = n56827 ^ n54200 ;
  assign n56830 = n56829 ^ n56828 ;
  assign n56802 = n56431 ^ n56406 ;
  assign n56779 = n56427 ^ n56424 ;
  assign n56803 = n56802 ^ n56779 ;
  assign n56726 = n56417 ^ n56416 ;
  assign n56688 = n54510 ^ n46777 ;
  assign n56689 = n56688 ^ n50798 ;
  assign n56690 = n56689 ^ n45408 ;
  assign n56691 = n56690 ^ n53152 ;
  assign n56638 = n54236 ^ n53300 ;
  assign n56639 = n56638 ^ n55277 ;
  assign n56686 = n56639 ^ n53231 ;
  assign n56684 = n55971 ^ n55920 ;
  assign n56682 = n55273 ^ n54234 ;
  assign n56683 = n56682 ^ n53295 ;
  assign n56685 = n56684 ^ n56683 ;
  assign n56687 = n56686 ^ n56685 ;
  assign n56692 = n56691 ^ n56687 ;
  assign n56649 = n54499 ^ n46781 ;
  assign n56650 = n56649 ^ n50803 ;
  assign n56651 = n56650 ^ n45429 ;
  assign n56693 = n56692 ^ n56651 ;
  assign n56587 = n55966 ^ n55928 ;
  assign n56636 = n56635 ^ n56587 ;
  assign n56585 = n55279 ^ n54596 ;
  assign n56586 = n56585 ^ n53843 ;
  assign n56588 = n56587 ^ n56586 ;
  assign n56539 = n55290 ^ n54548 ;
  assign n56540 = n56539 ^ n53847 ;
  assign n56542 = n56541 ^ n56540 ;
  assign n56513 = n54552 ^ n53851 ;
  assign n56514 = n56513 ^ n55287 ;
  assign n56516 = n56515 ^ n56514 ;
  assign n56102 = n55954 ^ n55949 ;
  assign n56106 = n56105 ^ n56102 ;
  assign n56099 = n55890 ^ n53855 ;
  assign n56100 = n56099 ^ n54556 ;
  assign n56096 = n56095 ^ n55653 ;
  assign n56097 = n55654 & n56096 ;
  assign n56098 = n56097 ^ n55653 ;
  assign n56101 = n56100 ^ n56098 ;
  assign n56103 = n56102 ^ n56098 ;
  assign n56104 = n56101 & n56103 ;
  assign n56107 = n56106 ^ n56104 ;
  assign n55103 = n55102 ^ n53860 ;
  assign n55104 = n55103 ^ n54562 ;
  assign n56510 = n56105 ^ n55104 ;
  assign n56511 = n56107 & ~n56510 ;
  assign n56512 = n56511 ^ n56105 ;
  assign n56543 = n56515 ^ n56512 ;
  assign n56544 = n56516 & n56543 ;
  assign n56545 = n56544 ^ n56515 ;
  assign n56582 = n56545 ^ n56541 ;
  assign n56583 = n56542 & n56582 ;
  assign n56584 = n56583 ^ n56541 ;
  assign n56633 = n56587 ^ n56584 ;
  assign n56634 = n56588 & ~n56633 ;
  assign n56637 = n56636 ^ n56634 ;
  assign n56680 = n56639 ^ n56635 ;
  assign n56681 = n56637 & n56680 ;
  assign n56694 = n56693 ^ n56681 ;
  assign n56110 = n56102 ^ n56101 ;
  assign n56111 = n56110 ^ n53093 ;
  assign n56235 = n56234 ^ n56233 ;
  assign n56237 = ~n56235 & n56236 ;
  assign n56238 = n56237 ^ n53833 ;
  assign n56239 = n56238 ^ n56110 ;
  assign n56240 = ~n56111 & n56239 ;
  assign n56241 = n56240 ^ n53093 ;
  assign n56108 = n56107 ^ n55104 ;
  assign n56109 = n56108 ^ n53096 ;
  assign n56242 = n56241 ^ n56109 ;
  assign n56294 = n56243 & n56293 ;
  assign n56295 = n56238 ^ n56111 ;
  assign n56296 = ~n56294 & n56295 ;
  assign n56509 = ~n56242 & ~n56296 ;
  assign n56519 = n56241 ^ n56108 ;
  assign n56520 = ~n56109 & n56519 ;
  assign n56521 = n56520 ^ n53096 ;
  assign n56517 = n56516 ^ n56512 ;
  assign n56518 = n56517 ^ n53084 ;
  assign n56522 = n56521 ^ n56518 ;
  assign n56537 = ~n56509 & n56522 ;
  assign n56538 = n56521 ^ n56517 ;
  assign n56546 = n56545 ^ n56542 ;
  assign n56547 = n56546 ^ n53084 ;
  assign n56548 = n56547 ^ n56517 ;
  assign n56549 = n56548 ^ n56546 ;
  assign n56550 = ~n56538 & ~n56549 ;
  assign n56551 = n56550 ^ n56547 ;
  assign n56552 = n56551 ^ n53080 ;
  assign n56581 = ~n56537 & n56552 ;
  assign n56589 = n56588 ^ n56584 ;
  assign n56591 = n56589 ^ n53080 ;
  assign n56590 = n56589 ^ n56546 ;
  assign n56592 = n56591 ^ n56590 ;
  assign n56593 = n56551 & ~n56592 ;
  assign n56594 = n56593 ^ n56591 ;
  assign n56595 = n56594 ^ n53129 ;
  assign n56629 = n56581 & n56595 ;
  assign n56640 = n56639 ^ n56637 ;
  assign n56641 = n56640 ^ n53152 ;
  assign n56630 = n56589 ^ n53129 ;
  assign n56631 = n56594 & ~n56630 ;
  assign n56632 = n56631 ^ n53129 ;
  assign n56642 = n56641 ^ n56632 ;
  assign n56679 = ~n56629 & ~n56642 ;
  assign n56695 = n56694 ^ n56679 ;
  assign n56677 = n56640 ^ n56632 ;
  assign n56678 = ~n56641 & ~n56677 ;
  assign n56696 = n56695 ^ n56678 ;
  assign n56523 = n56522 ^ n56509 ;
  assign n56506 = n54400 ^ n46797 ;
  assign n56507 = n56506 ^ n50807 ;
  assign n56508 = n56507 ^ n45294 ;
  assign n56524 = n56523 ^ n56508 ;
  assign n56553 = n56552 ^ n56537 ;
  assign n56554 = n56553 ^ n56508 ;
  assign n56555 = n56554 ^ n56553 ;
  assign n56297 = n56296 ^ n56242 ;
  assign n1401 = n1400 ^ n1334 ;
  assign n1438 = n1437 ^ n1401 ;
  assign n1448 = n1447 ^ n1438 ;
  assign n56298 = n56297 ^ n1448 ;
  assign n56302 = n56295 ^ n56294 ;
  assign n56502 = n56302 ^ n56297 ;
  assign n56299 = n54408 ^ n46803 ;
  assign n56300 = n56299 ^ n50818 ;
  assign n56301 = n56300 ^ n1429 ;
  assign n56303 = n56302 ^ n56301 ;
  assign n56498 = n56497 ^ n56306 ;
  assign n56499 = n56309 & n56498 ;
  assign n56307 = n56306 ^ n56302 ;
  assign n56500 = n56499 ^ n56307 ;
  assign n56501 = n56303 & n56500 ;
  assign n56503 = n56502 ^ n56501 ;
  assign n56504 = n56298 & n56503 ;
  assign n56505 = n56504 ^ n56297 ;
  assign n56556 = n56555 ^ n56505 ;
  assign n56557 = n56524 & n56556 ;
  assign n56558 = n56557 ^ n56554 ;
  assign n56596 = n56595 ^ n56581 ;
  assign n56598 = n56596 ^ n56553 ;
  assign n56559 = n54244 ^ n46792 ;
  assign n56560 = n56559 ^ n50984 ;
  assign n56561 = n56560 ^ n45440 ;
  assign n56597 = n56596 ^ n56561 ;
  assign n56599 = n56598 ^ n56597 ;
  assign n56600 = ~n56558 & ~n56599 ;
  assign n56601 = n56600 ^ n56598 ;
  assign n56643 = n56642 ^ n56629 ;
  assign n56645 = n56643 ^ n56596 ;
  assign n56602 = n54502 ^ n46786 ;
  assign n56603 = n56602 ^ n50992 ;
  assign n56604 = n56603 ^ n45434 ;
  assign n56644 = n56643 ^ n56604 ;
  assign n56646 = n56645 ^ n56644 ;
  assign n56647 = ~n56601 & n56646 ;
  assign n56648 = n56647 ^ n56645 ;
  assign n56675 = n56651 ^ n56643 ;
  assign n56676 = n56648 & ~n56675 ;
  assign n56697 = n56696 ^ n56676 ;
  assign n56727 = n56726 ^ n56697 ;
  assign n56701 = n55720 ^ n55134 ;
  assign n56702 = n56701 ^ n54214 ;
  assign n56652 = n56651 ^ n56648 ;
  assign n56605 = n56604 ^ n56601 ;
  assign n56653 = n56652 ^ n56605 ;
  assign n56525 = n56524 ^ n56505 ;
  assign n56526 = n55735 ^ n55145 ;
  assign n56527 = n56526 ^ n54229 ;
  assign n56565 = n56525 & ~n56527 ;
  assign n56563 = n55141 ^ n54220 ;
  assign n56564 = n56563 ^ n55731 ;
  assign n56566 = n56565 ^ n56564 ;
  assign n56606 = n56605 ^ n56564 ;
  assign n56607 = n56606 ^ n56605 ;
  assign n56562 = n56561 ^ n56558 ;
  assign n56608 = n56607 ^ n56562 ;
  assign n56609 = n56566 & ~n56608 ;
  assign n56610 = n56609 ^ n56606 ;
  assign n56611 = n55728 ^ n54616 ;
  assign n56612 = n56611 ^ n55139 ;
  assign n56627 = n56612 ^ n56605 ;
  assign n56628 = ~n56610 & ~n56627 ;
  assign n56654 = n56653 ^ n56628 ;
  assign n56655 = n55132 ^ n54218 ;
  assign n56656 = n56655 ^ n55722 ;
  assign n56698 = n56656 ^ n56652 ;
  assign n56699 = ~n56654 & n56698 ;
  assign n56700 = n56699 ^ n56656 ;
  assign n56703 = n56702 ^ n56700 ;
  assign n56724 = n56700 ^ n56697 ;
  assign n56725 = ~n56703 & ~n56724 ;
  assign n56728 = n56727 ^ n56725 ;
  assign n56729 = n55716 ^ n55321 ;
  assign n56730 = n56729 ^ n54210 ;
  assign n56758 = n56730 ^ n56726 ;
  assign n56759 = ~n56728 & n56758 ;
  assign n56755 = n56413 ^ n56245 ;
  assign n56756 = n56755 ^ n56418 ;
  assign n56757 = n56756 ^ n56726 ;
  assign n56760 = n56759 ^ n56757 ;
  assign n56780 = n56779 ^ n56756 ;
  assign n56781 = n56780 ^ n56779 ;
  assign n56753 = n55712 ^ n54205 ;
  assign n56754 = n56753 ^ n55128 ;
  assign n56782 = n56781 ^ n56754 ;
  assign n56783 = ~n56760 & ~n56782 ;
  assign n56784 = n56783 ^ n56780 ;
  assign n56785 = n55122 ^ n54631 ;
  assign n56786 = n56785 ^ n55708 ;
  assign n56800 = n56786 ^ n56779 ;
  assign n56801 = ~n56784 & ~n56800 ;
  assign n56804 = n56803 ^ n56801 ;
  assign n56805 = n55704 ^ n54638 ;
  assign n56806 = n56805 ^ n55118 ;
  assign n56824 = n56806 ^ n56802 ;
  assign n56825 = n56804 & ~n56824 ;
  assign n56826 = n56825 ^ n56806 ;
  assign n56849 = n56828 ^ n56826 ;
  assign n56850 = n56830 & ~n56849 ;
  assign n56851 = n56850 ^ n56829 ;
  assign n56877 = n56876 ^ n56851 ;
  assign n56878 = ~n56855 & n56877 ;
  assign n56879 = n56878 ^ n56875 ;
  assign n56905 = n56903 ^ n56874 ;
  assign n56880 = n55688 ^ n55445 ;
  assign n56881 = n56880 ^ n54190 ;
  assign n56904 = n56903 ^ n56881 ;
  assign n56906 = n56905 ^ n56904 ;
  assign n56907 = n56879 & ~n56906 ;
  assign n56908 = n56907 ^ n56905 ;
  assign n56909 = n55686 ^ n55646 ;
  assign n56910 = n56909 ^ n54182 ;
  assign n56921 = n56910 ^ n56903 ;
  assign n56922 = ~n56908 & ~n56921 ;
  assign n56926 = n56925 ^ n56922 ;
  assign n56927 = n56449 ^ n56389 ;
  assign n56946 = n56927 ^ n56924 ;
  assign n56947 = n56926 & n56946 ;
  assign n56948 = n56947 ^ n56927 ;
  assign n56976 = n56951 ^ n56948 ;
  assign n56977 = ~n56952 & ~n56976 ;
  assign n56980 = n56979 ^ n56977 ;
  assign n56981 = n55683 ^ n55675 ;
  assign n56982 = n56981 ^ n54667 ;
  assign n57000 = n56982 ^ n56978 ;
  assign n57001 = n56980 & n57000 ;
  assign n57002 = n57001 ^ n56982 ;
  assign n57021 = n57004 ^ n57002 ;
  assign n57022 = n57006 & ~n57021 ;
  assign n57023 = n57022 ^ n57005 ;
  assign n57042 = n57025 ^ n57023 ;
  assign n57043 = ~n57027 & n57042 ;
  assign n57044 = n57043 ^ n57026 ;
  assign n57067 = n57046 ^ n57044 ;
  assign n57068 = n57048 & n57067 ;
  assign n57069 = n57068 ^ n57047 ;
  assign n57097 = n57072 ^ n57069 ;
  assign n57098 = n57073 & n57097 ;
  assign n57101 = n57100 ^ n57098 ;
  assign n57102 = n56102 ^ n55173 ;
  assign n57103 = n57102 ^ n55661 ;
  assign n57120 = n57103 ^ n57099 ;
  assign n57121 = n57101 & ~n57120 ;
  assign n57122 = n57121 ^ n57103 ;
  assign n57137 = n57124 ^ n57122 ;
  assign n57138 = n57126 & ~n57137 ;
  assign n57139 = n57138 ^ n57125 ;
  assign n57163 = n57141 ^ n57139 ;
  assign n57164 = ~n57143 & n57163 ;
  assign n57165 = n57164 ^ n57142 ;
  assign n57192 = n57166 ^ n57165 ;
  assign n57193 = ~n57169 & ~n57192 ;
  assign n57196 = n57195 ^ n57193 ;
  assign n57197 = n56587 ^ n55106 ;
  assign n57198 = n57197 ^ n55102 ;
  assign n57214 = n57198 ^ n57194 ;
  assign n57215 = ~n57196 & n57214 ;
  assign n57216 = n57215 ^ n57198 ;
  assign n57247 = n57217 ^ n57216 ;
  assign n57248 = ~n57220 & ~n57247 ;
  assign n57251 = n57250 ^ n57248 ;
  assign n57252 = n56684 ^ n54562 ;
  assign n57253 = n57252 ^ n55290 ;
  assign n57273 = n57253 ^ n57249 ;
  assign n57274 = n57251 & n57273 ;
  assign n57275 = n57274 ^ n57253 ;
  assign n57294 = n57277 ^ n57275 ;
  assign n57295 = n57279 & ~n57294 ;
  assign n57296 = n57295 ^ n57278 ;
  assign n57315 = n57298 ^ n57296 ;
  assign n57316 = n57300 & n57315 ;
  assign n57317 = n57316 ^ n57299 ;
  assign n57322 = n57321 ^ n57317 ;
  assign n57323 = n57322 ^ n53843 ;
  assign n57301 = n57300 ^ n57296 ;
  assign n57302 = n57301 ^ n53847 ;
  assign n57280 = n57279 ^ n57275 ;
  assign n57281 = n57280 ^ n53851 ;
  assign n57254 = n57253 ^ n57251 ;
  assign n57255 = n57254 ^ n53860 ;
  assign n57127 = n57126 ^ n57122 ;
  assign n57128 = n57127 ^ n54484 ;
  assign n57104 = n57103 ^ n57101 ;
  assign n57105 = n57104 ^ n54315 ;
  assign n57074 = n57073 ^ n57069 ;
  assign n57075 = n57074 ^ n54174 ;
  assign n57049 = n57048 ^ n57044 ;
  assign n57050 = n57049 ^ n54179 ;
  assign n57028 = n57027 ^ n57023 ;
  assign n57029 = n57028 ^ n54183 ;
  assign n57007 = n57006 ^ n57002 ;
  assign n57008 = n57007 ^ n54187 ;
  assign n56983 = n56982 ^ n56980 ;
  assign n56984 = n56983 ^ n54192 ;
  assign n56953 = n56952 ^ n56948 ;
  assign n56954 = n56953 ^ n54197 ;
  assign n56928 = n56927 ^ n56926 ;
  assign n56929 = n56928 ^ n54264 ;
  assign n56882 = n56881 ^ n56879 ;
  assign n56883 = n56882 ^ n54202 ;
  assign n56787 = n56786 ^ n56784 ;
  assign n56788 = n56787 ^ n54006 ;
  assign n56704 = n56703 ^ n56697 ;
  assign n56613 = n56612 ^ n56610 ;
  assign n56614 = n56613 ^ n53279 ;
  assign n56528 = n56527 ^ n56525 ;
  assign n56568 = n53286 & ~n56528 ;
  assign n56569 = n56568 ^ n53284 ;
  assign n56567 = n56566 ^ n56562 ;
  assign n56615 = n56568 ^ n56567 ;
  assign n56616 = ~n56569 & n56615 ;
  assign n56617 = n56616 ^ n53284 ;
  assign n56623 = n56617 ^ n56613 ;
  assign n56624 = ~n56614 & ~n56623 ;
  assign n56625 = n56624 ^ n53279 ;
  assign n56626 = n56625 ^ n53271 ;
  assign n56657 = n56656 ^ n56654 ;
  assign n56671 = n56657 ^ n56625 ;
  assign n56672 = n56626 & n56671 ;
  assign n56673 = n56672 ^ n53271 ;
  assign n56723 = n56704 ^ n56673 ;
  assign n56731 = n56730 ^ n56728 ;
  assign n56732 = n56731 ^ n53239 ;
  assign n56733 = n56732 ^ n56731 ;
  assign n56734 = n56733 ^ n56704 ;
  assign n56735 = ~n56723 & n56734 ;
  assign n56736 = n56735 ^ n56732 ;
  assign n56749 = n56731 ^ n53268 ;
  assign n56750 = ~n56736 & n56749 ;
  assign n56751 = n56750 ^ n53268 ;
  assign n56752 = n56751 ^ n53967 ;
  assign n56761 = n56760 ^ n56754 ;
  assign n56776 = n56761 ^ n56751 ;
  assign n56777 = n56752 & ~n56776 ;
  assign n56778 = n56777 ^ n53967 ;
  assign n56808 = n56787 ^ n56778 ;
  assign n56809 = n56788 & n56808 ;
  assign n56810 = n56809 ^ n54006 ;
  assign n56811 = n56810 ^ n54141 ;
  assign n56807 = n56806 ^ n56804 ;
  assign n56833 = n56810 ^ n56807 ;
  assign n56834 = ~n56811 & n56833 ;
  assign n56835 = n56834 ^ n54141 ;
  assign n56831 = n56830 ^ n56826 ;
  assign n56848 = n56835 ^ n56831 ;
  assign n56856 = n56855 ^ n56851 ;
  assign n56857 = n56856 ^ n54164 ;
  assign n56858 = n56857 ^ n56856 ;
  assign n56859 = n56858 ^ n56831 ;
  assign n56860 = n56848 & n56859 ;
  assign n56861 = n56860 ^ n56857 ;
  assign n56884 = n56856 ^ n54208 ;
  assign n56885 = n56861 & n56884 ;
  assign n56886 = n56885 ^ n54208 ;
  assign n56899 = n56886 ^ n56882 ;
  assign n56900 = n56883 & ~n56899 ;
  assign n56901 = n56900 ^ n54202 ;
  assign n56902 = n56901 ^ n54268 ;
  assign n56911 = n56910 ^ n56908 ;
  assign n56918 = n56911 ^ n56901 ;
  assign n56919 = ~n56902 & ~n56918 ;
  assign n56920 = n56919 ^ n54268 ;
  assign n56955 = n56928 ^ n56920 ;
  assign n56956 = ~n56929 & n56955 ;
  assign n56957 = n56956 ^ n54264 ;
  assign n56973 = n56957 ^ n56953 ;
  assign n56974 = ~n56954 & n56973 ;
  assign n56975 = n56974 ^ n54197 ;
  assign n56997 = n56983 ^ n56975 ;
  assign n56998 = n56984 & n56997 ;
  assign n56999 = n56998 ^ n54192 ;
  assign n57030 = n57007 ^ n56999 ;
  assign n57031 = n57008 & n57030 ;
  assign n57032 = n57031 ^ n54187 ;
  assign n57039 = n57032 ^ n57028 ;
  assign n57040 = n57029 & n57039 ;
  assign n57041 = n57040 ^ n54183 ;
  assign n57076 = n57049 ^ n57041 ;
  assign n57077 = ~n57050 & n57076 ;
  assign n57078 = n57077 ^ n54179 ;
  assign n57094 = n57078 ^ n57074 ;
  assign n57095 = ~n57075 & ~n57094 ;
  assign n57096 = n57095 ^ n54174 ;
  assign n57129 = n57104 ^ n57096 ;
  assign n57130 = n57105 & ~n57129 ;
  assign n57131 = n57130 ^ n54315 ;
  assign n57146 = n57131 ^ n57127 ;
  assign n57147 = n57128 & n57146 ;
  assign n57148 = n57147 ^ n54484 ;
  assign n57144 = n57143 ^ n57139 ;
  assign n57162 = n57148 ^ n57144 ;
  assign n57170 = n57169 ^ n57165 ;
  assign n57171 = n57170 ^ n54524 ;
  assign n57172 = n57171 ^ n57170 ;
  assign n57173 = n57172 ^ n57144 ;
  assign n57174 = n57162 & n57173 ;
  assign n57175 = n57174 ^ n57171 ;
  assign n57201 = n57170 ^ n54533 ;
  assign n57202 = ~n57175 & n57201 ;
  assign n57203 = n57202 ^ n54533 ;
  assign n57199 = n57198 ^ n57196 ;
  assign n57213 = n57203 ^ n57199 ;
  assign n57221 = n57220 ^ n57216 ;
  assign n57222 = n57221 ^ n54585 ;
  assign n57223 = n57222 ^ n57221 ;
  assign n57224 = n57223 ^ n57199 ;
  assign n57225 = ~n57213 & n57224 ;
  assign n57226 = n57225 ^ n57222 ;
  assign n57256 = n57221 ^ n53855 ;
  assign n57257 = n57226 & ~n57256 ;
  assign n57258 = n57257 ^ n53855 ;
  assign n57270 = n57258 ^ n57254 ;
  assign n57271 = n57255 & n57270 ;
  assign n57272 = n57271 ^ n53860 ;
  assign n57303 = n57280 ^ n57272 ;
  assign n57304 = n57281 & n57303 ;
  assign n57305 = n57304 ^ n53851 ;
  assign n57312 = n57305 ^ n57301 ;
  assign n57313 = n57302 & ~n57312 ;
  assign n57314 = n57313 ^ n53847 ;
  assign n57354 = n57322 ^ n57314 ;
  assign n57355 = n57323 & ~n57354 ;
  assign n57356 = n57355 ^ n53843 ;
  assign n57350 = n56500 ^ n56301 ;
  assign n57348 = n56009 ^ n54236 ;
  assign n57349 = n57348 ^ n55156 ;
  assign n57351 = n57350 ^ n57349 ;
  assign n57345 = n57319 ^ n57317 ;
  assign n57346 = ~n57321 & n57345 ;
  assign n57347 = n57346 ^ n57320 ;
  assign n57352 = n57351 ^ n57347 ;
  assign n57378 = n57356 ^ n57352 ;
  assign n57324 = n57323 ^ n57314 ;
  assign n57306 = n57305 ^ n57302 ;
  assign n57282 = n57281 ^ n57272 ;
  assign n57259 = n57258 ^ n57255 ;
  assign n57227 = n57226 ^ n53855 ;
  assign n57200 = n57199 ^ n54585 ;
  assign n57204 = n57203 ^ n57200 ;
  assign n57176 = n57175 ^ n54533 ;
  assign n57145 = n57144 ^ n54524 ;
  assign n57149 = n57148 ^ n57145 ;
  assign n57132 = n57131 ^ n57128 ;
  assign n57106 = n57105 ^ n57096 ;
  assign n57079 = n57078 ^ n57075 ;
  assign n57051 = n57050 ^ n57041 ;
  assign n57033 = n57032 ^ n57029 ;
  assign n57009 = n57008 ^ n56999 ;
  assign n56985 = n56984 ^ n56975 ;
  assign n56958 = n56957 ^ n56954 ;
  assign n56930 = n56929 ^ n56920 ;
  assign n56912 = n56911 ^ n56902 ;
  assign n56887 = n56886 ^ n56883 ;
  assign n56862 = n56861 ^ n54208 ;
  assign n56832 = n56831 ^ n54164 ;
  assign n56836 = n56835 ^ n56832 ;
  assign n56812 = n56811 ^ n56807 ;
  assign n56789 = n56788 ^ n56778 ;
  assign n56762 = n56761 ^ n56752 ;
  assign n56737 = n56736 ^ n53268 ;
  assign n56674 = n56673 ^ n53239 ;
  assign n56705 = n56704 ^ n56674 ;
  assign n56658 = n56657 ^ n56626 ;
  assign n56570 = n56569 ^ n56567 ;
  assign n56618 = n56617 ^ n56614 ;
  assign n56659 = ~n56570 & ~n56618 ;
  assign n56706 = ~n56658 & ~n56659 ;
  assign n56738 = ~n56705 & ~n56706 ;
  assign n56763 = n56737 & ~n56738 ;
  assign n56790 = ~n56762 & ~n56763 ;
  assign n56813 = ~n56789 & n56790 ;
  assign n56837 = n56812 & n56813 ;
  assign n56863 = n56836 & ~n56837 ;
  assign n56888 = ~n56862 & n56863 ;
  assign n56913 = n56887 & n56888 ;
  assign n56931 = ~n56912 & n56913 ;
  assign n56959 = n56930 & n56931 ;
  assign n56986 = ~n56958 & ~n56959 ;
  assign n57010 = n56985 & n56986 ;
  assign n57034 = n57009 & ~n57010 ;
  assign n57052 = n57033 & ~n57034 ;
  assign n57080 = ~n57051 & ~n57052 ;
  assign n57107 = ~n57079 & n57080 ;
  assign n57133 = ~n57106 & n57107 ;
  assign n57150 = n57132 & ~n57133 ;
  assign n57177 = ~n57149 & n57150 ;
  assign n57205 = ~n57176 & ~n57177 ;
  assign n57228 = ~n57204 & n57205 ;
  assign n57260 = ~n57227 & ~n57228 ;
  assign n57283 = ~n57259 & ~n57260 ;
  assign n57307 = ~n57282 & ~n57283 ;
  assign n57325 = ~n57306 & ~n57307 ;
  assign n57358 = ~n57324 & n57325 ;
  assign n57381 = n57378 ^ n57358 ;
  assign n57382 = ~n53300 & n57381 ;
  assign n57379 = n57358 ^ n57352 ;
  assign n57380 = ~n57378 & n57379 ;
  assign n57383 = n57382 ^ n57380 ;
  assign n57375 = n53300 ^ n53295 ;
  assign n57372 = n56503 ^ n1448 ;
  assign n57370 = n56003 ^ n55152 ;
  assign n57371 = n57370 ^ n54234 ;
  assign n57373 = n57372 ^ n57371 ;
  assign n57374 = n57373 ^ n57349 ;
  assign n57376 = n57375 ^ n57374 ;
  assign n57368 = n57349 ^ n57347 ;
  assign n57369 = ~n57351 & ~n57368 ;
  assign n57377 = n57376 ^ n57369 ;
  assign n57384 = n57383 ^ n57377 ;
  assign n57365 = n55162 ^ n47501 ;
  assign n57366 = n57365 ^ n51587 ;
  assign n57367 = n57366 ^ n46091 ;
  assign n57385 = n57384 ^ n57367 ;
  assign n57340 = n55228 ^ n47456 ;
  assign n57341 = n57340 ^ n51592 ;
  assign n57342 = n57341 ^ n46095 ;
  assign n57308 = n57307 ^ n57306 ;
  assign n57291 = n55237 ^ n47397 ;
  assign n57292 = n57291 ^ n51601 ;
  assign n57293 = n57292 ^ n46105 ;
  assign n57309 = n57308 ^ n57293 ;
  assign n57326 = n57325 ^ n57324 ;
  assign n57327 = n57326 ^ n57293 ;
  assign n57328 = n57327 ^ n57326 ;
  assign n57284 = n57283 ^ n57282 ;
  assign n57267 = n55085 ^ n44026 ;
  assign n57268 = n57267 ^ n51606 ;
  assign n57269 = n57268 ^ n46110 ;
  assign n57285 = n57284 ^ n57269 ;
  assign n57233 = n54884 ^ n47182 ;
  assign n57234 = n57233 ^ n51616 ;
  assign n57235 = n57234 ^ n45940 ;
  assign n57206 = n57205 ^ n57204 ;
  assign n57189 = n54890 ^ n1740 ;
  assign n57190 = n57189 ^ n51621 ;
  assign n57191 = n57190 ^ n45301 ;
  assign n57207 = n57206 ^ n57191 ;
  assign n57108 = n57107 ^ n57106 ;
  assign n57091 = n54910 ^ n47205 ;
  assign n57092 = n57091 ^ n51641 ;
  assign n57093 = n57092 ^ n45760 ;
  assign n57109 = n57108 ^ n57093 ;
  assign n57112 = n54904 ^ n47201 ;
  assign n57113 = n57112 ^ n51636 ;
  assign n57114 = n57113 ^ n45755 ;
  assign n57115 = n57114 ^ n57108 ;
  assign n57116 = n57115 ^ n57114 ;
  assign n57081 = n57080 ^ n57079 ;
  assign n57064 = n54917 ^ n47210 ;
  assign n57065 = n57064 ^ n51646 ;
  assign n57066 = n57065 ^ n45766 ;
  assign n57082 = n57081 ^ n57066 ;
  assign n57035 = n57034 ^ n57033 ;
  assign n57018 = n54927 ^ n45775 ;
  assign n57019 = n57018 ^ n51656 ;
  assign n57020 = n57019 ^ n47222 ;
  assign n57036 = n57035 ^ n57020 ;
  assign n57053 = n57052 ^ n57051 ;
  assign n57054 = n57053 ^ n57020 ;
  assign n57055 = n57054 ^ n57053 ;
  assign n57011 = n57010 ^ n57009 ;
  assign n56994 = n54932 ^ n47228 ;
  assign n56995 = n56994 ^ n51661 ;
  assign n56996 = n56995 ^ n45780 ;
  assign n57012 = n57011 ^ n56996 ;
  assign n56987 = n56986 ^ n56985 ;
  assign n56970 = n54938 ^ n47233 ;
  assign n56971 = n56970 ^ n51666 ;
  assign n56972 = n56971 ^ n45787 ;
  assign n56988 = n56987 ^ n56972 ;
  assign n56960 = n56959 ^ n56958 ;
  assign n56943 = n54943 ^ n47238 ;
  assign n56944 = n56943 ^ n51298 ;
  assign n56945 = n56944 ^ n45791 ;
  assign n56961 = n56960 ^ n56945 ;
  assign n56914 = n56913 ^ n56912 ;
  assign n56896 = n54953 ^ n47247 ;
  assign n56897 = n56896 ^ n2441 ;
  assign n56898 = n56897 ^ n45801 ;
  assign n56915 = n56914 ^ n56898 ;
  assign n56932 = n56931 ^ n56930 ;
  assign n56933 = n56932 ^ n56898 ;
  assign n56934 = n56933 ^ n56932 ;
  assign n56889 = n56888 ^ n56887 ;
  assign n56871 = n54958 ^ n47253 ;
  assign n56872 = n56871 ^ n51165 ;
  assign n56873 = n56872 ^ n2430 ;
  assign n56890 = n56889 ^ n56873 ;
  assign n56864 = n56863 ^ n56862 ;
  assign n56845 = n54963 ^ n2279 ;
  assign n56846 = n56845 ^ n51171 ;
  assign n56847 = n56846 ^ n45809 ;
  assign n56865 = n56864 ^ n56847 ;
  assign n56838 = n56837 ^ n56836 ;
  assign n56821 = n54969 ^ n47261 ;
  assign n56822 = n56821 ^ n51176 ;
  assign n56823 = n56822 ^ n45813 ;
  assign n56839 = n56838 ^ n56823 ;
  assign n56814 = n56813 ^ n56812 ;
  assign n56797 = n54973 ^ n47265 ;
  assign n56798 = n56797 ^ n51181 ;
  assign n56799 = n56798 ^ n45819 ;
  assign n56815 = n56814 ^ n56799 ;
  assign n56764 = n56763 ^ n56762 ;
  assign n56746 = n54984 ^ n51187 ;
  assign n56747 = n56746 ^ n47276 ;
  assign n56748 = n56747 ^ n45828 ;
  assign n56765 = n56764 ^ n56748 ;
  assign n56768 = n54980 ^ n47271 ;
  assign n56769 = n56768 ^ n51192 ;
  assign n56770 = n56769 ^ n45824 ;
  assign n56771 = n56770 ^ n56764 ;
  assign n56739 = n56738 ^ n56737 ;
  assign n56720 = n55016 ^ n47281 ;
  assign n56721 = n56720 ^ n51197 ;
  assign n56722 = n56721 ^ n45833 ;
  assign n56740 = n56739 ^ n56722 ;
  assign n56619 = n56618 ^ n56570 ;
  assign n56578 = n54999 ^ n47300 ;
  assign n56579 = n56578 ^ n51214 ;
  assign n56580 = n56579 ^ n45848 ;
  assign n56620 = n56619 ^ n56580 ;
  assign n56660 = n56659 ^ n56658 ;
  assign n56661 = n56660 ^ n56580 ;
  assign n56534 = n55002 ^ n47296 ;
  assign n56535 = n56534 ^ n51218 ;
  assign n56536 = n56535 ^ n45852 ;
  assign n56571 = n56570 ^ n56536 ;
  assign n56529 = n56528 ^ n53286 ;
  assign n56530 = n55263 ^ n47535 ;
  assign n56531 = n56530 ^ n51737 ;
  assign n56532 = n56531 ^ n46154 ;
  assign n56572 = ~n56529 & n56532 ;
  assign n56575 = n56572 ^ n56570 ;
  assign n56576 = ~n56571 & ~n56575 ;
  assign n56577 = n56576 ^ n56570 ;
  assign n56662 = n56661 ^ n56577 ;
  assign n56663 = n56662 ^ n56660 ;
  assign n56664 = ~n56620 & ~n56663 ;
  assign n56665 = n56664 ^ n56661 ;
  assign n56666 = n54995 ^ n47290 ;
  assign n56667 = n56666 ^ n51207 ;
  assign n56668 = n56667 ^ n45844 ;
  assign n56711 = n56668 ^ n56660 ;
  assign n56712 = n56665 & n56711 ;
  assign n56713 = n56712 ^ n56660 ;
  assign n56708 = n54990 ^ n47285 ;
  assign n56709 = n56708 ^ n51203 ;
  assign n56710 = n56709 ^ n45838 ;
  assign n56714 = n56713 ^ n56710 ;
  assign n56707 = n56706 ^ n56705 ;
  assign n56717 = n56713 ^ n56707 ;
  assign n56718 = n56714 & ~n56717 ;
  assign n56719 = n56718 ^ n56713 ;
  assign n56743 = n56722 ^ n56719 ;
  assign n56744 = ~n56740 & n56743 ;
  assign n56745 = n56744 ^ n56722 ;
  assign n56772 = n56771 ^ n56745 ;
  assign n56773 = n56772 ^ n56770 ;
  assign n56774 = ~n56765 & ~n56773 ;
  assign n56775 = n56774 ^ n56771 ;
  assign n56791 = n56790 ^ n56789 ;
  assign n56794 = n56791 ^ n56770 ;
  assign n56795 = ~n56775 & n56794 ;
  assign n56796 = n56795 ^ n56770 ;
  assign n56818 = n56799 ^ n56796 ;
  assign n56819 = ~n56815 & n56818 ;
  assign n56820 = n56819 ^ n56799 ;
  assign n56842 = n56823 ^ n56820 ;
  assign n56843 = ~n56839 & ~n56842 ;
  assign n56844 = n56843 ^ n56838 ;
  assign n56868 = n56847 ^ n56844 ;
  assign n56869 = ~n56865 & n56868 ;
  assign n56870 = n56869 ^ n56864 ;
  assign n56893 = n56873 ^ n56870 ;
  assign n56894 = n56890 & n56893 ;
  assign n56895 = n56894 ^ n56889 ;
  assign n56935 = n56934 ^ n56895 ;
  assign n56936 = ~n56915 & n56935 ;
  assign n56937 = n56936 ^ n56933 ;
  assign n56938 = n54948 ^ n47243 ;
  assign n56939 = n56938 ^ n51255 ;
  assign n56940 = n56939 ^ n45796 ;
  assign n56962 = n56940 ^ n56932 ;
  assign n56963 = n56937 & n56962 ;
  assign n56964 = n56963 ^ n56932 ;
  assign n56967 = n56964 ^ n56945 ;
  assign n56968 = n56961 & n56967 ;
  assign n56969 = n56968 ^ n56964 ;
  assign n56991 = n56972 ^ n56969 ;
  assign n56992 = ~n56988 & n56991 ;
  assign n56993 = n56992 ^ n56972 ;
  assign n57015 = n56996 ^ n56993 ;
  assign n57016 = ~n57012 & n57015 ;
  assign n57017 = n57016 ^ n56996 ;
  assign n57056 = n57055 ^ n57017 ;
  assign n57057 = n57036 & n57056 ;
  assign n57058 = n57057 ^ n57054 ;
  assign n57059 = n54923 ^ n47216 ;
  assign n57060 = n57059 ^ n51651 ;
  assign n57061 = n57060 ^ n45771 ;
  assign n57083 = n57061 ^ n57053 ;
  assign n57084 = n57058 & n57083 ;
  assign n57085 = n57084 ^ n57053 ;
  assign n57088 = n57085 ^ n57066 ;
  assign n57089 = n57082 & n57088 ;
  assign n57090 = n57089 ^ n57085 ;
  assign n57117 = n57116 ^ n57090 ;
  assign n57118 = ~n57109 & ~n57117 ;
  assign n57119 = n57118 ^ n57115 ;
  assign n57151 = n57150 ^ n57149 ;
  assign n57153 = n57151 ^ n57114 ;
  assign n57134 = n57133 ^ n57132 ;
  assign n57152 = n57151 ^ n57134 ;
  assign n57154 = n57153 ^ n57152 ;
  assign n57155 = ~n57119 & n57154 ;
  assign n57156 = n57155 ^ n57153 ;
  assign n57178 = n57177 ^ n57176 ;
  assign n57180 = n57178 ^ n57151 ;
  assign n57157 = n54900 ^ n47195 ;
  assign n57158 = n57157 ^ n51632 ;
  assign n57159 = n57158 ^ n965 ;
  assign n57179 = n57178 ^ n57159 ;
  assign n57181 = n57180 ^ n57179 ;
  assign n57182 = n57156 & n57181 ;
  assign n57183 = n57182 ^ n57180 ;
  assign n57184 = n54894 ^ n47190 ;
  assign n57185 = n57184 ^ n51626 ;
  assign n57186 = n57185 ^ n45747 ;
  assign n57208 = n57186 ^ n57178 ;
  assign n57209 = n57183 & n57208 ;
  assign n57210 = n57209 ^ n57178 ;
  assign n57230 = n57210 ^ n57191 ;
  assign n57231 = n57207 & n57230 ;
  assign n57232 = n57231 ^ n57210 ;
  assign n57236 = n57235 ^ n57232 ;
  assign n57239 = n47177 ^ n1775 ;
  assign n57240 = n57239 ^ n51611 ;
  assign n57241 = n57240 ^ n46116 ;
  assign n57229 = n57228 ^ n57227 ;
  assign n57242 = n57241 ^ n57229 ;
  assign n57243 = n57242 ^ n57241 ;
  assign n57244 = n57243 ^ n57232 ;
  assign n57245 = ~n57236 & ~n57244 ;
  assign n57246 = n57245 ^ n57242 ;
  assign n57261 = n57260 ^ n57259 ;
  assign n57264 = n57261 ^ n57241 ;
  assign n57265 = ~n57246 & n57264 ;
  assign n57266 = n57265 ^ n57241 ;
  assign n57288 = n57284 ^ n57266 ;
  assign n57289 = ~n57285 & ~n57288 ;
  assign n57290 = n57289 ^ n57284 ;
  assign n57329 = n57328 ^ n57290 ;
  assign n57330 = n57309 & ~n57329 ;
  assign n57331 = n57330 ^ n57327 ;
  assign n57332 = n55232 ^ n47410 ;
  assign n57333 = n57332 ^ n51596 ;
  assign n57334 = n57333 ^ n46101 ;
  assign n57337 = n57334 ^ n57326 ;
  assign n57338 = ~n57331 & ~n57337 ;
  assign n57339 = n57338 ^ n57326 ;
  assign n57343 = n57342 ^ n57339 ;
  assign n57353 = n57352 ^ n53300 ;
  assign n57357 = n57356 ^ n57353 ;
  assign n57359 = n57358 ^ n57357 ;
  assign n57360 = n57359 ^ n57339 ;
  assign n57363 = n57343 & n57360 ;
  assign n56533 = n56532 ^ n56529 ;
  assign n56573 = n56572 ^ n56571 ;
  assign n56574 = ~n56533 & ~n56573 ;
  assign n56621 = n56620 ^ n56577 ;
  assign n56622 = n56574 & n56621 ;
  assign n56669 = n56668 ^ n56665 ;
  assign n56670 = n56622 & n56669 ;
  assign n56715 = n56714 ^ n56707 ;
  assign n56716 = n56670 & ~n56715 ;
  assign n56741 = n56740 ^ n56719 ;
  assign n56742 = n56716 & ~n56741 ;
  assign n56766 = n56765 ^ n56745 ;
  assign n56767 = n56742 & ~n56766 ;
  assign n56792 = n56791 ^ n56775 ;
  assign n56793 = n56767 & ~n56792 ;
  assign n56816 = n56815 ^ n56796 ;
  assign n56817 = ~n56793 & n56816 ;
  assign n56840 = n56839 ^ n56820 ;
  assign n56841 = n56817 & n56840 ;
  assign n56866 = n56865 ^ n56844 ;
  assign n56867 = ~n56841 & n56866 ;
  assign n56891 = n56890 ^ n56870 ;
  assign n56892 = n56867 & ~n56891 ;
  assign n56916 = n56915 ^ n56895 ;
  assign n56917 = n56892 & ~n56916 ;
  assign n56941 = n56940 ^ n56937 ;
  assign n56942 = ~n56917 & ~n56941 ;
  assign n56965 = n56964 ^ n56961 ;
  assign n56966 = ~n56942 & ~n56965 ;
  assign n56989 = n56988 ^ n56969 ;
  assign n56990 = n56966 & ~n56989 ;
  assign n57013 = n57012 ^ n56993 ;
  assign n57014 = ~n56990 & n57013 ;
  assign n57037 = n57036 ^ n57017 ;
  assign n57038 = ~n57014 & n57037 ;
  assign n57062 = n57061 ^ n57058 ;
  assign n57063 = ~n57038 & ~n57062 ;
  assign n57086 = n57085 ^ n57082 ;
  assign n57087 = ~n57063 & ~n57086 ;
  assign n57110 = n57109 ^ n57090 ;
  assign n57111 = n57087 & ~n57110 ;
  assign n57135 = n57134 ^ n57119 ;
  assign n57136 = n57111 & ~n57135 ;
  assign n57160 = n57159 ^ n57156 ;
  assign n57161 = ~n57136 & ~n57160 ;
  assign n57187 = n57186 ^ n57183 ;
  assign n57188 = ~n57161 & n57187 ;
  assign n57211 = n57210 ^ n57207 ;
  assign n57212 = ~n57188 & n57211 ;
  assign n57237 = n57236 ^ n57229 ;
  assign n57238 = n57212 & n57237 ;
  assign n57262 = n57261 ^ n57246 ;
  assign n57263 = n57238 & n57262 ;
  assign n57286 = n57285 ^ n57266 ;
  assign n57287 = ~n57263 & ~n57286 ;
  assign n57310 = n57309 ^ n57290 ;
  assign n57311 = n57287 & ~n57310 ;
  assign n57335 = n57334 ^ n57331 ;
  assign n57336 = ~n57311 & n57335 ;
  assign n57344 = n57343 ^ n57339 ;
  assign n57361 = n57360 ^ n57344 ;
  assign n57362 = ~n57336 & n57361 ;
  assign n57364 = n57363 ^ n57362 ;
  assign n57386 = n57385 ^ n57364 ;
  assign n57387 = n57359 ^ n57343 ;
  assign n57388 = n57387 ^ n57336 ;
  assign n57389 = n57335 ^ n57311 ;
  assign n57390 = n57310 ^ n57287 ;
  assign n57391 = n57286 ^ n57263 ;
  assign n57392 = n57262 ^ n57238 ;
  assign n57393 = n57237 ^ n57212 ;
  assign n57394 = n57211 ^ n57188 ;
  assign n57395 = n57187 ^ n57161 ;
  assign n57396 = n57160 ^ n57136 ;
  assign n57397 = n57135 ^ n57111 ;
  assign n57398 = n57110 ^ n57087 ;
  assign n57399 = n57086 ^ n57063 ;
  assign n57400 = n57062 ^ n57038 ;
  assign n57401 = n57037 ^ n57014 ;
  assign n57402 = n57013 ^ n56990 ;
  assign n57403 = n56989 ^ n56966 ;
  assign n57404 = n56965 ^ n56942 ;
  assign n57405 = n56941 ^ n56917 ;
  assign n57406 = n56916 ^ n56892 ;
  assign n57407 = n56891 ^ n56867 ;
  assign n57408 = n56866 ^ n56841 ;
  assign n57409 = n56840 ^ n56817 ;
  assign n57410 = n56816 ^ n56793 ;
  assign n57411 = n56792 ^ n56767 ;
  assign n57412 = n56766 ^ n56742 ;
  assign n57413 = n56741 ^ n56716 ;
  assign n57414 = n56715 ^ n56670 ;
  assign n57415 = n56669 ^ n56622 ;
  assign n57416 = n56621 ^ n56574 ;
  assign n57417 = n56573 ^ n56533 ;
  assign n57418 = ~n56726 & n56756 ;
  assign n57419 = ~n56779 & n57418 ;
  assign n57420 = ~n56802 & ~n57419 ;
  assign n57421 = ~n56829 & ~n57420 ;
  assign n57422 = ~n56854 & n57421 ;
  assign n57423 = ~n56874 & n57422 ;
  assign n57424 = ~n56903 & ~n57423 ;
  assign n57425 = n56927 & n57424 ;
  assign n57426 = ~n56951 & n57425 ;
  assign n57427 = ~n56978 & ~n57426 ;
  assign n57428 = n57005 & ~n57427 ;
  assign n57429 = ~n57026 & ~n57428 ;
  assign n57430 = ~n57047 & ~n57429 ;
  assign n57431 = n57072 & ~n57430 ;
  assign n57432 = n57099 & ~n57431 ;
  assign n57433 = ~n57125 & n57432 ;
  assign n57434 = n57142 & ~n57433 ;
  assign n57435 = n57166 & ~n57434 ;
  assign n57436 = n57194 & n57435 ;
  assign n57437 = n57217 & ~n57436 ;
  assign n57438 = ~n57249 & n57437 ;
  assign n57439 = n57278 & ~n57438 ;
  assign n57440 = ~n57299 & n57439 ;
  assign n57441 = ~n57320 & n57440 ;
  assign n57442 = ~n57350 & n57441 ;
  assign n57443 = ~n57372 & n57442 ;
  assign n57444 = ~n56525 & n57443 ;
  assign n57445 = ~n56562 & ~n57444 ;
  assign n57446 = n56605 & ~n57445 ;
  assign n57447 = n56652 & n57446 ;
  assign n57448 = n57447 ^ n56697 ;
  assign n57449 = n57446 ^ n56652 ;
  assign n57450 = n57445 ^ n56605 ;
  assign n57451 = n57444 ^ n56562 ;
  assign n57452 = n57443 ^ n56525 ;
  assign n57453 = n57442 ^ n57372 ;
  assign n57454 = n57441 ^ n57350 ;
  assign n57455 = n57440 ^ n57320 ;
  assign n57456 = n57439 ^ n57299 ;
  assign n57457 = n57438 ^ n57278 ;
  assign n57458 = n57437 ^ n57249 ;
  assign n57459 = n57436 ^ n57217 ;
  assign n57460 = n57435 ^ n57194 ;
  assign n57461 = n57434 ^ n57166 ;
  assign n57462 = n57433 ^ n57142 ;
  assign n57463 = n57432 ^ n57125 ;
  assign n57464 = n57431 ^ n57099 ;
  assign n57465 = n57430 ^ n57072 ;
  assign n57466 = n57429 ^ n57047 ;
  assign n57467 = n57428 ^ n57026 ;
  assign n57468 = n57427 ^ n57005 ;
  assign n57469 = n57426 ^ n56978 ;
  assign n57470 = n57425 ^ n56951 ;
  assign n57471 = n57424 ^ n56927 ;
  assign n57472 = n57423 ^ n56903 ;
  assign n57473 = n57422 ^ n56874 ;
  assign n57474 = n57421 ^ n56854 ;
  assign n57475 = n57420 ^ n56829 ;
  assign n57476 = n57419 ^ n56802 ;
  assign n57477 = n57418 ^ n56779 ;
  assign n57478 = ~n55720 & ~n55722 ;
  assign n57479 = n55716 & n57478 ;
  assign n57480 = n55712 & n57479 ;
  assign n57481 = n55708 & n57480 ;
  assign n57482 = n55704 & n57481 ;
  assign n57483 = ~n55700 & n57482 ;
  assign n57484 = n55696 & ~n57483 ;
  assign n57485 = ~n55688 & n57484 ;
  assign n57486 = ~n55686 & ~n57485 ;
  assign n57487 = n55681 & n57486 ;
  assign n57488 = n55670 & n57487 ;
  assign n57489 = ~n55675 & ~n57488 ;
  assign n57490 = ~n55665 & ~n57489 ;
  assign n57491 = n55663 & n57490 ;
  assign n57492 = n55655 & ~n57491 ;
  assign n57493 = ~n55653 & ~n57492 ;
  assign n57494 = n56102 & ~n57493 ;
  assign n57495 = ~n56105 & ~n57494 ;
  assign n57496 = ~n56515 & n57495 ;
  assign n57497 = ~n56541 & n57496 ;
  assign n57498 = ~n56587 & ~n57497 ;
  assign n57499 = ~n56635 & ~n57498 ;
  assign n57500 = ~n56684 & ~n57499 ;
  assign n57501 = n56017 & n57500 ;
  assign n57502 = ~n56022 & n57501 ;
  assign n57503 = ~n56013 & ~n57502 ;
  assign n57504 = n56009 & n57503 ;
  assign n57505 = ~n56003 & ~n57504 ;
  assign n57506 = n55735 & n57505 ;
  assign n57507 = n57506 ^ n55731 ;
  assign n57508 = n57505 ^ n55735 ;
  assign n57509 = n57504 ^ n56003 ;
  assign n57510 = n57503 ^ n56009 ;
  assign n57511 = n57502 ^ n56013 ;
  assign n57512 = n57501 ^ n56022 ;
  assign n57513 = n57500 ^ n56017 ;
  assign n57514 = n57499 ^ n56684 ;
  assign n57515 = n57498 ^ n56635 ;
  assign n57516 = n57497 ^ n56587 ;
  assign n57517 = n57496 ^ n56541 ;
  assign n57518 = n57495 ^ n56515 ;
  assign n57519 = n57494 ^ n56105 ;
  assign n57520 = n57493 ^ n56102 ;
  assign n57521 = n57492 ^ n55653 ;
  assign n57522 = n57491 ^ n55655 ;
  assign n57523 = n57490 ^ n55663 ;
  assign n57524 = n57489 ^ n55665 ;
  assign n57525 = n57488 ^ n55675 ;
  assign n57526 = n57487 ^ n55670 ;
  assign n57527 = n57486 ^ n55681 ;
  assign n57528 = n57485 ^ n55686 ;
  assign n57529 = n57484 ^ n55688 ;
  assign n57530 = n57483 ^ n55696 ;
  assign n57531 = n57482 ^ n55700 ;
  assign n57532 = n57481 ^ n55704 ;
  assign n57533 = n57480 ^ n55708 ;
  assign n57534 = n57479 ^ n55712 ;
  assign n57535 = n57478 ^ n55716 ;
  assign n57536 = n55722 ^ n55720 ;
  assign n57537 = n55139 & ~n55141 ;
  assign n57538 = n55132 & ~n57537 ;
  assign n57539 = ~n55134 & ~n57538 ;
  assign n57540 = ~n55321 & n57539 ;
  assign n57541 = n55128 & n57540 ;
  assign n57542 = n55122 & ~n57541 ;
  assign n57543 = ~n55118 & n57542 ;
  assign n57544 = ~n55114 & n57543 ;
  assign n57545 = n55345 & ~n57544 ;
  assign n57546 = ~n55445 & ~n57545 ;
  assign n57547 = n55646 & ~n57546 ;
  assign n57548 = ~n55693 & ~n57547 ;
  assign n57549 = ~n55689 & ~n57548 ;
  assign n57550 = ~n55683 & ~n57549 ;
  assign n57551 = n55678 & n57550 ;
  assign n57552 = ~n55671 & ~n57551 ;
  assign n57553 = n55750 & ~n57552 ;
  assign n57554 = ~n55666 & n57553 ;
  assign n57555 = n55661 & ~n57554 ;
  assign n57556 = n55657 & n57555 ;
  assign n57557 = n55105 & ~n57556 ;
  assign n57558 = n55890 & n57557 ;
  assign n57559 = ~n55102 & n57558 ;
  assign n57560 = ~n55287 & n57559 ;
  assign n57561 = n55290 & n57560 ;
  assign n57562 = ~n55279 & n57561 ;
  assign n57563 = ~n55277 & ~n57562 ;
  assign n57564 = n55273 & ~n57563 ;
  assign n57565 = ~n55156 & n57564 ;
  assign n57566 = n57565 ^ n55152 ;
  assign n57567 = n57564 ^ n55156 ;
  assign n57568 = n57563 ^ n55273 ;
  assign n57569 = n57562 ^ n55277 ;
  assign n57570 = n57561 ^ n55279 ;
  assign n57571 = n57560 ^ n55290 ;
  assign n57572 = n57559 ^ n55287 ;
  assign n57573 = n57558 ^ n55102 ;
  assign n57574 = n57557 ^ n55890 ;
  assign n57575 = n57556 ^ n55105 ;
  assign n57576 = n57555 ^ n55657 ;
  assign n57577 = n57554 ^ n55661 ;
  assign n57578 = n57553 ^ n55666 ;
  assign n57579 = n57552 ^ n55750 ;
  assign n57580 = n57551 ^ n55671 ;
  assign n57581 = n57550 ^ n55678 ;
  assign n57582 = n57549 ^ n55683 ;
  assign n57583 = n57548 ^ n55689 ;
  assign n57584 = n57547 ^ n55693 ;
  assign n57585 = n57546 ^ n55646 ;
  assign n57586 = n57545 ^ n55445 ;
  assign n57587 = n57544 ^ n55345 ;
  assign n57588 = n57543 ^ n55114 ;
  assign n57589 = n57542 ^ n55118 ;
  assign n57590 = n57541 ^ n55122 ;
  assign n57591 = n57540 ^ n55128 ;
  assign n57592 = n57539 ^ n55321 ;
  assign n57593 = n57538 ^ n55134 ;
  assign n57594 = n57537 ^ n55132 ;
  assign n57595 = n55141 ^ n55139 ;
  assign n57596 = ~n54210 & n54214 ;
  assign n57597 = n54205 & n57596 ;
  assign n57598 = n54631 & n57597 ;
  assign n57599 = n54638 & n57598 ;
  assign n57600 = n54200 & ~n57599 ;
  assign n57601 = ~n54195 & n57600 ;
  assign n57602 = n54190 & n57601 ;
  assign n57603 = n54182 & n57602 ;
  assign n57604 = n54177 & ~n57603 ;
  assign n57605 = ~n54172 & n57604 ;
  assign n57606 = n54667 & n57605 ;
  assign n57607 = ~n54791 & ~n57606 ;
  assign n57608 = n54795 & ~n57607 ;
  assign n57609 = n54809 & ~n57608 ;
  assign n57610 = ~n55095 & n57609 ;
  assign n57611 = n55173 & ~n57610 ;
  assign n57612 = ~n55169 & ~n57611 ;
  assign n57613 = n55165 & ~n57612 ;
  assign n57614 = ~n55209 & n57613 ;
  assign n57615 = n55106 & n57614 ;
  assign n57616 = ~n54556 & n57615 ;
  assign n57617 = n54562 & ~n57616 ;
  assign n57618 = n54552 & n57617 ;
  assign n57619 = ~n54548 & n57618 ;
  assign n57620 = ~n54596 & n57619 ;
  assign n57621 = n54236 & ~n57620 ;
  assign n57622 = n57621 ^ n54234 ;
  assign n57623 = n57620 ^ n54236 ;
  assign n57624 = n57619 ^ n54596 ;
  assign n57625 = n57618 ^ n54548 ;
  assign n57626 = n57617 ^ n54552 ;
  assign n57627 = n57616 ^ n54562 ;
  assign n57628 = n57615 ^ n54556 ;
  assign n57629 = n57614 ^ n55106 ;
  assign n57630 = n57613 ^ n55209 ;
  assign n57631 = n57612 ^ n55165 ;
  assign n57632 = n57611 ^ n55169 ;
  assign n57633 = n57610 ^ n55173 ;
  assign n57634 = n57609 ^ n55095 ;
  assign n57635 = n57608 ^ n54809 ;
  assign n57636 = n57607 ^ n54795 ;
  assign n57637 = n57606 ^ n54791 ;
  assign n57638 = n57605 ^ n54667 ;
  assign n57639 = n57604 ^ n54172 ;
  assign n57640 = n57603 ^ n54177 ;
  assign n57641 = n57602 ^ n54182 ;
  assign n57642 = n57601 ^ n54190 ;
  assign n57643 = n57600 ^ n54195 ;
  assign n57644 = n57599 ^ n54200 ;
  assign n57645 = n57598 ^ n54638 ;
  assign n57646 = n57597 ^ n54631 ;
  assign n57647 = n57596 ^ n54205 ;
  assign n57648 = n54214 ^ n54210 ;
  assign y0 = ~n57386 ;
  assign y1 = ~n57388 ;
  assign y2 = n57389 ;
  assign y3 = ~n57390 ;
  assign y4 = n57391 ;
  assign y5 = ~n57392 ;
  assign y6 = ~n57393 ;
  assign y7 = n57394 ;
  assign y8 = ~n57395 ;
  assign y9 = ~n57396 ;
  assign y10 = ~n57397 ;
  assign y11 = ~n57398 ;
  assign y12 = n57399 ;
  assign y13 = ~n57400 ;
  assign y14 = ~n57401 ;
  assign y15 = n57402 ;
  assign y16 = ~n57403 ;
  assign y17 = n57404 ;
  assign y18 = ~n57405 ;
  assign y19 = ~n57406 ;
  assign y20 = ~n57407 ;
  assign y21 = ~n57408 ;
  assign y22 = ~n57409 ;
  assign y23 = n57410 ;
  assign y24 = ~n57411 ;
  assign y25 = ~n57412 ;
  assign y26 = ~n57413 ;
  assign y27 = ~n57414 ;
  assign y28 = n57415 ;
  assign y29 = n57416 ;
  assign y30 = n57417 ;
  assign y31 = n56533 ;
  assign y32 = n57448 ;
  assign y33 = ~n57449 ;
  assign y34 = n57450 ;
  assign y35 = n57451 ;
  assign y36 = n57452 ;
  assign y37 = n57453 ;
  assign y38 = n57454 ;
  assign y39 = n57455 ;
  assign y40 = n57456 ;
  assign y41 = n57457 ;
  assign y42 = ~n57458 ;
  assign y43 = ~n57459 ;
  assign y44 = ~n57460 ;
  assign y45 = n57461 ;
  assign y46 = ~n57462 ;
  assign y47 = n57463 ;
  assign y48 = n57464 ;
  assign y49 = ~n57465 ;
  assign y50 = ~n57466 ;
  assign y51 = n57467 ;
  assign y52 = n57468 ;
  assign y53 = n57469 ;
  assign y54 = n57470 ;
  assign y55 = ~n57471 ;
  assign y56 = ~n57472 ;
  assign y57 = ~n57473 ;
  assign y58 = ~n57474 ;
  assign y59 = n57475 ;
  assign y60 = ~n57476 ;
  assign y61 = ~n57477 ;
  assign y62 = ~n56757 ;
  assign y63 = n56726 ;
  assign y64 = n57507 ;
  assign y65 = n57508 ;
  assign y66 = n57509 ;
  assign y67 = ~n57510 ;
  assign y68 = ~n57511 ;
  assign y69 = ~n57512 ;
  assign y70 = n57513 ;
  assign y71 = n57514 ;
  assign y72 = ~n57515 ;
  assign y73 = n57516 ;
  assign y74 = n57517 ;
  assign y75 = n57518 ;
  assign y76 = ~n57519 ;
  assign y77 = ~n57520 ;
  assign y78 = ~n57521 ;
  assign y79 = ~n57522 ;
  assign y80 = ~n57523 ;
  assign y81 = ~n57524 ;
  assign y82 = n57525 ;
  assign y83 = ~n57526 ;
  assign y84 = ~n57527 ;
  assign y85 = ~n57528 ;
  assign y86 = ~n57529 ;
  assign y87 = ~n57530 ;
  assign y88 = n57531 ;
  assign y89 = ~n57532 ;
  assign y90 = ~n57533 ;
  assign y91 = ~n57534 ;
  assign y92 = ~n57535 ;
  assign y93 = ~n57536 ;
  assign y94 = ~n55722 ;
  assign y95 = n55728 ;
  assign y96 = ~n57566 ;
  assign y97 = ~n57567 ;
  assign y98 = ~n57568 ;
  assign y99 = ~n57569 ;
  assign y100 = ~n57570 ;
  assign y101 = n57571 ;
  assign y102 = ~n57572 ;
  assign y103 = ~n57573 ;
  assign y104 = n57574 ;
  assign y105 = ~n57575 ;
  assign y106 = ~n57576 ;
  assign y107 = n57577 ;
  assign y108 = ~n57578 ;
  assign y109 = ~n57579 ;
  assign y110 = ~n57580 ;
  assign y111 = n57581 ;
  assign y112 = n57582 ;
  assign y113 = ~n57583 ;
  assign y114 = n57584 ;
  assign y115 = n57585 ;
  assign y116 = n57586 ;
  assign y117 = n57587 ;
  assign y118 = ~n57588 ;
  assign y119 = ~n57589 ;
  assign y120 = ~n57590 ;
  assign y121 = ~n57591 ;
  assign y122 = n57592 ;
  assign y123 = ~n57593 ;
  assign y124 = ~n57594 ;
  assign y125 = n57595 ;
  assign y126 = ~n55141 ;
  assign y127 = ~n55145 ;
  assign y128 = ~n57622 ;
  assign y129 = n57623 ;
  assign y130 = ~n57624 ;
  assign y131 = ~n57625 ;
  assign y132 = n57626 ;
  assign y133 = ~n57627 ;
  assign y134 = n57628 ;
  assign y135 = ~n57629 ;
  assign y136 = n57630 ;
  assign y137 = n57631 ;
  assign y138 = n57632 ;
  assign y139 = n57633 ;
  assign y140 = ~n57634 ;
  assign y141 = ~n57635 ;
  assign y142 = n57636 ;
  assign y143 = n57637 ;
  assign y144 = ~n57638 ;
  assign y145 = n57639 ;
  assign y146 = n57640 ;
  assign y147 = n57641 ;
  assign y148 = n57642 ;
  assign y149 = ~n57643 ;
  assign y150 = ~n57644 ;
  assign y151 = ~n57645 ;
  assign y152 = ~n57646 ;
  assign y153 = ~n57647 ;
  assign y154 = n57648 ;
  assign y155 = n54214 ;
  assign y156 = ~n54218 ;
  assign y157 = ~n54616 ;
  assign y158 = ~n54220 ;
  assign y159 = n54229 ;
endmodule
