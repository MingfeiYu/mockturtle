module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n135 , n136 , n137 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n157 , n158 , n161 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n187 , n188 , n189 , n191 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n204 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n253 , n254 , n255 , n258 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n271 , n272 , n273 , n274 , n275 , n277 , n278 , n279 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n312 , n313 , n314 , n315 , n316 , n318 , n319 , n320 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n358 , n359 , n360 , n362 , n363 , n364 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n426 , n427 , n428 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n480 , n481 , n482 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n539 , n540 , n541 , n542 , n543 , n544 , n546 , n547 , n548 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n583 , n584 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n614 , n615 , n616 , n617 , n618 , n620 , n621 , n622 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n683 , n684 , n685 , n686 , n687 , n689 , n690 , n691 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n755 , n756 , n757 , n758 , n759 , n761 , n762 , n763 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n839 , n840 , n841 , n843 , n844 , n845 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n920 , n921 , n922 , n923 , n924 , n926 , n927 , n928 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n956 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1011 , n1012 , n1013 , n1015 , n1016 , n1017 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1101 , n1102 , n1103 , n1105 , n1106 , n1107 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1240 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1543 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1890 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2021 , n2022 , n2023 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3208 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3719 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4283 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4873 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6198 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6937 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7673 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7938 , n7939 , n7940 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8384 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8480 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8744 , n8745 , n8746 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8905 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8952 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9270 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9372 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9635 , n9636 , n9637 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9839 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15661 , n15662 , n15663 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16680 , n16681 , n16682 , n16683 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18085 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19132 , n19133 , n19134 , n19135 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19555 , n19556 , n19557 , n19558 , n19559 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19986 , n19988 , n19989 , n19990 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20014 , n20015 , n20016 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20065 , n20066 , n20067 , n20068 , n20069 , n20075 , n20076 , n20077 , n20078 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20092 , n20093 , n20094 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20103 , n20104 , n20105 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20229 , n20231 , n20233 , n20234 , n20235 , n20236 , n20240 , n20241 , n20242 , n20243 , n20245 , n20247 , n20248 , n20250 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20273 , n20279 , n20280 , n20281 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20433 , n20434 , n20435 , n20436 , n20437 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20498 , n20499 , n20500 , n20504 , n20505 , n20506 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 ;
  assign n129 = x0 & x64 ;
  assign n131 = x0 & x65 ;
  assign n130 = x1 & x64 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = x66 ^ x2 ;
  assign n146 = n129 & ~n133 ;
  assign n135 = x1 & x65 ;
  assign n143 = n135 ^ x66 ;
  assign n144 = ~x64 & ~n143 ;
  assign n136 = n135 ^ x2 ;
  assign n137 = n136 ^ x66 ;
  assign n140 = x64 & ~n137 ;
  assign n141 = n140 ^ x66 ;
  assign n142 = ~x0 & n141 ;
  assign n145 = n144 ^ n142 ;
  assign n147 = n146 ^ n145 ;
  assign n170 = x2 & ~x64 ;
  assign n171 = ~x65 & ~x66 ;
  assign n172 = n170 & n171 ;
  assign n173 = n172 ^ n170 ;
  assign n177 = ~x0 & ~n135 ;
  assign n178 = n173 & n177 ;
  assign n175 = x3 & x64 ;
  assign n174 = n173 ^ x2 ;
  assign n176 = n175 ^ n174 ;
  assign n179 = n178 ^ n176 ;
  assign n164 = x2 & x65 ;
  assign n165 = n164 ^ x66 ;
  assign n166 = ~x1 & n165 ;
  assign n149 = ~x64 & ~x65 ;
  assign n150 = n149 ^ x64 ;
  assign n151 = n150 ^ x65 ;
  assign n152 = ~x66 & n151 ;
  assign n148 = x65 & x66 ;
  assign n153 = n152 ^ n148 ;
  assign n10129 = x2 ^ x1 ;
  assign n157 = n153 & n10129 ;
  assign n155 = x67 ^ x1 ;
  assign n158 = n157 ^ n155 ;
  assign n161 = n158 ^ n133 ;
  assign n167 = n166 ^ n161 ;
  assign n168 = ~x0 & n167 ;
  assign n169 = n168 ^ n158 ;
  assign n180 = n179 ^ n169 ;
  assign n213 = n169 & n179 ;
  assign n207 = x2 & x66 ;
  assign n208 = n207 ^ x67 ;
  assign n209 = ~x1 & n208 ;
  assign n182 = x67 & ~n152 ;
  assign n181 = ~x67 & ~n148 ;
  assign n183 = n182 ^ n181 ;
  assign n187 = n183 & n10129 ;
  assign n185 = x68 ^ x1 ;
  assign n188 = n187 ^ n185 ;
  assign n154 = x67 ^ x2 ;
  assign n204 = n188 ^ n154 ;
  assign n210 = n209 ^ n204 ;
  assign n211 = ~x0 & n210 ;
  assign n197 = x65 ^ x3 ;
  assign n198 = x3 ^ x2 ;
  assign n199 = ~n197 & n198 ;
  assign n193 = x2 & x3 ;
  assign n194 = n193 ^ x4 ;
  assign n195 = ~x64 & n194 ;
  assign n189 = x4 ^ x2 ;
  assign n196 = n195 ^ n189 ;
  assign n200 = n199 ^ n196 ;
  assign n201 = n200 ^ n188 ;
  assign n212 = n211 ^ n201 ;
  assign n214 = n213 ^ n212 ;
  assign n255 = x1 ^ x0 ;
  assign n261 = x2 & x67 ;
  assign n262 = n261 ^ x68 ;
  assign n263 = ~n255 & n262 ;
  assign n248 = ~x68 & ~n182 ;
  assign n247 = x68 & ~n181 ;
  assign n249 = n248 ^ n247 ;
  assign n253 = n249 & n10129 ;
  assign n251 = x69 ^ x1 ;
  assign n254 = n253 ^ n251 ;
  assign n184 = x68 ^ x2 ;
  assign n258 = n254 ^ n184 ;
  assign n264 = n263 ^ n258 ;
  assign n265 = ~x0 & n264 ;
  assign n266 = n265 ^ n254 ;
  assign n243 = x66 & n198 ;
  assign n229 = x5 ^ x4 ;
  assign n230 = n198 & ~n229 ;
  assign n231 = n230 ^ n198 ;
  assign n239 = x65 & n231 ;
  assign n232 = x5 ^ x3 ;
  assign n233 = ~n198 & n232 ;
  assign n234 = n229 & n233 ;
  assign n240 = n239 ^ n234 ;
  assign n241 = ~x64 & n240 ;
  assign n242 = n241 ^ n234 ;
  assign n244 = n243 ^ n242 ;
  assign n191 = x4 ^ x3 ;
  assign n227 = n191 & ~n198 ;
  assign n228 = x65 & n227 ;
  assign n245 = n244 ^ n228 ;
  assign n218 = n189 ^ x65 ;
  assign n219 = ~x64 & ~n218 ;
  assign n220 = n219 ^ n189 ;
  assign n221 = n198 ^ x64 ;
  assign n222 = n221 ^ x5 ;
  assign n223 = ~n220 & ~n222 ;
  assign n224 = n223 ^ x64 ;
  assign n225 = x5 & ~n224 ;
  assign n226 = n225 ^ x5 ;
  assign n246 = n245 ^ n226 ;
  assign n267 = n266 ^ n246 ;
  assign n215 = n213 ^ n200 ;
  assign n216 = n212 & n215 ;
  assign n217 = n216 ^ n200 ;
  assign n268 = n267 ^ n217 ;
  assign n303 = n266 ^ n217 ;
  assign n304 = n267 & n303 ;
  assign n305 = n304 ^ n266 ;
  assign n294 = x65 & n234 ;
  assign n293 = x67 & n230 ;
  assign n295 = n294 ^ n293 ;
  assign n296 = n295 ^ x5 ;
  assign n291 = n153 ^ x67 ;
  assign n292 = n231 & ~n291 ;
  assign n297 = n296 ^ n292 ;
  assign n290 = x66 & n227 ;
  assign n298 = n297 ^ n290 ;
  assign n289 = n225 & ~n245 ;
  assign n299 = n298 ^ n289 ;
  assign n287 = x6 ^ x5 ;
  assign n288 = x64 & n287 ;
  assign n300 = n299 ^ n288 ;
  assign n272 = x69 & ~n248 ;
  assign n271 = ~x69 & ~n247 ;
  assign n273 = n272 ^ n271 ;
  assign n277 = n273 & n10129 ;
  assign n275 = x70 ^ x1 ;
  assign n278 = n277 ^ n275 ;
  assign n301 = n300 ^ n278 ;
  assign n282 = x2 & x68 ;
  assign n283 = n282 ^ x69 ;
  assign n284 = ~x1 & n283 ;
  assign n250 = x69 ^ x2 ;
  assign n279 = n278 ^ n250 ;
  assign n285 = n284 ^ n279 ;
  assign n286 = ~x0 & n285 ;
  assign n302 = n301 ^ n286 ;
  assign n306 = n305 ^ n302 ;
  assign n349 = ~n289 & n298 ;
  assign n350 = ~n288 & n349 ;
  assign n351 = n350 ^ n298 ;
  assign n343 = x66 & n234 ;
  assign n342 = x68 & n230 ;
  assign n344 = n343 ^ n342 ;
  assign n345 = n344 ^ x5 ;
  assign n340 = n183 ^ x68 ;
  assign n341 = n231 & ~n340 ;
  assign n346 = n345 ^ n341 ;
  assign n339 = x67 & n227 ;
  assign n347 = n346 ^ n339 ;
  assign n337 = ~x7 & x64 ;
  assign n328 = ~x5 & ~x6 ;
  assign n329 = n328 ^ n287 ;
  assign n334 = x65 & ~n328 ;
  assign n335 = n334 ^ x64 ;
  assign n336 = n329 & n335 ;
  assign n338 = n337 ^ n336 ;
  assign n348 = n347 ^ n338 ;
  assign n352 = n351 ^ n348 ;
  assign n313 = ~x70 & ~n272 ;
  assign n312 = x70 & ~n271 ;
  assign n314 = n313 ^ n312 ;
  assign n318 = n314 & n10129 ;
  assign n316 = x71 ^ x1 ;
  assign n319 = n318 ^ n316 ;
  assign n353 = n352 ^ n319 ;
  assign n323 = x2 & x69 ;
  assign n324 = n323 ^ x70 ;
  assign n325 = ~x1 & n324 ;
  assign n274 = x70 ^ x2 ;
  assign n320 = n319 ^ n274 ;
  assign n326 = n325 ^ n320 ;
  assign n327 = ~x0 & n326 ;
  assign n354 = n353 ^ n327 ;
  assign n307 = n305 ^ n300 ;
  assign n308 = ~n302 & n307 ;
  assign n309 = n308 ^ n305 ;
  assign n355 = n354 ^ n309 ;
  assign n409 = n352 ^ n309 ;
  assign n410 = n354 & n409 ;
  assign n411 = n410 ^ n352 ;
  assign n404 = x68 & n227 ;
  assign n394 = ~n288 & ~n338 ;
  assign n389 = x7 ^ x6 ;
  assign n390 = ~n287 & n389 ;
  assign n391 = x65 & n390 ;
  assign n382 = x8 ^ x7 ;
  assign n383 = n287 & ~n382 ;
  assign n384 = n383 ^ n287 ;
  assign n387 = ~n150 & n384 ;
  assign n386 = x66 & n287 ;
  assign n388 = n387 ^ n386 ;
  assign n392 = n391 ^ n388 ;
  assign n381 = n328 & n337 ;
  assign n393 = n392 ^ n381 ;
  assign n395 = n394 ^ n393 ;
  assign n396 = n395 ^ n392 ;
  assign n379 = n337 ^ x64 ;
  assign n380 = ~n329 & n379 ;
  assign n397 = n396 ^ n380 ;
  assign n398 = ~x8 & ~n397 ;
  assign n399 = n398 ^ n395 ;
  assign n400 = n399 ^ x5 ;
  assign n378 = x67 & n234 ;
  assign n401 = n400 ^ n378 ;
  assign n377 = x69 & n230 ;
  assign n402 = n401 ^ n377 ;
  assign n375 = n249 ^ x69 ;
  assign n376 = n231 & ~n375 ;
  assign n403 = n402 ^ n376 ;
  assign n405 = n404 ^ n403 ;
  assign n372 = n351 ^ n347 ;
  assign n373 = ~n348 & n372 ;
  assign n374 = n373 ^ n351 ;
  assign n406 = n405 ^ n374 ;
  assign n356 = x71 ^ x70 ;
  assign n358 = n314 & n356 ;
  assign n362 = ~n358 & n10129 ;
  assign n360 = x72 ^ x1 ;
  assign n363 = n362 ^ n360 ;
  assign n407 = n406 ^ n363 ;
  assign n367 = x2 & x70 ;
  assign n368 = n367 ^ x71 ;
  assign n369 = ~x1 & n368 ;
  assign n315 = x71 ^ x2 ;
  assign n364 = n363 ^ n315 ;
  assign n370 = n369 ^ n364 ;
  assign n371 = ~x0 & n370 ;
  assign n408 = n407 ^ n371 ;
  assign n412 = n411 ^ n408 ;
  assign n462 = n399 ^ n374 ;
  assign n463 = ~n405 & ~n462 ;
  assign n464 = n463 ^ n399 ;
  assign n460 = x69 & n227 ;
  assign n453 = x8 & ~n393 ;
  assign n454 = n395 & n453 ;
  assign n445 = ~n287 & n382 ;
  assign n446 = ~n389 & n445 ;
  assign n447 = x65 & n446 ;
  assign n444 = x67 & n383 ;
  assign n448 = n447 ^ n444 ;
  assign n449 = n448 ^ x8 ;
  assign n443 = ~n291 & n384 ;
  assign n450 = n449 ^ n443 ;
  assign n442 = x66 & n390 ;
  assign n451 = n450 ^ n442 ;
  assign n440 = x9 ^ x8 ;
  assign n441 = x64 & n440 ;
  assign n452 = n451 ^ n441 ;
  assign n455 = n454 ^ n452 ;
  assign n456 = n455 ^ x5 ;
  assign n439 = x68 & n234 ;
  assign n457 = n456 ^ n439 ;
  assign n438 = x70 & n230 ;
  assign n458 = n457 ^ n438 ;
  assign n436 = n273 ^ x70 ;
  assign n437 = n231 & ~n436 ;
  assign n459 = n458 ^ n437 ;
  assign n461 = n460 ^ n459 ;
  assign n465 = n464 ^ n461 ;
  assign n418 = x71 & ~x72 ;
  assign n421 = ~n313 & n418 ;
  assign n416 = x72 ^ x71 ;
  assign n419 = n418 ^ n416 ;
  assign n420 = ~n312 & n419 ;
  assign n422 = n421 ^ n420 ;
  assign n426 = ~n422 & n10129 ;
  assign n424 = x73 ^ x1 ;
  assign n427 = n426 ^ n424 ;
  assign n466 = n465 ^ n427 ;
  assign n431 = x2 & x71 ;
  assign n432 = n431 ^ x72 ;
  assign n433 = ~x1 & n432 ;
  assign n359 = x72 ^ x2 ;
  assign n428 = n427 ^ n359 ;
  assign n434 = n433 ^ n428 ;
  assign n435 = ~x0 & n434 ;
  assign n467 = n466 ^ n435 ;
  assign n413 = n411 ^ n406 ;
  assign n414 = n408 & ~n413 ;
  assign n415 = n414 ^ n411 ;
  assign n468 = n467 ^ n415 ;
  assign n530 = n465 ^ n415 ;
  assign n531 = ~n467 & ~n530 ;
  assign n532 = n531 ^ n465 ;
  assign n525 = x70 & n227 ;
  assign n515 = x66 & n446 ;
  assign n514 = x68 & n383 ;
  assign n516 = n515 ^ n514 ;
  assign n517 = n516 ^ x8 ;
  assign n513 = ~n340 & n384 ;
  assign n518 = n517 ^ n513 ;
  assign n512 = x67 & n390 ;
  assign n519 = n518 ^ n512 ;
  assign n508 = n451 & ~n454 ;
  assign n509 = ~n441 & n508 ;
  assign n510 = n509 ^ n451 ;
  assign n503 = ~x8 & ~x9 ;
  assign n504 = n503 ^ n440 ;
  assign n505 = n504 ^ x10 ;
  assign n506 = ~x64 & ~n505 ;
  assign n497 = x65 ^ x9 ;
  assign n500 = x65 ^ x8 ;
  assign n501 = ~n497 & n500 ;
  assign n498 = x10 ^ x8 ;
  assign n502 = n501 ^ n498 ;
  assign n507 = n506 ^ n502 ;
  assign n511 = n510 ^ n507 ;
  assign n520 = n519 ^ n511 ;
  assign n521 = n520 ^ x5 ;
  assign n496 = x69 & n234 ;
  assign n522 = n521 ^ n496 ;
  assign n495 = x71 & n230 ;
  assign n523 = n522 ^ n495 ;
  assign n493 = n314 ^ x71 ;
  assign n494 = n231 & ~n493 ;
  assign n524 = n523 ^ n494 ;
  assign n526 = n525 ^ n524 ;
  assign n490 = n464 ^ n455 ;
  assign n491 = ~n461 & ~n490 ;
  assign n492 = n491 ^ n464 ;
  assign n527 = n526 ^ n492 ;
  assign n473 = n421 ^ x72 ;
  assign n474 = x73 & n473 ;
  assign n475 = n474 ^ x73 ;
  assign n471 = x72 & ~x73 ;
  assign n472 = ~n420 & n471 ;
  assign n476 = n475 ^ n472 ;
  assign n480 = ~n476 & n10129 ;
  assign n478 = x74 ^ x1 ;
  assign n481 = n480 ^ n478 ;
  assign n528 = n527 ^ n481 ;
  assign n485 = x2 & x72 ;
  assign n486 = n485 ^ x73 ;
  assign n487 = ~x1 & n486 ;
  assign n423 = x73 ^ x2 ;
  assign n482 = n481 ^ n423 ;
  assign n488 = n487 ^ n482 ;
  assign n489 = ~x0 & n488 ;
  assign n529 = n528 ^ n489 ;
  assign n533 = n532 ^ n529 ;
  assign n605 = n520 ^ n492 ;
  assign n606 = n526 & ~n605 ;
  assign n607 = n606 ^ n520 ;
  assign n603 = x71 & n227 ;
  assign n596 = x68 & n390 ;
  assign n593 = x69 & n383 ;
  assign n591 = x67 & n446 ;
  assign n570 = ~x10 & ~n440 ;
  assign n578 = n570 ^ n503 ;
  assign n586 = n578 ^ n440 ;
  assign n587 = x64 & ~n586 ;
  assign n588 = ~x11 & n587 ;
  assign n579 = x65 & n578 ;
  assign n569 = x11 ^ x10 ;
  assign n571 = n570 ^ n569 ;
  assign n568 = x11 & ~n440 ;
  assign n572 = n571 ^ n568 ;
  assign n573 = n572 ^ n440 ;
  assign n576 = ~n150 & ~n573 ;
  assign n575 = x66 & n440 ;
  assign n577 = n576 ^ n575 ;
  assign n580 = n579 ^ n577 ;
  assign n566 = ~x10 & x64 ;
  assign n567 = n503 & n566 ;
  assign n581 = n580 ^ n567 ;
  assign n583 = n581 ^ x11 ;
  assign n564 = x11 & ~n441 ;
  assign n565 = ~n507 & n564 ;
  assign n584 = n583 ^ n565 ;
  assign n589 = n588 ^ n584 ;
  assign n590 = n589 ^ x8 ;
  assign n592 = n591 ^ n590 ;
  assign n594 = n593 ^ n592 ;
  assign n563 = ~n375 & n384 ;
  assign n595 = n594 ^ n563 ;
  assign n597 = n596 ^ n595 ;
  assign n560 = n519 ^ n510 ;
  assign n561 = ~n511 & n560 ;
  assign n562 = n561 ^ n519 ;
  assign n598 = n597 ^ n562 ;
  assign n599 = n598 ^ x5 ;
  assign n559 = x70 & n234 ;
  assign n600 = n599 ^ n559 ;
  assign n558 = x72 & n230 ;
  assign n601 = n600 ^ n558 ;
  assign n556 = n358 ^ x72 ;
  assign n557 = n231 & n556 ;
  assign n602 = n601 ^ n557 ;
  assign n604 = n603 ^ n602 ;
  assign n608 = n607 ^ n604 ;
  assign n541 = ~x74 & ~n474 ;
  assign n539 = n472 ^ x73 ;
  assign n540 = x74 & n539 ;
  assign n542 = n541 ^ n540 ;
  assign n546 = n542 & n10129 ;
  assign n544 = x75 ^ x1 ;
  assign n547 = n546 ^ n544 ;
  assign n609 = n608 ^ n547 ;
  assign n551 = x2 & x73 ;
  assign n552 = n551 ^ x74 ;
  assign n553 = ~x1 & n552 ;
  assign n477 = x74 ^ x2 ;
  assign n548 = n547 ^ n477 ;
  assign n554 = n553 ^ n548 ;
  assign n555 = ~x0 & n554 ;
  assign n610 = n609 ^ n555 ;
  assign n534 = n532 ^ n527 ;
  assign n535 = n529 & n534 ;
  assign n536 = n535 ^ n532 ;
  assign n611 = n610 ^ n536 ;
  assign n674 = n608 ^ n536 ;
  assign n675 = n610 & ~n674 ;
  assign n676 = n675 ^ n608 ;
  assign n669 = x72 & n227 ;
  assign n658 = x68 & n446 ;
  assign n657 = x70 & n383 ;
  assign n659 = n658 ^ n657 ;
  assign n660 = n659 ^ x8 ;
  assign n656 = n384 & ~n436 ;
  assign n661 = n660 ^ n656 ;
  assign n655 = x69 & n390 ;
  assign n662 = n661 ^ n655 ;
  assign n646 = n568 ^ n504 ;
  assign n647 = n569 & ~n646 ;
  assign n648 = x65 & n647 ;
  assign n645 = x67 & ~n572 ;
  assign n649 = n648 ^ n645 ;
  assign n650 = n649 ^ x11 ;
  assign n644 = ~n291 & ~n573 ;
  assign n651 = n650 ^ n644 ;
  assign n643 = x66 & n578 ;
  assign n652 = n651 ^ n643 ;
  assign n641 = x12 ^ x11 ;
  assign n642 = x64 & n641 ;
  assign n653 = n652 ^ n642 ;
  assign n640 = n565 & ~n581 ;
  assign n654 = n653 ^ n640 ;
  assign n663 = n662 ^ n654 ;
  assign n637 = n589 ^ n562 ;
  assign n638 = ~n597 & n637 ;
  assign n639 = n638 ^ n562 ;
  assign n664 = n663 ^ n639 ;
  assign n665 = n664 ^ x5 ;
  assign n636 = x71 & n234 ;
  assign n666 = n665 ^ n636 ;
  assign n635 = x73 & n230 ;
  assign n667 = n666 ^ n635 ;
  assign n633 = n422 ^ x73 ;
  assign n634 = n231 & n633 ;
  assign n668 = n667 ^ n634 ;
  assign n670 = n669 ^ n668 ;
  assign n630 = n607 ^ n598 ;
  assign n631 = ~n604 & n630 ;
  assign n632 = n631 ^ n607 ;
  assign n671 = n670 ^ n632 ;
  assign n615 = x75 & ~n541 ;
  assign n614 = ~x75 & ~n540 ;
  assign n616 = n615 ^ n614 ;
  assign n620 = n616 & n10129 ;
  assign n618 = x76 ^ x1 ;
  assign n621 = n620 ^ n618 ;
  assign n672 = n671 ^ n621 ;
  assign n625 = x2 & x74 ;
  assign n626 = n625 ^ x75 ;
  assign n627 = ~x1 & n626 ;
  assign n543 = x75 ^ x2 ;
  assign n622 = n621 ^ n543 ;
  assign n628 = n627 ^ n622 ;
  assign n629 = ~x0 & n628 ;
  assign n673 = n672 ^ n629 ;
  assign n677 = n676 ^ n673 ;
  assign n746 = n664 ^ n632 ;
  assign n747 = n670 & n746 ;
  assign n748 = n747 ^ n664 ;
  assign n744 = x73 & n227 ;
  assign n737 = x70 & n390 ;
  assign n727 = ~n642 & n652 ;
  assign n728 = ~n640 & n727 ;
  assign n729 = n728 ^ n652 ;
  assign n726 = ~n150 & n641 ;
  assign n730 = n729 ^ n726 ;
  assign n717 = x13 ^ x12 ;
  assign n718 = n717 ^ x65 ;
  assign n719 = n718 ^ x12 ;
  assign n720 = n719 ^ n717 ;
  assign n723 = n641 & n720 ;
  assign n724 = n723 ^ n717 ;
  assign n725 = x64 & n724 ;
  assign n731 = n730 ^ n725 ;
  assign n712 = x66 & n647 ;
  assign n711 = x68 & ~n572 ;
  assign n713 = n712 ^ n711 ;
  assign n714 = n713 ^ x11 ;
  assign n710 = ~n340 & ~n573 ;
  assign n715 = n714 ^ n710 ;
  assign n709 = x67 & n578 ;
  assign n716 = n715 ^ n709 ;
  assign n732 = n731 ^ n716 ;
  assign n733 = n732 ^ x8 ;
  assign n708 = x69 & n446 ;
  assign n734 = n733 ^ n708 ;
  assign n707 = x71 & n383 ;
  assign n735 = n734 ^ n707 ;
  assign n706 = n384 & ~n493 ;
  assign n736 = n735 ^ n706 ;
  assign n738 = n737 ^ n736 ;
  assign n703 = n662 ^ n639 ;
  assign n704 = n663 & n703 ;
  assign n705 = n704 ^ n662 ;
  assign n739 = n738 ^ n705 ;
  assign n740 = n739 ^ x5 ;
  assign n702 = x72 & n234 ;
  assign n741 = n740 ^ n702 ;
  assign n701 = x74 & n230 ;
  assign n742 = n741 ^ n701 ;
  assign n699 = n476 ^ x74 ;
  assign n700 = n231 & n699 ;
  assign n743 = n742 ^ n700 ;
  assign n745 = n744 ^ n743 ;
  assign n749 = n748 ^ n745 ;
  assign n684 = ~x76 & ~n615 ;
  assign n683 = x76 & ~n614 ;
  assign n685 = n684 ^ n683 ;
  assign n689 = n685 & n10129 ;
  assign n687 = x77 ^ x1 ;
  assign n690 = n689 ^ n687 ;
  assign n750 = n749 ^ n690 ;
  assign n694 = x2 & x75 ;
  assign n695 = n694 ^ x76 ;
  assign n696 = ~x1 & n695 ;
  assign n617 = x76 ^ x2 ;
  assign n691 = n690 ^ n617 ;
  assign n697 = n696 ^ n691 ;
  assign n698 = ~x0 & n697 ;
  assign n751 = n750 ^ n698 ;
  assign n678 = n676 ^ n671 ;
  assign n679 = ~n673 & n678 ;
  assign n680 = n679 ^ n676 ;
  assign n752 = n751 ^ n680 ;
  assign n830 = n749 ^ n680 ;
  assign n831 = n751 & n830 ;
  assign n832 = n831 ^ n749 ;
  assign n825 = x74 & n227 ;
  assign n817 = n732 ^ n705 ;
  assign n818 = n738 & n817 ;
  assign n819 = n818 ^ n732 ;
  assign n815 = x71 & n390 ;
  assign n807 = n729 ^ n716 ;
  assign n808 = n731 & n807 ;
  assign n809 = n808 ^ n729 ;
  assign n804 = n726 ^ x64 ;
  assign n805 = x14 & n804 ;
  assign n800 = x11 & x12 ;
  assign n801 = x13 & x64 ;
  assign n802 = n800 & n801 ;
  assign n794 = x67 & n647 ;
  assign n793 = x69 & ~n572 ;
  assign n795 = n794 ^ n793 ;
  assign n796 = n795 ^ x11 ;
  assign n792 = ~n375 & ~n573 ;
  assign n797 = n796 ^ n792 ;
  assign n791 = x68 & n578 ;
  assign n798 = n797 ^ n791 ;
  assign n788 = ~n641 & n717 ;
  assign n789 = x65 & n788 ;
  assign n781 = x14 ^ x13 ;
  assign n782 = n641 & ~n781 ;
  assign n783 = n782 ^ n641 ;
  assign n786 = ~n150 & n783 ;
  assign n785 = x66 & n641 ;
  assign n787 = n786 ^ n785 ;
  assign n790 = n789 ^ n787 ;
  assign n799 = n798 ^ n790 ;
  assign n803 = n802 ^ n799 ;
  assign n806 = n805 ^ n803 ;
  assign n810 = n809 ^ n806 ;
  assign n811 = n810 ^ x8 ;
  assign n780 = x70 & n446 ;
  assign n812 = n811 ^ n780 ;
  assign n779 = x72 & n383 ;
  assign n813 = n812 ^ n779 ;
  assign n778 = n384 & n556 ;
  assign n814 = n813 ^ n778 ;
  assign n816 = n815 ^ n814 ;
  assign n820 = n819 ^ n816 ;
  assign n821 = n820 ^ x5 ;
  assign n777 = x73 & n234 ;
  assign n822 = n821 ^ n777 ;
  assign n776 = x75 & n230 ;
  assign n823 = n822 ^ n776 ;
  assign n774 = n542 ^ x75 ;
  assign n775 = n231 & ~n774 ;
  assign n824 = n823 ^ n775 ;
  assign n826 = n825 ^ n824 ;
  assign n771 = n748 ^ n739 ;
  assign n772 = ~n745 & n771 ;
  assign n773 = n772 ^ n748 ;
  assign n827 = n826 ^ n773 ;
  assign n756 = x77 & ~n684 ;
  assign n755 = ~x77 & ~n683 ;
  assign n757 = n756 ^ n755 ;
  assign n761 = n757 & n10129 ;
  assign n759 = x78 ^ x1 ;
  assign n762 = n761 ^ n759 ;
  assign n828 = n827 ^ n762 ;
  assign n766 = x2 & x76 ;
  assign n767 = n766 ^ x77 ;
  assign n768 = ~x1 & n767 ;
  assign n686 = x77 ^ x2 ;
  assign n763 = n762 ^ n686 ;
  assign n769 = n768 ^ n763 ;
  assign n770 = ~x0 & n769 ;
  assign n829 = n828 ^ n770 ;
  assign n833 = n832 ^ n829 ;
  assign n907 = n820 ^ n773 ;
  assign n908 = n826 & n907 ;
  assign n909 = n908 ^ n820 ;
  assign n905 = x75 & n227 ;
  assign n898 = x72 & n390 ;
  assign n887 = x68 & n647 ;
  assign n886 = x70 & ~n572 ;
  assign n888 = n887 ^ n886 ;
  assign n889 = n888 ^ x11 ;
  assign n885 = ~n436 & ~n573 ;
  assign n890 = n889 ^ n885 ;
  assign n884 = x69 & n578 ;
  assign n891 = n890 ^ n884 ;
  assign n875 = x14 ^ x12 ;
  assign n876 = ~n641 & n875 ;
  assign n877 = n781 & n876 ;
  assign n878 = x65 & n877 ;
  assign n874 = x67 & n782 ;
  assign n879 = n878 ^ n874 ;
  assign n880 = n879 ^ x14 ;
  assign n873 = ~n291 & n783 ;
  assign n881 = n880 ^ n873 ;
  assign n872 = x66 & n788 ;
  assign n882 = n881 ^ n872 ;
  assign n869 = x15 ^ x14 ;
  assign n870 = x64 & n869 ;
  assign n866 = x14 & ~n790 ;
  assign n867 = n804 ^ n802 ;
  assign n868 = n866 & ~n867 ;
  assign n871 = n870 ^ n868 ;
  assign n883 = n882 ^ n871 ;
  assign n892 = n891 ^ n883 ;
  assign n863 = n809 ^ n798 ;
  assign n864 = ~n806 & n863 ;
  assign n865 = n864 ^ n809 ;
  assign n893 = n892 ^ n865 ;
  assign n894 = n893 ^ x8 ;
  assign n862 = x71 & n446 ;
  assign n895 = n894 ^ n862 ;
  assign n861 = x73 & n383 ;
  assign n896 = n895 ^ n861 ;
  assign n860 = n384 & n633 ;
  assign n897 = n896 ^ n860 ;
  assign n899 = n898 ^ n897 ;
  assign n857 = n819 ^ n810 ;
  assign n858 = ~n816 & n857 ;
  assign n859 = n858 ^ n819 ;
  assign n900 = n899 ^ n859 ;
  assign n901 = n900 ^ x5 ;
  assign n856 = x74 & n234 ;
  assign n902 = n901 ^ n856 ;
  assign n855 = x76 & n230 ;
  assign n903 = n902 ^ n855 ;
  assign n853 = n616 ^ x76 ;
  assign n854 = n231 & ~n853 ;
  assign n904 = n903 ^ n854 ;
  assign n906 = n905 ^ n904 ;
  assign n910 = n909 ^ n906 ;
  assign n837 = x78 ^ x77 ;
  assign n839 = n757 & n837 ;
  assign n843 = ~n839 & n10129 ;
  assign n841 = x79 ^ x1 ;
  assign n844 = n843 ^ n841 ;
  assign n911 = n910 ^ n844 ;
  assign n848 = x2 & x77 ;
  assign n849 = n848 ^ x78 ;
  assign n850 = ~x1 & n849 ;
  assign n758 = x78 ^ x2 ;
  assign n845 = n844 ^ n758 ;
  assign n851 = n850 ^ n845 ;
  assign n852 = ~x0 & n851 ;
  assign n912 = n911 ^ n852 ;
  assign n834 = n832 ^ n827 ;
  assign n835 = ~n829 & n834 ;
  assign n836 = n835 ^ n832 ;
  assign n913 = n912 ^ n836 ;
  assign n1002 = n910 ^ n836 ;
  assign n1003 = n912 & n1002 ;
  assign n1004 = n1003 ^ n910 ;
  assign n997 = x76 & n227 ;
  assign n989 = n893 ^ n859 ;
  assign n990 = n899 & n989 ;
  assign n991 = n990 ^ n893 ;
  assign n987 = x73 & n390 ;
  assign n979 = n891 ^ n865 ;
  assign n980 = n892 & n979 ;
  assign n981 = n980 ^ n891 ;
  assign n977 = x70 & n578 ;
  assign n967 = x66 & n877 ;
  assign n966 = x68 & n782 ;
  assign n968 = n967 ^ n966 ;
  assign n969 = n968 ^ x14 ;
  assign n965 = ~n340 & n783 ;
  assign n970 = n969 ^ n965 ;
  assign n964 = x67 & n788 ;
  assign n971 = n970 ^ n964 ;
  assign n958 = x14 & x15 ;
  assign n959 = n958 ^ x16 ;
  assign n960 = ~x64 & n959 ;
  assign n954 = x16 ^ x14 ;
  assign n961 = n960 ^ n954 ;
  assign n952 = x65 ^ x15 ;
  assign n953 = n869 & ~n952 ;
  assign n962 = n961 ^ n953 ;
  assign n949 = ~n870 & n882 ;
  assign n950 = ~n868 & n949 ;
  assign n951 = n950 ^ n882 ;
  assign n963 = n962 ^ n951 ;
  assign n972 = n971 ^ n963 ;
  assign n973 = n972 ^ x11 ;
  assign n948 = x69 & n647 ;
  assign n974 = n973 ^ n948 ;
  assign n947 = x71 & ~n572 ;
  assign n975 = n974 ^ n947 ;
  assign n946 = ~n493 & ~n573 ;
  assign n976 = n975 ^ n946 ;
  assign n978 = n977 ^ n976 ;
  assign n982 = n981 ^ n978 ;
  assign n983 = n982 ^ x8 ;
  assign n945 = x72 & n446 ;
  assign n984 = n983 ^ n945 ;
  assign n944 = x74 & n383 ;
  assign n985 = n984 ^ n944 ;
  assign n943 = n384 & n699 ;
  assign n986 = n985 ^ n943 ;
  assign n988 = n987 ^ n986 ;
  assign n992 = n991 ^ n988 ;
  assign n993 = n992 ^ x5 ;
  assign n942 = x75 & n234 ;
  assign n994 = n993 ^ n942 ;
  assign n941 = x77 & n230 ;
  assign n995 = n994 ^ n941 ;
  assign n939 = n685 ^ x77 ;
  assign n940 = n231 & ~n939 ;
  assign n996 = n995 ^ n940 ;
  assign n998 = n997 ^ n996 ;
  assign n936 = n909 ^ n900 ;
  assign n937 = ~n906 & n936 ;
  assign n938 = n937 ^ n909 ;
  assign n999 = n998 ^ n938 ;
  assign n914 = x79 ^ x78 ;
  assign n920 = ~x79 & n757 ;
  assign n921 = n920 ^ n756 ;
  assign n922 = n914 & ~n921 ;
  assign n926 = ~n922 & n10129 ;
  assign n924 = x80 ^ x1 ;
  assign n927 = n926 ^ n924 ;
  assign n1000 = n999 ^ n927 ;
  assign n931 = x2 & x78 ;
  assign n932 = n931 ^ x79 ;
  assign n933 = ~x1 & n932 ;
  assign n840 = x79 ^ x2 ;
  assign n928 = n927 ^ n840 ;
  assign n934 = n933 ^ n928 ;
  assign n935 = ~x0 & n934 ;
  assign n1001 = n1000 ^ n935 ;
  assign n1005 = n1004 ^ n1001 ;
  assign n1092 = n992 ^ n938 ;
  assign n1093 = n998 & n1092 ;
  assign n1094 = n1093 ^ n992 ;
  assign n1090 = x77 & n227 ;
  assign n1083 = x74 & n390 ;
  assign n1076 = x71 & n578 ;
  assign n1069 = x68 & n788 ;
  assign n1062 = x17 & ~n870 ;
  assign n1063 = ~n962 & n1062 ;
  assign n956 = x16 ^ x15 ;
  assign n1058 = ~n869 & n956 ;
  assign n1059 = x65 & n1058 ;
  assign n1047 = x17 ^ x16 ;
  assign n1053 = n869 & ~n1047 ;
  assign n1054 = n1053 ^ n869 ;
  assign n1055 = ~n150 & n1054 ;
  assign n1052 = x66 & n869 ;
  assign n1056 = n1055 ^ n1052 ;
  assign n1057 = n1056 ^ x17 ;
  assign n1060 = n1059 ^ n1057 ;
  assign n1048 = x17 ^ x15 ;
  assign n1049 = ~n869 & n1048 ;
  assign n1050 = n1047 & n1049 ;
  assign n1051 = x64 & n1050 ;
  assign n1061 = n1060 ^ n1051 ;
  assign n1064 = n1063 ^ n1061 ;
  assign n1065 = n1064 ^ x14 ;
  assign n1046 = x67 & n877 ;
  assign n1066 = n1065 ^ n1046 ;
  assign n1045 = x69 & n782 ;
  assign n1067 = n1066 ^ n1045 ;
  assign n1044 = ~n375 & n783 ;
  assign n1068 = n1067 ^ n1044 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1041 = n971 ^ n962 ;
  assign n1042 = ~n963 & n1041 ;
  assign n1043 = n1042 ^ n971 ;
  assign n1071 = n1070 ^ n1043 ;
  assign n1072 = n1071 ^ x11 ;
  assign n1040 = x70 & n647 ;
  assign n1073 = n1072 ^ n1040 ;
  assign n1039 = x72 & ~n572 ;
  assign n1074 = n1073 ^ n1039 ;
  assign n1038 = n556 & ~n573 ;
  assign n1075 = n1074 ^ n1038 ;
  assign n1077 = n1076 ^ n1075 ;
  assign n1035 = n981 ^ n972 ;
  assign n1036 = ~n978 & n1035 ;
  assign n1037 = n1036 ^ n981 ;
  assign n1078 = n1077 ^ n1037 ;
  assign n1079 = n1078 ^ x8 ;
  assign n1034 = x73 & n446 ;
  assign n1080 = n1079 ^ n1034 ;
  assign n1033 = x75 & n383 ;
  assign n1081 = n1080 ^ n1033 ;
  assign n1032 = n384 & ~n774 ;
  assign n1082 = n1081 ^ n1032 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1029 = n991 ^ n982 ;
  assign n1030 = ~n988 & n1029 ;
  assign n1031 = n1030 ^ n991 ;
  assign n1085 = n1084 ^ n1031 ;
  assign n1086 = n1085 ^ x5 ;
  assign n1028 = x76 & n234 ;
  assign n1087 = n1086 ^ n1028 ;
  assign n1027 = x78 & n230 ;
  assign n1088 = n1087 ^ n1027 ;
  assign n1025 = n757 ^ x78 ;
  assign n1026 = n231 & ~n1025 ;
  assign n1089 = n1088 ^ n1026 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1095 = n1094 ^ n1091 ;
  assign n1009 = x80 ^ x79 ;
  assign n1011 = ~n922 & n1009 ;
  assign n1015 = ~n1011 & n10129 ;
  assign n1013 = x81 ^ x1 ;
  assign n1016 = n1015 ^ n1013 ;
  assign n1096 = n1095 ^ n1016 ;
  assign n1020 = x2 & x79 ;
  assign n1021 = n1020 ^ x80 ;
  assign n1022 = ~n255 & n1021 ;
  assign n923 = x80 ^ x2 ;
  assign n1017 = n1016 ^ n923 ;
  assign n1023 = n1022 ^ n1017 ;
  assign n1024 = ~x0 & n1023 ;
  assign n1097 = n1096 ^ n1024 ;
  assign n1006 = n1004 ^ n999 ;
  assign n1007 = ~n1001 & n1006 ;
  assign n1008 = n1007 ^ n1004 ;
  assign n1098 = n1097 ^ n1008 ;
  assign n1183 = n1095 ^ n1008 ;
  assign n1184 = n1097 & n1183 ;
  assign n1185 = n1184 ^ n1095 ;
  assign n1178 = x78 & n227 ;
  assign n1170 = n1078 ^ n1031 ;
  assign n1171 = n1084 & n1170 ;
  assign n1172 = n1171 ^ n1078 ;
  assign n1168 = x75 & n390 ;
  assign n1160 = n1071 ^ n1037 ;
  assign n1161 = n1077 & n1160 ;
  assign n1162 = n1161 ^ n1071 ;
  assign n1158 = x72 & n578 ;
  assign n1150 = n1064 ^ n1043 ;
  assign n1151 = n1070 & n1150 ;
  assign n1152 = n1151 ^ n1064 ;
  assign n1148 = x69 & n788 ;
  assign n1137 = x65 & n1050 ;
  assign n1136 = x67 & n1053 ;
  assign n1138 = n1137 ^ n1136 ;
  assign n1139 = n1138 ^ x17 ;
  assign n1135 = ~n291 & n1054 ;
  assign n1140 = n1139 ^ n1135 ;
  assign n1134 = x66 & n1058 ;
  assign n1141 = n1140 ^ n1134 ;
  assign n1132 = x18 ^ x17 ;
  assign n1133 = x64 & n1132 ;
  assign n1142 = n1141 ^ n1133 ;
  assign n1131 = n1061 & n1063 ;
  assign n1143 = n1142 ^ n1131 ;
  assign n1144 = n1143 ^ x14 ;
  assign n1130 = x68 & n877 ;
  assign n1145 = n1144 ^ n1130 ;
  assign n1129 = x70 & n782 ;
  assign n1146 = n1145 ^ n1129 ;
  assign n1128 = ~n436 & n783 ;
  assign n1147 = n1146 ^ n1128 ;
  assign n1149 = n1148 ^ n1147 ;
  assign n1153 = n1152 ^ n1149 ;
  assign n1154 = n1153 ^ x11 ;
  assign n1127 = x71 & n647 ;
  assign n1155 = n1154 ^ n1127 ;
  assign n1126 = x73 & ~n572 ;
  assign n1156 = n1155 ^ n1126 ;
  assign n1125 = ~n573 & n633 ;
  assign n1157 = n1156 ^ n1125 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1163 = n1162 ^ n1159 ;
  assign n1164 = n1163 ^ x8 ;
  assign n1124 = x74 & n446 ;
  assign n1165 = n1164 ^ n1124 ;
  assign n1123 = x76 & n383 ;
  assign n1166 = n1165 ^ n1123 ;
  assign n1122 = n384 & ~n853 ;
  assign n1167 = n1166 ^ n1122 ;
  assign n1169 = n1168 ^ n1167 ;
  assign n1173 = n1172 ^ n1169 ;
  assign n1174 = n1173 ^ x5 ;
  assign n1121 = x77 & n234 ;
  assign n1175 = n1174 ^ n1121 ;
  assign n1120 = x79 & n230 ;
  assign n1176 = n1175 ^ n1120 ;
  assign n1118 = n839 ^ x79 ;
  assign n1119 = n231 & n1118 ;
  assign n1177 = n1176 ^ n1119 ;
  assign n1179 = n1178 ^ n1177 ;
  assign n1115 = n1094 ^ n1085 ;
  assign n1116 = ~n1091 & n1115 ;
  assign n1117 = n1116 ^ n1094 ;
  assign n1180 = n1179 ^ n1117 ;
  assign n1099 = x81 ^ x80 ;
  assign n1101 = ~n1011 & n1099 ;
  assign n1105 = ~n1101 & n10129 ;
  assign n1103 = x82 ^ x1 ;
  assign n1106 = n1105 ^ n1103 ;
  assign n1181 = n1180 ^ n1106 ;
  assign n1110 = x2 & x80 ;
  assign n1111 = n1110 ^ x81 ;
  assign n1112 = ~x1 & n1111 ;
  assign n1012 = x81 ^ x2 ;
  assign n1107 = n1106 ^ n1012 ;
  assign n1113 = n1112 ^ n1107 ;
  assign n1114 = ~x0 & n1113 ;
  assign n1182 = n1181 ^ n1114 ;
  assign n1186 = n1185 ^ n1182 ;
  assign n1279 = n1173 ^ n1117 ;
  assign n1280 = n1179 & n1279 ;
  assign n1281 = n1280 ^ n1173 ;
  assign n1277 = x79 & n227 ;
  assign n1270 = x76 & n390 ;
  assign n1263 = x73 & n578 ;
  assign n1256 = x70 & n788 ;
  assign n1248 = ~n1133 & n1141 ;
  assign n1249 = ~n1131 & n1248 ;
  assign n1250 = n1249 ^ n1141 ;
  assign n1242 = x17 & x18 ;
  assign n1243 = n1242 ^ x19 ;
  assign n1244 = ~x64 & n1243 ;
  assign n1238 = x19 ^ x17 ;
  assign n1245 = n1244 ^ n1238 ;
  assign n1236 = x65 ^ x18 ;
  assign n1237 = n1132 & ~n1236 ;
  assign n1246 = n1245 ^ n1237 ;
  assign n1231 = x66 & n1050 ;
  assign n1230 = x68 & n1053 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1233 = n1232 ^ x17 ;
  assign n1229 = ~n340 & n1054 ;
  assign n1234 = n1233 ^ n1229 ;
  assign n1228 = x67 & n1058 ;
  assign n1235 = n1234 ^ n1228 ;
  assign n1247 = n1246 ^ n1235 ;
  assign n1251 = n1250 ^ n1247 ;
  assign n1252 = n1251 ^ x14 ;
  assign n1227 = x69 & n877 ;
  assign n1253 = n1252 ^ n1227 ;
  assign n1226 = x71 & n782 ;
  assign n1254 = n1253 ^ n1226 ;
  assign n1225 = ~n493 & n783 ;
  assign n1255 = n1254 ^ n1225 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1222 = n1152 ^ n1143 ;
  assign n1223 = ~n1149 & n1222 ;
  assign n1224 = n1223 ^ n1152 ;
  assign n1258 = n1257 ^ n1224 ;
  assign n1259 = n1258 ^ x11 ;
  assign n1221 = x72 & n647 ;
  assign n1260 = n1259 ^ n1221 ;
  assign n1220 = x74 & ~n572 ;
  assign n1261 = n1260 ^ n1220 ;
  assign n1219 = ~n573 & n699 ;
  assign n1262 = n1261 ^ n1219 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1216 = n1162 ^ n1153 ;
  assign n1217 = ~n1159 & n1216 ;
  assign n1218 = n1217 ^ n1162 ;
  assign n1265 = n1264 ^ n1218 ;
  assign n1266 = n1265 ^ x8 ;
  assign n1215 = x75 & n446 ;
  assign n1267 = n1266 ^ n1215 ;
  assign n1214 = x77 & n383 ;
  assign n1268 = n1267 ^ n1214 ;
  assign n1213 = n384 & ~n939 ;
  assign n1269 = n1268 ^ n1213 ;
  assign n1271 = n1270 ^ n1269 ;
  assign n1210 = n1172 ^ n1163 ;
  assign n1211 = ~n1169 & n1210 ;
  assign n1212 = n1211 ^ n1172 ;
  assign n1272 = n1271 ^ n1212 ;
  assign n1273 = n1272 ^ x5 ;
  assign n1209 = x78 & n234 ;
  assign n1274 = n1273 ^ n1209 ;
  assign n1208 = x80 & n230 ;
  assign n1275 = n1274 ^ n1208 ;
  assign n1206 = n922 ^ x80 ;
  assign n1207 = n231 & n1206 ;
  assign n1276 = n1275 ^ n1207 ;
  assign n1278 = n1277 ^ n1276 ;
  assign n1282 = n1281 ^ n1278 ;
  assign n1190 = x82 ^ x81 ;
  assign n1192 = ~n1101 & n1190 ;
  assign n1194 = x83 ^ x1 ;
  assign n1193 = x83 ^ x2 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1196 = ~n1192 & n1195 ;
  assign n1197 = n1196 ^ n1194 ;
  assign n1283 = n1282 ^ n1197 ;
  assign n1201 = x2 & x81 ;
  assign n1202 = n1201 ^ x82 ;
  assign n1203 = ~x1 & n1202 ;
  assign n1102 = x82 ^ x2 ;
  assign n1198 = n1197 ^ n1102 ;
  assign n1204 = n1203 ^ n1198 ;
  assign n1205 = ~x0 & n1204 ;
  assign n1284 = n1283 ^ n1205 ;
  assign n1187 = n1185 ^ n1180 ;
  assign n1188 = ~n1182 & n1187 ;
  assign n1189 = n1188 ^ n1185 ;
  assign n1285 = n1284 ^ n1189 ;
  assign n1388 = n1282 ^ n1189 ;
  assign n1389 = n1284 & n1388 ;
  assign n1390 = n1389 ^ n1282 ;
  assign n1383 = x80 & n227 ;
  assign n1375 = n1265 ^ n1212 ;
  assign n1376 = n1271 & n1375 ;
  assign n1377 = n1376 ^ n1265 ;
  assign n1373 = x77 & n390 ;
  assign n1365 = n1258 ^ n1218 ;
  assign n1366 = n1264 & n1365 ;
  assign n1367 = n1366 ^ n1258 ;
  assign n1363 = x74 & n578 ;
  assign n1355 = n1251 ^ n1224 ;
  assign n1356 = n1257 & n1355 ;
  assign n1357 = n1356 ^ n1251 ;
  assign n1353 = x71 & n788 ;
  assign n1346 = x68 & n1058 ;
  assign n1339 = x20 & ~n1133 ;
  assign n1340 = ~n1246 & n1339 ;
  assign n1240 = x19 ^ x18 ;
  assign n1335 = ~n1132 & n1240 ;
  assign n1336 = x65 & n1335 ;
  assign n1324 = x20 ^ x19 ;
  assign n1330 = n1132 & ~n1324 ;
  assign n1331 = n1330 ^ n1132 ;
  assign n1332 = ~n150 & n1331 ;
  assign n1329 = x66 & n1132 ;
  assign n1333 = n1332 ^ n1329 ;
  assign n1334 = n1333 ^ x20 ;
  assign n1337 = n1336 ^ n1334 ;
  assign n1325 = x20 ^ x18 ;
  assign n1326 = ~n1132 & n1325 ;
  assign n1327 = n1324 & n1326 ;
  assign n1328 = x64 & n1327 ;
  assign n1338 = n1337 ^ n1328 ;
  assign n1341 = n1340 ^ n1338 ;
  assign n1342 = n1341 ^ x17 ;
  assign n1323 = x67 & n1050 ;
  assign n1343 = n1342 ^ n1323 ;
  assign n1322 = x69 & n1053 ;
  assign n1344 = n1343 ^ n1322 ;
  assign n1321 = ~n375 & n1054 ;
  assign n1345 = n1344 ^ n1321 ;
  assign n1347 = n1346 ^ n1345 ;
  assign n1318 = n1250 ^ n1246 ;
  assign n1319 = ~n1247 & n1318 ;
  assign n1320 = n1319 ^ n1250 ;
  assign n1348 = n1347 ^ n1320 ;
  assign n1349 = n1348 ^ x14 ;
  assign n1317 = x70 & n877 ;
  assign n1350 = n1349 ^ n1317 ;
  assign n1316 = x72 & n782 ;
  assign n1351 = n1350 ^ n1316 ;
  assign n1315 = n556 & n783 ;
  assign n1352 = n1351 ^ n1315 ;
  assign n1354 = n1353 ^ n1352 ;
  assign n1358 = n1357 ^ n1354 ;
  assign n1359 = n1358 ^ x11 ;
  assign n1314 = x73 & n647 ;
  assign n1360 = n1359 ^ n1314 ;
  assign n1313 = x75 & ~n572 ;
  assign n1361 = n1360 ^ n1313 ;
  assign n1312 = ~n573 & ~n774 ;
  assign n1362 = n1361 ^ n1312 ;
  assign n1364 = n1363 ^ n1362 ;
  assign n1368 = n1367 ^ n1364 ;
  assign n1369 = n1368 ^ x8 ;
  assign n1311 = x76 & n446 ;
  assign n1370 = n1369 ^ n1311 ;
  assign n1310 = x78 & n383 ;
  assign n1371 = n1370 ^ n1310 ;
  assign n1309 = n384 & ~n1025 ;
  assign n1372 = n1371 ^ n1309 ;
  assign n1374 = n1373 ^ n1372 ;
  assign n1378 = n1377 ^ n1374 ;
  assign n1379 = n1378 ^ x5 ;
  assign n1308 = x79 & n234 ;
  assign n1380 = n1379 ^ n1308 ;
  assign n1307 = x81 & n230 ;
  assign n1381 = n1380 ^ n1307 ;
  assign n1305 = n1011 ^ x81 ;
  assign n1306 = n231 & n1305 ;
  assign n1382 = n1381 ^ n1306 ;
  assign n1384 = n1383 ^ n1382 ;
  assign n1302 = n1281 ^ n1272 ;
  assign n1303 = ~n1278 & n1302 ;
  assign n1304 = n1303 ^ n1281 ;
  assign n1385 = n1384 ^ n1304 ;
  assign n1286 = x83 ^ x82 ;
  assign n1288 = ~n1192 & n1286 ;
  assign n1290 = x84 ^ x1 ;
  assign n1289 = x84 ^ x2 ;
  assign n1291 = n1290 ^ n1289 ;
  assign n1292 = ~n1288 & n1291 ;
  assign n1293 = n1292 ^ n1290 ;
  assign n1386 = n1385 ^ n1293 ;
  assign n1297 = x2 & x82 ;
  assign n1298 = n1297 ^ x83 ;
  assign n1299 = ~n255 & n1298 ;
  assign n1294 = n1293 ^ n1193 ;
  assign n1300 = n1299 ^ n1294 ;
  assign n1301 = ~x0 & n1300 ;
  assign n1387 = n1386 ^ n1301 ;
  assign n1391 = n1390 ^ n1387 ;
  assign n1486 = n1378 ^ n1304 ;
  assign n1487 = n1384 & n1486 ;
  assign n1488 = n1487 ^ n1378 ;
  assign n1484 = x81 & n227 ;
  assign n1477 = x78 & n390 ;
  assign n1470 = x75 & n578 ;
  assign n1463 = x72 & n788 ;
  assign n1455 = n1341 ^ n1320 ;
  assign n1456 = n1347 & n1455 ;
  assign n1457 = n1456 ^ n1341 ;
  assign n1453 = x69 & n1058 ;
  assign n1442 = x65 & n1327 ;
  assign n1441 = x67 & n1330 ;
  assign n1443 = n1442 ^ n1441 ;
  assign n1444 = n1443 ^ x20 ;
  assign n1440 = ~n291 & n1331 ;
  assign n1445 = n1444 ^ n1440 ;
  assign n1439 = x66 & n1335 ;
  assign n1446 = n1445 ^ n1439 ;
  assign n1437 = x21 ^ x20 ;
  assign n1438 = x64 & n1437 ;
  assign n1447 = n1446 ^ n1438 ;
  assign n1436 = n1338 & n1340 ;
  assign n1448 = n1447 ^ n1436 ;
  assign n1449 = n1448 ^ x17 ;
  assign n1435 = x68 & n1050 ;
  assign n1450 = n1449 ^ n1435 ;
  assign n1434 = x70 & n1053 ;
  assign n1451 = n1450 ^ n1434 ;
  assign n1433 = ~n436 & n1054 ;
  assign n1452 = n1451 ^ n1433 ;
  assign n1454 = n1453 ^ n1452 ;
  assign n1458 = n1457 ^ n1454 ;
  assign n1459 = n1458 ^ x14 ;
  assign n1432 = x71 & n877 ;
  assign n1460 = n1459 ^ n1432 ;
  assign n1431 = x73 & n782 ;
  assign n1461 = n1460 ^ n1431 ;
  assign n1430 = n633 & n783 ;
  assign n1462 = n1461 ^ n1430 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1427 = n1357 ^ n1348 ;
  assign n1428 = ~n1354 & n1427 ;
  assign n1429 = n1428 ^ n1357 ;
  assign n1465 = n1464 ^ n1429 ;
  assign n1466 = n1465 ^ x11 ;
  assign n1426 = x74 & n647 ;
  assign n1467 = n1466 ^ n1426 ;
  assign n1425 = x76 & ~n572 ;
  assign n1468 = n1467 ^ n1425 ;
  assign n1424 = ~n573 & ~n853 ;
  assign n1469 = n1468 ^ n1424 ;
  assign n1471 = n1470 ^ n1469 ;
  assign n1421 = n1367 ^ n1358 ;
  assign n1422 = ~n1364 & n1421 ;
  assign n1423 = n1422 ^ n1367 ;
  assign n1472 = n1471 ^ n1423 ;
  assign n1473 = n1472 ^ x8 ;
  assign n1420 = x77 & n446 ;
  assign n1474 = n1473 ^ n1420 ;
  assign n1419 = x79 & n383 ;
  assign n1475 = n1474 ^ n1419 ;
  assign n1418 = n384 & n1118 ;
  assign n1476 = n1475 ^ n1418 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1415 = n1377 ^ n1368 ;
  assign n1416 = ~n1374 & n1415 ;
  assign n1417 = n1416 ^ n1377 ;
  assign n1479 = n1478 ^ n1417 ;
  assign n1480 = n1479 ^ x5 ;
  assign n1414 = x80 & n234 ;
  assign n1481 = n1480 ^ n1414 ;
  assign n1413 = x82 & n230 ;
  assign n1482 = n1481 ^ n1413 ;
  assign n1411 = n1101 ^ x82 ;
  assign n1412 = n231 & n1411 ;
  assign n1483 = n1482 ^ n1412 ;
  assign n1485 = n1484 ^ n1483 ;
  assign n1489 = n1488 ^ n1485 ;
  assign n1395 = x84 ^ x83 ;
  assign n1397 = ~n1288 & n1395 ;
  assign n1399 = x85 ^ x1 ;
  assign n1398 = x85 ^ x2 ;
  assign n1400 = n1399 ^ n1398 ;
  assign n1401 = ~n1397 & n1400 ;
  assign n1402 = n1401 ^ n1399 ;
  assign n1490 = n1489 ^ n1402 ;
  assign n1406 = x2 & x83 ;
  assign n1407 = n1406 ^ x84 ;
  assign n1408 = ~x1 & n1407 ;
  assign n1403 = n1402 ^ n1289 ;
  assign n1409 = n1408 ^ n1403 ;
  assign n1410 = ~x0 & n1409 ;
  assign n1491 = n1490 ^ n1410 ;
  assign n1392 = n1390 ^ n1385 ;
  assign n1393 = ~n1387 & n1392 ;
  assign n1394 = n1393 ^ n1390 ;
  assign n1492 = n1491 ^ n1394 ;
  assign n1601 = n1489 ^ n1394 ;
  assign n1602 = n1491 & n1601 ;
  assign n1603 = n1602 ^ n1489 ;
  assign n1596 = x82 & n227 ;
  assign n1588 = n1472 ^ n1417 ;
  assign n1589 = n1478 & n1588 ;
  assign n1590 = n1589 ^ n1472 ;
  assign n1586 = x79 & n390 ;
  assign n1578 = n1465 ^ n1423 ;
  assign n1579 = n1471 & n1578 ;
  assign n1580 = n1579 ^ n1465 ;
  assign n1576 = x76 & n578 ;
  assign n1568 = n1458 ^ n1429 ;
  assign n1569 = n1464 & n1568 ;
  assign n1570 = n1569 ^ n1458 ;
  assign n1566 = x73 & n788 ;
  assign n1559 = x70 & n1058 ;
  assign n1551 = ~n1438 & n1446 ;
  assign n1552 = ~n1436 & n1551 ;
  assign n1553 = n1552 ^ n1446 ;
  assign n1545 = x20 & x21 ;
  assign n1546 = n1545 ^ x22 ;
  assign n1547 = ~x64 & n1546 ;
  assign n1541 = x22 ^ x20 ;
  assign n1548 = n1547 ^ n1541 ;
  assign n1539 = x65 ^ x21 ;
  assign n1540 = n1437 & ~n1539 ;
  assign n1549 = n1548 ^ n1540 ;
  assign n1534 = x66 & n1327 ;
  assign n1533 = x68 & n1330 ;
  assign n1535 = n1534 ^ n1533 ;
  assign n1536 = n1535 ^ x20 ;
  assign n1532 = ~n340 & n1331 ;
  assign n1537 = n1536 ^ n1532 ;
  assign n1531 = x67 & n1335 ;
  assign n1538 = n1537 ^ n1531 ;
  assign n1550 = n1549 ^ n1538 ;
  assign n1554 = n1553 ^ n1550 ;
  assign n1555 = n1554 ^ x17 ;
  assign n1530 = x69 & n1050 ;
  assign n1556 = n1555 ^ n1530 ;
  assign n1529 = x71 & n1053 ;
  assign n1557 = n1556 ^ n1529 ;
  assign n1528 = ~n493 & n1054 ;
  assign n1558 = n1557 ^ n1528 ;
  assign n1560 = n1559 ^ n1558 ;
  assign n1525 = n1457 ^ n1448 ;
  assign n1526 = ~n1454 & n1525 ;
  assign n1527 = n1526 ^ n1457 ;
  assign n1561 = n1560 ^ n1527 ;
  assign n1562 = n1561 ^ x14 ;
  assign n1524 = x72 & n877 ;
  assign n1563 = n1562 ^ n1524 ;
  assign n1523 = x74 & n782 ;
  assign n1564 = n1563 ^ n1523 ;
  assign n1522 = n699 & n783 ;
  assign n1565 = n1564 ^ n1522 ;
  assign n1567 = n1566 ^ n1565 ;
  assign n1571 = n1570 ^ n1567 ;
  assign n1572 = n1571 ^ x11 ;
  assign n1521 = x75 & n647 ;
  assign n1573 = n1572 ^ n1521 ;
  assign n1520 = x77 & ~n572 ;
  assign n1574 = n1573 ^ n1520 ;
  assign n1519 = ~n573 & ~n939 ;
  assign n1575 = n1574 ^ n1519 ;
  assign n1577 = n1576 ^ n1575 ;
  assign n1581 = n1580 ^ n1577 ;
  assign n1582 = n1581 ^ x8 ;
  assign n1518 = x78 & n446 ;
  assign n1583 = n1582 ^ n1518 ;
  assign n1517 = x80 & n383 ;
  assign n1584 = n1583 ^ n1517 ;
  assign n1516 = n384 & n1206 ;
  assign n1585 = n1584 ^ n1516 ;
  assign n1587 = n1586 ^ n1585 ;
  assign n1591 = n1590 ^ n1587 ;
  assign n1592 = n1591 ^ x5 ;
  assign n1515 = x81 & n234 ;
  assign n1593 = n1592 ^ n1515 ;
  assign n1514 = x83 & n230 ;
  assign n1594 = n1593 ^ n1514 ;
  assign n1512 = n1192 ^ x83 ;
  assign n1513 = n231 & n1512 ;
  assign n1595 = n1594 ^ n1513 ;
  assign n1597 = n1596 ^ n1595 ;
  assign n1509 = n1488 ^ n1479 ;
  assign n1510 = ~n1485 & n1509 ;
  assign n1511 = n1510 ^ n1488 ;
  assign n1598 = n1597 ^ n1511 ;
  assign n1493 = x85 ^ x84 ;
  assign n1495 = ~n1397 & n1493 ;
  assign n1497 = x86 ^ x1 ;
  assign n1496 = x86 ^ x2 ;
  assign n1498 = n1497 ^ n1496 ;
  assign n1499 = ~n1495 & n1498 ;
  assign n1500 = n1499 ^ n1497 ;
  assign n1599 = n1598 ^ n1500 ;
  assign n1504 = x2 & x84 ;
  assign n1505 = n1504 ^ x85 ;
  assign n1506 = ~x1 & n1505 ;
  assign n1501 = n1500 ^ n1398 ;
  assign n1507 = n1506 ^ n1501 ;
  assign n1508 = ~x0 & n1507 ;
  assign n1600 = n1599 ^ n1508 ;
  assign n1604 = n1603 ^ n1600 ;
  assign n1717 = n1591 ^ n1511 ;
  assign n1718 = n1597 & n1717 ;
  assign n1719 = n1718 ^ n1591 ;
  assign n1715 = x83 & n227 ;
  assign n1708 = x80 & n390 ;
  assign n1701 = x77 & n578 ;
  assign n1694 = x74 & n788 ;
  assign n1686 = n1554 ^ n1527 ;
  assign n1687 = n1560 & n1686 ;
  assign n1688 = n1687 ^ n1554 ;
  assign n1684 = x71 & n1058 ;
  assign n1677 = x68 & n1335 ;
  assign n1670 = x23 & ~n1438 ;
  assign n1671 = ~n1549 & n1670 ;
  assign n1543 = x22 ^ x21 ;
  assign n1666 = ~n1437 & n1543 ;
  assign n1667 = x65 & n1666 ;
  assign n1655 = x23 ^ x22 ;
  assign n1661 = n1437 & ~n1655 ;
  assign n1662 = n1661 ^ n1437 ;
  assign n1663 = ~n150 & n1662 ;
  assign n1660 = x66 & n1437 ;
  assign n1664 = n1663 ^ n1660 ;
  assign n1665 = n1664 ^ x23 ;
  assign n1668 = n1667 ^ n1665 ;
  assign n1656 = x23 ^ x21 ;
  assign n1657 = ~n1437 & n1656 ;
  assign n1658 = n1655 & n1657 ;
  assign n1659 = x64 & n1658 ;
  assign n1669 = n1668 ^ n1659 ;
  assign n1672 = n1671 ^ n1669 ;
  assign n1673 = n1672 ^ x20 ;
  assign n1654 = x67 & n1327 ;
  assign n1674 = n1673 ^ n1654 ;
  assign n1653 = x69 & n1330 ;
  assign n1675 = n1674 ^ n1653 ;
  assign n1652 = ~n375 & n1331 ;
  assign n1676 = n1675 ^ n1652 ;
  assign n1678 = n1677 ^ n1676 ;
  assign n1649 = n1553 ^ n1549 ;
  assign n1650 = ~n1550 & n1649 ;
  assign n1651 = n1650 ^ n1553 ;
  assign n1679 = n1678 ^ n1651 ;
  assign n1680 = n1679 ^ x17 ;
  assign n1648 = x70 & n1050 ;
  assign n1681 = n1680 ^ n1648 ;
  assign n1647 = x72 & n1053 ;
  assign n1682 = n1681 ^ n1647 ;
  assign n1646 = n556 & n1054 ;
  assign n1683 = n1682 ^ n1646 ;
  assign n1685 = n1684 ^ n1683 ;
  assign n1689 = n1688 ^ n1685 ;
  assign n1690 = n1689 ^ x14 ;
  assign n1645 = x73 & n877 ;
  assign n1691 = n1690 ^ n1645 ;
  assign n1644 = x75 & n782 ;
  assign n1692 = n1691 ^ n1644 ;
  assign n1643 = ~n774 & n783 ;
  assign n1693 = n1692 ^ n1643 ;
  assign n1695 = n1694 ^ n1693 ;
  assign n1640 = n1570 ^ n1561 ;
  assign n1641 = ~n1567 & n1640 ;
  assign n1642 = n1641 ^ n1570 ;
  assign n1696 = n1695 ^ n1642 ;
  assign n1697 = n1696 ^ x11 ;
  assign n1639 = x76 & n647 ;
  assign n1698 = n1697 ^ n1639 ;
  assign n1638 = x78 & ~n572 ;
  assign n1699 = n1698 ^ n1638 ;
  assign n1637 = ~n573 & ~n1025 ;
  assign n1700 = n1699 ^ n1637 ;
  assign n1702 = n1701 ^ n1700 ;
  assign n1634 = n1580 ^ n1571 ;
  assign n1635 = ~n1577 & n1634 ;
  assign n1636 = n1635 ^ n1580 ;
  assign n1703 = n1702 ^ n1636 ;
  assign n1704 = n1703 ^ x8 ;
  assign n1633 = x79 & n446 ;
  assign n1705 = n1704 ^ n1633 ;
  assign n1632 = x81 & n383 ;
  assign n1706 = n1705 ^ n1632 ;
  assign n1631 = n384 & n1305 ;
  assign n1707 = n1706 ^ n1631 ;
  assign n1709 = n1708 ^ n1707 ;
  assign n1628 = n1590 ^ n1581 ;
  assign n1629 = ~n1587 & n1628 ;
  assign n1630 = n1629 ^ n1590 ;
  assign n1710 = n1709 ^ n1630 ;
  assign n1711 = n1710 ^ x5 ;
  assign n1627 = x82 & n234 ;
  assign n1712 = n1711 ^ n1627 ;
  assign n1626 = x84 & n230 ;
  assign n1713 = n1712 ^ n1626 ;
  assign n1624 = n1288 ^ x84 ;
  assign n1625 = n231 & n1624 ;
  assign n1714 = n1713 ^ n1625 ;
  assign n1716 = n1715 ^ n1714 ;
  assign n1720 = n1719 ^ n1716 ;
  assign n1608 = x86 ^ x85 ;
  assign n1610 = ~n1495 & n1608 ;
  assign n1612 = x87 ^ x1 ;
  assign n1611 = x87 ^ x2 ;
  assign n1613 = n1612 ^ n1611 ;
  assign n1614 = ~n1610 & n1613 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1721 = n1720 ^ n1615 ;
  assign n1619 = x2 & x85 ;
  assign n1620 = n1619 ^ x86 ;
  assign n1621 = ~x1 & n1620 ;
  assign n1616 = n1615 ^ n1496 ;
  assign n1622 = n1621 ^ n1616 ;
  assign n1623 = ~x0 & n1622 ;
  assign n1722 = n1721 ^ n1623 ;
  assign n1605 = n1603 ^ n1598 ;
  assign n1606 = ~n1600 & n1605 ;
  assign n1607 = n1606 ^ n1603 ;
  assign n1723 = n1722 ^ n1607 ;
  assign n1834 = n1720 ^ n1607 ;
  assign n1835 = n1722 & n1834 ;
  assign n1836 = n1835 ^ n1720 ;
  assign n1829 = x84 & n227 ;
  assign n1821 = n1703 ^ n1630 ;
  assign n1822 = n1709 & n1821 ;
  assign n1823 = n1822 ^ n1703 ;
  assign n1819 = x81 & n390 ;
  assign n1811 = n1696 ^ n1636 ;
  assign n1812 = n1702 & n1811 ;
  assign n1813 = n1812 ^ n1696 ;
  assign n1809 = x78 & n578 ;
  assign n1801 = n1689 ^ n1642 ;
  assign n1802 = n1695 & n1801 ;
  assign n1803 = n1802 ^ n1689 ;
  assign n1799 = x75 & n788 ;
  assign n1792 = x72 & n1058 ;
  assign n1784 = n1672 ^ n1651 ;
  assign n1785 = n1678 & n1784 ;
  assign n1786 = n1785 ^ n1672 ;
  assign n1782 = x69 & n1335 ;
  assign n1771 = x65 & n1658 ;
  assign n1770 = x67 & n1661 ;
  assign n1772 = n1771 ^ n1770 ;
  assign n1773 = n1772 ^ x23 ;
  assign n1769 = ~n291 & n1662 ;
  assign n1774 = n1773 ^ n1769 ;
  assign n1768 = x66 & n1666 ;
  assign n1775 = n1774 ^ n1768 ;
  assign n1766 = x24 ^ x23 ;
  assign n1767 = x64 & n1766 ;
  assign n1776 = n1775 ^ n1767 ;
  assign n1765 = n1669 & n1671 ;
  assign n1777 = n1776 ^ n1765 ;
  assign n1778 = n1777 ^ x20 ;
  assign n1764 = x68 & n1327 ;
  assign n1779 = n1778 ^ n1764 ;
  assign n1763 = x70 & n1330 ;
  assign n1780 = n1779 ^ n1763 ;
  assign n1762 = ~n436 & n1331 ;
  assign n1781 = n1780 ^ n1762 ;
  assign n1783 = n1782 ^ n1781 ;
  assign n1787 = n1786 ^ n1783 ;
  assign n1788 = n1787 ^ x17 ;
  assign n1761 = x71 & n1050 ;
  assign n1789 = n1788 ^ n1761 ;
  assign n1760 = x73 & n1053 ;
  assign n1790 = n1789 ^ n1760 ;
  assign n1759 = n633 & n1054 ;
  assign n1791 = n1790 ^ n1759 ;
  assign n1793 = n1792 ^ n1791 ;
  assign n1756 = n1688 ^ n1679 ;
  assign n1757 = ~n1685 & n1756 ;
  assign n1758 = n1757 ^ n1688 ;
  assign n1794 = n1793 ^ n1758 ;
  assign n1795 = n1794 ^ x14 ;
  assign n1755 = x74 & n877 ;
  assign n1796 = n1795 ^ n1755 ;
  assign n1754 = x76 & n782 ;
  assign n1797 = n1796 ^ n1754 ;
  assign n1753 = n783 & ~n853 ;
  assign n1798 = n1797 ^ n1753 ;
  assign n1800 = n1799 ^ n1798 ;
  assign n1804 = n1803 ^ n1800 ;
  assign n1805 = n1804 ^ x11 ;
  assign n1752 = x77 & n647 ;
  assign n1806 = n1805 ^ n1752 ;
  assign n1751 = x79 & ~n572 ;
  assign n1807 = n1806 ^ n1751 ;
  assign n1750 = ~n573 & n1118 ;
  assign n1808 = n1807 ^ n1750 ;
  assign n1810 = n1809 ^ n1808 ;
  assign n1814 = n1813 ^ n1810 ;
  assign n1815 = n1814 ^ x8 ;
  assign n1749 = x80 & n446 ;
  assign n1816 = n1815 ^ n1749 ;
  assign n1748 = x82 & n383 ;
  assign n1817 = n1816 ^ n1748 ;
  assign n1747 = n384 & n1411 ;
  assign n1818 = n1817 ^ n1747 ;
  assign n1820 = n1819 ^ n1818 ;
  assign n1824 = n1823 ^ n1820 ;
  assign n1825 = n1824 ^ x5 ;
  assign n1746 = x83 & n234 ;
  assign n1826 = n1825 ^ n1746 ;
  assign n1745 = x85 & n230 ;
  assign n1827 = n1826 ^ n1745 ;
  assign n1743 = n1397 ^ x85 ;
  assign n1744 = n231 & n1743 ;
  assign n1828 = n1827 ^ n1744 ;
  assign n1830 = n1829 ^ n1828 ;
  assign n1740 = n1719 ^ n1710 ;
  assign n1741 = ~n1716 & n1740 ;
  assign n1742 = n1741 ^ n1719 ;
  assign n1831 = n1830 ^ n1742 ;
  assign n1724 = x87 ^ x86 ;
  assign n1726 = ~n1610 & n1724 ;
  assign n1728 = x88 ^ x1 ;
  assign n1727 = x88 ^ x2 ;
  assign n1729 = n1728 ^ n1727 ;
  assign n1730 = ~n1726 & n1729 ;
  assign n1731 = n1730 ^ n1728 ;
  assign n1832 = n1831 ^ n1731 ;
  assign n1735 = x2 & x86 ;
  assign n1736 = n1735 ^ x87 ;
  assign n1737 = ~x1 & n1736 ;
  assign n1732 = n1731 ^ n1611 ;
  assign n1738 = n1737 ^ n1732 ;
  assign n1739 = ~x0 & n1738 ;
  assign n1833 = n1832 ^ n1739 ;
  assign n1837 = n1836 ^ n1833 ;
  assign n1956 = n1824 ^ n1742 ;
  assign n1957 = n1830 & n1956 ;
  assign n1958 = n1957 ^ n1824 ;
  assign n1954 = x85 & n227 ;
  assign n1947 = x82 & n390 ;
  assign n1940 = x79 & n578 ;
  assign n1933 = x76 & n788 ;
  assign n1925 = n1787 ^ n1758 ;
  assign n1926 = n1793 & n1925 ;
  assign n1927 = n1926 ^ n1787 ;
  assign n1923 = x73 & n1058 ;
  assign n1916 = x70 & n1335 ;
  assign n1908 = ~n1767 & n1775 ;
  assign n1909 = ~n1765 & n1908 ;
  assign n1910 = n1909 ^ n1775 ;
  assign n1902 = x66 & n1658 ;
  assign n1901 = x68 & n1661 ;
  assign n1903 = n1902 ^ n1901 ;
  assign n1904 = n1903 ^ x23 ;
  assign n1900 = ~n340 & n1662 ;
  assign n1905 = n1904 ^ n1900 ;
  assign n1899 = x67 & n1666 ;
  assign n1906 = n1905 ^ n1899 ;
  assign n1896 = x65 ^ x24 ;
  assign n1897 = n1766 & ~n1896 ;
  assign n1892 = x23 & x24 ;
  assign n1893 = n1892 ^ x25 ;
  assign n1894 = ~x64 & n1893 ;
  assign n1888 = x25 ^ x23 ;
  assign n1895 = n1894 ^ n1888 ;
  assign n1898 = n1897 ^ n1895 ;
  assign n1907 = n1906 ^ n1898 ;
  assign n1911 = n1910 ^ n1907 ;
  assign n1912 = n1911 ^ x20 ;
  assign n1887 = x69 & n1327 ;
  assign n1913 = n1912 ^ n1887 ;
  assign n1886 = x71 & n1330 ;
  assign n1914 = n1913 ^ n1886 ;
  assign n1885 = ~n493 & n1331 ;
  assign n1915 = n1914 ^ n1885 ;
  assign n1917 = n1916 ^ n1915 ;
  assign n1882 = n1786 ^ n1777 ;
  assign n1883 = ~n1783 & n1882 ;
  assign n1884 = n1883 ^ n1786 ;
  assign n1918 = n1917 ^ n1884 ;
  assign n1919 = n1918 ^ x17 ;
  assign n1881 = x72 & n1050 ;
  assign n1920 = n1919 ^ n1881 ;
  assign n1880 = x74 & n1053 ;
  assign n1921 = n1920 ^ n1880 ;
  assign n1879 = n699 & n1054 ;
  assign n1922 = n1921 ^ n1879 ;
  assign n1924 = n1923 ^ n1922 ;
  assign n1928 = n1927 ^ n1924 ;
  assign n1929 = n1928 ^ x14 ;
  assign n1878 = x75 & n877 ;
  assign n1930 = n1929 ^ n1878 ;
  assign n1877 = x77 & n782 ;
  assign n1931 = n1930 ^ n1877 ;
  assign n1876 = n783 & ~n939 ;
  assign n1932 = n1931 ^ n1876 ;
  assign n1934 = n1933 ^ n1932 ;
  assign n1873 = n1803 ^ n1794 ;
  assign n1874 = ~n1800 & n1873 ;
  assign n1875 = n1874 ^ n1803 ;
  assign n1935 = n1934 ^ n1875 ;
  assign n1936 = n1935 ^ x11 ;
  assign n1872 = x78 & n647 ;
  assign n1937 = n1936 ^ n1872 ;
  assign n1871 = x80 & ~n572 ;
  assign n1938 = n1937 ^ n1871 ;
  assign n1870 = ~n573 & n1206 ;
  assign n1939 = n1938 ^ n1870 ;
  assign n1941 = n1940 ^ n1939 ;
  assign n1867 = n1813 ^ n1804 ;
  assign n1868 = ~n1810 & n1867 ;
  assign n1869 = n1868 ^ n1813 ;
  assign n1942 = n1941 ^ n1869 ;
  assign n1943 = n1942 ^ x8 ;
  assign n1866 = x81 & n446 ;
  assign n1944 = n1943 ^ n1866 ;
  assign n1865 = x83 & n383 ;
  assign n1945 = n1944 ^ n1865 ;
  assign n1864 = n384 & n1512 ;
  assign n1946 = n1945 ^ n1864 ;
  assign n1948 = n1947 ^ n1946 ;
  assign n1861 = n1823 ^ n1814 ;
  assign n1862 = ~n1820 & n1861 ;
  assign n1863 = n1862 ^ n1823 ;
  assign n1949 = n1948 ^ n1863 ;
  assign n1950 = n1949 ^ x5 ;
  assign n1860 = x84 & n234 ;
  assign n1951 = n1950 ^ n1860 ;
  assign n1859 = x86 & n230 ;
  assign n1952 = n1951 ^ n1859 ;
  assign n1857 = n1495 ^ x86 ;
  assign n1858 = n231 & n1857 ;
  assign n1953 = n1952 ^ n1858 ;
  assign n1955 = n1954 ^ n1953 ;
  assign n1959 = n1958 ^ n1955 ;
  assign n1841 = x88 ^ x87 ;
  assign n1843 = ~n1726 & n1841 ;
  assign n1845 = x89 ^ x1 ;
  assign n1844 = x89 ^ x2 ;
  assign n1846 = n1845 ^ n1844 ;
  assign n1847 = ~n1843 & n1846 ;
  assign n1848 = n1847 ^ n1845 ;
  assign n1960 = n1959 ^ n1848 ;
  assign n1852 = x2 & x87 ;
  assign n1853 = n1852 ^ x88 ;
  assign n1854 = ~x1 & n1853 ;
  assign n1849 = n1848 ^ n1727 ;
  assign n1855 = n1854 ^ n1849 ;
  assign n1856 = ~x0 & n1855 ;
  assign n1961 = n1960 ^ n1856 ;
  assign n1838 = n1836 ^ n1831 ;
  assign n1839 = ~n1833 & n1838 ;
  assign n1840 = n1839 ^ n1836 ;
  assign n1962 = n1961 ^ n1840 ;
  assign n2096 = n1959 ^ n1840 ;
  assign n2097 = n1961 & n2096 ;
  assign n2098 = n2097 ^ n1959 ;
  assign n2091 = x86 & n227 ;
  assign n2083 = n1942 ^ n1863 ;
  assign n2084 = n1948 & n2083 ;
  assign n2085 = n2084 ^ n1942 ;
  assign n2081 = x83 & n390 ;
  assign n2073 = n1935 ^ n1869 ;
  assign n2074 = n1941 & n2073 ;
  assign n2075 = n2074 ^ n1935 ;
  assign n2071 = x80 & n578 ;
  assign n2063 = n1928 ^ n1875 ;
  assign n2064 = n1934 & n2063 ;
  assign n2065 = n2064 ^ n1928 ;
  assign n2061 = x77 & n788 ;
  assign n2052 = n1911 ^ n1884 ;
  assign n2053 = n1917 & n2052 ;
  assign n2054 = n2053 ^ n1911 ;
  assign n2050 = x71 & n1335 ;
  assign n2039 = x67 & n1658 ;
  assign n2038 = x69 & n1661 ;
  assign n2040 = n2039 ^ n2038 ;
  assign n2041 = n2040 ^ x23 ;
  assign n2037 = ~n375 & n1662 ;
  assign n2042 = n2041 ^ n2037 ;
  assign n2036 = x68 & n1666 ;
  assign n2043 = n2042 ^ n2036 ;
  assign n2032 = x26 & ~n1767 ;
  assign n2033 = ~n1898 & n2032 ;
  assign n2034 = n2033 ^ x26 ;
  assign n2029 = x66 & n1766 ;
  assign n2016 = x26 ^ x25 ;
  assign n2021 = n1766 & ~n2016 ;
  assign n2022 = n2021 ^ n1766 ;
  assign n2025 = x65 & n2022 ;
  assign n1890 = x25 ^ x24 ;
  assign n2017 = ~n1766 & ~n1890 ;
  assign n2018 = n2016 & n2017 ;
  assign n2026 = n2025 ^ n2018 ;
  assign n2027 = ~x64 & n2026 ;
  assign n2028 = n2027 ^ n2018 ;
  assign n2030 = n2029 ^ n2028 ;
  assign n2014 = ~n1766 & n1890 ;
  assign n2015 = x65 & n2014 ;
  assign n2031 = n2030 ^ n2015 ;
  assign n2035 = n2034 ^ n2031 ;
  assign n2044 = n2043 ^ n2035 ;
  assign n2011 = n1910 ^ n1906 ;
  assign n2012 = ~n1907 & n2011 ;
  assign n2013 = n2012 ^ n1910 ;
  assign n2045 = n2044 ^ n2013 ;
  assign n2046 = n2045 ^ x20 ;
  assign n2010 = x70 & n1327 ;
  assign n2047 = n2046 ^ n2010 ;
  assign n2009 = x72 & n1330 ;
  assign n2048 = n2047 ^ n2009 ;
  assign n2008 = n556 & n1331 ;
  assign n2049 = n2048 ^ n2008 ;
  assign n2051 = n2050 ^ n2049 ;
  assign n2055 = n2054 ^ n2051 ;
  assign n1998 = x73 & n1050 ;
  assign n1997 = x75 & n1053 ;
  assign n1999 = n1998 ^ n1997 ;
  assign n2000 = n1999 ^ x17 ;
  assign n1996 = ~n774 & n1054 ;
  assign n2001 = n2000 ^ n1996 ;
  assign n1995 = x74 & n1058 ;
  assign n2002 = n2001 ^ n1995 ;
  assign n2003 = n2002 ^ n1927 ;
  assign n2004 = n2003 ^ n1918 ;
  assign n2005 = n2004 ^ n2002 ;
  assign n2006 = ~n1924 & n2005 ;
  assign n2007 = n2006 ^ n2003 ;
  assign n2056 = n2055 ^ n2007 ;
  assign n2057 = n2056 ^ x14 ;
  assign n1994 = x76 & n877 ;
  assign n2058 = n2057 ^ n1994 ;
  assign n1993 = x78 & n782 ;
  assign n2059 = n2058 ^ n1993 ;
  assign n1992 = n783 & ~n1025 ;
  assign n2060 = n2059 ^ n1992 ;
  assign n2062 = n2061 ^ n2060 ;
  assign n2066 = n2065 ^ n2062 ;
  assign n2067 = n2066 ^ x11 ;
  assign n1991 = x79 & n647 ;
  assign n2068 = n2067 ^ n1991 ;
  assign n1990 = x81 & ~n572 ;
  assign n2069 = n2068 ^ n1990 ;
  assign n1989 = ~n573 & n1305 ;
  assign n2070 = n2069 ^ n1989 ;
  assign n2072 = n2071 ^ n2070 ;
  assign n2076 = n2075 ^ n2072 ;
  assign n2077 = n2076 ^ x8 ;
  assign n1988 = x82 & n446 ;
  assign n2078 = n2077 ^ n1988 ;
  assign n1987 = x84 & n383 ;
  assign n2079 = n2078 ^ n1987 ;
  assign n1986 = n384 & n1624 ;
  assign n2080 = n2079 ^ n1986 ;
  assign n2082 = n2081 ^ n2080 ;
  assign n2086 = n2085 ^ n2082 ;
  assign n2087 = n2086 ^ x5 ;
  assign n1985 = x85 & n234 ;
  assign n2088 = n2087 ^ n1985 ;
  assign n1984 = x87 & n230 ;
  assign n2089 = n2088 ^ n1984 ;
  assign n1982 = n1610 ^ x87 ;
  assign n1983 = n231 & n1982 ;
  assign n2090 = n2089 ^ n1983 ;
  assign n2092 = n2091 ^ n2090 ;
  assign n1979 = n1958 ^ n1949 ;
  assign n1980 = ~n1955 & n1979 ;
  assign n1981 = n1980 ^ n1958 ;
  assign n2093 = n2092 ^ n1981 ;
  assign n1963 = x89 ^ x88 ;
  assign n1965 = ~n1843 & n1963 ;
  assign n1967 = x90 ^ x1 ;
  assign n1966 = x90 ^ x2 ;
  assign n1968 = n1967 ^ n1966 ;
  assign n1969 = ~n1965 & n1968 ;
  assign n1970 = n1969 ^ n1967 ;
  assign n2094 = n2093 ^ n1970 ;
  assign n1974 = x2 & x88 ;
  assign n1975 = n1974 ^ x89 ;
  assign n1976 = ~x1 & n1975 ;
  assign n1971 = n1970 ^ n1844 ;
  assign n1977 = n1976 ^ n1971 ;
  assign n1978 = ~x0 & n1977 ;
  assign n2095 = n2094 ^ n1978 ;
  assign n2099 = n2098 ^ n2095 ;
  assign n2223 = n2086 ^ n1981 ;
  assign n2224 = n2092 & n2223 ;
  assign n2225 = n2224 ^ n2086 ;
  assign n2221 = x87 & n227 ;
  assign n2214 = x84 & n390 ;
  assign n2207 = x81 & n578 ;
  assign n2200 = x78 & n788 ;
  assign n2193 = x75 & n1058 ;
  assign n2186 = x72 & n1335 ;
  assign n2178 = n2043 ^ n2013 ;
  assign n2179 = n2044 & n2178 ;
  assign n2180 = n2179 ^ n2043 ;
  assign n2172 = x68 & n1658 ;
  assign n2171 = x70 & n1661 ;
  assign n2173 = n2172 ^ n2171 ;
  assign n2174 = n2173 ^ x23 ;
  assign n2170 = ~n436 & n1662 ;
  assign n2175 = n2174 ^ n2170 ;
  assign n2169 = x69 & n1666 ;
  assign n2176 = n2175 ^ n2169 ;
  assign n2166 = ~n2031 & n2033 ;
  assign n2164 = x27 ^ x26 ;
  assign n2165 = x64 & n2164 ;
  assign n2167 = n2166 ^ n2165 ;
  assign n2160 = x65 & n2018 ;
  assign n2159 = x66 & n2014 ;
  assign n2161 = n2160 ^ n2159 ;
  assign n2162 = n2161 ^ x26 ;
  assign n2156 = ~n153 & ~n2016 ;
  assign n2157 = n2156 ^ n291 ;
  assign n2158 = n1766 & ~n2157 ;
  assign n2163 = n2162 ^ n2158 ;
  assign n2168 = n2167 ^ n2163 ;
  assign n2177 = n2176 ^ n2168 ;
  assign n2181 = n2180 ^ n2177 ;
  assign n2182 = n2181 ^ x20 ;
  assign n2152 = x71 & n1327 ;
  assign n2183 = n2182 ^ n2152 ;
  assign n2151 = x73 & n1330 ;
  assign n2184 = n2183 ^ n2151 ;
  assign n2150 = n633 & n1331 ;
  assign n2185 = n2184 ^ n2150 ;
  assign n2187 = n2186 ^ n2185 ;
  assign n2147 = n2054 ^ n2045 ;
  assign n2148 = ~n2051 & n2147 ;
  assign n2149 = n2148 ^ n2054 ;
  assign n2188 = n2187 ^ n2149 ;
  assign n2189 = n2188 ^ x17 ;
  assign n2146 = x74 & n1050 ;
  assign n2190 = n2189 ^ n2146 ;
  assign n2145 = x76 & n1053 ;
  assign n2191 = n2190 ^ n2145 ;
  assign n2144 = ~n853 & n1054 ;
  assign n2192 = n2191 ^ n2144 ;
  assign n2194 = n2193 ^ n2192 ;
  assign n2141 = n2055 ^ n2002 ;
  assign n2142 = n2007 & n2141 ;
  assign n2143 = n2142 ^ n2002 ;
  assign n2195 = n2194 ^ n2143 ;
  assign n2196 = n2195 ^ x14 ;
  assign n2140 = x77 & n877 ;
  assign n2197 = n2196 ^ n2140 ;
  assign n2139 = x79 & n782 ;
  assign n2198 = n2197 ^ n2139 ;
  assign n2138 = n783 & n1118 ;
  assign n2199 = n2198 ^ n2138 ;
  assign n2201 = n2200 ^ n2199 ;
  assign n2135 = n2065 ^ n2056 ;
  assign n2136 = ~n2062 & n2135 ;
  assign n2137 = n2136 ^ n2065 ;
  assign n2202 = n2201 ^ n2137 ;
  assign n2203 = n2202 ^ x11 ;
  assign n2134 = x80 & n647 ;
  assign n2204 = n2203 ^ n2134 ;
  assign n2133 = x82 & ~n572 ;
  assign n2205 = n2204 ^ n2133 ;
  assign n2132 = ~n573 & n1411 ;
  assign n2206 = n2205 ^ n2132 ;
  assign n2208 = n2207 ^ n2206 ;
  assign n2129 = n2075 ^ n2066 ;
  assign n2130 = ~n2072 & n2129 ;
  assign n2131 = n2130 ^ n2075 ;
  assign n2209 = n2208 ^ n2131 ;
  assign n2210 = n2209 ^ x8 ;
  assign n2128 = x83 & n446 ;
  assign n2211 = n2210 ^ n2128 ;
  assign n2127 = x85 & n383 ;
  assign n2212 = n2211 ^ n2127 ;
  assign n2126 = n384 & n1743 ;
  assign n2213 = n2212 ^ n2126 ;
  assign n2215 = n2214 ^ n2213 ;
  assign n2123 = n2085 ^ n2076 ;
  assign n2124 = ~n2082 & n2123 ;
  assign n2125 = n2124 ^ n2085 ;
  assign n2216 = n2215 ^ n2125 ;
  assign n2217 = n2216 ^ x5 ;
  assign n2122 = x86 & n234 ;
  assign n2218 = n2217 ^ n2122 ;
  assign n2121 = x88 & n230 ;
  assign n2219 = n2218 ^ n2121 ;
  assign n2119 = n1726 ^ x88 ;
  assign n2120 = n231 & n2119 ;
  assign n2220 = n2219 ^ n2120 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2226 = n2225 ^ n2222 ;
  assign n2103 = x90 ^ x89 ;
  assign n2105 = ~n1965 & n2103 ;
  assign n2107 = x91 ^ x1 ;
  assign n2106 = x91 ^ x2 ;
  assign n2108 = n2107 ^ n2106 ;
  assign n2109 = ~n2105 & n2108 ;
  assign n2110 = n2109 ^ n2107 ;
  assign n2227 = n2226 ^ n2110 ;
  assign n2114 = x2 & x89 ;
  assign n2115 = n2114 ^ x90 ;
  assign n2116 = ~x1 & n2115 ;
  assign n2111 = n2110 ^ n1966 ;
  assign n2117 = n2116 ^ n2111 ;
  assign n2118 = ~x0 & n2117 ;
  assign n2228 = n2227 ^ n2118 ;
  assign n2100 = n2098 ^ n2093 ;
  assign n2101 = ~n2095 & n2100 ;
  assign n2102 = n2101 ^ n2098 ;
  assign n2229 = n2228 ^ n2102 ;
  assign n2363 = n2226 ^ n2102 ;
  assign n2364 = n2228 & n2363 ;
  assign n2365 = n2364 ^ n2226 ;
  assign n2358 = x88 & n227 ;
  assign n2350 = n2209 ^ n2125 ;
  assign n2351 = n2215 & n2350 ;
  assign n2352 = n2351 ^ n2209 ;
  assign n2348 = x85 & n390 ;
  assign n2340 = n2202 ^ n2131 ;
  assign n2341 = n2208 & n2340 ;
  assign n2342 = n2341 ^ n2202 ;
  assign n2338 = x82 & n578 ;
  assign n2330 = n2195 ^ n2137 ;
  assign n2331 = n2201 & n2330 ;
  assign n2332 = n2331 ^ n2195 ;
  assign n2328 = x79 & n788 ;
  assign n2321 = x76 & n1058 ;
  assign n2313 = n2181 ^ n2149 ;
  assign n2314 = n2187 & n2313 ;
  assign n2315 = n2314 ^ n2181 ;
  assign n2311 = x73 & n1335 ;
  assign n2300 = x69 & n1658 ;
  assign n2299 = x71 & n1661 ;
  assign n2301 = n2300 ^ n2299 ;
  assign n2302 = n2301 ^ x23 ;
  assign n2298 = ~n493 & n1662 ;
  assign n2303 = n2302 ^ n2298 ;
  assign n2297 = x70 & n1666 ;
  assign n2304 = n2303 ^ n2297 ;
  assign n2293 = ~n2165 & ~n2166 ;
  assign n2294 = n2163 & n2293 ;
  assign n2295 = n2294 ^ n2163 ;
  assign n2287 = x66 & n2018 ;
  assign n2286 = x68 & n2021 ;
  assign n2288 = n2287 ^ n2286 ;
  assign n2289 = n2288 ^ x26 ;
  assign n2285 = ~n340 & n2022 ;
  assign n2290 = n2289 ^ n2285 ;
  assign n2284 = x67 & n2014 ;
  assign n2291 = n2290 ^ n2284 ;
  assign n2280 = x26 & x27 ;
  assign n2281 = n2280 ^ x28 ;
  assign n2282 = ~x64 & n2281 ;
  assign n2274 = x65 ^ x27 ;
  assign n2277 = x65 ^ x26 ;
  assign n2278 = ~n2274 & n2277 ;
  assign n2275 = x28 ^ x26 ;
  assign n2279 = n2278 ^ n2275 ;
  assign n2283 = n2282 ^ n2279 ;
  assign n2292 = n2291 ^ n2283 ;
  assign n2296 = n2295 ^ n2292 ;
  assign n2305 = n2304 ^ n2296 ;
  assign n2271 = n2180 ^ n2176 ;
  assign n2272 = ~n2177 & n2271 ;
  assign n2273 = n2272 ^ n2180 ;
  assign n2306 = n2305 ^ n2273 ;
  assign n2307 = n2306 ^ x20 ;
  assign n2270 = x72 & n1327 ;
  assign n2308 = n2307 ^ n2270 ;
  assign n2269 = x74 & n1330 ;
  assign n2309 = n2308 ^ n2269 ;
  assign n2268 = n699 & n1331 ;
  assign n2310 = n2309 ^ n2268 ;
  assign n2312 = n2311 ^ n2310 ;
  assign n2316 = n2315 ^ n2312 ;
  assign n2317 = n2316 ^ x17 ;
  assign n2267 = x75 & n1050 ;
  assign n2318 = n2317 ^ n2267 ;
  assign n2266 = x77 & n1053 ;
  assign n2319 = n2318 ^ n2266 ;
  assign n2265 = ~n939 & n1054 ;
  assign n2320 = n2319 ^ n2265 ;
  assign n2322 = n2321 ^ n2320 ;
  assign n2262 = n2188 ^ n2143 ;
  assign n2263 = n2194 & n2262 ;
  assign n2264 = n2263 ^ n2188 ;
  assign n2323 = n2322 ^ n2264 ;
  assign n2324 = n2323 ^ x14 ;
  assign n2261 = x78 & n877 ;
  assign n2325 = n2324 ^ n2261 ;
  assign n2260 = x80 & n782 ;
  assign n2326 = n2325 ^ n2260 ;
  assign n2259 = n783 & n1206 ;
  assign n2327 = n2326 ^ n2259 ;
  assign n2329 = n2328 ^ n2327 ;
  assign n2333 = n2332 ^ n2329 ;
  assign n2334 = n2333 ^ x11 ;
  assign n2258 = x81 & n647 ;
  assign n2335 = n2334 ^ n2258 ;
  assign n2257 = x83 & ~n572 ;
  assign n2336 = n2335 ^ n2257 ;
  assign n2256 = ~n573 & n1512 ;
  assign n2337 = n2336 ^ n2256 ;
  assign n2339 = n2338 ^ n2337 ;
  assign n2343 = n2342 ^ n2339 ;
  assign n2344 = n2343 ^ x8 ;
  assign n2255 = x84 & n446 ;
  assign n2345 = n2344 ^ n2255 ;
  assign n2254 = x86 & n383 ;
  assign n2346 = n2345 ^ n2254 ;
  assign n2253 = n384 & n1857 ;
  assign n2347 = n2346 ^ n2253 ;
  assign n2349 = n2348 ^ n2347 ;
  assign n2353 = n2352 ^ n2349 ;
  assign n2354 = n2353 ^ x5 ;
  assign n2252 = x87 & n234 ;
  assign n2355 = n2354 ^ n2252 ;
  assign n2251 = x89 & n230 ;
  assign n2356 = n2355 ^ n2251 ;
  assign n2249 = n1843 ^ x89 ;
  assign n2250 = n231 & n2249 ;
  assign n2357 = n2356 ^ n2250 ;
  assign n2359 = n2358 ^ n2357 ;
  assign n2246 = n2225 ^ n2216 ;
  assign n2247 = ~n2222 & n2246 ;
  assign n2248 = n2247 ^ n2225 ;
  assign n2360 = n2359 ^ n2248 ;
  assign n2230 = x91 ^ x90 ;
  assign n2232 = ~n2105 & n2230 ;
  assign n2234 = x92 ^ x1 ;
  assign n2233 = x92 ^ x2 ;
  assign n2235 = n2234 ^ n2233 ;
  assign n2236 = ~n2232 & n2235 ;
  assign n2237 = n2236 ^ n2234 ;
  assign n2361 = n2360 ^ n2237 ;
  assign n2241 = x2 & x90 ;
  assign n2242 = n2241 ^ x91 ;
  assign n2243 = ~n255 & n2242 ;
  assign n2238 = n2237 ^ n2106 ;
  assign n2244 = n2243 ^ n2238 ;
  assign n2245 = ~x0 & n2244 ;
  assign n2362 = n2361 ^ n2245 ;
  assign n2366 = n2365 ^ n2362 ;
  assign n2513 = n2353 ^ n2248 ;
  assign n2514 = n2359 & n2513 ;
  assign n2515 = n2514 ^ n2353 ;
  assign n2511 = x89 & n227 ;
  assign n2504 = x86 & n390 ;
  assign n2497 = x83 & n578 ;
  assign n2490 = x80 & n788 ;
  assign n2482 = n2316 ^ n2264 ;
  assign n2483 = n2322 & n2482 ;
  assign n2484 = n2483 ^ n2316 ;
  assign n2480 = x77 & n1058 ;
  assign n2473 = x74 & n1335 ;
  assign n2465 = n2304 ^ n2273 ;
  assign n2466 = n2305 & n2465 ;
  assign n2467 = n2466 ^ n2304 ;
  assign n2459 = x70 & n1658 ;
  assign n2458 = x72 & n1661 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2461 = n2460 ^ x23 ;
  assign n2457 = n556 & n1662 ;
  assign n2462 = n2461 ^ n2457 ;
  assign n2456 = x71 & n1666 ;
  assign n2463 = n2462 ^ n2456 ;
  assign n2453 = x68 & n2014 ;
  assign n2450 = x69 & n2021 ;
  assign n2448 = x67 & n2018 ;
  assign n2428 = x28 ^ x27 ;
  assign n2429 = ~n2164 & n2428 ;
  assign n2430 = x65 & n2429 ;
  assign n2421 = x29 ^ x28 ;
  assign n2422 = n2164 & ~n2421 ;
  assign n2423 = n2422 ^ n2164 ;
  assign n2426 = ~n150 & n2423 ;
  assign n2425 = x66 & n2164 ;
  assign n2427 = n2426 ^ n2425 ;
  assign n2431 = n2430 ^ n2427 ;
  assign n2442 = x29 & ~n2431 ;
  assign n2433 = ~n2165 & ~n2283 ;
  assign n2436 = x28 & x64 ;
  assign n2443 = n2436 ^ x64 ;
  assign n2444 = n2433 & ~n2443 ;
  assign n2445 = n2442 & n2444 ;
  assign n2432 = n2431 ^ x29 ;
  assign n2437 = n2280 & n2436 ;
  assign n2438 = n2437 ^ n2433 ;
  assign n2439 = ~n2431 & n2438 ;
  assign n2440 = n2439 ^ n2433 ;
  assign n2441 = ~n2432 & ~n2440 ;
  assign n2446 = n2445 ^ n2441 ;
  assign n2447 = n2446 ^ x26 ;
  assign n2449 = n2448 ^ n2447 ;
  assign n2451 = n2450 ^ n2449 ;
  assign n2420 = ~n375 & n2022 ;
  assign n2452 = n2451 ^ n2420 ;
  assign n2454 = n2453 ^ n2452 ;
  assign n2417 = n2295 ^ n2291 ;
  assign n2418 = ~n2292 & n2417 ;
  assign n2419 = n2418 ^ n2295 ;
  assign n2455 = n2454 ^ n2419 ;
  assign n2464 = n2463 ^ n2455 ;
  assign n2468 = n2467 ^ n2464 ;
  assign n2469 = n2468 ^ x20 ;
  assign n2416 = x73 & n1327 ;
  assign n2470 = n2469 ^ n2416 ;
  assign n2415 = x75 & n1330 ;
  assign n2471 = n2470 ^ n2415 ;
  assign n2414 = ~n774 & n1331 ;
  assign n2472 = n2471 ^ n2414 ;
  assign n2474 = n2473 ^ n2472 ;
  assign n2411 = n2315 ^ n2306 ;
  assign n2412 = ~n2312 & n2411 ;
  assign n2413 = n2412 ^ n2315 ;
  assign n2475 = n2474 ^ n2413 ;
  assign n2476 = n2475 ^ x17 ;
  assign n2410 = x76 & n1050 ;
  assign n2477 = n2476 ^ n2410 ;
  assign n2409 = x78 & n1053 ;
  assign n2478 = n2477 ^ n2409 ;
  assign n2408 = ~n1025 & n1054 ;
  assign n2479 = n2478 ^ n2408 ;
  assign n2481 = n2480 ^ n2479 ;
  assign n2485 = n2484 ^ n2481 ;
  assign n2486 = n2485 ^ x14 ;
  assign n2407 = x79 & n877 ;
  assign n2487 = n2486 ^ n2407 ;
  assign n2406 = x81 & n782 ;
  assign n2488 = n2487 ^ n2406 ;
  assign n2405 = n783 & n1305 ;
  assign n2489 = n2488 ^ n2405 ;
  assign n2491 = n2490 ^ n2489 ;
  assign n2402 = n2332 ^ n2323 ;
  assign n2403 = ~n2329 & n2402 ;
  assign n2404 = n2403 ^ n2332 ;
  assign n2492 = n2491 ^ n2404 ;
  assign n2493 = n2492 ^ x11 ;
  assign n2401 = x82 & n647 ;
  assign n2494 = n2493 ^ n2401 ;
  assign n2400 = x84 & ~n572 ;
  assign n2495 = n2494 ^ n2400 ;
  assign n2399 = ~n573 & n1624 ;
  assign n2496 = n2495 ^ n2399 ;
  assign n2498 = n2497 ^ n2496 ;
  assign n2396 = n2342 ^ n2333 ;
  assign n2397 = ~n2339 & n2396 ;
  assign n2398 = n2397 ^ n2342 ;
  assign n2499 = n2498 ^ n2398 ;
  assign n2500 = n2499 ^ x8 ;
  assign n2395 = x85 & n446 ;
  assign n2501 = n2500 ^ n2395 ;
  assign n2394 = x87 & n383 ;
  assign n2502 = n2501 ^ n2394 ;
  assign n2393 = n384 & n1982 ;
  assign n2503 = n2502 ^ n2393 ;
  assign n2505 = n2504 ^ n2503 ;
  assign n2390 = n2352 ^ n2343 ;
  assign n2391 = ~n2349 & n2390 ;
  assign n2392 = n2391 ^ n2352 ;
  assign n2506 = n2505 ^ n2392 ;
  assign n2507 = n2506 ^ x5 ;
  assign n2389 = x88 & n234 ;
  assign n2508 = n2507 ^ n2389 ;
  assign n2388 = x90 & n230 ;
  assign n2509 = n2508 ^ n2388 ;
  assign n2386 = n1965 ^ x90 ;
  assign n2387 = n231 & n2386 ;
  assign n2510 = n2509 ^ n2387 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2516 = n2515 ^ n2512 ;
  assign n2370 = x92 ^ x91 ;
  assign n2372 = ~n2232 & n2370 ;
  assign n2374 = x93 ^ x1 ;
  assign n2373 = x93 ^ x2 ;
  assign n2375 = n2374 ^ n2373 ;
  assign n2376 = ~n2372 & n2375 ;
  assign n2377 = n2376 ^ n2374 ;
  assign n2517 = n2516 ^ n2377 ;
  assign n2381 = x2 & x91 ;
  assign n2382 = n2381 ^ x92 ;
  assign n2383 = ~n255 & n2382 ;
  assign n2378 = n2377 ^ n2233 ;
  assign n2384 = n2383 ^ n2378 ;
  assign n2385 = ~x0 & n2384 ;
  assign n2518 = n2517 ^ n2385 ;
  assign n2367 = n2365 ^ n2360 ;
  assign n2368 = ~n2362 & n2367 ;
  assign n2369 = n2368 ^ n2365 ;
  assign n2519 = n2518 ^ n2369 ;
  assign n2661 = n2516 ^ n2369 ;
  assign n2662 = ~n2518 & ~n2661 ;
  assign n2663 = n2662 ^ n2516 ;
  assign n2656 = x90 & n227 ;
  assign n2648 = n2499 ^ n2392 ;
  assign n2649 = ~n2505 & ~n2648 ;
  assign n2650 = n2649 ^ n2499 ;
  assign n2646 = x87 & n390 ;
  assign n2638 = n2492 ^ n2398 ;
  assign n2639 = ~n2498 & ~n2638 ;
  assign n2640 = n2639 ^ n2492 ;
  assign n2636 = x84 & n578 ;
  assign n2628 = n2485 ^ n2404 ;
  assign n2629 = ~n2491 & ~n2628 ;
  assign n2630 = n2629 ^ n2485 ;
  assign n2626 = x81 & n788 ;
  assign n2619 = x78 & n1058 ;
  assign n2611 = n2468 ^ n2413 ;
  assign n2612 = ~n2474 & ~n2611 ;
  assign n2613 = n2612 ^ n2468 ;
  assign n2609 = x75 & n1335 ;
  assign n2602 = x72 & n1666 ;
  assign n2591 = x68 & n2018 ;
  assign n2590 = x70 & n2021 ;
  assign n2592 = n2591 ^ n2590 ;
  assign n2593 = n2592 ^ x26 ;
  assign n2589 = ~n436 & n2022 ;
  assign n2594 = n2593 ^ n2589 ;
  assign n2588 = x69 & n2014 ;
  assign n2595 = n2594 ^ n2588 ;
  assign n2579 = x29 ^ x27 ;
  assign n2580 = ~n2164 & n2579 ;
  assign n2581 = n2421 & n2580 ;
  assign n2582 = x65 & n2581 ;
  assign n2578 = x67 & n2422 ;
  assign n2583 = n2582 ^ n2578 ;
  assign n2584 = n2583 ^ x29 ;
  assign n2577 = ~n291 & n2423 ;
  assign n2585 = n2584 ^ n2577 ;
  assign n2576 = x66 & n2429 ;
  assign n2586 = n2585 ^ n2576 ;
  assign n2573 = x30 ^ x29 ;
  assign n2574 = x64 & n2573 ;
  assign n2575 = n2574 ^ n2445 ;
  assign n2587 = n2586 ^ n2575 ;
  assign n2596 = n2595 ^ n2587 ;
  assign n2570 = n2446 ^ n2419 ;
  assign n2571 = n2454 & ~n2570 ;
  assign n2572 = n2571 ^ n2419 ;
  assign n2597 = n2596 ^ n2572 ;
  assign n2598 = n2597 ^ x23 ;
  assign n2569 = x71 & n1658 ;
  assign n2599 = n2598 ^ n2569 ;
  assign n2568 = x73 & n1661 ;
  assign n2600 = n2599 ^ n2568 ;
  assign n2567 = n633 & n1662 ;
  assign n2601 = n2600 ^ n2567 ;
  assign n2603 = n2602 ^ n2601 ;
  assign n2564 = n2467 ^ n2463 ;
  assign n2565 = n2464 & n2564 ;
  assign n2566 = n2565 ^ n2467 ;
  assign n2604 = n2603 ^ n2566 ;
  assign n2605 = n2604 ^ x20 ;
  assign n2563 = x74 & n1327 ;
  assign n2606 = n2605 ^ n2563 ;
  assign n2562 = x76 & n1330 ;
  assign n2607 = n2606 ^ n2562 ;
  assign n2561 = ~n853 & n1331 ;
  assign n2608 = n2607 ^ n2561 ;
  assign n2610 = n2609 ^ n2608 ;
  assign n2614 = n2613 ^ n2610 ;
  assign n2615 = n2614 ^ x17 ;
  assign n2560 = x77 & n1050 ;
  assign n2616 = n2615 ^ n2560 ;
  assign n2559 = x79 & n1053 ;
  assign n2617 = n2616 ^ n2559 ;
  assign n2558 = n1054 & n1118 ;
  assign n2618 = n2617 ^ n2558 ;
  assign n2620 = n2619 ^ n2618 ;
  assign n2555 = n2484 ^ n2475 ;
  assign n2556 = n2481 & ~n2555 ;
  assign n2557 = n2556 ^ n2484 ;
  assign n2621 = n2620 ^ n2557 ;
  assign n2622 = n2621 ^ x14 ;
  assign n2554 = x80 & n877 ;
  assign n2623 = n2622 ^ n2554 ;
  assign n2553 = x82 & n782 ;
  assign n2624 = n2623 ^ n2553 ;
  assign n2552 = n783 & n1411 ;
  assign n2625 = n2624 ^ n2552 ;
  assign n2627 = n2626 ^ n2625 ;
  assign n2631 = n2630 ^ n2627 ;
  assign n2632 = n2631 ^ x11 ;
  assign n2551 = x83 & n647 ;
  assign n2633 = n2632 ^ n2551 ;
  assign n2550 = x85 & ~n572 ;
  assign n2634 = n2633 ^ n2550 ;
  assign n2549 = ~n573 & n1743 ;
  assign n2635 = n2634 ^ n2549 ;
  assign n2637 = n2636 ^ n2635 ;
  assign n2641 = n2640 ^ n2637 ;
  assign n2642 = n2641 ^ x8 ;
  assign n2548 = x86 & n446 ;
  assign n2643 = n2642 ^ n2548 ;
  assign n2547 = x88 & n383 ;
  assign n2644 = n2643 ^ n2547 ;
  assign n2546 = n384 & n2119 ;
  assign n2645 = n2644 ^ n2546 ;
  assign n2647 = n2646 ^ n2645 ;
  assign n2651 = n2650 ^ n2647 ;
  assign n2652 = n2651 ^ x5 ;
  assign n2545 = x89 & n234 ;
  assign n2653 = n2652 ^ n2545 ;
  assign n2544 = x91 & n230 ;
  assign n2654 = n2653 ^ n2544 ;
  assign n2542 = n2105 ^ x91 ;
  assign n2543 = n231 & n2542 ;
  assign n2655 = n2654 ^ n2543 ;
  assign n2657 = n2656 ^ n2655 ;
  assign n2539 = n2515 ^ n2506 ;
  assign n2540 = n2512 & ~n2539 ;
  assign n2541 = n2540 ^ n2515 ;
  assign n2658 = n2657 ^ n2541 ;
  assign n2522 = x93 ^ x91 ;
  assign n2520 = x93 ^ x92 ;
  assign n2523 = ~n2232 & n2520 ;
  assign n2524 = ~n2522 & n2523 ;
  assign n2525 = n2524 ^ n2520 ;
  assign n2527 = x94 ^ x1 ;
  assign n2526 = x94 ^ x2 ;
  assign n2528 = n2527 ^ n2526 ;
  assign n2529 = ~n2525 & n2528 ;
  assign n2530 = n2529 ^ n2527 ;
  assign n2659 = n2658 ^ n2530 ;
  assign n2534 = x2 & x92 ;
  assign n2535 = n2534 ^ x93 ;
  assign n2536 = ~x1 & n2535 ;
  assign n2531 = n2530 ^ n2373 ;
  assign n2537 = n2536 ^ n2531 ;
  assign n2538 = ~x0 & n2537 ;
  assign n2660 = n2659 ^ n2538 ;
  assign n2664 = n2663 ^ n2660 ;
  assign n2810 = n2651 ^ n2541 ;
  assign n2811 = n2657 & n2810 ;
  assign n2812 = n2811 ^ n2651 ;
  assign n2808 = x91 & n227 ;
  assign n2801 = x88 & n390 ;
  assign n2794 = x85 & n578 ;
  assign n2787 = x82 & n788 ;
  assign n2779 = n2614 ^ n2557 ;
  assign n2780 = ~n2620 & ~n2779 ;
  assign n2781 = n2780 ^ n2614 ;
  assign n2777 = x79 & n1058 ;
  assign n2770 = x76 & n1335 ;
  assign n2762 = n2597 ^ n2566 ;
  assign n2763 = n2603 & n2762 ;
  assign n2764 = n2763 ^ n2597 ;
  assign n2760 = x73 & n1666 ;
  assign n2751 = ~n2445 & n2586 ;
  assign n2752 = ~n2574 & n2751 ;
  assign n2753 = n2752 ^ n2586 ;
  assign n2745 = x66 & n2581 ;
  assign n2744 = x68 & n2422 ;
  assign n2746 = n2745 ^ n2744 ;
  assign n2747 = n2746 ^ x29 ;
  assign n2743 = ~n340 & n2423 ;
  assign n2748 = n2747 ^ n2743 ;
  assign n2742 = x67 & n2429 ;
  assign n2749 = n2748 ^ n2742 ;
  assign n2737 = ~x29 & ~x30 ;
  assign n2738 = n2737 ^ n2573 ;
  assign n2739 = n2738 ^ x31 ;
  assign n2740 = ~x64 & ~n2739 ;
  assign n2731 = x65 ^ x30 ;
  assign n2734 = x65 ^ x29 ;
  assign n2735 = ~n2731 & n2734 ;
  assign n2732 = x31 ^ x29 ;
  assign n2736 = n2735 ^ n2732 ;
  assign n2741 = n2740 ^ n2736 ;
  assign n2750 = n2749 ^ n2741 ;
  assign n2754 = n2753 ^ n2750 ;
  assign n2721 = x69 & n2018 ;
  assign n2720 = x71 & n2021 ;
  assign n2722 = n2721 ^ n2720 ;
  assign n2723 = n2722 ^ x26 ;
  assign n2719 = ~n493 & n2022 ;
  assign n2724 = n2723 ^ n2719 ;
  assign n2718 = x70 & n2014 ;
  assign n2725 = n2724 ^ n2718 ;
  assign n2726 = n2725 ^ n2595 ;
  assign n2727 = n2726 ^ n2572 ;
  assign n2728 = n2727 ^ n2725 ;
  assign n2729 = n2596 & n2728 ;
  assign n2730 = n2729 ^ n2726 ;
  assign n2755 = n2754 ^ n2730 ;
  assign n2756 = n2755 ^ x23 ;
  assign n2717 = x72 & n1658 ;
  assign n2757 = n2756 ^ n2717 ;
  assign n2716 = x74 & n1661 ;
  assign n2758 = n2757 ^ n2716 ;
  assign n2715 = n699 & n1662 ;
  assign n2759 = n2758 ^ n2715 ;
  assign n2761 = n2760 ^ n2759 ;
  assign n2765 = n2764 ^ n2761 ;
  assign n2766 = n2765 ^ x20 ;
  assign n2714 = x75 & n1327 ;
  assign n2767 = n2766 ^ n2714 ;
  assign n2713 = x77 & n1330 ;
  assign n2768 = n2767 ^ n2713 ;
  assign n2712 = ~n939 & n1331 ;
  assign n2769 = n2768 ^ n2712 ;
  assign n2771 = n2770 ^ n2769 ;
  assign n2709 = n2613 ^ n2604 ;
  assign n2710 = ~n2610 & ~n2709 ;
  assign n2711 = n2710 ^ n2613 ;
  assign n2772 = n2771 ^ n2711 ;
  assign n2773 = n2772 ^ x17 ;
  assign n2708 = x78 & n1050 ;
  assign n2774 = n2773 ^ n2708 ;
  assign n2707 = x80 & n1053 ;
  assign n2775 = n2774 ^ n2707 ;
  assign n2706 = n1054 & n1206 ;
  assign n2776 = n2775 ^ n2706 ;
  assign n2778 = n2777 ^ n2776 ;
  assign n2782 = n2781 ^ n2778 ;
  assign n2783 = n2782 ^ x14 ;
  assign n2705 = x81 & n877 ;
  assign n2784 = n2783 ^ n2705 ;
  assign n2704 = x83 & n782 ;
  assign n2785 = n2784 ^ n2704 ;
  assign n2703 = n783 & n1512 ;
  assign n2786 = n2785 ^ n2703 ;
  assign n2788 = n2787 ^ n2786 ;
  assign n2700 = n2630 ^ n2621 ;
  assign n2701 = n2627 & n2700 ;
  assign n2702 = n2701 ^ n2630 ;
  assign n2789 = n2788 ^ n2702 ;
  assign n2790 = n2789 ^ x11 ;
  assign n2699 = x84 & n647 ;
  assign n2791 = n2790 ^ n2699 ;
  assign n2698 = x86 & ~n572 ;
  assign n2792 = n2791 ^ n2698 ;
  assign n2697 = ~n573 & n1857 ;
  assign n2793 = n2792 ^ n2697 ;
  assign n2795 = n2794 ^ n2793 ;
  assign n2694 = n2640 ^ n2631 ;
  assign n2695 = ~n2637 & ~n2694 ;
  assign n2696 = n2695 ^ n2640 ;
  assign n2796 = n2795 ^ n2696 ;
  assign n2797 = n2796 ^ x8 ;
  assign n2693 = x87 & n446 ;
  assign n2798 = n2797 ^ n2693 ;
  assign n2692 = x89 & n383 ;
  assign n2799 = n2798 ^ n2692 ;
  assign n2691 = n384 & n2249 ;
  assign n2800 = n2799 ^ n2691 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2688 = n2650 ^ n2641 ;
  assign n2689 = n2647 & n2688 ;
  assign n2690 = n2689 ^ n2650 ;
  assign n2803 = n2802 ^ n2690 ;
  assign n2804 = n2803 ^ x5 ;
  assign n2687 = x90 & n234 ;
  assign n2805 = n2804 ^ n2687 ;
  assign n2686 = x92 & n230 ;
  assign n2806 = n2805 ^ n2686 ;
  assign n2684 = n2232 ^ x92 ;
  assign n2685 = n231 & n2684 ;
  assign n2807 = n2806 ^ n2685 ;
  assign n2809 = n2808 ^ n2807 ;
  assign n2813 = n2812 ^ n2809 ;
  assign n2668 = x94 ^ x93 ;
  assign n2670 = ~n2525 & n2668 ;
  assign n2672 = x95 ^ x1 ;
  assign n2671 = x95 ^ x2 ;
  assign n2673 = n2672 ^ n2671 ;
  assign n2674 = ~n2670 & n2673 ;
  assign n2675 = n2674 ^ n2672 ;
  assign n2814 = n2813 ^ n2675 ;
  assign n2679 = x2 & x93 ;
  assign n2680 = n2679 ^ x94 ;
  assign n2681 = ~n255 & n2680 ;
  assign n2676 = n2675 ^ n2526 ;
  assign n2682 = n2681 ^ n2676 ;
  assign n2683 = ~x0 & n2682 ;
  assign n2815 = n2814 ^ n2683 ;
  assign n2665 = n2663 ^ n2658 ;
  assign n2666 = ~n2660 & ~n2665 ;
  assign n2667 = n2666 ^ n2663 ;
  assign n2816 = n2815 ^ n2667 ;
  assign n2971 = n2813 ^ n2667 ;
  assign n2972 = ~n2815 & n2971 ;
  assign n2973 = n2972 ^ n2813 ;
  assign n2966 = x92 & n227 ;
  assign n2958 = n2796 ^ n2690 ;
  assign n2959 = n2802 & ~n2958 ;
  assign n2960 = n2959 ^ n2796 ;
  assign n2956 = x89 & n390 ;
  assign n2948 = n2789 ^ n2696 ;
  assign n2949 = ~n2795 & n2948 ;
  assign n2950 = n2949 ^ n2789 ;
  assign n2946 = x86 & n578 ;
  assign n2938 = n2782 ^ n2702 ;
  assign n2939 = n2788 & ~n2938 ;
  assign n2940 = n2939 ^ n2782 ;
  assign n2936 = x83 & n788 ;
  assign n2929 = x80 & n1058 ;
  assign n2921 = n2765 ^ n2711 ;
  assign n2922 = n2771 & ~n2921 ;
  assign n2923 = n2922 ^ n2765 ;
  assign n2919 = x77 & n1335 ;
  assign n2912 = x74 & n1666 ;
  assign n2905 = x71 & n2014 ;
  assign n2898 = x68 & n2429 ;
  assign n2891 = x32 & ~n2574 ;
  assign n2892 = ~n2741 & n2891 ;
  assign n2876 = x31 ^ x30 ;
  assign n2887 = ~n2573 & n2876 ;
  assign n2888 = x65 & n2887 ;
  assign n2877 = x32 ^ x31 ;
  assign n2882 = n2573 & ~n2877 ;
  assign n2883 = n2882 ^ n2573 ;
  assign n2884 = ~n150 & n2883 ;
  assign n2881 = x66 & n2573 ;
  assign n2885 = n2884 ^ n2881 ;
  assign n2886 = n2885 ^ x32 ;
  assign n2889 = n2888 ^ n2886 ;
  assign n2878 = ~n2573 & n2877 ;
  assign n2879 = ~n2876 & n2878 ;
  assign n2880 = x64 & n2879 ;
  assign n2890 = n2889 ^ n2880 ;
  assign n2893 = n2892 ^ n2890 ;
  assign n2894 = n2893 ^ x29 ;
  assign n2875 = x67 & n2581 ;
  assign n2895 = n2894 ^ n2875 ;
  assign n2874 = x69 & n2422 ;
  assign n2896 = n2895 ^ n2874 ;
  assign n2873 = ~n375 & n2423 ;
  assign n2897 = n2896 ^ n2873 ;
  assign n2899 = n2898 ^ n2897 ;
  assign n2870 = n2753 ^ n2749 ;
  assign n2871 = ~n2750 & n2870 ;
  assign n2872 = n2871 ^ n2753 ;
  assign n2900 = n2899 ^ n2872 ;
  assign n2901 = n2900 ^ x26 ;
  assign n2869 = x70 & n2018 ;
  assign n2902 = n2901 ^ n2869 ;
  assign n2868 = x72 & n2021 ;
  assign n2903 = n2902 ^ n2868 ;
  assign n2867 = n556 & n2022 ;
  assign n2904 = n2903 ^ n2867 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n2864 = n2754 ^ n2725 ;
  assign n2865 = n2730 & n2864 ;
  assign n2866 = n2865 ^ n2725 ;
  assign n2907 = n2906 ^ n2866 ;
  assign n2908 = n2907 ^ x23 ;
  assign n2863 = x73 & n1658 ;
  assign n2909 = n2908 ^ n2863 ;
  assign n2862 = x75 & n1661 ;
  assign n2910 = n2909 ^ n2862 ;
  assign n2861 = ~n774 & n1662 ;
  assign n2911 = n2910 ^ n2861 ;
  assign n2913 = n2912 ^ n2911 ;
  assign n2858 = n2764 ^ n2755 ;
  assign n2859 = ~n2761 & n2858 ;
  assign n2860 = n2859 ^ n2764 ;
  assign n2914 = n2913 ^ n2860 ;
  assign n2915 = n2914 ^ x20 ;
  assign n2857 = x76 & n1327 ;
  assign n2916 = n2915 ^ n2857 ;
  assign n2856 = x78 & n1330 ;
  assign n2917 = n2916 ^ n2856 ;
  assign n2855 = ~n1025 & n1331 ;
  assign n2918 = n2917 ^ n2855 ;
  assign n2920 = n2919 ^ n2918 ;
  assign n2924 = n2923 ^ n2920 ;
  assign n2925 = n2924 ^ x17 ;
  assign n2854 = x79 & n1050 ;
  assign n2926 = n2925 ^ n2854 ;
  assign n2853 = x81 & n1053 ;
  assign n2927 = n2926 ^ n2853 ;
  assign n2852 = n1054 & n1305 ;
  assign n2928 = n2927 ^ n2852 ;
  assign n2930 = n2929 ^ n2928 ;
  assign n2849 = n2781 ^ n2772 ;
  assign n2850 = n2778 & n2849 ;
  assign n2851 = n2850 ^ n2781 ;
  assign n2931 = n2930 ^ n2851 ;
  assign n2932 = n2931 ^ x14 ;
  assign n2848 = x82 & n877 ;
  assign n2933 = n2932 ^ n2848 ;
  assign n2847 = x84 & n782 ;
  assign n2934 = n2933 ^ n2847 ;
  assign n2846 = n783 & n1624 ;
  assign n2935 = n2934 ^ n2846 ;
  assign n2937 = n2936 ^ n2935 ;
  assign n2941 = n2940 ^ n2937 ;
  assign n2942 = n2941 ^ x11 ;
  assign n2845 = x85 & n647 ;
  assign n2943 = n2942 ^ n2845 ;
  assign n2844 = x87 & ~n572 ;
  assign n2944 = n2943 ^ n2844 ;
  assign n2843 = ~n573 & n1982 ;
  assign n2945 = n2944 ^ n2843 ;
  assign n2947 = n2946 ^ n2945 ;
  assign n2951 = n2950 ^ n2947 ;
  assign n2952 = n2951 ^ x8 ;
  assign n2842 = x88 & n446 ;
  assign n2953 = n2952 ^ n2842 ;
  assign n2841 = x90 & n383 ;
  assign n2954 = n2953 ^ n2841 ;
  assign n2840 = n384 & n2386 ;
  assign n2955 = n2954 ^ n2840 ;
  assign n2957 = n2956 ^ n2955 ;
  assign n2961 = n2960 ^ n2957 ;
  assign n2962 = n2961 ^ x5 ;
  assign n2839 = x91 & n234 ;
  assign n2963 = n2962 ^ n2839 ;
  assign n2838 = x93 & n230 ;
  assign n2964 = n2963 ^ n2838 ;
  assign n2836 = n2372 ^ x93 ;
  assign n2837 = n231 & n2836 ;
  assign n2965 = n2964 ^ n2837 ;
  assign n2967 = n2966 ^ n2965 ;
  assign n2833 = n2812 ^ n2803 ;
  assign n2834 = n2809 & ~n2833 ;
  assign n2835 = n2834 ^ n2812 ;
  assign n2968 = n2967 ^ n2835 ;
  assign n2817 = x95 ^ x94 ;
  assign n2819 = ~n2670 & n2817 ;
  assign n2821 = x96 ^ x1 ;
  assign n2820 = x96 ^ x2 ;
  assign n2822 = n2821 ^ n2820 ;
  assign n2823 = ~n2819 & n2822 ;
  assign n2824 = n2823 ^ n2821 ;
  assign n2969 = n2968 ^ n2824 ;
  assign n2828 = x2 & x94 ;
  assign n2829 = n2828 ^ x95 ;
  assign n2830 = ~x1 & n2829 ;
  assign n2825 = n2824 ^ n2671 ;
  assign n2831 = n2830 ^ n2825 ;
  assign n2832 = ~x0 & n2831 ;
  assign n2970 = n2969 ^ n2832 ;
  assign n2974 = n2973 ^ n2970 ;
  assign n3124 = n2961 ^ n2835 ;
  assign n3125 = n2967 & n3124 ;
  assign n3126 = n3125 ^ n2961 ;
  assign n3122 = x93 & n227 ;
  assign n3115 = x90 & n390 ;
  assign n3108 = x87 & n578 ;
  assign n3101 = x84 & n788 ;
  assign n3093 = n2924 ^ n2851 ;
  assign n3094 = n2930 & ~n3093 ;
  assign n3095 = n3094 ^ n2924 ;
  assign n3091 = x81 & n1058 ;
  assign n3084 = x78 & n1335 ;
  assign n3076 = n2907 ^ n2860 ;
  assign n3077 = n2913 & n3076 ;
  assign n3078 = n3077 ^ n2907 ;
  assign n3074 = x75 & n1666 ;
  assign n3067 = x72 & n2014 ;
  assign n3059 = n2893 ^ n2872 ;
  assign n3060 = n2899 & n3059 ;
  assign n3061 = n3060 ^ n2893 ;
  assign n3057 = x69 & n2429 ;
  assign n3046 = x65 & n2879 ;
  assign n3045 = x67 & n2882 ;
  assign n3047 = n3046 ^ n3045 ;
  assign n3048 = n3047 ^ x32 ;
  assign n3044 = ~n291 & n2883 ;
  assign n3049 = n3048 ^ n3044 ;
  assign n3043 = x66 & n2887 ;
  assign n3050 = n3049 ^ n3043 ;
  assign n3041 = x33 ^ x32 ;
  assign n3042 = x64 & n3041 ;
  assign n3051 = n3050 ^ n3042 ;
  assign n3040 = n2890 & n2892 ;
  assign n3052 = n3051 ^ n3040 ;
  assign n3053 = n3052 ^ x29 ;
  assign n3039 = x68 & n2581 ;
  assign n3054 = n3053 ^ n3039 ;
  assign n3038 = x70 & n2422 ;
  assign n3055 = n3054 ^ n3038 ;
  assign n3037 = ~n436 & n2423 ;
  assign n3056 = n3055 ^ n3037 ;
  assign n3058 = n3057 ^ n3056 ;
  assign n3062 = n3061 ^ n3058 ;
  assign n3063 = n3062 ^ x26 ;
  assign n3036 = x71 & n2018 ;
  assign n3064 = n3063 ^ n3036 ;
  assign n3035 = x73 & n2021 ;
  assign n3065 = n3064 ^ n3035 ;
  assign n3034 = n633 & n2022 ;
  assign n3066 = n3065 ^ n3034 ;
  assign n3068 = n3067 ^ n3066 ;
  assign n3031 = n2900 ^ n2866 ;
  assign n3032 = n2906 & n3031 ;
  assign n3033 = n3032 ^ n2900 ;
  assign n3069 = n3068 ^ n3033 ;
  assign n3070 = n3069 ^ x23 ;
  assign n3030 = x74 & n1658 ;
  assign n3071 = n3070 ^ n3030 ;
  assign n3029 = x76 & n1661 ;
  assign n3072 = n3071 ^ n3029 ;
  assign n3028 = ~n853 & n1662 ;
  assign n3073 = n3072 ^ n3028 ;
  assign n3075 = n3074 ^ n3073 ;
  assign n3079 = n3078 ^ n3075 ;
  assign n3080 = n3079 ^ x20 ;
  assign n3027 = x77 & n1327 ;
  assign n3081 = n3080 ^ n3027 ;
  assign n3026 = x79 & n1330 ;
  assign n3082 = n3081 ^ n3026 ;
  assign n3025 = n1118 & n1331 ;
  assign n3083 = n3082 ^ n3025 ;
  assign n3085 = n3084 ^ n3083 ;
  assign n3022 = n2923 ^ n2914 ;
  assign n3023 = ~n2920 & n3022 ;
  assign n3024 = n3023 ^ n2923 ;
  assign n3086 = n3085 ^ n3024 ;
  assign n3087 = n3086 ^ x17 ;
  assign n3021 = x80 & n1050 ;
  assign n3088 = n3087 ^ n3021 ;
  assign n3020 = x82 & n1053 ;
  assign n3089 = n3088 ^ n3020 ;
  assign n3019 = n1054 & n1411 ;
  assign n3090 = n3089 ^ n3019 ;
  assign n3092 = n3091 ^ n3090 ;
  assign n3096 = n3095 ^ n3092 ;
  assign n3097 = n3096 ^ x14 ;
  assign n3018 = x83 & n877 ;
  assign n3098 = n3097 ^ n3018 ;
  assign n3017 = x85 & n782 ;
  assign n3099 = n3098 ^ n3017 ;
  assign n3016 = n783 & n1743 ;
  assign n3100 = n3099 ^ n3016 ;
  assign n3102 = n3101 ^ n3100 ;
  assign n3013 = n2940 ^ n2931 ;
  assign n3014 = n2937 & ~n3013 ;
  assign n3015 = n3014 ^ n2940 ;
  assign n3103 = n3102 ^ n3015 ;
  assign n3104 = n3103 ^ x11 ;
  assign n3012 = x86 & n647 ;
  assign n3105 = n3104 ^ n3012 ;
  assign n3011 = x88 & ~n572 ;
  assign n3106 = n3105 ^ n3011 ;
  assign n3010 = ~n573 & n2119 ;
  assign n3107 = n3106 ^ n3010 ;
  assign n3109 = n3108 ^ n3107 ;
  assign n3007 = n2950 ^ n2941 ;
  assign n3008 = n2947 & n3007 ;
  assign n3009 = n3008 ^ n2950 ;
  assign n3110 = n3109 ^ n3009 ;
  assign n3111 = n3110 ^ x8 ;
  assign n3006 = x89 & n446 ;
  assign n3112 = n3111 ^ n3006 ;
  assign n3005 = x91 & n383 ;
  assign n3113 = n3112 ^ n3005 ;
  assign n3004 = n384 & n2542 ;
  assign n3114 = n3113 ^ n3004 ;
  assign n3116 = n3115 ^ n3114 ;
  assign n3001 = n2960 ^ n2951 ;
  assign n3002 = ~n2957 & n3001 ;
  assign n3003 = n3002 ^ n2960 ;
  assign n3117 = n3116 ^ n3003 ;
  assign n3118 = n3117 ^ x5 ;
  assign n3000 = x92 & n234 ;
  assign n3119 = n3118 ^ n3000 ;
  assign n2999 = x94 & n230 ;
  assign n3120 = n3119 ^ n2999 ;
  assign n2997 = n2525 ^ x94 ;
  assign n2998 = n231 & n2997 ;
  assign n3121 = n3120 ^ n2998 ;
  assign n3123 = n3122 ^ n3121 ;
  assign n3127 = n3126 ^ n3123 ;
  assign n2980 = x96 ^ x94 ;
  assign n2978 = x96 ^ x95 ;
  assign n2981 = ~n2670 & n2978 ;
  assign n2982 = ~n2980 & n2981 ;
  assign n2983 = n2982 ^ n2978 ;
  assign n2985 = x97 ^ x1 ;
  assign n2984 = x97 ^ x2 ;
  assign n2986 = n2985 ^ n2984 ;
  assign n2987 = ~n2983 & n2986 ;
  assign n2988 = n2987 ^ n2985 ;
  assign n3128 = n3127 ^ n2988 ;
  assign n2992 = x2 & x95 ;
  assign n2993 = n2992 ^ x96 ;
  assign n2994 = ~x1 & n2993 ;
  assign n2989 = n2988 ^ n2820 ;
  assign n2995 = n2994 ^ n2989 ;
  assign n2996 = ~x0 & n2995 ;
  assign n3129 = n3128 ^ n2996 ;
  assign n2975 = n2973 ^ n2968 ;
  assign n2976 = ~n2970 & ~n2975 ;
  assign n2977 = n2976 ^ n2973 ;
  assign n3130 = n3129 ^ n2977 ;
  assign n3300 = n3127 ^ n2977 ;
  assign n3301 = ~n3129 & n3300 ;
  assign n3302 = n3301 ^ n3127 ;
  assign n3295 = x94 & n227 ;
  assign n3287 = n3110 ^ n3003 ;
  assign n3288 = ~n3116 & ~n3287 ;
  assign n3289 = n3288 ^ n3110 ;
  assign n3285 = x91 & n390 ;
  assign n3277 = n3103 ^ n3009 ;
  assign n3278 = n3109 & ~n3277 ;
  assign n3279 = n3278 ^ n3103 ;
  assign n3275 = x88 & n578 ;
  assign n3267 = n3096 ^ n3015 ;
  assign n3268 = n3102 & n3267 ;
  assign n3269 = n3268 ^ n3096 ;
  assign n3265 = x85 & n788 ;
  assign n3258 = x82 & n1058 ;
  assign n3250 = n3079 ^ n3024 ;
  assign n3251 = n3085 & n3250 ;
  assign n3252 = n3251 ^ n3079 ;
  assign n3248 = x79 & n1335 ;
  assign n3241 = x76 & n1666 ;
  assign n3233 = n3062 ^ n3033 ;
  assign n3234 = n3068 & n3233 ;
  assign n3235 = n3234 ^ n3062 ;
  assign n3231 = x73 & n2014 ;
  assign n3224 = x70 & n2429 ;
  assign n3216 = ~n3042 & n3050 ;
  assign n3217 = ~n3040 & n3216 ;
  assign n3218 = n3217 ^ n3050 ;
  assign n3210 = x32 & x33 ;
  assign n3211 = n3210 ^ x34 ;
  assign n3212 = ~x64 & n3211 ;
  assign n3206 = x34 ^ x32 ;
  assign n3213 = n3212 ^ n3206 ;
  assign n3204 = x65 ^ x33 ;
  assign n3205 = n3041 & ~n3204 ;
  assign n3214 = n3213 ^ n3205 ;
  assign n3199 = x66 & n2879 ;
  assign n3198 = x68 & n2882 ;
  assign n3200 = n3199 ^ n3198 ;
  assign n3201 = n3200 ^ x32 ;
  assign n3197 = ~n340 & n2883 ;
  assign n3202 = n3201 ^ n3197 ;
  assign n3196 = x67 & n2887 ;
  assign n3203 = n3202 ^ n3196 ;
  assign n3215 = n3214 ^ n3203 ;
  assign n3219 = n3218 ^ n3215 ;
  assign n3220 = n3219 ^ x29 ;
  assign n3195 = x69 & n2581 ;
  assign n3221 = n3220 ^ n3195 ;
  assign n3194 = x71 & n2422 ;
  assign n3222 = n3221 ^ n3194 ;
  assign n3193 = ~n493 & n2423 ;
  assign n3223 = n3222 ^ n3193 ;
  assign n3225 = n3224 ^ n3223 ;
  assign n3190 = n3061 ^ n3052 ;
  assign n3191 = ~n3058 & n3190 ;
  assign n3192 = n3191 ^ n3061 ;
  assign n3226 = n3225 ^ n3192 ;
  assign n3227 = n3226 ^ x26 ;
  assign n3189 = x72 & n2018 ;
  assign n3228 = n3227 ^ n3189 ;
  assign n3188 = x74 & n2021 ;
  assign n3229 = n3228 ^ n3188 ;
  assign n3187 = n699 & n2022 ;
  assign n3230 = n3229 ^ n3187 ;
  assign n3232 = n3231 ^ n3230 ;
  assign n3236 = n3235 ^ n3232 ;
  assign n3237 = n3236 ^ x23 ;
  assign n3186 = x75 & n1658 ;
  assign n3238 = n3237 ^ n3186 ;
  assign n3185 = x77 & n1661 ;
  assign n3239 = n3238 ^ n3185 ;
  assign n3184 = ~n939 & n1662 ;
  assign n3240 = n3239 ^ n3184 ;
  assign n3242 = n3241 ^ n3240 ;
  assign n3181 = n3078 ^ n3069 ;
  assign n3182 = ~n3075 & n3181 ;
  assign n3183 = n3182 ^ n3078 ;
  assign n3243 = n3242 ^ n3183 ;
  assign n3244 = n3243 ^ x20 ;
  assign n3180 = x78 & n1327 ;
  assign n3245 = n3244 ^ n3180 ;
  assign n3179 = x80 & n1330 ;
  assign n3246 = n3245 ^ n3179 ;
  assign n3178 = n1206 & n1331 ;
  assign n3247 = n3246 ^ n3178 ;
  assign n3249 = n3248 ^ n3247 ;
  assign n3253 = n3252 ^ n3249 ;
  assign n3254 = n3253 ^ x17 ;
  assign n3177 = x81 & n1050 ;
  assign n3255 = n3254 ^ n3177 ;
  assign n3176 = x83 & n1053 ;
  assign n3256 = n3255 ^ n3176 ;
  assign n3175 = n1054 & n1512 ;
  assign n3257 = n3256 ^ n3175 ;
  assign n3259 = n3258 ^ n3257 ;
  assign n3172 = n3095 ^ n3086 ;
  assign n3173 = ~n3092 & n3172 ;
  assign n3174 = n3173 ^ n3095 ;
  assign n3260 = n3259 ^ n3174 ;
  assign n3261 = n3260 ^ x14 ;
  assign n3171 = x84 & n877 ;
  assign n3262 = n3261 ^ n3171 ;
  assign n3170 = x86 & n782 ;
  assign n3263 = n3262 ^ n3170 ;
  assign n3169 = n783 & n1857 ;
  assign n3264 = n3263 ^ n3169 ;
  assign n3266 = n3265 ^ n3264 ;
  assign n3270 = n3269 ^ n3266 ;
  assign n3271 = n3270 ^ x11 ;
  assign n3168 = x87 & n647 ;
  assign n3272 = n3271 ^ n3168 ;
  assign n3167 = x89 & ~n572 ;
  assign n3273 = n3272 ^ n3167 ;
  assign n3166 = ~n573 & n2249 ;
  assign n3274 = n3273 ^ n3166 ;
  assign n3276 = n3275 ^ n3274 ;
  assign n3280 = n3279 ^ n3276 ;
  assign n3281 = n3280 ^ x8 ;
  assign n3165 = x90 & n446 ;
  assign n3282 = n3281 ^ n3165 ;
  assign n3164 = x92 & n383 ;
  assign n3283 = n3282 ^ n3164 ;
  assign n3163 = n384 & n2684 ;
  assign n3284 = n3283 ^ n3163 ;
  assign n3286 = n3285 ^ n3284 ;
  assign n3290 = n3289 ^ n3286 ;
  assign n3291 = n3290 ^ x5 ;
  assign n3162 = x93 & n234 ;
  assign n3292 = n3291 ^ n3162 ;
  assign n3161 = x95 & n230 ;
  assign n3293 = n3292 ^ n3161 ;
  assign n3159 = n2670 ^ x95 ;
  assign n3160 = n231 & n3159 ;
  assign n3294 = n3293 ^ n3160 ;
  assign n3296 = n3295 ^ n3294 ;
  assign n3156 = n3126 ^ n3117 ;
  assign n3157 = n3123 & ~n3156 ;
  assign n3158 = n3157 ^ n3126 ;
  assign n3297 = n3296 ^ n3158 ;
  assign n3131 = x97 ^ x96 ;
  assign n3135 = n2978 ^ x94 ;
  assign n3136 = n3135 ^ x97 ;
  assign n3137 = n3136 ^ n2978 ;
  assign n3138 = n2981 & n3137 ;
  assign n3139 = n3138 ^ n2978 ;
  assign n3140 = n3131 & n3139 ;
  assign n3141 = n3140 ^ x96 ;
  assign n3142 = n3141 ^ x97 ;
  assign n3144 = x98 ^ x1 ;
  assign n3143 = x98 ^ x2 ;
  assign n3145 = n3144 ^ n3143 ;
  assign n3146 = ~n3142 & n3145 ;
  assign n3147 = n3146 ^ n3144 ;
  assign n3298 = n3297 ^ n3147 ;
  assign n3151 = x2 & x96 ;
  assign n3152 = n3151 ^ x97 ;
  assign n3153 = ~x1 & n3152 ;
  assign n3148 = n3147 ^ n2984 ;
  assign n3154 = n3153 ^ n3148 ;
  assign n3155 = ~x0 & n3154 ;
  assign n3299 = n3298 ^ n3155 ;
  assign n3303 = n3302 ^ n3299 ;
  assign n3468 = n3290 ^ n3158 ;
  assign n3469 = ~n3296 & ~n3468 ;
  assign n3470 = n3469 ^ n3290 ;
  assign n3466 = x95 & n227 ;
  assign n3459 = x92 & n390 ;
  assign n3452 = x89 & n578 ;
  assign n3445 = x86 & n788 ;
  assign n3437 = n3253 ^ n3174 ;
  assign n3438 = n3259 & n3437 ;
  assign n3439 = n3438 ^ n3253 ;
  assign n3435 = x83 & n1058 ;
  assign n3428 = x80 & n1335 ;
  assign n3420 = n3236 ^ n3183 ;
  assign n3421 = n3242 & n3420 ;
  assign n3422 = n3421 ^ n3236 ;
  assign n3418 = x77 & n1666 ;
  assign n3411 = x74 & n2014 ;
  assign n3403 = n3219 ^ n3192 ;
  assign n3404 = n3225 & n3403 ;
  assign n3405 = n3404 ^ n3219 ;
  assign n3401 = x71 & n2429 ;
  assign n3394 = x68 & n2887 ;
  assign n3387 = x35 & ~n3042 ;
  assign n3388 = ~n3214 & n3387 ;
  assign n3208 = x34 ^ x33 ;
  assign n3383 = ~n3041 & n3208 ;
  assign n3384 = x65 & n3383 ;
  assign n3372 = x35 ^ x34 ;
  assign n3378 = n3041 & ~n3372 ;
  assign n3379 = n3378 ^ n3041 ;
  assign n3380 = ~n150 & n3379 ;
  assign n3377 = x66 & n3041 ;
  assign n3381 = n3380 ^ n3377 ;
  assign n3382 = n3381 ^ x35 ;
  assign n3385 = n3384 ^ n3382 ;
  assign n3373 = x35 ^ x33 ;
  assign n3374 = ~n3041 & n3373 ;
  assign n3375 = n3372 & n3374 ;
  assign n3376 = x64 & n3375 ;
  assign n3386 = n3385 ^ n3376 ;
  assign n3389 = n3388 ^ n3386 ;
  assign n3390 = n3389 ^ x32 ;
  assign n3371 = x67 & n2879 ;
  assign n3391 = n3390 ^ n3371 ;
  assign n3370 = x69 & n2882 ;
  assign n3392 = n3391 ^ n3370 ;
  assign n3369 = ~n375 & n2883 ;
  assign n3393 = n3392 ^ n3369 ;
  assign n3395 = n3394 ^ n3393 ;
  assign n3366 = n3218 ^ n3214 ;
  assign n3367 = ~n3215 & n3366 ;
  assign n3368 = n3367 ^ n3218 ;
  assign n3396 = n3395 ^ n3368 ;
  assign n3397 = n3396 ^ x29 ;
  assign n3365 = x70 & n2581 ;
  assign n3398 = n3397 ^ n3365 ;
  assign n3364 = x72 & n2422 ;
  assign n3399 = n3398 ^ n3364 ;
  assign n3363 = n556 & n2423 ;
  assign n3400 = n3399 ^ n3363 ;
  assign n3402 = n3401 ^ n3400 ;
  assign n3406 = n3405 ^ n3402 ;
  assign n3407 = n3406 ^ x26 ;
  assign n3362 = x73 & n2018 ;
  assign n3408 = n3407 ^ n3362 ;
  assign n3361 = x75 & n2021 ;
  assign n3409 = n3408 ^ n3361 ;
  assign n3360 = ~n774 & n2022 ;
  assign n3410 = n3409 ^ n3360 ;
  assign n3412 = n3411 ^ n3410 ;
  assign n3357 = n3235 ^ n3226 ;
  assign n3358 = ~n3232 & n3357 ;
  assign n3359 = n3358 ^ n3235 ;
  assign n3413 = n3412 ^ n3359 ;
  assign n3414 = n3413 ^ x23 ;
  assign n3356 = x76 & n1658 ;
  assign n3415 = n3414 ^ n3356 ;
  assign n3355 = x78 & n1661 ;
  assign n3416 = n3415 ^ n3355 ;
  assign n3354 = ~n1025 & n1662 ;
  assign n3417 = n3416 ^ n3354 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n3423 = n3422 ^ n3419 ;
  assign n3424 = n3423 ^ x20 ;
  assign n3353 = x79 & n1327 ;
  assign n3425 = n3424 ^ n3353 ;
  assign n3352 = x81 & n1330 ;
  assign n3426 = n3425 ^ n3352 ;
  assign n3351 = n1305 & n1331 ;
  assign n3427 = n3426 ^ n3351 ;
  assign n3429 = n3428 ^ n3427 ;
  assign n3348 = n3252 ^ n3243 ;
  assign n3349 = ~n3249 & n3348 ;
  assign n3350 = n3349 ^ n3252 ;
  assign n3430 = n3429 ^ n3350 ;
  assign n3431 = n3430 ^ x17 ;
  assign n3347 = x82 & n1050 ;
  assign n3432 = n3431 ^ n3347 ;
  assign n3346 = x84 & n1053 ;
  assign n3433 = n3432 ^ n3346 ;
  assign n3345 = n1054 & n1624 ;
  assign n3434 = n3433 ^ n3345 ;
  assign n3436 = n3435 ^ n3434 ;
  assign n3440 = n3439 ^ n3436 ;
  assign n3441 = n3440 ^ x14 ;
  assign n3344 = x85 & n877 ;
  assign n3442 = n3441 ^ n3344 ;
  assign n3343 = x87 & n782 ;
  assign n3443 = n3442 ^ n3343 ;
  assign n3342 = n783 & n1982 ;
  assign n3444 = n3443 ^ n3342 ;
  assign n3446 = n3445 ^ n3444 ;
  assign n3339 = n3269 ^ n3260 ;
  assign n3340 = ~n3266 & n3339 ;
  assign n3341 = n3340 ^ n3269 ;
  assign n3447 = n3446 ^ n3341 ;
  assign n3448 = n3447 ^ x11 ;
  assign n3338 = x88 & n647 ;
  assign n3449 = n3448 ^ n3338 ;
  assign n3337 = x90 & ~n572 ;
  assign n3450 = n3449 ^ n3337 ;
  assign n3336 = ~n573 & n2386 ;
  assign n3451 = n3450 ^ n3336 ;
  assign n3453 = n3452 ^ n3451 ;
  assign n3333 = n3279 ^ n3270 ;
  assign n3334 = ~n3276 & n3333 ;
  assign n3335 = n3334 ^ n3279 ;
  assign n3454 = n3453 ^ n3335 ;
  assign n3455 = n3454 ^ x8 ;
  assign n3332 = x91 & n446 ;
  assign n3456 = n3455 ^ n3332 ;
  assign n3331 = x93 & n383 ;
  assign n3457 = n3456 ^ n3331 ;
  assign n3330 = n384 & n2836 ;
  assign n3458 = n3457 ^ n3330 ;
  assign n3460 = n3459 ^ n3458 ;
  assign n3327 = n3289 ^ n3280 ;
  assign n3328 = ~n3286 & ~n3327 ;
  assign n3329 = n3328 ^ n3289 ;
  assign n3461 = n3460 ^ n3329 ;
  assign n3462 = n3461 ^ x5 ;
  assign n3326 = x94 & n234 ;
  assign n3463 = n3462 ^ n3326 ;
  assign n3325 = x96 & n230 ;
  assign n3464 = n3463 ^ n3325 ;
  assign n3323 = n2819 ^ x96 ;
  assign n3324 = n231 & n3323 ;
  assign n3465 = n3464 ^ n3324 ;
  assign n3467 = n3466 ^ n3465 ;
  assign n3471 = n3470 ^ n3467 ;
  assign n3307 = x98 ^ x97 ;
  assign n3309 = ~n3142 & n3307 ;
  assign n3311 = x99 ^ x1 ;
  assign n3310 = x99 ^ x2 ;
  assign n3312 = n3311 ^ n3310 ;
  assign n3313 = ~n3309 & n3312 ;
  assign n3314 = n3313 ^ n3311 ;
  assign n3472 = n3471 ^ n3314 ;
  assign n3318 = x2 & x97 ;
  assign n3319 = n3318 ^ x98 ;
  assign n3320 = ~x1 & n3319 ;
  assign n3315 = n3314 ^ n3143 ;
  assign n3321 = n3320 ^ n3315 ;
  assign n3322 = ~x0 & n3321 ;
  assign n3473 = n3472 ^ n3322 ;
  assign n3304 = n3302 ^ n3297 ;
  assign n3305 = n3299 & n3304 ;
  assign n3306 = n3305 ^ n3302 ;
  assign n3474 = n3473 ^ n3306 ;
  assign n3637 = n3471 ^ n3306 ;
  assign n3638 = n3473 & ~n3637 ;
  assign n3639 = n3638 ^ n3471 ;
  assign n3632 = x96 & n227 ;
  assign n3624 = n3454 ^ n3329 ;
  assign n3625 = n3460 & ~n3624 ;
  assign n3626 = n3625 ^ n3454 ;
  assign n3622 = x93 & n390 ;
  assign n3614 = n3447 ^ n3335 ;
  assign n3615 = n3453 & n3614 ;
  assign n3616 = n3615 ^ n3447 ;
  assign n3612 = x90 & n578 ;
  assign n3604 = n3440 ^ n3341 ;
  assign n3605 = n3446 & n3604 ;
  assign n3606 = n3605 ^ n3440 ;
  assign n3602 = x87 & n788 ;
  assign n3595 = x84 & n1058 ;
  assign n3587 = n3423 ^ n3350 ;
  assign n3588 = n3429 & n3587 ;
  assign n3589 = n3588 ^ n3423 ;
  assign n3585 = x81 & n1335 ;
  assign n3578 = x78 & n1666 ;
  assign n3570 = n3406 ^ n3359 ;
  assign n3571 = n3412 & n3570 ;
  assign n3572 = n3571 ^ n3406 ;
  assign n3568 = x75 & n2014 ;
  assign n3557 = x71 & n2581 ;
  assign n3556 = x73 & n2422 ;
  assign n3558 = n3557 ^ n3556 ;
  assign n3559 = n3558 ^ x29 ;
  assign n3555 = n633 & n2423 ;
  assign n3560 = n3559 ^ n3555 ;
  assign n3554 = x72 & n2429 ;
  assign n3561 = n3560 ^ n3554 ;
  assign n3550 = n3389 ^ n3368 ;
  assign n3551 = n3395 & n3550 ;
  assign n3552 = n3551 ^ n3389 ;
  assign n3548 = x69 & n2887 ;
  assign n3537 = x65 & n3375 ;
  assign n3536 = x67 & n3378 ;
  assign n3538 = n3537 ^ n3536 ;
  assign n3539 = n3538 ^ x35 ;
  assign n3535 = ~n291 & n3379 ;
  assign n3540 = n3539 ^ n3535 ;
  assign n3534 = x66 & n3383 ;
  assign n3541 = n3540 ^ n3534 ;
  assign n3532 = x36 ^ x35 ;
  assign n3533 = x64 & n3532 ;
  assign n3542 = n3541 ^ n3533 ;
  assign n3531 = n3386 & n3388 ;
  assign n3543 = n3542 ^ n3531 ;
  assign n3544 = n3543 ^ x32 ;
  assign n3530 = x68 & n2879 ;
  assign n3545 = n3544 ^ n3530 ;
  assign n3529 = x70 & n2882 ;
  assign n3546 = n3545 ^ n3529 ;
  assign n3528 = ~n436 & n2883 ;
  assign n3547 = n3546 ^ n3528 ;
  assign n3549 = n3548 ^ n3547 ;
  assign n3553 = n3552 ^ n3549 ;
  assign n3562 = n3561 ^ n3553 ;
  assign n3525 = n3405 ^ n3396 ;
  assign n3526 = ~n3402 & n3525 ;
  assign n3527 = n3526 ^ n3405 ;
  assign n3563 = n3562 ^ n3527 ;
  assign n3564 = n3563 ^ x26 ;
  assign n3524 = x74 & n2018 ;
  assign n3565 = n3564 ^ n3524 ;
  assign n3523 = x76 & n2021 ;
  assign n3566 = n3565 ^ n3523 ;
  assign n3522 = ~n853 & n2022 ;
  assign n3567 = n3566 ^ n3522 ;
  assign n3569 = n3568 ^ n3567 ;
  assign n3573 = n3572 ^ n3569 ;
  assign n3574 = n3573 ^ x23 ;
  assign n3521 = x77 & n1658 ;
  assign n3575 = n3574 ^ n3521 ;
  assign n3520 = x79 & n1661 ;
  assign n3576 = n3575 ^ n3520 ;
  assign n3519 = n1118 & n1662 ;
  assign n3577 = n3576 ^ n3519 ;
  assign n3579 = n3578 ^ n3577 ;
  assign n3516 = n3422 ^ n3413 ;
  assign n3517 = ~n3419 & n3516 ;
  assign n3518 = n3517 ^ n3422 ;
  assign n3580 = n3579 ^ n3518 ;
  assign n3581 = n3580 ^ x20 ;
  assign n3515 = x80 & n1327 ;
  assign n3582 = n3581 ^ n3515 ;
  assign n3514 = x82 & n1330 ;
  assign n3583 = n3582 ^ n3514 ;
  assign n3513 = n1331 & n1411 ;
  assign n3584 = n3583 ^ n3513 ;
  assign n3586 = n3585 ^ n3584 ;
  assign n3590 = n3589 ^ n3586 ;
  assign n3591 = n3590 ^ x17 ;
  assign n3512 = x83 & n1050 ;
  assign n3592 = n3591 ^ n3512 ;
  assign n3511 = x85 & n1053 ;
  assign n3593 = n3592 ^ n3511 ;
  assign n3510 = n1054 & n1743 ;
  assign n3594 = n3593 ^ n3510 ;
  assign n3596 = n3595 ^ n3594 ;
  assign n3507 = n3439 ^ n3430 ;
  assign n3508 = ~n3436 & n3507 ;
  assign n3509 = n3508 ^ n3439 ;
  assign n3597 = n3596 ^ n3509 ;
  assign n3598 = n3597 ^ x14 ;
  assign n3506 = x86 & n877 ;
  assign n3599 = n3598 ^ n3506 ;
  assign n3505 = x88 & n782 ;
  assign n3600 = n3599 ^ n3505 ;
  assign n3504 = n783 & n2119 ;
  assign n3601 = n3600 ^ n3504 ;
  assign n3603 = n3602 ^ n3601 ;
  assign n3607 = n3606 ^ n3603 ;
  assign n3608 = n3607 ^ x11 ;
  assign n3503 = x89 & n647 ;
  assign n3609 = n3608 ^ n3503 ;
  assign n3502 = x91 & ~n572 ;
  assign n3610 = n3609 ^ n3502 ;
  assign n3501 = ~n573 & n2542 ;
  assign n3611 = n3610 ^ n3501 ;
  assign n3613 = n3612 ^ n3611 ;
  assign n3617 = n3616 ^ n3613 ;
  assign n3618 = n3617 ^ x8 ;
  assign n3500 = x92 & n446 ;
  assign n3619 = n3618 ^ n3500 ;
  assign n3499 = x94 & n383 ;
  assign n3620 = n3619 ^ n3499 ;
  assign n3498 = n384 & n2997 ;
  assign n3621 = n3620 ^ n3498 ;
  assign n3623 = n3622 ^ n3621 ;
  assign n3627 = n3626 ^ n3623 ;
  assign n3628 = n3627 ^ x5 ;
  assign n3497 = x95 & n234 ;
  assign n3629 = n3628 ^ n3497 ;
  assign n3496 = x97 & n230 ;
  assign n3630 = n3629 ^ n3496 ;
  assign n3494 = n2983 ^ x97 ;
  assign n3495 = n231 & n3494 ;
  assign n3631 = n3630 ^ n3495 ;
  assign n3633 = n3632 ^ n3631 ;
  assign n3491 = n3470 ^ n3461 ;
  assign n3492 = n3467 & n3491 ;
  assign n3493 = n3492 ^ n3470 ;
  assign n3634 = n3633 ^ n3493 ;
  assign n3475 = x99 ^ x98 ;
  assign n3477 = ~n3309 & n3475 ;
  assign n3479 = x100 ^ x1 ;
  assign n3478 = x100 ^ x2 ;
  assign n3480 = n3479 ^ n3478 ;
  assign n3481 = ~n3477 & n3480 ;
  assign n3482 = n3481 ^ n3479 ;
  assign n3635 = n3634 ^ n3482 ;
  assign n3486 = x2 & x98 ;
  assign n3487 = n3486 ^ x99 ;
  assign n3488 = ~x1 & n3487 ;
  assign n3483 = n3482 ^ n3310 ;
  assign n3489 = n3488 ^ n3483 ;
  assign n3490 = ~x0 & n3489 ;
  assign n3636 = n3635 ^ n3490 ;
  assign n3640 = n3639 ^ n3636 ;
  assign n3811 = n3627 ^ n3493 ;
  assign n3812 = n3633 & ~n3811 ;
  assign n3813 = n3812 ^ n3627 ;
  assign n3809 = x97 & n227 ;
  assign n3802 = x94 & n390 ;
  assign n3795 = x91 & n578 ;
  assign n3788 = x88 & n788 ;
  assign n3780 = n3590 ^ n3509 ;
  assign n3781 = n3596 & n3780 ;
  assign n3782 = n3781 ^ n3590 ;
  assign n3778 = x85 & n1058 ;
  assign n3771 = x82 & n1335 ;
  assign n3763 = n3573 ^ n3518 ;
  assign n3764 = n3579 & n3763 ;
  assign n3765 = n3764 ^ n3573 ;
  assign n3761 = x79 & n1666 ;
  assign n3754 = x76 & n2014 ;
  assign n3747 = x73 & n2429 ;
  assign n3740 = x70 & n2887 ;
  assign n3730 = x66 & n3375 ;
  assign n3729 = x68 & n3378 ;
  assign n3731 = n3730 ^ n3729 ;
  assign n3732 = n3731 ^ x35 ;
  assign n3728 = ~n340 & n3379 ;
  assign n3733 = n3732 ^ n3728 ;
  assign n3727 = x67 & n3383 ;
  assign n3734 = n3733 ^ n3727 ;
  assign n3721 = x35 & x36 ;
  assign n3722 = n3721 ^ x37 ;
  assign n3723 = ~x64 & n3722 ;
  assign n3717 = x37 ^ x35 ;
  assign n3724 = n3723 ^ n3717 ;
  assign n3715 = x65 ^ x36 ;
  assign n3716 = n3532 & ~n3715 ;
  assign n3725 = n3724 ^ n3716 ;
  assign n3712 = ~n3533 & n3541 ;
  assign n3713 = ~n3531 & n3712 ;
  assign n3714 = n3713 ^ n3541 ;
  assign n3726 = n3725 ^ n3714 ;
  assign n3735 = n3734 ^ n3726 ;
  assign n3736 = n3735 ^ x32 ;
  assign n3711 = x69 & n2879 ;
  assign n3737 = n3736 ^ n3711 ;
  assign n3710 = x71 & n2882 ;
  assign n3738 = n3737 ^ n3710 ;
  assign n3709 = ~n493 & n2883 ;
  assign n3739 = n3738 ^ n3709 ;
  assign n3741 = n3740 ^ n3739 ;
  assign n3706 = n3552 ^ n3543 ;
  assign n3707 = ~n3549 & n3706 ;
  assign n3708 = n3707 ^ n3552 ;
  assign n3742 = n3741 ^ n3708 ;
  assign n3743 = n3742 ^ x29 ;
  assign n3705 = x72 & n2581 ;
  assign n3744 = n3743 ^ n3705 ;
  assign n3704 = x74 & n2422 ;
  assign n3745 = n3744 ^ n3704 ;
  assign n3703 = n699 & n2423 ;
  assign n3746 = n3745 ^ n3703 ;
  assign n3748 = n3747 ^ n3746 ;
  assign n3700 = n3553 ^ n3527 ;
  assign n3701 = n3562 & ~n3700 ;
  assign n3702 = n3701 ^ n3561 ;
  assign n3749 = n3748 ^ n3702 ;
  assign n3750 = n3749 ^ x26 ;
  assign n3699 = x75 & n2018 ;
  assign n3751 = n3750 ^ n3699 ;
  assign n3698 = x77 & n2021 ;
  assign n3752 = n3751 ^ n3698 ;
  assign n3697 = ~n939 & n2022 ;
  assign n3753 = n3752 ^ n3697 ;
  assign n3755 = n3754 ^ n3753 ;
  assign n3694 = n3572 ^ n3563 ;
  assign n3695 = ~n3569 & n3694 ;
  assign n3696 = n3695 ^ n3572 ;
  assign n3756 = n3755 ^ n3696 ;
  assign n3757 = n3756 ^ x23 ;
  assign n3693 = x78 & n1658 ;
  assign n3758 = n3757 ^ n3693 ;
  assign n3692 = x80 & n1661 ;
  assign n3759 = n3758 ^ n3692 ;
  assign n3691 = n1206 & n1662 ;
  assign n3760 = n3759 ^ n3691 ;
  assign n3762 = n3761 ^ n3760 ;
  assign n3766 = n3765 ^ n3762 ;
  assign n3767 = n3766 ^ x20 ;
  assign n3690 = x81 & n1327 ;
  assign n3768 = n3767 ^ n3690 ;
  assign n3689 = x83 & n1330 ;
  assign n3769 = n3768 ^ n3689 ;
  assign n3688 = n1331 & n1512 ;
  assign n3770 = n3769 ^ n3688 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3685 = n3589 ^ n3580 ;
  assign n3686 = ~n3586 & n3685 ;
  assign n3687 = n3686 ^ n3589 ;
  assign n3773 = n3772 ^ n3687 ;
  assign n3774 = n3773 ^ x17 ;
  assign n3684 = x84 & n1050 ;
  assign n3775 = n3774 ^ n3684 ;
  assign n3683 = x86 & n1053 ;
  assign n3776 = n3775 ^ n3683 ;
  assign n3682 = n1054 & n1857 ;
  assign n3777 = n3776 ^ n3682 ;
  assign n3779 = n3778 ^ n3777 ;
  assign n3783 = n3782 ^ n3779 ;
  assign n3784 = n3783 ^ x14 ;
  assign n3681 = x87 & n877 ;
  assign n3785 = n3784 ^ n3681 ;
  assign n3680 = x89 & n782 ;
  assign n3786 = n3785 ^ n3680 ;
  assign n3679 = n783 & n2249 ;
  assign n3787 = n3786 ^ n3679 ;
  assign n3789 = n3788 ^ n3787 ;
  assign n3676 = n3606 ^ n3597 ;
  assign n3677 = ~n3603 & n3676 ;
  assign n3678 = n3677 ^ n3606 ;
  assign n3790 = n3789 ^ n3678 ;
  assign n3791 = n3790 ^ x11 ;
  assign n3675 = x90 & n647 ;
  assign n3792 = n3791 ^ n3675 ;
  assign n3674 = x92 & ~n572 ;
  assign n3793 = n3792 ^ n3674 ;
  assign n3673 = ~n573 & n2684 ;
  assign n3794 = n3793 ^ n3673 ;
  assign n3796 = n3795 ^ n3794 ;
  assign n3670 = n3616 ^ n3607 ;
  assign n3671 = ~n3613 & n3670 ;
  assign n3672 = n3671 ^ n3616 ;
  assign n3797 = n3796 ^ n3672 ;
  assign n3798 = n3797 ^ x8 ;
  assign n3669 = x93 & n446 ;
  assign n3799 = n3798 ^ n3669 ;
  assign n3668 = x95 & n383 ;
  assign n3800 = n3799 ^ n3668 ;
  assign n3667 = n384 & n3159 ;
  assign n3801 = n3800 ^ n3667 ;
  assign n3803 = n3802 ^ n3801 ;
  assign n3664 = n3626 ^ n3617 ;
  assign n3665 = ~n3623 & n3664 ;
  assign n3666 = n3665 ^ n3626 ;
  assign n3804 = n3803 ^ n3666 ;
  assign n3805 = n3804 ^ x5 ;
  assign n3663 = x96 & n234 ;
  assign n3806 = n3805 ^ n3663 ;
  assign n3662 = x98 & n230 ;
  assign n3807 = n3806 ^ n3662 ;
  assign n3660 = n3307 ^ n3141 ;
  assign n3661 = n231 & n3660 ;
  assign n3808 = n3807 ^ n3661 ;
  assign n3810 = n3809 ^ n3808 ;
  assign n3814 = n3813 ^ n3810 ;
  assign n3644 = x100 ^ x99 ;
  assign n3646 = ~n3477 & n3644 ;
  assign n3648 = x101 ^ x1 ;
  assign n3647 = x101 ^ x2 ;
  assign n3649 = n3648 ^ n3647 ;
  assign n3650 = ~n3646 & n3649 ;
  assign n3651 = n3650 ^ n3648 ;
  assign n3815 = n3814 ^ n3651 ;
  assign n3655 = x2 & x99 ;
  assign n3656 = n3655 ^ x100 ;
  assign n3657 = ~n255 & n3656 ;
  assign n3652 = n3651 ^ n3478 ;
  assign n3658 = n3657 ^ n3652 ;
  assign n3659 = ~x0 & n3658 ;
  assign n3816 = n3815 ^ n3659 ;
  assign n3641 = n3639 ^ n3634 ;
  assign n3642 = n3636 & ~n3641 ;
  assign n3643 = n3642 ^ n3639 ;
  assign n3817 = n3816 ^ n3643 ;
  assign n4007 = n3814 ^ n3643 ;
  assign n4008 = n3816 & n4007 ;
  assign n4009 = n4008 ^ n3814 ;
  assign n4002 = x98 & n227 ;
  assign n3994 = n3797 ^ n3666 ;
  assign n3995 = n3803 & n3994 ;
  assign n3996 = n3995 ^ n3797 ;
  assign n3992 = x95 & n390 ;
  assign n3984 = n3790 ^ n3672 ;
  assign n3985 = n3796 & n3984 ;
  assign n3986 = n3985 ^ n3790 ;
  assign n3982 = x92 & n578 ;
  assign n3974 = n3783 ^ n3678 ;
  assign n3975 = n3789 & n3974 ;
  assign n3976 = n3975 ^ n3783 ;
  assign n3972 = x89 & n788 ;
  assign n3965 = x86 & n1058 ;
  assign n3957 = n3766 ^ n3687 ;
  assign n3958 = n3772 & n3957 ;
  assign n3959 = n3958 ^ n3766 ;
  assign n3955 = x83 & n1335 ;
  assign n3944 = n3735 ^ n3708 ;
  assign n3945 = n3741 & n3944 ;
  assign n3946 = n3945 ^ n3735 ;
  assign n3942 = x71 & n2887 ;
  assign n3935 = x68 & n3383 ;
  assign n3928 = x38 & ~n3533 ;
  assign n3929 = ~n3725 & n3928 ;
  assign n3719 = x37 ^ x36 ;
  assign n3924 = ~n3532 & n3719 ;
  assign n3925 = x65 & n3924 ;
  assign n3913 = x38 ^ x37 ;
  assign n3919 = n3532 & ~n3913 ;
  assign n3920 = n3919 ^ n3532 ;
  assign n3921 = ~n150 & n3920 ;
  assign n3918 = x66 & n3532 ;
  assign n3922 = n3921 ^ n3918 ;
  assign n3923 = n3922 ^ x38 ;
  assign n3926 = n3925 ^ n3923 ;
  assign n3914 = x38 ^ x36 ;
  assign n3915 = ~n3532 & n3914 ;
  assign n3916 = n3913 & n3915 ;
  assign n3917 = x64 & n3916 ;
  assign n3927 = n3926 ^ n3917 ;
  assign n3930 = n3929 ^ n3927 ;
  assign n3931 = n3930 ^ x35 ;
  assign n3912 = x67 & n3375 ;
  assign n3932 = n3931 ^ n3912 ;
  assign n3911 = x69 & n3378 ;
  assign n3933 = n3932 ^ n3911 ;
  assign n3910 = ~n375 & n3379 ;
  assign n3934 = n3933 ^ n3910 ;
  assign n3936 = n3935 ^ n3934 ;
  assign n3907 = n3734 ^ n3725 ;
  assign n3908 = ~n3726 & n3907 ;
  assign n3909 = n3908 ^ n3734 ;
  assign n3937 = n3936 ^ n3909 ;
  assign n3938 = n3937 ^ x32 ;
  assign n3906 = x70 & n2879 ;
  assign n3939 = n3938 ^ n3906 ;
  assign n3905 = x72 & n2882 ;
  assign n3940 = n3939 ^ n3905 ;
  assign n3904 = n556 & n2883 ;
  assign n3941 = n3940 ^ n3904 ;
  assign n3943 = n3942 ^ n3941 ;
  assign n3947 = n3946 ^ n3943 ;
  assign n3901 = n3742 ^ n3702 ;
  assign n3902 = n3748 & n3901 ;
  assign n3894 = x73 & n2581 ;
  assign n3893 = x75 & n2422 ;
  assign n3895 = n3894 ^ n3893 ;
  assign n3896 = n3895 ^ x29 ;
  assign n3892 = ~n774 & n2423 ;
  assign n3897 = n3896 ^ n3892 ;
  assign n3891 = x74 & n2429 ;
  assign n3898 = n3897 ^ n3891 ;
  assign n3899 = n3898 ^ n3742 ;
  assign n3903 = n3902 ^ n3899 ;
  assign n3948 = n3947 ^ n3903 ;
  assign n3888 = n3749 ^ n3696 ;
  assign n3889 = n3755 & n3888 ;
  assign n3881 = x76 & n2018 ;
  assign n3880 = x78 & n2021 ;
  assign n3882 = n3881 ^ n3880 ;
  assign n3883 = n3882 ^ x26 ;
  assign n3879 = ~n1025 & n2022 ;
  assign n3884 = n3883 ^ n3879 ;
  assign n3878 = x77 & n2014 ;
  assign n3885 = n3884 ^ n3878 ;
  assign n3886 = n3885 ^ n3749 ;
  assign n3890 = n3889 ^ n3886 ;
  assign n3949 = n3948 ^ n3890 ;
  assign n3868 = x79 & n1658 ;
  assign n3867 = x81 & n1661 ;
  assign n3869 = n3868 ^ n3867 ;
  assign n3870 = n3869 ^ x23 ;
  assign n3866 = n1305 & n1662 ;
  assign n3871 = n3870 ^ n3866 ;
  assign n3865 = x80 & n1666 ;
  assign n3872 = n3871 ^ n3865 ;
  assign n3873 = n3872 ^ n3765 ;
  assign n3874 = n3873 ^ n3756 ;
  assign n3875 = n3874 ^ n3872 ;
  assign n3876 = ~n3762 & n3875 ;
  assign n3877 = n3876 ^ n3873 ;
  assign n3950 = n3949 ^ n3877 ;
  assign n3951 = n3950 ^ x20 ;
  assign n3864 = x82 & n1327 ;
  assign n3952 = n3951 ^ n3864 ;
  assign n3863 = x84 & n1330 ;
  assign n3953 = n3952 ^ n3863 ;
  assign n3862 = n1331 & n1624 ;
  assign n3954 = n3953 ^ n3862 ;
  assign n3956 = n3955 ^ n3954 ;
  assign n3960 = n3959 ^ n3956 ;
  assign n3961 = n3960 ^ x17 ;
  assign n3861 = x85 & n1050 ;
  assign n3962 = n3961 ^ n3861 ;
  assign n3860 = x87 & n1053 ;
  assign n3963 = n3962 ^ n3860 ;
  assign n3859 = n1054 & n1982 ;
  assign n3964 = n3963 ^ n3859 ;
  assign n3966 = n3965 ^ n3964 ;
  assign n3856 = n3782 ^ n3773 ;
  assign n3857 = ~n3779 & n3856 ;
  assign n3858 = n3857 ^ n3782 ;
  assign n3967 = n3966 ^ n3858 ;
  assign n3968 = n3967 ^ x14 ;
  assign n3855 = x88 & n877 ;
  assign n3969 = n3968 ^ n3855 ;
  assign n3854 = x90 & n782 ;
  assign n3970 = n3969 ^ n3854 ;
  assign n3853 = n783 & n2386 ;
  assign n3971 = n3970 ^ n3853 ;
  assign n3973 = n3972 ^ n3971 ;
  assign n3977 = n3976 ^ n3973 ;
  assign n3978 = n3977 ^ x11 ;
  assign n3852 = x91 & n647 ;
  assign n3979 = n3978 ^ n3852 ;
  assign n3851 = x93 & ~n572 ;
  assign n3980 = n3979 ^ n3851 ;
  assign n3850 = ~n573 & n2836 ;
  assign n3981 = n3980 ^ n3850 ;
  assign n3983 = n3982 ^ n3981 ;
  assign n3987 = n3986 ^ n3983 ;
  assign n3988 = n3987 ^ x8 ;
  assign n3849 = x94 & n446 ;
  assign n3989 = n3988 ^ n3849 ;
  assign n3848 = x96 & n383 ;
  assign n3990 = n3989 ^ n3848 ;
  assign n3847 = n384 & n3323 ;
  assign n3991 = n3990 ^ n3847 ;
  assign n3993 = n3992 ^ n3991 ;
  assign n3997 = n3996 ^ n3993 ;
  assign n3998 = n3997 ^ x5 ;
  assign n3846 = x97 & n234 ;
  assign n3999 = n3998 ^ n3846 ;
  assign n3845 = x99 & n230 ;
  assign n4000 = n3999 ^ n3845 ;
  assign n3843 = n3309 ^ x99 ;
  assign n3844 = n231 & n3843 ;
  assign n4001 = n4000 ^ n3844 ;
  assign n4003 = n4002 ^ n4001 ;
  assign n3840 = n3813 ^ n3804 ;
  assign n3841 = ~n3810 & n3840 ;
  assign n3842 = n3841 ^ n3813 ;
  assign n4004 = n4003 ^ n3842 ;
  assign n3820 = x101 ^ x98 ;
  assign n3818 = x101 ^ x100 ;
  assign n3821 = n3644 & n3818 ;
  assign n3822 = ~n3309 & n3821 ;
  assign n3823 = n3820 & n3822 ;
  assign n3824 = n3823 ^ n3821 ;
  assign n3825 = n3824 ^ x100 ;
  assign n3826 = n3825 ^ x101 ;
  assign n3828 = x102 ^ x1 ;
  assign n3827 = x102 ^ x2 ;
  assign n3829 = n3828 ^ n3827 ;
  assign n3830 = ~n3826 & n3829 ;
  assign n3831 = n3830 ^ n3828 ;
  assign n4005 = n4004 ^ n3831 ;
  assign n3835 = x2 & x100 ;
  assign n3836 = n3835 ^ x101 ;
  assign n3837 = ~x1 & n3836 ;
  assign n3832 = n3831 ^ n3647 ;
  assign n3838 = n3837 ^ n3832 ;
  assign n3839 = ~x0 & n3838 ;
  assign n4006 = n4005 ^ n3839 ;
  assign n4010 = n4009 ^ n4006 ;
  assign n4187 = n3997 ^ n3842 ;
  assign n4188 = n4003 & n4187 ;
  assign n4189 = n4188 ^ n3997 ;
  assign n4185 = x99 & n227 ;
  assign n4178 = x96 & n390 ;
  assign n4171 = x93 & n578 ;
  assign n4164 = x90 & n788 ;
  assign n4156 = n3960 ^ n3858 ;
  assign n4157 = n3966 & n4156 ;
  assign n4158 = n4157 ^ n3960 ;
  assign n4154 = x87 & n1058 ;
  assign n4147 = x84 & n1335 ;
  assign n4140 = x81 & n1666 ;
  assign n4133 = x78 & n2014 ;
  assign n4126 = x75 & n2429 ;
  assign n4119 = x72 & n2887 ;
  assign n4111 = n3930 ^ n3909 ;
  assign n4112 = n3936 & n4111 ;
  assign n4113 = n4112 ^ n3930 ;
  assign n4109 = x69 & n3383 ;
  assign n4098 = x65 & n3916 ;
  assign n4097 = x67 & n3919 ;
  assign n4099 = n4098 ^ n4097 ;
  assign n4100 = n4099 ^ x38 ;
  assign n4096 = ~n291 & n3920 ;
  assign n4101 = n4100 ^ n4096 ;
  assign n4095 = x66 & n3924 ;
  assign n4102 = n4101 ^ n4095 ;
  assign n4093 = x39 ^ x38 ;
  assign n4094 = x64 & n4093 ;
  assign n4103 = n4102 ^ n4094 ;
  assign n4092 = n3927 & n3929 ;
  assign n4104 = n4103 ^ n4092 ;
  assign n4105 = n4104 ^ x35 ;
  assign n4091 = x68 & n3375 ;
  assign n4106 = n4105 ^ n4091 ;
  assign n4090 = x70 & n3378 ;
  assign n4107 = n4106 ^ n4090 ;
  assign n4089 = ~n436 & n3379 ;
  assign n4108 = n4107 ^ n4089 ;
  assign n4110 = n4109 ^ n4108 ;
  assign n4114 = n4113 ^ n4110 ;
  assign n4115 = n4114 ^ x32 ;
  assign n4088 = x71 & n2879 ;
  assign n4116 = n4115 ^ n4088 ;
  assign n4087 = x73 & n2882 ;
  assign n4117 = n4116 ^ n4087 ;
  assign n4086 = n633 & n2883 ;
  assign n4118 = n4117 ^ n4086 ;
  assign n4120 = n4119 ^ n4118 ;
  assign n4083 = n3946 ^ n3937 ;
  assign n4084 = ~n3943 & n4083 ;
  assign n4085 = n4084 ^ n3946 ;
  assign n4121 = n4120 ^ n4085 ;
  assign n4122 = n4121 ^ x29 ;
  assign n4082 = x74 & n2581 ;
  assign n4123 = n4122 ^ n4082 ;
  assign n4081 = x76 & n2422 ;
  assign n4124 = n4123 ^ n4081 ;
  assign n4080 = ~n853 & n2423 ;
  assign n4125 = n4124 ^ n4080 ;
  assign n4127 = n4126 ^ n4125 ;
  assign n4077 = n3947 ^ n3898 ;
  assign n4078 = n3903 & n4077 ;
  assign n4079 = n4078 ^ n3898 ;
  assign n4128 = n4127 ^ n4079 ;
  assign n4129 = n4128 ^ x26 ;
  assign n4076 = x77 & n2018 ;
  assign n4130 = n4129 ^ n4076 ;
  assign n4075 = x79 & n2021 ;
  assign n4131 = n4130 ^ n4075 ;
  assign n4074 = n1118 & n2022 ;
  assign n4132 = n4131 ^ n4074 ;
  assign n4134 = n4133 ^ n4132 ;
  assign n4071 = n3948 ^ n3885 ;
  assign n4072 = n3890 & n4071 ;
  assign n4073 = n4072 ^ n3885 ;
  assign n4135 = n4134 ^ n4073 ;
  assign n4136 = n4135 ^ x23 ;
  assign n4070 = x80 & n1658 ;
  assign n4137 = n4136 ^ n4070 ;
  assign n4069 = x82 & n1661 ;
  assign n4138 = n4137 ^ n4069 ;
  assign n4068 = n1411 & n1662 ;
  assign n4139 = n4138 ^ n4068 ;
  assign n4141 = n4140 ^ n4139 ;
  assign n4065 = n3949 ^ n3872 ;
  assign n4066 = n3877 & n4065 ;
  assign n4067 = n4066 ^ n3872 ;
  assign n4142 = n4141 ^ n4067 ;
  assign n4143 = n4142 ^ x20 ;
  assign n4064 = x83 & n1327 ;
  assign n4144 = n4143 ^ n4064 ;
  assign n4063 = x85 & n1330 ;
  assign n4145 = n4144 ^ n4063 ;
  assign n4062 = n1331 & n1743 ;
  assign n4146 = n4145 ^ n4062 ;
  assign n4148 = n4147 ^ n4146 ;
  assign n4059 = n3959 ^ n3950 ;
  assign n4060 = ~n3956 & n4059 ;
  assign n4061 = n4060 ^ n3959 ;
  assign n4149 = n4148 ^ n4061 ;
  assign n4150 = n4149 ^ x17 ;
  assign n4058 = x86 & n1050 ;
  assign n4151 = n4150 ^ n4058 ;
  assign n4057 = x88 & n1053 ;
  assign n4152 = n4151 ^ n4057 ;
  assign n4056 = n1054 & n2119 ;
  assign n4153 = n4152 ^ n4056 ;
  assign n4155 = n4154 ^ n4153 ;
  assign n4159 = n4158 ^ n4155 ;
  assign n4160 = n4159 ^ x14 ;
  assign n4055 = x89 & n877 ;
  assign n4161 = n4160 ^ n4055 ;
  assign n4054 = x91 & n782 ;
  assign n4162 = n4161 ^ n4054 ;
  assign n4053 = n783 & n2542 ;
  assign n4163 = n4162 ^ n4053 ;
  assign n4165 = n4164 ^ n4163 ;
  assign n4050 = n3976 ^ n3967 ;
  assign n4051 = ~n3973 & n4050 ;
  assign n4052 = n4051 ^ n3976 ;
  assign n4166 = n4165 ^ n4052 ;
  assign n4167 = n4166 ^ x11 ;
  assign n4049 = x92 & n647 ;
  assign n4168 = n4167 ^ n4049 ;
  assign n4048 = x94 & ~n572 ;
  assign n4169 = n4168 ^ n4048 ;
  assign n4047 = ~n573 & n2997 ;
  assign n4170 = n4169 ^ n4047 ;
  assign n4172 = n4171 ^ n4170 ;
  assign n4044 = n3986 ^ n3977 ;
  assign n4045 = ~n3983 & n4044 ;
  assign n4046 = n4045 ^ n3986 ;
  assign n4173 = n4172 ^ n4046 ;
  assign n4174 = n4173 ^ x8 ;
  assign n4043 = x95 & n446 ;
  assign n4175 = n4174 ^ n4043 ;
  assign n4042 = x97 & n383 ;
  assign n4176 = n4175 ^ n4042 ;
  assign n4041 = n384 & n3494 ;
  assign n4177 = n4176 ^ n4041 ;
  assign n4179 = n4178 ^ n4177 ;
  assign n4038 = n3996 ^ n3987 ;
  assign n4039 = ~n3993 & n4038 ;
  assign n4040 = n4039 ^ n3996 ;
  assign n4180 = n4179 ^ n4040 ;
  assign n4181 = n4180 ^ x5 ;
  assign n4037 = x98 & n234 ;
  assign n4182 = n4181 ^ n4037 ;
  assign n4036 = x100 & n230 ;
  assign n4183 = n4182 ^ n4036 ;
  assign n4034 = n3477 ^ x100 ;
  assign n4035 = n231 & n4034 ;
  assign n4184 = n4183 ^ n4035 ;
  assign n4186 = n4185 ^ n4184 ;
  assign n4190 = n4189 ^ n4186 ;
  assign n4016 = x101 & n3825 ;
  assign n4018 = n4016 ^ n3826 ;
  assign n4019 = x102 & n4018 ;
  assign n4017 = ~x102 & ~n4016 ;
  assign n4020 = n4019 ^ n4017 ;
  assign n4022 = x103 ^ x1 ;
  assign n4021 = x103 ^ x2 ;
  assign n4023 = n4022 ^ n4021 ;
  assign n4024 = n4020 & n4023 ;
  assign n4025 = n4024 ^ n4022 ;
  assign n4191 = n4190 ^ n4025 ;
  assign n4029 = x2 & x101 ;
  assign n4030 = n4029 ^ x102 ;
  assign n4031 = ~x1 & n4030 ;
  assign n4026 = n4025 ^ n3827 ;
  assign n4032 = n4031 ^ n4026 ;
  assign n4033 = ~x0 & n4032 ;
  assign n4192 = n4191 ^ n4033 ;
  assign n4011 = n4009 ^ n4004 ;
  assign n4012 = ~n4006 & n4011 ;
  assign n4013 = n4012 ^ n4009 ;
  assign n4193 = n4192 ^ n4013 ;
  assign n4385 = n4190 ^ n4013 ;
  assign n4386 = n4192 & n4385 ;
  assign n4387 = n4386 ^ n4190 ;
  assign n4380 = x100 & n227 ;
  assign n4372 = n4173 ^ n4040 ;
  assign n4373 = n4179 & n4372 ;
  assign n4374 = n4373 ^ n4173 ;
  assign n4370 = x97 & n390 ;
  assign n4362 = n4166 ^ n4046 ;
  assign n4363 = n4172 & n4362 ;
  assign n4364 = n4363 ^ n4166 ;
  assign n4360 = x94 & n578 ;
  assign n4352 = n4159 ^ n4052 ;
  assign n4353 = n4165 & n4352 ;
  assign n4354 = n4353 ^ n4159 ;
  assign n4350 = x91 & n788 ;
  assign n4343 = x88 & n1058 ;
  assign n4335 = n4142 ^ n4061 ;
  assign n4336 = n4148 & n4335 ;
  assign n4337 = n4336 ^ n4142 ;
  assign n4333 = x85 & n1335 ;
  assign n4326 = x82 & n1666 ;
  assign n4319 = x79 & n2014 ;
  assign n4312 = x76 & n2429 ;
  assign n4304 = n4114 ^ n4085 ;
  assign n4305 = n4120 & n4304 ;
  assign n4306 = n4305 ^ n4114 ;
  assign n4302 = x73 & n2887 ;
  assign n4291 = ~n4094 & n4102 ;
  assign n4292 = ~n4092 & n4291 ;
  assign n4293 = n4292 ^ n4102 ;
  assign n4285 = ~x38 & ~x39 ;
  assign n4286 = n4285 ^ x40 ;
  assign n4287 = ~x64 & ~n4286 ;
  assign n4288 = n4287 ^ n4093 ;
  assign n4289 = n4288 ^ n4094 ;
  assign n4281 = x40 ^ x38 ;
  assign n4290 = n4289 ^ n4281 ;
  assign n4294 = n4293 ^ n4290 ;
  assign n4279 = x65 ^ x39 ;
  assign n4280 = n4093 & ~n4279 ;
  assign n4295 = n4294 ^ n4280 ;
  assign n4274 = x66 & n3916 ;
  assign n4273 = x68 & n3919 ;
  assign n4275 = n4274 ^ n4273 ;
  assign n4276 = n4275 ^ x38 ;
  assign n4272 = ~n340 & n3920 ;
  assign n4277 = n4276 ^ n4272 ;
  assign n4271 = x67 & n3924 ;
  assign n4278 = n4277 ^ n4271 ;
  assign n4296 = n4295 ^ n4278 ;
  assign n4261 = x69 & n3375 ;
  assign n4260 = x71 & n3378 ;
  assign n4262 = n4261 ^ n4260 ;
  assign n4263 = n4262 ^ x35 ;
  assign n4259 = ~n493 & n3379 ;
  assign n4264 = n4263 ^ n4259 ;
  assign n4258 = x70 & n3383 ;
  assign n4265 = n4264 ^ n4258 ;
  assign n4266 = n4265 ^ n4113 ;
  assign n4267 = n4266 ^ n4104 ;
  assign n4268 = n4267 ^ n4265 ;
  assign n4269 = ~n4110 & n4268 ;
  assign n4270 = n4269 ^ n4266 ;
  assign n4297 = n4296 ^ n4270 ;
  assign n4298 = n4297 ^ x32 ;
  assign n4257 = x72 & n2879 ;
  assign n4299 = n4298 ^ n4257 ;
  assign n4256 = x74 & n2882 ;
  assign n4300 = n4299 ^ n4256 ;
  assign n4255 = n699 & n2883 ;
  assign n4301 = n4300 ^ n4255 ;
  assign n4303 = n4302 ^ n4301 ;
  assign n4307 = n4306 ^ n4303 ;
  assign n4308 = n4307 ^ x29 ;
  assign n4254 = x75 & n2581 ;
  assign n4309 = n4308 ^ n4254 ;
  assign n4253 = x77 & n2422 ;
  assign n4310 = n4309 ^ n4253 ;
  assign n4252 = ~n939 & n2423 ;
  assign n4311 = n4310 ^ n4252 ;
  assign n4313 = n4312 ^ n4311 ;
  assign n4249 = n4121 ^ n4079 ;
  assign n4250 = n4127 & n4249 ;
  assign n4251 = n4250 ^ n4121 ;
  assign n4314 = n4313 ^ n4251 ;
  assign n4315 = n4314 ^ x26 ;
  assign n4248 = x78 & n2018 ;
  assign n4316 = n4315 ^ n4248 ;
  assign n4247 = x80 & n2021 ;
  assign n4317 = n4316 ^ n4247 ;
  assign n4246 = n1206 & n2022 ;
  assign n4318 = n4317 ^ n4246 ;
  assign n4320 = n4319 ^ n4318 ;
  assign n4243 = n4128 ^ n4073 ;
  assign n4244 = n4134 & n4243 ;
  assign n4245 = n4244 ^ n4128 ;
  assign n4321 = n4320 ^ n4245 ;
  assign n4322 = n4321 ^ x23 ;
  assign n4242 = x81 & n1658 ;
  assign n4323 = n4322 ^ n4242 ;
  assign n4241 = x83 & n1661 ;
  assign n4324 = n4323 ^ n4241 ;
  assign n4240 = n1512 & n1662 ;
  assign n4325 = n4324 ^ n4240 ;
  assign n4327 = n4326 ^ n4325 ;
  assign n4237 = n4135 ^ n4067 ;
  assign n4238 = n4141 & n4237 ;
  assign n4239 = n4238 ^ n4135 ;
  assign n4328 = n4327 ^ n4239 ;
  assign n4329 = n4328 ^ x20 ;
  assign n4236 = x84 & n1327 ;
  assign n4330 = n4329 ^ n4236 ;
  assign n4235 = x86 & n1330 ;
  assign n4331 = n4330 ^ n4235 ;
  assign n4234 = n1331 & n1857 ;
  assign n4332 = n4331 ^ n4234 ;
  assign n4334 = n4333 ^ n4332 ;
  assign n4338 = n4337 ^ n4334 ;
  assign n4339 = n4338 ^ x17 ;
  assign n4233 = x87 & n1050 ;
  assign n4340 = n4339 ^ n4233 ;
  assign n4232 = x89 & n1053 ;
  assign n4341 = n4340 ^ n4232 ;
  assign n4231 = n1054 & n2249 ;
  assign n4342 = n4341 ^ n4231 ;
  assign n4344 = n4343 ^ n4342 ;
  assign n4228 = n4158 ^ n4149 ;
  assign n4229 = ~n4155 & n4228 ;
  assign n4230 = n4229 ^ n4158 ;
  assign n4345 = n4344 ^ n4230 ;
  assign n4346 = n4345 ^ x14 ;
  assign n4227 = x90 & n877 ;
  assign n4347 = n4346 ^ n4227 ;
  assign n4226 = x92 & n782 ;
  assign n4348 = n4347 ^ n4226 ;
  assign n4225 = n783 & n2684 ;
  assign n4349 = n4348 ^ n4225 ;
  assign n4351 = n4350 ^ n4349 ;
  assign n4355 = n4354 ^ n4351 ;
  assign n4356 = n4355 ^ x11 ;
  assign n4224 = x93 & n647 ;
  assign n4357 = n4356 ^ n4224 ;
  assign n4223 = x95 & ~n572 ;
  assign n4358 = n4357 ^ n4223 ;
  assign n4222 = ~n573 & n3159 ;
  assign n4359 = n4358 ^ n4222 ;
  assign n4361 = n4360 ^ n4359 ;
  assign n4365 = n4364 ^ n4361 ;
  assign n4366 = n4365 ^ x8 ;
  assign n4221 = x96 & n446 ;
  assign n4367 = n4366 ^ n4221 ;
  assign n4220 = x98 & n383 ;
  assign n4368 = n4367 ^ n4220 ;
  assign n4219 = n384 & n3660 ;
  assign n4369 = n4368 ^ n4219 ;
  assign n4371 = n4370 ^ n4369 ;
  assign n4375 = n4374 ^ n4371 ;
  assign n4376 = n4375 ^ x5 ;
  assign n4218 = x99 & n234 ;
  assign n4377 = n4376 ^ n4218 ;
  assign n4217 = x101 & n230 ;
  assign n4378 = n4377 ^ n4217 ;
  assign n4215 = n3646 ^ x101 ;
  assign n4216 = n231 & n4215 ;
  assign n4379 = n4378 ^ n4216 ;
  assign n4381 = n4380 ^ n4379 ;
  assign n4212 = n4189 ^ n4180 ;
  assign n4213 = ~n4186 & n4212 ;
  assign n4214 = n4213 ^ n4189 ;
  assign n4382 = n4381 ^ n4214 ;
  assign n4197 = ~x103 & ~n4019 ;
  assign n4196 = x103 & ~n4017 ;
  assign n4198 = n4197 ^ n4196 ;
  assign n4200 = x104 ^ x1 ;
  assign n4199 = x104 ^ x2 ;
  assign n4201 = n4200 ^ n4199 ;
  assign n4202 = n4198 & n4201 ;
  assign n4203 = n4202 ^ n4200 ;
  assign n4383 = n4382 ^ n4203 ;
  assign n4207 = x2 & x102 ;
  assign n4208 = n4207 ^ x103 ;
  assign n4209 = ~x1 & n4208 ;
  assign n4204 = n4203 ^ n4021 ;
  assign n4210 = n4209 ^ n4204 ;
  assign n4211 = ~x0 & n4210 ;
  assign n4384 = n4383 ^ n4211 ;
  assign n4388 = n4387 ^ n4384 ;
  assign n4587 = n4375 ^ n4214 ;
  assign n4588 = n4381 & n4587 ;
  assign n4589 = n4588 ^ n4375 ;
  assign n4585 = x101 & n227 ;
  assign n4578 = x98 & n390 ;
  assign n4571 = x95 & n578 ;
  assign n4564 = x92 & n788 ;
  assign n4556 = n4338 ^ n4230 ;
  assign n4557 = n4344 & n4556 ;
  assign n4558 = n4557 ^ n4338 ;
  assign n4554 = x89 & n1058 ;
  assign n4547 = x86 & n1335 ;
  assign n4539 = n4321 ^ n4239 ;
  assign n4540 = n4327 & n4539 ;
  assign n4541 = n4540 ^ n4321 ;
  assign n4537 = x83 & n1666 ;
  assign n4529 = n4314 ^ n4245 ;
  assign n4530 = n4320 & n4529 ;
  assign n4531 = n4530 ^ n4314 ;
  assign n4527 = x80 & n2014 ;
  assign n4519 = n4307 ^ n4251 ;
  assign n4520 = n4313 & n4519 ;
  assign n4521 = n4520 ^ n4307 ;
  assign n4517 = x77 & n2429 ;
  assign n4510 = x74 & n2887 ;
  assign n4503 = x71 & n3383 ;
  assign n4495 = n4293 ^ n4278 ;
  assign n4496 = n4295 & n4495 ;
  assign n4497 = n4496 ^ n4293 ;
  assign n4489 = x67 & n3916 ;
  assign n4488 = x69 & n3919 ;
  assign n4490 = n4489 ^ n4488 ;
  assign n4491 = n4490 ^ x38 ;
  assign n4487 = ~n375 & n3920 ;
  assign n4492 = n4491 ^ n4487 ;
  assign n4486 = x68 & n3924 ;
  assign n4493 = n4492 ^ n4486 ;
  assign n4470 = x41 ^ x40 ;
  assign n4471 = n4093 & ~n4470 ;
  assign n4472 = n4471 ^ n4093 ;
  assign n4479 = x65 & n4472 ;
  assign n4283 = x40 ^ x39 ;
  assign n4473 = ~n4093 & ~n4283 ;
  assign n4474 = n4470 & n4473 ;
  assign n4480 = n4479 ^ n4474 ;
  assign n4481 = ~x64 & n4480 ;
  assign n4482 = n4481 ^ n4474 ;
  assign n4469 = x66 & n4093 ;
  assign n4483 = n4482 ^ n4469 ;
  assign n4467 = ~n4093 & n4283 ;
  assign n4468 = x65 & n4467 ;
  assign n4484 = n4483 ^ n4468 ;
  assign n4462 = n4287 ^ n4283 ;
  assign n4463 = x41 & ~n149 ;
  assign n4464 = ~n4093 & n4463 ;
  assign n4465 = ~n4462 & n4464 ;
  assign n4466 = n4465 ^ n4463 ;
  assign n4485 = n4484 ^ n4466 ;
  assign n4494 = n4493 ^ n4485 ;
  assign n4498 = n4497 ^ n4494 ;
  assign n4499 = n4498 ^ x35 ;
  assign n4461 = x70 & n3375 ;
  assign n4500 = n4499 ^ n4461 ;
  assign n4460 = x72 & n3378 ;
  assign n4501 = n4500 ^ n4460 ;
  assign n4459 = n556 & n3379 ;
  assign n4502 = n4501 ^ n4459 ;
  assign n4504 = n4503 ^ n4502 ;
  assign n4456 = n4296 ^ n4265 ;
  assign n4457 = n4270 & n4456 ;
  assign n4458 = n4457 ^ n4265 ;
  assign n4505 = n4504 ^ n4458 ;
  assign n4506 = n4505 ^ x32 ;
  assign n4455 = x73 & n2879 ;
  assign n4507 = n4506 ^ n4455 ;
  assign n4454 = x75 & n2882 ;
  assign n4508 = n4507 ^ n4454 ;
  assign n4453 = ~n774 & n2883 ;
  assign n4509 = n4508 ^ n4453 ;
  assign n4511 = n4510 ^ n4509 ;
  assign n4450 = n4306 ^ n4297 ;
  assign n4451 = ~n4303 & n4450 ;
  assign n4452 = n4451 ^ n4306 ;
  assign n4512 = n4511 ^ n4452 ;
  assign n4513 = n4512 ^ x29 ;
  assign n4449 = x76 & n2581 ;
  assign n4514 = n4513 ^ n4449 ;
  assign n4448 = x78 & n2422 ;
  assign n4515 = n4514 ^ n4448 ;
  assign n4447 = ~n1025 & n2423 ;
  assign n4516 = n4515 ^ n4447 ;
  assign n4518 = n4517 ^ n4516 ;
  assign n4522 = n4521 ^ n4518 ;
  assign n4523 = n4522 ^ x26 ;
  assign n4446 = x79 & n2018 ;
  assign n4524 = n4523 ^ n4446 ;
  assign n4445 = x81 & n2021 ;
  assign n4525 = n4524 ^ n4445 ;
  assign n4444 = n1305 & n2022 ;
  assign n4526 = n4525 ^ n4444 ;
  assign n4528 = n4527 ^ n4526 ;
  assign n4532 = n4531 ^ n4528 ;
  assign n4533 = n4532 ^ x23 ;
  assign n4443 = x82 & n1658 ;
  assign n4534 = n4533 ^ n4443 ;
  assign n4442 = x84 & n1661 ;
  assign n4535 = n4534 ^ n4442 ;
  assign n4441 = n1624 & n1662 ;
  assign n4536 = n4535 ^ n4441 ;
  assign n4538 = n4537 ^ n4536 ;
  assign n4542 = n4541 ^ n4538 ;
  assign n4543 = n4542 ^ x20 ;
  assign n4440 = x85 & n1327 ;
  assign n4544 = n4543 ^ n4440 ;
  assign n4439 = x87 & n1330 ;
  assign n4545 = n4544 ^ n4439 ;
  assign n4438 = n1331 & n1982 ;
  assign n4546 = n4545 ^ n4438 ;
  assign n4548 = n4547 ^ n4546 ;
  assign n4435 = n4337 ^ n4328 ;
  assign n4436 = ~n4334 & n4435 ;
  assign n4437 = n4436 ^ n4337 ;
  assign n4549 = n4548 ^ n4437 ;
  assign n4550 = n4549 ^ x17 ;
  assign n4434 = x88 & n1050 ;
  assign n4551 = n4550 ^ n4434 ;
  assign n4433 = x90 & n1053 ;
  assign n4552 = n4551 ^ n4433 ;
  assign n4432 = n1054 & n2386 ;
  assign n4553 = n4552 ^ n4432 ;
  assign n4555 = n4554 ^ n4553 ;
  assign n4559 = n4558 ^ n4555 ;
  assign n4560 = n4559 ^ x14 ;
  assign n4431 = x91 & n877 ;
  assign n4561 = n4560 ^ n4431 ;
  assign n4430 = x93 & n782 ;
  assign n4562 = n4561 ^ n4430 ;
  assign n4429 = n783 & n2836 ;
  assign n4563 = n4562 ^ n4429 ;
  assign n4565 = n4564 ^ n4563 ;
  assign n4426 = n4354 ^ n4345 ;
  assign n4427 = ~n4351 & n4426 ;
  assign n4428 = n4427 ^ n4354 ;
  assign n4566 = n4565 ^ n4428 ;
  assign n4567 = n4566 ^ x11 ;
  assign n4425 = x94 & n647 ;
  assign n4568 = n4567 ^ n4425 ;
  assign n4424 = x96 & ~n572 ;
  assign n4569 = n4568 ^ n4424 ;
  assign n4423 = ~n573 & n3323 ;
  assign n4570 = n4569 ^ n4423 ;
  assign n4572 = n4571 ^ n4570 ;
  assign n4420 = n4364 ^ n4355 ;
  assign n4421 = ~n4361 & n4420 ;
  assign n4422 = n4421 ^ n4364 ;
  assign n4573 = n4572 ^ n4422 ;
  assign n4574 = n4573 ^ x8 ;
  assign n4419 = x97 & n446 ;
  assign n4575 = n4574 ^ n4419 ;
  assign n4418 = x99 & n383 ;
  assign n4576 = n4575 ^ n4418 ;
  assign n4417 = n384 & n3843 ;
  assign n4577 = n4576 ^ n4417 ;
  assign n4579 = n4578 ^ n4577 ;
  assign n4414 = n4374 ^ n4365 ;
  assign n4415 = ~n4371 & n4414 ;
  assign n4416 = n4415 ^ n4374 ;
  assign n4580 = n4579 ^ n4416 ;
  assign n4581 = n4580 ^ x5 ;
  assign n4413 = x100 & n234 ;
  assign n4582 = n4581 ^ n4413 ;
  assign n4412 = x102 & n230 ;
  assign n4583 = n4582 ^ n4412 ;
  assign n4410 = n3826 ^ x102 ;
  assign n4411 = n231 & n4410 ;
  assign n4584 = n4583 ^ n4411 ;
  assign n4586 = n4585 ^ n4584 ;
  assign n4590 = n4589 ^ n4586 ;
  assign n4395 = x104 & ~n4197 ;
  assign n4394 = ~x104 & ~n4196 ;
  assign n4396 = n4395 ^ n4394 ;
  assign n4398 = x105 ^ x1 ;
  assign n4397 = x105 ^ x2 ;
  assign n4399 = n4398 ^ n4397 ;
  assign n4400 = n4396 & n4399 ;
  assign n4401 = n4400 ^ n4398 ;
  assign n4591 = n4590 ^ n4401 ;
  assign n4405 = x2 & x103 ;
  assign n4406 = n4405 ^ x104 ;
  assign n4407 = ~x1 & n4406 ;
  assign n4402 = n4401 ^ n4199 ;
  assign n4408 = n4407 ^ n4402 ;
  assign n4409 = ~x0 & n4408 ;
  assign n4592 = n4591 ^ n4409 ;
  assign n4389 = n4387 ^ n4382 ;
  assign n4390 = ~n4384 & n4389 ;
  assign n4391 = n4390 ^ n4387 ;
  assign n4593 = n4592 ^ n4391 ;
  assign n4789 = n4590 ^ n4391 ;
  assign n4790 = n4592 & n4789 ;
  assign n4791 = n4790 ^ n4590 ;
  assign n4784 = x102 & n227 ;
  assign n4776 = n4573 ^ n4416 ;
  assign n4777 = n4579 & n4776 ;
  assign n4778 = n4777 ^ n4573 ;
  assign n4774 = x99 & n390 ;
  assign n4766 = n4566 ^ n4422 ;
  assign n4767 = n4572 & n4766 ;
  assign n4768 = n4767 ^ n4566 ;
  assign n4764 = x96 & n578 ;
  assign n4756 = n4559 ^ n4428 ;
  assign n4757 = n4565 & n4756 ;
  assign n4758 = n4757 ^ n4559 ;
  assign n4754 = x93 & n788 ;
  assign n4747 = x90 & n1058 ;
  assign n4739 = n4542 ^ n4437 ;
  assign n4740 = n4548 & n4739 ;
  assign n4741 = n4740 ^ n4542 ;
  assign n4737 = x87 & n1335 ;
  assign n4730 = x84 & n1666 ;
  assign n4723 = x81 & n2014 ;
  assign n4716 = x78 & n2429 ;
  assign n4708 = n4505 ^ n4452 ;
  assign n4709 = n4511 & n4708 ;
  assign n4710 = n4709 ^ n4505 ;
  assign n4706 = x75 & n2887 ;
  assign n4699 = x72 & n3383 ;
  assign n4692 = x69 & n3924 ;
  assign n4684 = x66 & n4467 ;
  assign n4682 = x65 & n4474 ;
  assign n4678 = ~n153 & n4470 ;
  assign n4679 = n4678 ^ x67 ;
  assign n4680 = n4093 & n4679 ;
  assign n4681 = n4680 ^ x41 ;
  assign n4683 = n4682 ^ n4681 ;
  assign n4685 = n4684 ^ n4683 ;
  assign n4672 = x41 & ~n4484 ;
  assign n4673 = ~n4466 & n4672 ;
  assign n4686 = n4685 ^ n4673 ;
  assign n4670 = x42 ^ x41 ;
  assign n4671 = x64 & n4670 ;
  assign n4687 = n4686 ^ n4671 ;
  assign n4688 = n4687 ^ x38 ;
  assign n4669 = x68 & n3916 ;
  assign n4689 = n4688 ^ n4669 ;
  assign n4668 = x70 & n3919 ;
  assign n4690 = n4689 ^ n4668 ;
  assign n4667 = ~n436 & n3920 ;
  assign n4691 = n4690 ^ n4667 ;
  assign n4693 = n4692 ^ n4691 ;
  assign n4664 = n4497 ^ n4493 ;
  assign n4665 = ~n4494 & n4664 ;
  assign n4666 = n4665 ^ n4497 ;
  assign n4694 = n4693 ^ n4666 ;
  assign n4695 = n4694 ^ x35 ;
  assign n4663 = x71 & n3375 ;
  assign n4696 = n4695 ^ n4663 ;
  assign n4662 = x73 & n3378 ;
  assign n4697 = n4696 ^ n4662 ;
  assign n4661 = n633 & n3379 ;
  assign n4698 = n4697 ^ n4661 ;
  assign n4700 = n4699 ^ n4698 ;
  assign n4658 = n4498 ^ n4458 ;
  assign n4659 = n4504 & n4658 ;
  assign n4660 = n4659 ^ n4498 ;
  assign n4701 = n4700 ^ n4660 ;
  assign n4702 = n4701 ^ x32 ;
  assign n4657 = x74 & n2879 ;
  assign n4703 = n4702 ^ n4657 ;
  assign n4656 = x76 & n2882 ;
  assign n4704 = n4703 ^ n4656 ;
  assign n4655 = ~n853 & n2883 ;
  assign n4705 = n4704 ^ n4655 ;
  assign n4707 = n4706 ^ n4705 ;
  assign n4711 = n4710 ^ n4707 ;
  assign n4712 = n4711 ^ x29 ;
  assign n4654 = x77 & n2581 ;
  assign n4713 = n4712 ^ n4654 ;
  assign n4653 = x79 & n2422 ;
  assign n4714 = n4713 ^ n4653 ;
  assign n4652 = n1118 & n2423 ;
  assign n4715 = n4714 ^ n4652 ;
  assign n4717 = n4716 ^ n4715 ;
  assign n4649 = n4521 ^ n4512 ;
  assign n4650 = ~n4518 & n4649 ;
  assign n4651 = n4650 ^ n4521 ;
  assign n4718 = n4717 ^ n4651 ;
  assign n4719 = n4718 ^ x26 ;
  assign n4648 = x80 & n2018 ;
  assign n4720 = n4719 ^ n4648 ;
  assign n4647 = x82 & n2021 ;
  assign n4721 = n4720 ^ n4647 ;
  assign n4646 = n1411 & n2022 ;
  assign n4722 = n4721 ^ n4646 ;
  assign n4724 = n4723 ^ n4722 ;
  assign n4643 = n4531 ^ n4522 ;
  assign n4644 = ~n4528 & n4643 ;
  assign n4645 = n4644 ^ n4531 ;
  assign n4725 = n4724 ^ n4645 ;
  assign n4726 = n4725 ^ x23 ;
  assign n4642 = x83 & n1658 ;
  assign n4727 = n4726 ^ n4642 ;
  assign n4641 = x85 & n1661 ;
  assign n4728 = n4727 ^ n4641 ;
  assign n4640 = n1662 & n1743 ;
  assign n4729 = n4728 ^ n4640 ;
  assign n4731 = n4730 ^ n4729 ;
  assign n4637 = n4541 ^ n4532 ;
  assign n4638 = ~n4538 & n4637 ;
  assign n4639 = n4638 ^ n4541 ;
  assign n4732 = n4731 ^ n4639 ;
  assign n4733 = n4732 ^ x20 ;
  assign n4636 = x86 & n1327 ;
  assign n4734 = n4733 ^ n4636 ;
  assign n4635 = x88 & n1330 ;
  assign n4735 = n4734 ^ n4635 ;
  assign n4634 = n1331 & n2119 ;
  assign n4736 = n4735 ^ n4634 ;
  assign n4738 = n4737 ^ n4736 ;
  assign n4742 = n4741 ^ n4738 ;
  assign n4743 = n4742 ^ x17 ;
  assign n4633 = x89 & n1050 ;
  assign n4744 = n4743 ^ n4633 ;
  assign n4632 = x91 & n1053 ;
  assign n4745 = n4744 ^ n4632 ;
  assign n4631 = n1054 & n2542 ;
  assign n4746 = n4745 ^ n4631 ;
  assign n4748 = n4747 ^ n4746 ;
  assign n4628 = n4558 ^ n4549 ;
  assign n4629 = ~n4555 & n4628 ;
  assign n4630 = n4629 ^ n4558 ;
  assign n4749 = n4748 ^ n4630 ;
  assign n4750 = n4749 ^ x14 ;
  assign n4627 = x92 & n877 ;
  assign n4751 = n4750 ^ n4627 ;
  assign n4626 = x94 & n782 ;
  assign n4752 = n4751 ^ n4626 ;
  assign n4625 = n783 & n2997 ;
  assign n4753 = n4752 ^ n4625 ;
  assign n4755 = n4754 ^ n4753 ;
  assign n4759 = n4758 ^ n4755 ;
  assign n4760 = n4759 ^ x11 ;
  assign n4624 = x95 & n647 ;
  assign n4761 = n4760 ^ n4624 ;
  assign n4623 = x97 & ~n572 ;
  assign n4762 = n4761 ^ n4623 ;
  assign n4622 = ~n573 & n3494 ;
  assign n4763 = n4762 ^ n4622 ;
  assign n4765 = n4764 ^ n4763 ;
  assign n4769 = n4768 ^ n4765 ;
  assign n4770 = n4769 ^ x8 ;
  assign n4621 = x98 & n446 ;
  assign n4771 = n4770 ^ n4621 ;
  assign n4620 = x100 & n383 ;
  assign n4772 = n4771 ^ n4620 ;
  assign n4619 = n384 & n4034 ;
  assign n4773 = n4772 ^ n4619 ;
  assign n4775 = n4774 ^ n4773 ;
  assign n4779 = n4778 ^ n4775 ;
  assign n4780 = n4779 ^ x5 ;
  assign n4618 = x101 & n234 ;
  assign n4781 = n4780 ^ n4618 ;
  assign n4617 = x103 & n230 ;
  assign n4782 = n4781 ^ n4617 ;
  assign n4615 = n4020 ^ x103 ;
  assign n4616 = n231 & ~n4615 ;
  assign n4783 = n4782 ^ n4616 ;
  assign n4785 = n4784 ^ n4783 ;
  assign n4612 = n4589 ^ n4580 ;
  assign n4613 = ~n4586 & n4612 ;
  assign n4614 = n4613 ^ n4589 ;
  assign n4786 = n4785 ^ n4614 ;
  assign n4597 = ~x105 & ~n4395 ;
  assign n4596 = x105 & ~n4394 ;
  assign n4598 = n4597 ^ n4596 ;
  assign n4600 = x106 ^ x1 ;
  assign n4599 = x106 ^ x2 ;
  assign n4601 = n4600 ^ n4599 ;
  assign n4602 = n4598 & n4601 ;
  assign n4603 = n4602 ^ n4600 ;
  assign n4787 = n4786 ^ n4603 ;
  assign n4607 = x2 & x104 ;
  assign n4608 = n4607 ^ x105 ;
  assign n4609 = ~x1 & n4608 ;
  assign n4604 = n4603 ^ n4397 ;
  assign n4610 = n4609 ^ n4604 ;
  assign n4611 = ~x0 & n4610 ;
  assign n4788 = n4787 ^ n4611 ;
  assign n4792 = n4791 ^ n4788 ;
  assign n4991 = n4779 ^ n4614 ;
  assign n4992 = n4785 & n4991 ;
  assign n4993 = n4992 ^ n4779 ;
  assign n4989 = x103 & n227 ;
  assign n4982 = x100 & n390 ;
  assign n4975 = x97 & n578 ;
  assign n4968 = x94 & n788 ;
  assign n4960 = n4742 ^ n4630 ;
  assign n4961 = n4748 & n4960 ;
  assign n4962 = n4961 ^ n4742 ;
  assign n4958 = x91 & n1058 ;
  assign n4951 = x88 & n1335 ;
  assign n4943 = n4725 ^ n4639 ;
  assign n4944 = n4731 & n4943 ;
  assign n4945 = n4944 ^ n4725 ;
  assign n4941 = x85 & n1666 ;
  assign n4933 = n4718 ^ n4645 ;
  assign n4934 = n4724 & n4933 ;
  assign n4935 = n4934 ^ n4718 ;
  assign n4931 = x82 & n2014 ;
  assign n4923 = n4711 ^ n4651 ;
  assign n4924 = n4717 & n4923 ;
  assign n4925 = n4924 ^ n4711 ;
  assign n4921 = x79 & n2429 ;
  assign n4914 = x76 & n2887 ;
  assign n4906 = n4694 ^ n4660 ;
  assign n4907 = n4700 & n4906 ;
  assign n4908 = n4907 ^ n4694 ;
  assign n4904 = x73 & n3383 ;
  assign n4896 = n4687 ^ n4666 ;
  assign n4897 = n4693 & n4896 ;
  assign n4898 = n4897 ^ n4687 ;
  assign n4894 = x70 & n3924 ;
  assign n4884 = x66 & n4474 ;
  assign n4883 = x68 & n4471 ;
  assign n4885 = n4884 ^ n4883 ;
  assign n4886 = n4885 ^ x41 ;
  assign n4882 = ~n340 & n4472 ;
  assign n4887 = n4886 ^ n4882 ;
  assign n4881 = x67 & n4467 ;
  assign n4888 = n4887 ^ n4881 ;
  assign n4875 = x41 & x42 ;
  assign n4876 = n4875 ^ x43 ;
  assign n4877 = ~x64 & n4876 ;
  assign n4871 = x43 ^ x41 ;
  assign n4878 = n4877 ^ n4871 ;
  assign n4869 = x65 ^ x42 ;
  assign n4870 = n4670 & ~n4869 ;
  assign n4879 = n4878 ^ n4870 ;
  assign n4866 = n4685 & n4686 ;
  assign n4867 = ~n4671 & n4866 ;
  assign n4868 = n4867 ^ n4685 ;
  assign n4880 = n4879 ^ n4868 ;
  assign n4889 = n4888 ^ n4880 ;
  assign n4890 = n4889 ^ x38 ;
  assign n4865 = x69 & n3916 ;
  assign n4891 = n4890 ^ n4865 ;
  assign n4864 = x71 & n3919 ;
  assign n4892 = n4891 ^ n4864 ;
  assign n4863 = ~n493 & n3920 ;
  assign n4893 = n4892 ^ n4863 ;
  assign n4895 = n4894 ^ n4893 ;
  assign n4899 = n4898 ^ n4895 ;
  assign n4900 = n4899 ^ x35 ;
  assign n4862 = x72 & n3375 ;
  assign n4901 = n4900 ^ n4862 ;
  assign n4861 = x74 & n3378 ;
  assign n4902 = n4901 ^ n4861 ;
  assign n4860 = n699 & n3379 ;
  assign n4903 = n4902 ^ n4860 ;
  assign n4905 = n4904 ^ n4903 ;
  assign n4909 = n4908 ^ n4905 ;
  assign n4910 = n4909 ^ x32 ;
  assign n4859 = x75 & n2879 ;
  assign n4911 = n4910 ^ n4859 ;
  assign n4858 = x77 & n2882 ;
  assign n4912 = n4911 ^ n4858 ;
  assign n4857 = ~n939 & n2883 ;
  assign n4913 = n4912 ^ n4857 ;
  assign n4915 = n4914 ^ n4913 ;
  assign n4854 = n4710 ^ n4701 ;
  assign n4855 = ~n4707 & n4854 ;
  assign n4856 = n4855 ^ n4710 ;
  assign n4916 = n4915 ^ n4856 ;
  assign n4917 = n4916 ^ x29 ;
  assign n4853 = x78 & n2581 ;
  assign n4918 = n4917 ^ n4853 ;
  assign n4852 = x80 & n2422 ;
  assign n4919 = n4918 ^ n4852 ;
  assign n4851 = n1206 & n2423 ;
  assign n4920 = n4919 ^ n4851 ;
  assign n4922 = n4921 ^ n4920 ;
  assign n4926 = n4925 ^ n4922 ;
  assign n4927 = n4926 ^ x26 ;
  assign n4850 = x81 & n2018 ;
  assign n4928 = n4927 ^ n4850 ;
  assign n4849 = x83 & n2021 ;
  assign n4929 = n4928 ^ n4849 ;
  assign n4848 = n1512 & n2022 ;
  assign n4930 = n4929 ^ n4848 ;
  assign n4932 = n4931 ^ n4930 ;
  assign n4936 = n4935 ^ n4932 ;
  assign n4937 = n4936 ^ x23 ;
  assign n4847 = x84 & n1658 ;
  assign n4938 = n4937 ^ n4847 ;
  assign n4846 = x86 & n1661 ;
  assign n4939 = n4938 ^ n4846 ;
  assign n4845 = n1662 & n1857 ;
  assign n4940 = n4939 ^ n4845 ;
  assign n4942 = n4941 ^ n4940 ;
  assign n4946 = n4945 ^ n4942 ;
  assign n4947 = n4946 ^ x20 ;
  assign n4844 = x87 & n1327 ;
  assign n4948 = n4947 ^ n4844 ;
  assign n4843 = x89 & n1330 ;
  assign n4949 = n4948 ^ n4843 ;
  assign n4842 = n1331 & n2249 ;
  assign n4950 = n4949 ^ n4842 ;
  assign n4952 = n4951 ^ n4950 ;
  assign n4839 = n4741 ^ n4732 ;
  assign n4840 = ~n4738 & n4839 ;
  assign n4841 = n4840 ^ n4741 ;
  assign n4953 = n4952 ^ n4841 ;
  assign n4954 = n4953 ^ x17 ;
  assign n4838 = x90 & n1050 ;
  assign n4955 = n4954 ^ n4838 ;
  assign n4837 = x92 & n1053 ;
  assign n4956 = n4955 ^ n4837 ;
  assign n4836 = n1054 & n2684 ;
  assign n4957 = n4956 ^ n4836 ;
  assign n4959 = n4958 ^ n4957 ;
  assign n4963 = n4962 ^ n4959 ;
  assign n4964 = n4963 ^ x14 ;
  assign n4835 = x93 & n877 ;
  assign n4965 = n4964 ^ n4835 ;
  assign n4834 = x95 & n782 ;
  assign n4966 = n4965 ^ n4834 ;
  assign n4833 = n783 & n3159 ;
  assign n4967 = n4966 ^ n4833 ;
  assign n4969 = n4968 ^ n4967 ;
  assign n4830 = n4758 ^ n4749 ;
  assign n4831 = ~n4755 & n4830 ;
  assign n4832 = n4831 ^ n4758 ;
  assign n4970 = n4969 ^ n4832 ;
  assign n4971 = n4970 ^ x11 ;
  assign n4829 = x96 & n647 ;
  assign n4972 = n4971 ^ n4829 ;
  assign n4828 = x98 & ~n572 ;
  assign n4973 = n4972 ^ n4828 ;
  assign n4827 = ~n573 & n3660 ;
  assign n4974 = n4973 ^ n4827 ;
  assign n4976 = n4975 ^ n4974 ;
  assign n4824 = n4768 ^ n4759 ;
  assign n4825 = ~n4765 & n4824 ;
  assign n4826 = n4825 ^ n4768 ;
  assign n4977 = n4976 ^ n4826 ;
  assign n4978 = n4977 ^ x8 ;
  assign n4823 = x99 & n446 ;
  assign n4979 = n4978 ^ n4823 ;
  assign n4822 = x101 & n383 ;
  assign n4980 = n4979 ^ n4822 ;
  assign n4821 = n384 & n4215 ;
  assign n4981 = n4980 ^ n4821 ;
  assign n4983 = n4982 ^ n4981 ;
  assign n4818 = n4778 ^ n4769 ;
  assign n4819 = ~n4775 & n4818 ;
  assign n4820 = n4819 ^ n4778 ;
  assign n4984 = n4983 ^ n4820 ;
  assign n4985 = n4984 ^ x5 ;
  assign n4817 = x102 & n234 ;
  assign n4986 = n4985 ^ n4817 ;
  assign n4816 = x104 & n230 ;
  assign n4987 = n4986 ^ n4816 ;
  assign n4814 = n4198 ^ x104 ;
  assign n4815 = n231 & ~n4814 ;
  assign n4988 = n4987 ^ n4815 ;
  assign n4990 = n4989 ^ n4988 ;
  assign n4994 = n4993 ^ n4990 ;
  assign n4799 = x106 & ~n4597 ;
  assign n4798 = ~x106 & ~n4596 ;
  assign n4800 = n4799 ^ n4798 ;
  assign n4802 = x107 ^ x1 ;
  assign n4801 = x107 ^ x2 ;
  assign n4803 = n4802 ^ n4801 ;
  assign n4804 = n4800 & n4803 ;
  assign n4805 = n4804 ^ n4802 ;
  assign n4995 = n4994 ^ n4805 ;
  assign n4809 = x2 & x105 ;
  assign n4810 = n4809 ^ x106 ;
  assign n4811 = ~x1 & n4810 ;
  assign n4806 = n4805 ^ n4599 ;
  assign n4812 = n4811 ^ n4806 ;
  assign n4813 = ~x0 & n4812 ;
  assign n4996 = n4995 ^ n4813 ;
  assign n4793 = n4791 ^ n4786 ;
  assign n4794 = ~n4788 & n4793 ;
  assign n4795 = n4794 ^ n4791 ;
  assign n4997 = n4996 ^ n4795 ;
  assign n5211 = n4994 ^ n4795 ;
  assign n5212 = n4996 & n5211 ;
  assign n5213 = n5212 ^ n4994 ;
  assign n5206 = x104 & n227 ;
  assign n5198 = n4977 ^ n4820 ;
  assign n5199 = n4983 & n5198 ;
  assign n5200 = n5199 ^ n4977 ;
  assign n5196 = x101 & n390 ;
  assign n5188 = n4970 ^ n4826 ;
  assign n5189 = n4976 & n5188 ;
  assign n5190 = n5189 ^ n4970 ;
  assign n5186 = x98 & n578 ;
  assign n5178 = n4963 ^ n4832 ;
  assign n5179 = n4969 & n5178 ;
  assign n5180 = n5179 ^ n4963 ;
  assign n5176 = x95 & n788 ;
  assign n5169 = x92 & n1058 ;
  assign n5161 = n4946 ^ n4841 ;
  assign n5162 = n4952 & n5161 ;
  assign n5163 = n5162 ^ n4946 ;
  assign n5159 = x89 & n1335 ;
  assign n5152 = x86 & n1666 ;
  assign n5145 = x83 & n2014 ;
  assign n5138 = x80 & n2429 ;
  assign n5130 = n4909 ^ n4856 ;
  assign n5131 = n4915 & n5130 ;
  assign n5132 = n5131 ^ n4909 ;
  assign n5128 = x77 & n2887 ;
  assign n5120 = x71 & n3924 ;
  assign n5113 = x68 & n4467 ;
  assign n5106 = x44 & ~n4671 ;
  assign n5107 = ~n4879 & n5106 ;
  assign n4873 = x43 ^ x42 ;
  assign n5102 = ~n4670 & n4873 ;
  assign n5103 = x65 & n5102 ;
  assign n5091 = x44 ^ x43 ;
  assign n5097 = n4670 & ~n5091 ;
  assign n5098 = n5097 ^ n4670 ;
  assign n5099 = ~n150 & n5098 ;
  assign n5096 = x66 & n4670 ;
  assign n5100 = n5099 ^ n5096 ;
  assign n5101 = n5100 ^ x44 ;
  assign n5104 = n5103 ^ n5101 ;
  assign n5092 = x44 ^ x42 ;
  assign n5093 = ~n4670 & n5092 ;
  assign n5094 = n5091 & n5093 ;
  assign n5095 = x64 & n5094 ;
  assign n5105 = n5104 ^ n5095 ;
  assign n5108 = n5107 ^ n5105 ;
  assign n5109 = n5108 ^ x41 ;
  assign n5090 = x67 & n4474 ;
  assign n5110 = n5109 ^ n5090 ;
  assign n5089 = x69 & n4471 ;
  assign n5111 = n5110 ^ n5089 ;
  assign n5088 = ~n375 & n4472 ;
  assign n5112 = n5111 ^ n5088 ;
  assign n5114 = n5113 ^ n5112 ;
  assign n5085 = n4888 ^ n4879 ;
  assign n5086 = ~n4880 & n5085 ;
  assign n5087 = n5086 ^ n4888 ;
  assign n5115 = n5114 ^ n5087 ;
  assign n5116 = n5115 ^ x38 ;
  assign n5084 = x70 & n3916 ;
  assign n5117 = n5116 ^ n5084 ;
  assign n5083 = x72 & n3919 ;
  assign n5118 = n5117 ^ n5083 ;
  assign n5082 = n556 & n3920 ;
  assign n5119 = n5118 ^ n5082 ;
  assign n5121 = n5120 ^ n5119 ;
  assign n5079 = n4898 ^ n4889 ;
  assign n5080 = ~n4895 & n5079 ;
  assign n5081 = n5080 ^ n4898 ;
  assign n5122 = n5121 ^ n5081 ;
  assign n5069 = x73 & n3375 ;
  assign n5068 = x75 & n3378 ;
  assign n5070 = n5069 ^ n5068 ;
  assign n5071 = n5070 ^ x35 ;
  assign n5067 = ~n774 & n3379 ;
  assign n5072 = n5071 ^ n5067 ;
  assign n5066 = x74 & n3383 ;
  assign n5073 = n5072 ^ n5066 ;
  assign n5074 = n5073 ^ n4908 ;
  assign n5075 = n5074 ^ n4899 ;
  assign n5076 = n5075 ^ n5073 ;
  assign n5077 = ~n4905 & n5076 ;
  assign n5078 = n5077 ^ n5074 ;
  assign n5123 = n5122 ^ n5078 ;
  assign n5124 = n5123 ^ x32 ;
  assign n5065 = x76 & n2879 ;
  assign n5125 = n5124 ^ n5065 ;
  assign n5064 = x78 & n2882 ;
  assign n5126 = n5125 ^ n5064 ;
  assign n5063 = ~n1025 & n2883 ;
  assign n5127 = n5126 ^ n5063 ;
  assign n5129 = n5128 ^ n5127 ;
  assign n5133 = n5132 ^ n5129 ;
  assign n5134 = n5133 ^ x29 ;
  assign n5062 = x79 & n2581 ;
  assign n5135 = n5134 ^ n5062 ;
  assign n5061 = x81 & n2422 ;
  assign n5136 = n5135 ^ n5061 ;
  assign n5060 = n1305 & n2423 ;
  assign n5137 = n5136 ^ n5060 ;
  assign n5139 = n5138 ^ n5137 ;
  assign n5057 = n4925 ^ n4916 ;
  assign n5058 = ~n4922 & n5057 ;
  assign n5059 = n5058 ^ n4925 ;
  assign n5140 = n5139 ^ n5059 ;
  assign n5141 = n5140 ^ x26 ;
  assign n5056 = x82 & n2018 ;
  assign n5142 = n5141 ^ n5056 ;
  assign n5055 = x84 & n2021 ;
  assign n5143 = n5142 ^ n5055 ;
  assign n5054 = n1624 & n2022 ;
  assign n5144 = n5143 ^ n5054 ;
  assign n5146 = n5145 ^ n5144 ;
  assign n5051 = n4935 ^ n4926 ;
  assign n5052 = ~n4932 & n5051 ;
  assign n5053 = n5052 ^ n4935 ;
  assign n5147 = n5146 ^ n5053 ;
  assign n5148 = n5147 ^ x23 ;
  assign n5050 = x85 & n1658 ;
  assign n5149 = n5148 ^ n5050 ;
  assign n5049 = x87 & n1661 ;
  assign n5150 = n5149 ^ n5049 ;
  assign n5048 = n1662 & n1982 ;
  assign n5151 = n5150 ^ n5048 ;
  assign n5153 = n5152 ^ n5151 ;
  assign n5045 = n4945 ^ n4936 ;
  assign n5046 = ~n4942 & n5045 ;
  assign n5047 = n5046 ^ n4945 ;
  assign n5154 = n5153 ^ n5047 ;
  assign n5155 = n5154 ^ x20 ;
  assign n5044 = x88 & n1327 ;
  assign n5156 = n5155 ^ n5044 ;
  assign n5043 = x90 & n1330 ;
  assign n5157 = n5156 ^ n5043 ;
  assign n5042 = n1331 & n2386 ;
  assign n5158 = n5157 ^ n5042 ;
  assign n5160 = n5159 ^ n5158 ;
  assign n5164 = n5163 ^ n5160 ;
  assign n5165 = n5164 ^ x17 ;
  assign n5041 = x91 & n1050 ;
  assign n5166 = n5165 ^ n5041 ;
  assign n5040 = x93 & n1053 ;
  assign n5167 = n5166 ^ n5040 ;
  assign n5039 = n1054 & n2836 ;
  assign n5168 = n5167 ^ n5039 ;
  assign n5170 = n5169 ^ n5168 ;
  assign n5036 = n4962 ^ n4953 ;
  assign n5037 = ~n4959 & n5036 ;
  assign n5038 = n5037 ^ n4962 ;
  assign n5171 = n5170 ^ n5038 ;
  assign n5172 = n5171 ^ x14 ;
  assign n5035 = x94 & n877 ;
  assign n5173 = n5172 ^ n5035 ;
  assign n5034 = x96 & n782 ;
  assign n5174 = n5173 ^ n5034 ;
  assign n5033 = n783 & n3323 ;
  assign n5175 = n5174 ^ n5033 ;
  assign n5177 = n5176 ^ n5175 ;
  assign n5181 = n5180 ^ n5177 ;
  assign n5182 = n5181 ^ x11 ;
  assign n5032 = x97 & n647 ;
  assign n5183 = n5182 ^ n5032 ;
  assign n5031 = x99 & ~n572 ;
  assign n5184 = n5183 ^ n5031 ;
  assign n5030 = ~n573 & n3843 ;
  assign n5185 = n5184 ^ n5030 ;
  assign n5187 = n5186 ^ n5185 ;
  assign n5191 = n5190 ^ n5187 ;
  assign n5192 = n5191 ^ x8 ;
  assign n5029 = x100 & n446 ;
  assign n5193 = n5192 ^ n5029 ;
  assign n5028 = x102 & n383 ;
  assign n5194 = n5193 ^ n5028 ;
  assign n5027 = n384 & n4410 ;
  assign n5195 = n5194 ^ n5027 ;
  assign n5197 = n5196 ^ n5195 ;
  assign n5201 = n5200 ^ n5197 ;
  assign n5202 = n5201 ^ x5 ;
  assign n5026 = x103 & n234 ;
  assign n5203 = n5202 ^ n5026 ;
  assign n5025 = x105 & n230 ;
  assign n5204 = n5203 ^ n5025 ;
  assign n5023 = n4396 ^ x105 ;
  assign n5024 = n231 & ~n5023 ;
  assign n5205 = n5204 ^ n5024 ;
  assign n5207 = n5206 ^ n5205 ;
  assign n5020 = n4993 ^ n4984 ;
  assign n5021 = ~n4990 & n5020 ;
  assign n5022 = n5021 ^ n4993 ;
  assign n5208 = n5207 ^ n5022 ;
  assign n4998 = x107 ^ x106 ;
  assign n5004 = x107 & n4598 ;
  assign n5005 = n5004 ^ n4597 ;
  assign n5006 = n4998 & ~n5005 ;
  assign n5008 = x108 ^ x1 ;
  assign n5007 = x108 ^ x2 ;
  assign n5009 = n5008 ^ n5007 ;
  assign n5010 = ~n5006 & n5009 ;
  assign n5011 = n5010 ^ n5008 ;
  assign n5209 = n5208 ^ n5011 ;
  assign n5015 = x2 & x106 ;
  assign n5016 = n5015 ^ x107 ;
  assign n5017 = ~x1 & n5016 ;
  assign n5012 = n5011 ^ n4801 ;
  assign n5018 = n5017 ^ n5012 ;
  assign n5019 = ~x0 & n5018 ;
  assign n5210 = n5209 ^ n5019 ;
  assign n5214 = n5213 ^ n5210 ;
  assign n5420 = n5201 ^ n5022 ;
  assign n5421 = n5207 & n5420 ;
  assign n5422 = n5421 ^ n5201 ;
  assign n5418 = x105 & n227 ;
  assign n5411 = x102 & n390 ;
  assign n5404 = x99 & n578 ;
  assign n5397 = x96 & n788 ;
  assign n5389 = n5164 ^ n5038 ;
  assign n5390 = n5170 & n5389 ;
  assign n5391 = n5390 ^ n5164 ;
  assign n5387 = x93 & n1058 ;
  assign n5380 = x90 & n1335 ;
  assign n5372 = n5147 ^ n5047 ;
  assign n5373 = n5153 & n5372 ;
  assign n5374 = n5373 ^ n5147 ;
  assign n5370 = x87 & n1666 ;
  assign n5362 = n5140 ^ n5053 ;
  assign n5363 = n5146 & n5362 ;
  assign n5364 = n5363 ^ n5140 ;
  assign n5360 = x84 & n2014 ;
  assign n5352 = n5133 ^ n5059 ;
  assign n5353 = n5139 & n5352 ;
  assign n5354 = n5353 ^ n5133 ;
  assign n5350 = x81 & n2429 ;
  assign n5343 = x78 & n2887 ;
  assign n5336 = x75 & n3383 ;
  assign n5327 = n5108 ^ n5087 ;
  assign n5328 = n5114 & n5327 ;
  assign n5329 = n5328 ^ n5108 ;
  assign n5325 = x69 & n4467 ;
  assign n5314 = x65 & n5094 ;
  assign n5313 = x67 & n5097 ;
  assign n5315 = n5314 ^ n5313 ;
  assign n5316 = n5315 ^ x44 ;
  assign n5312 = ~n291 & n5098 ;
  assign n5317 = n5316 ^ n5312 ;
  assign n5311 = x66 & n5102 ;
  assign n5318 = n5317 ^ n5311 ;
  assign n5309 = x45 ^ x44 ;
  assign n5310 = x64 & n5309 ;
  assign n5319 = n5318 ^ n5310 ;
  assign n5308 = n5105 & n5107 ;
  assign n5320 = n5319 ^ n5308 ;
  assign n5321 = n5320 ^ x41 ;
  assign n5307 = x68 & n4474 ;
  assign n5322 = n5321 ^ n5307 ;
  assign n5306 = x70 & n4471 ;
  assign n5323 = n5322 ^ n5306 ;
  assign n5305 = ~n436 & n4472 ;
  assign n5324 = n5323 ^ n5305 ;
  assign n5326 = n5325 ^ n5324 ;
  assign n5330 = n5329 ^ n5326 ;
  assign n5302 = n5115 ^ n5081 ;
  assign n5303 = n5121 & n5302 ;
  assign n5295 = x71 & n3916 ;
  assign n5294 = x73 & n3919 ;
  assign n5296 = n5295 ^ n5294 ;
  assign n5297 = n5296 ^ x38 ;
  assign n5293 = n633 & n3920 ;
  assign n5298 = n5297 ^ n5293 ;
  assign n5292 = x72 & n3924 ;
  assign n5299 = n5298 ^ n5292 ;
  assign n5300 = n5299 ^ n5115 ;
  assign n5304 = n5303 ^ n5300 ;
  assign n5331 = n5330 ^ n5304 ;
  assign n5332 = n5331 ^ x35 ;
  assign n5291 = x74 & n3375 ;
  assign n5333 = n5332 ^ n5291 ;
  assign n5290 = x76 & n3378 ;
  assign n5334 = n5333 ^ n5290 ;
  assign n5289 = ~n853 & n3379 ;
  assign n5335 = n5334 ^ n5289 ;
  assign n5337 = n5336 ^ n5335 ;
  assign n5286 = n5122 ^ n5073 ;
  assign n5287 = n5078 & n5286 ;
  assign n5288 = n5287 ^ n5073 ;
  assign n5338 = n5337 ^ n5288 ;
  assign n5339 = n5338 ^ x32 ;
  assign n5285 = x77 & n2879 ;
  assign n5340 = n5339 ^ n5285 ;
  assign n5284 = x79 & n2882 ;
  assign n5341 = n5340 ^ n5284 ;
  assign n5283 = n1118 & n2883 ;
  assign n5342 = n5341 ^ n5283 ;
  assign n5344 = n5343 ^ n5342 ;
  assign n5280 = n5132 ^ n5123 ;
  assign n5281 = ~n5129 & n5280 ;
  assign n5282 = n5281 ^ n5132 ;
  assign n5345 = n5344 ^ n5282 ;
  assign n5346 = n5345 ^ x29 ;
  assign n5279 = x80 & n2581 ;
  assign n5347 = n5346 ^ n5279 ;
  assign n5278 = x82 & n2422 ;
  assign n5348 = n5347 ^ n5278 ;
  assign n5277 = n1411 & n2423 ;
  assign n5349 = n5348 ^ n5277 ;
  assign n5351 = n5350 ^ n5349 ;
  assign n5355 = n5354 ^ n5351 ;
  assign n5356 = n5355 ^ x26 ;
  assign n5276 = x83 & n2018 ;
  assign n5357 = n5356 ^ n5276 ;
  assign n5275 = x85 & n2021 ;
  assign n5358 = n5357 ^ n5275 ;
  assign n5274 = n1743 & n2022 ;
  assign n5359 = n5358 ^ n5274 ;
  assign n5361 = n5360 ^ n5359 ;
  assign n5365 = n5364 ^ n5361 ;
  assign n5366 = n5365 ^ x23 ;
  assign n5273 = x86 & n1658 ;
  assign n5367 = n5366 ^ n5273 ;
  assign n5272 = x88 & n1661 ;
  assign n5368 = n5367 ^ n5272 ;
  assign n5271 = n1662 & n2119 ;
  assign n5369 = n5368 ^ n5271 ;
  assign n5371 = n5370 ^ n5369 ;
  assign n5375 = n5374 ^ n5371 ;
  assign n5376 = n5375 ^ x20 ;
  assign n5270 = x89 & n1327 ;
  assign n5377 = n5376 ^ n5270 ;
  assign n5269 = x91 & n1330 ;
  assign n5378 = n5377 ^ n5269 ;
  assign n5268 = n1331 & n2542 ;
  assign n5379 = n5378 ^ n5268 ;
  assign n5381 = n5380 ^ n5379 ;
  assign n5265 = n5163 ^ n5154 ;
  assign n5266 = ~n5160 & n5265 ;
  assign n5267 = n5266 ^ n5163 ;
  assign n5382 = n5381 ^ n5267 ;
  assign n5383 = n5382 ^ x17 ;
  assign n5264 = x92 & n1050 ;
  assign n5384 = n5383 ^ n5264 ;
  assign n5263 = x94 & n1053 ;
  assign n5385 = n5384 ^ n5263 ;
  assign n5262 = n1054 & n2997 ;
  assign n5386 = n5385 ^ n5262 ;
  assign n5388 = n5387 ^ n5386 ;
  assign n5392 = n5391 ^ n5388 ;
  assign n5393 = n5392 ^ x14 ;
  assign n5261 = x95 & n877 ;
  assign n5394 = n5393 ^ n5261 ;
  assign n5260 = x97 & n782 ;
  assign n5395 = n5394 ^ n5260 ;
  assign n5259 = n783 & n3494 ;
  assign n5396 = n5395 ^ n5259 ;
  assign n5398 = n5397 ^ n5396 ;
  assign n5256 = n5180 ^ n5171 ;
  assign n5257 = ~n5177 & n5256 ;
  assign n5258 = n5257 ^ n5180 ;
  assign n5399 = n5398 ^ n5258 ;
  assign n5400 = n5399 ^ x11 ;
  assign n5255 = x98 & n647 ;
  assign n5401 = n5400 ^ n5255 ;
  assign n5254 = x100 & ~n572 ;
  assign n5402 = n5401 ^ n5254 ;
  assign n5253 = ~n573 & n4034 ;
  assign n5403 = n5402 ^ n5253 ;
  assign n5405 = n5404 ^ n5403 ;
  assign n5250 = n5190 ^ n5181 ;
  assign n5251 = ~n5187 & n5250 ;
  assign n5252 = n5251 ^ n5190 ;
  assign n5406 = n5405 ^ n5252 ;
  assign n5407 = n5406 ^ x8 ;
  assign n5249 = x101 & n446 ;
  assign n5408 = n5407 ^ n5249 ;
  assign n5248 = x103 & n383 ;
  assign n5409 = n5408 ^ n5248 ;
  assign n5247 = n384 & ~n4615 ;
  assign n5410 = n5409 ^ n5247 ;
  assign n5412 = n5411 ^ n5410 ;
  assign n5244 = n5200 ^ n5191 ;
  assign n5245 = ~n5197 & n5244 ;
  assign n5246 = n5245 ^ n5200 ;
  assign n5413 = n5412 ^ n5246 ;
  assign n5414 = n5413 ^ x5 ;
  assign n5243 = x104 & n234 ;
  assign n5415 = n5414 ^ n5243 ;
  assign n5242 = x106 & n230 ;
  assign n5416 = n5415 ^ n5242 ;
  assign n5240 = n4598 ^ x106 ;
  assign n5241 = n231 & ~n5240 ;
  assign n5417 = n5416 ^ n5241 ;
  assign n5419 = n5418 ^ n5417 ;
  assign n5423 = n5422 ^ n5419 ;
  assign n5218 = x108 ^ x107 ;
  assign n5224 = x108 & n4800 ;
  assign n5225 = n5224 ^ n4798 ;
  assign n5226 = n5218 & ~n5225 ;
  assign n5228 = x109 ^ x1 ;
  assign n5227 = x109 ^ x2 ;
  assign n5229 = n5228 ^ n5227 ;
  assign n5230 = ~n5226 & n5229 ;
  assign n5231 = n5230 ^ n5228 ;
  assign n5424 = n5423 ^ n5231 ;
  assign n5235 = x2 & x107 ;
  assign n5236 = n5235 ^ x108 ;
  assign n5237 = ~n255 & n5236 ;
  assign n5232 = n5231 ^ n5007 ;
  assign n5238 = n5237 ^ n5232 ;
  assign n5239 = ~x0 & n5238 ;
  assign n5425 = n5424 ^ n5239 ;
  assign n5215 = n5213 ^ n5208 ;
  assign n5216 = ~n5210 & n5215 ;
  assign n5217 = n5216 ^ n5213 ;
  assign n5426 = n5425 ^ n5217 ;
  assign n5643 = n5423 ^ n5217 ;
  assign n5644 = n5425 & n5643 ;
  assign n5645 = n5644 ^ n5423 ;
  assign n5638 = x106 & n227 ;
  assign n5630 = n5406 ^ n5246 ;
  assign n5631 = n5412 & n5630 ;
  assign n5632 = n5631 ^ n5406 ;
  assign n5628 = x103 & n390 ;
  assign n5620 = n5399 ^ n5252 ;
  assign n5621 = n5405 & n5620 ;
  assign n5622 = n5621 ^ n5399 ;
  assign n5618 = x100 & n578 ;
  assign n5610 = n5392 ^ n5258 ;
  assign n5611 = n5398 & n5610 ;
  assign n5612 = n5611 ^ n5392 ;
  assign n5608 = x97 & n788 ;
  assign n5601 = x94 & n1058 ;
  assign n5593 = n5375 ^ n5267 ;
  assign n5594 = n5381 & n5593 ;
  assign n5595 = n5594 ^ n5375 ;
  assign n5591 = x91 & n1335 ;
  assign n5584 = x88 & n1666 ;
  assign n5577 = x85 & n2014 ;
  assign n5570 = x82 & n2429 ;
  assign n5562 = n5338 ^ n5282 ;
  assign n5563 = n5344 & n5562 ;
  assign n5564 = n5563 ^ n5338 ;
  assign n5560 = x79 & n2887 ;
  assign n5552 = x73 & n3924 ;
  assign n5543 = ~n5310 & n5318 ;
  assign n5544 = ~n5308 & n5543 ;
  assign n5545 = n5544 ^ n5318 ;
  assign n5537 = x66 & n5094 ;
  assign n5536 = x68 & n5097 ;
  assign n5538 = n5537 ^ n5536 ;
  assign n5539 = n5538 ^ x44 ;
  assign n5535 = ~n340 & n5098 ;
  assign n5540 = n5539 ^ n5535 ;
  assign n5534 = x67 & n5102 ;
  assign n5541 = n5540 ^ n5534 ;
  assign n5529 = ~x44 & ~x45 ;
  assign n5530 = n5529 ^ n5309 ;
  assign n5531 = n5530 ^ x46 ;
  assign n5532 = ~x64 & ~n5531 ;
  assign n5523 = x65 ^ x45 ;
  assign n5526 = x65 ^ x44 ;
  assign n5527 = ~n5523 & n5526 ;
  assign n5524 = x46 ^ x44 ;
  assign n5528 = n5527 ^ n5524 ;
  assign n5533 = n5532 ^ n5528 ;
  assign n5542 = n5541 ^ n5533 ;
  assign n5546 = n5545 ^ n5542 ;
  assign n5513 = x69 & n4474 ;
  assign n5512 = x71 & n4471 ;
  assign n5514 = n5513 ^ n5512 ;
  assign n5515 = n5514 ^ x41 ;
  assign n5511 = ~n493 & n4472 ;
  assign n5516 = n5515 ^ n5511 ;
  assign n5510 = x70 & n4467 ;
  assign n5517 = n5516 ^ n5510 ;
  assign n5518 = n5517 ^ n5329 ;
  assign n5519 = n5518 ^ n5320 ;
  assign n5520 = n5519 ^ n5517 ;
  assign n5521 = ~n5326 & n5520 ;
  assign n5522 = n5521 ^ n5518 ;
  assign n5547 = n5546 ^ n5522 ;
  assign n5548 = n5547 ^ x38 ;
  assign n5509 = x72 & n3916 ;
  assign n5549 = n5548 ^ n5509 ;
  assign n5508 = x74 & n3919 ;
  assign n5550 = n5549 ^ n5508 ;
  assign n5507 = n699 & n3920 ;
  assign n5551 = n5550 ^ n5507 ;
  assign n5553 = n5552 ^ n5551 ;
  assign n5504 = n5330 ^ n5299 ;
  assign n5505 = n5304 & n5504 ;
  assign n5506 = n5505 ^ n5299 ;
  assign n5554 = n5553 ^ n5506 ;
  assign n5494 = x75 & n3375 ;
  assign n5493 = x77 & n3378 ;
  assign n5495 = n5494 ^ n5493 ;
  assign n5496 = n5495 ^ x35 ;
  assign n5492 = ~n939 & n3379 ;
  assign n5497 = n5496 ^ n5492 ;
  assign n5491 = x76 & n3383 ;
  assign n5498 = n5497 ^ n5491 ;
  assign n5499 = n5498 ^ n5331 ;
  assign n5500 = n5499 ^ n5288 ;
  assign n5501 = n5500 ^ n5498 ;
  assign n5502 = n5337 & n5501 ;
  assign n5503 = n5502 ^ n5499 ;
  assign n5555 = n5554 ^ n5503 ;
  assign n5556 = n5555 ^ x32 ;
  assign n5490 = x78 & n2879 ;
  assign n5557 = n5556 ^ n5490 ;
  assign n5489 = x80 & n2882 ;
  assign n5558 = n5557 ^ n5489 ;
  assign n5488 = n1206 & n2883 ;
  assign n5559 = n5558 ^ n5488 ;
  assign n5561 = n5560 ^ n5559 ;
  assign n5565 = n5564 ^ n5561 ;
  assign n5566 = n5565 ^ x29 ;
  assign n5487 = x81 & n2581 ;
  assign n5567 = n5566 ^ n5487 ;
  assign n5486 = x83 & n2422 ;
  assign n5568 = n5567 ^ n5486 ;
  assign n5485 = n1512 & n2423 ;
  assign n5569 = n5568 ^ n5485 ;
  assign n5571 = n5570 ^ n5569 ;
  assign n5482 = n5354 ^ n5345 ;
  assign n5483 = ~n5351 & n5482 ;
  assign n5484 = n5483 ^ n5354 ;
  assign n5572 = n5571 ^ n5484 ;
  assign n5573 = n5572 ^ x26 ;
  assign n5481 = x84 & n2018 ;
  assign n5574 = n5573 ^ n5481 ;
  assign n5480 = x86 & n2021 ;
  assign n5575 = n5574 ^ n5480 ;
  assign n5479 = n1857 & n2022 ;
  assign n5576 = n5575 ^ n5479 ;
  assign n5578 = n5577 ^ n5576 ;
  assign n5476 = n5364 ^ n5355 ;
  assign n5477 = ~n5361 & n5476 ;
  assign n5478 = n5477 ^ n5364 ;
  assign n5579 = n5578 ^ n5478 ;
  assign n5580 = n5579 ^ x23 ;
  assign n5475 = x87 & n1658 ;
  assign n5581 = n5580 ^ n5475 ;
  assign n5474 = x89 & n1661 ;
  assign n5582 = n5581 ^ n5474 ;
  assign n5473 = n1662 & n2249 ;
  assign n5583 = n5582 ^ n5473 ;
  assign n5585 = n5584 ^ n5583 ;
  assign n5470 = n5374 ^ n5365 ;
  assign n5471 = ~n5371 & n5470 ;
  assign n5472 = n5471 ^ n5374 ;
  assign n5586 = n5585 ^ n5472 ;
  assign n5587 = n5586 ^ x20 ;
  assign n5469 = x90 & n1327 ;
  assign n5588 = n5587 ^ n5469 ;
  assign n5468 = x92 & n1330 ;
  assign n5589 = n5588 ^ n5468 ;
  assign n5467 = n1331 & n2684 ;
  assign n5590 = n5589 ^ n5467 ;
  assign n5592 = n5591 ^ n5590 ;
  assign n5596 = n5595 ^ n5592 ;
  assign n5597 = n5596 ^ x17 ;
  assign n5466 = x93 & n1050 ;
  assign n5598 = n5597 ^ n5466 ;
  assign n5465 = x95 & n1053 ;
  assign n5599 = n5598 ^ n5465 ;
  assign n5464 = n1054 & n3159 ;
  assign n5600 = n5599 ^ n5464 ;
  assign n5602 = n5601 ^ n5600 ;
  assign n5461 = n5391 ^ n5382 ;
  assign n5462 = ~n5388 & n5461 ;
  assign n5463 = n5462 ^ n5391 ;
  assign n5603 = n5602 ^ n5463 ;
  assign n5604 = n5603 ^ x14 ;
  assign n5460 = x96 & n877 ;
  assign n5605 = n5604 ^ n5460 ;
  assign n5459 = x98 & n782 ;
  assign n5606 = n5605 ^ n5459 ;
  assign n5458 = n783 & n3660 ;
  assign n5607 = n5606 ^ n5458 ;
  assign n5609 = n5608 ^ n5607 ;
  assign n5613 = n5612 ^ n5609 ;
  assign n5614 = n5613 ^ x11 ;
  assign n5457 = x99 & n647 ;
  assign n5615 = n5614 ^ n5457 ;
  assign n5456 = x101 & ~n572 ;
  assign n5616 = n5615 ^ n5456 ;
  assign n5455 = ~n573 & n4215 ;
  assign n5617 = n5616 ^ n5455 ;
  assign n5619 = n5618 ^ n5617 ;
  assign n5623 = n5622 ^ n5619 ;
  assign n5624 = n5623 ^ x8 ;
  assign n5454 = x102 & n446 ;
  assign n5625 = n5624 ^ n5454 ;
  assign n5453 = x104 & n383 ;
  assign n5626 = n5625 ^ n5453 ;
  assign n5452 = n384 & ~n4814 ;
  assign n5627 = n5626 ^ n5452 ;
  assign n5629 = n5628 ^ n5627 ;
  assign n5633 = n5632 ^ n5629 ;
  assign n5634 = n5633 ^ x5 ;
  assign n5451 = x105 & n234 ;
  assign n5635 = n5634 ^ n5451 ;
  assign n5450 = x107 & n230 ;
  assign n5636 = n5635 ^ n5450 ;
  assign n5448 = n4800 ^ x107 ;
  assign n5449 = n231 & ~n5448 ;
  assign n5637 = n5636 ^ n5449 ;
  assign n5639 = n5638 ^ n5637 ;
  assign n5445 = n5422 ^ n5413 ;
  assign n5446 = ~n5419 & n5445 ;
  assign n5447 = n5446 ^ n5422 ;
  assign n5640 = n5639 ^ n5447 ;
  assign n5427 = x109 ^ x108 ;
  assign n5429 = n5226 & n5427 ;
  assign n5430 = n5429 ^ x108 ;
  assign n5431 = n5430 ^ x109 ;
  assign n5433 = x110 ^ x1 ;
  assign n5432 = x110 ^ x2 ;
  assign n5434 = n5433 ^ n5432 ;
  assign n5435 = ~n5431 & n5434 ;
  assign n5436 = n5435 ^ n5433 ;
  assign n5641 = n5640 ^ n5436 ;
  assign n5440 = x2 & x108 ;
  assign n5441 = n5440 ^ x109 ;
  assign n5442 = ~n255 & n5441 ;
  assign n5437 = n5436 ^ n5227 ;
  assign n5443 = n5442 ^ n5437 ;
  assign n5444 = ~x0 & n5443 ;
  assign n5642 = n5641 ^ n5444 ;
  assign n5646 = n5645 ^ n5642 ;
  assign n5874 = n5633 ^ n5447 ;
  assign n5875 = n5639 & n5874 ;
  assign n5876 = n5875 ^ n5633 ;
  assign n5872 = x107 & n227 ;
  assign n5865 = x104 & n390 ;
  assign n5858 = x101 & n578 ;
  assign n5851 = x98 & n788 ;
  assign n5843 = n5596 ^ n5463 ;
  assign n5844 = n5602 & n5843 ;
  assign n5845 = n5844 ^ n5596 ;
  assign n5841 = x95 & n1058 ;
  assign n5834 = x92 & n1335 ;
  assign n5826 = n5579 ^ n5472 ;
  assign n5827 = n5585 & n5826 ;
  assign n5828 = n5827 ^ n5579 ;
  assign n5824 = x89 & n1666 ;
  assign n5816 = n5572 ^ n5478 ;
  assign n5817 = n5578 & n5816 ;
  assign n5818 = n5817 ^ n5572 ;
  assign n5814 = x86 & n2014 ;
  assign n5806 = n5565 ^ n5484 ;
  assign n5807 = n5571 & n5806 ;
  assign n5808 = n5807 ^ n5565 ;
  assign n5804 = x83 & n2429 ;
  assign n5797 = x80 & n2887 ;
  assign n5790 = x77 & n3383 ;
  assign n5780 = x73 & n3916 ;
  assign n5779 = x75 & n3919 ;
  assign n5781 = n5780 ^ n5779 ;
  assign n5782 = n5781 ^ x38 ;
  assign n5778 = ~n774 & n3920 ;
  assign n5783 = n5782 ^ n5778 ;
  assign n5777 = x74 & n3924 ;
  assign n5784 = n5783 ^ n5777 ;
  assign n5770 = x70 & n4474 ;
  assign n5769 = x72 & n4471 ;
  assign n5771 = n5770 ^ n5769 ;
  assign n5772 = n5771 ^ x41 ;
  assign n5768 = n556 & n4472 ;
  assign n5773 = n5772 ^ n5768 ;
  assign n5767 = x71 & n4467 ;
  assign n5774 = n5773 ^ n5767 ;
  assign n5756 = x67 & n5094 ;
  assign n5755 = x69 & n5097 ;
  assign n5757 = n5756 ^ n5755 ;
  assign n5758 = n5757 ^ x44 ;
  assign n5754 = ~n375 & n5098 ;
  assign n5759 = n5758 ^ n5754 ;
  assign n5753 = x68 & n5102 ;
  assign n5760 = n5759 ^ n5753 ;
  assign n5739 = ~x46 & x47 ;
  assign n5740 = x64 & n5529 ;
  assign n5741 = n5739 & n5740 ;
  assign n5735 = x46 ^ x45 ;
  assign n5736 = ~n5309 & n5735 ;
  assign n5737 = x65 & n5736 ;
  assign n5728 = x47 ^ x46 ;
  assign n5729 = n5309 & ~n5728 ;
  assign n5730 = n5729 ^ n5309 ;
  assign n5733 = ~n150 & n5730 ;
  assign n5732 = x66 & n5309 ;
  assign n5734 = n5733 ^ n5732 ;
  assign n5738 = n5737 ^ n5734 ;
  assign n5742 = n5741 ^ n5738 ;
  assign n5727 = ~n5310 & ~n5533 ;
  assign n5743 = n5742 ^ n5727 ;
  assign n5744 = n5743 ^ n5738 ;
  assign n5725 = x46 & x64 ;
  assign n5726 = ~n5530 & n5725 ;
  assign n5745 = n5744 ^ n5726 ;
  assign n5746 = ~x47 & ~n5745 ;
  assign n5747 = n5746 ^ n5743 ;
  assign n5748 = n5747 ^ n5545 ;
  assign n5749 = n5748 ^ n5533 ;
  assign n5750 = n5749 ^ n5747 ;
  assign n5751 = ~n5542 & n5750 ;
  assign n5752 = n5751 ^ n5748 ;
  assign n5761 = n5760 ^ n5752 ;
  assign n5763 = n5761 ^ n5517 ;
  assign n5762 = n5761 ^ n5546 ;
  assign n5764 = n5763 ^ n5762 ;
  assign n5765 = n5522 & n5764 ;
  assign n5766 = n5765 ^ n5763 ;
  assign n5775 = n5774 ^ n5766 ;
  assign n5722 = n5547 ^ n5506 ;
  assign n5723 = n5553 & n5722 ;
  assign n5724 = n5723 ^ n5547 ;
  assign n5776 = n5775 ^ n5724 ;
  assign n5785 = n5784 ^ n5776 ;
  assign n5786 = n5785 ^ x35 ;
  assign n5721 = x76 & n3375 ;
  assign n5787 = n5786 ^ n5721 ;
  assign n5720 = x78 & n3378 ;
  assign n5788 = n5787 ^ n5720 ;
  assign n5719 = ~n1025 & n3379 ;
  assign n5789 = n5788 ^ n5719 ;
  assign n5791 = n5790 ^ n5789 ;
  assign n5716 = n5554 ^ n5498 ;
  assign n5717 = n5503 & n5716 ;
  assign n5718 = n5717 ^ n5498 ;
  assign n5792 = n5791 ^ n5718 ;
  assign n5793 = n5792 ^ x32 ;
  assign n5715 = x79 & n2879 ;
  assign n5794 = n5793 ^ n5715 ;
  assign n5714 = x81 & n2882 ;
  assign n5795 = n5794 ^ n5714 ;
  assign n5713 = n1305 & n2883 ;
  assign n5796 = n5795 ^ n5713 ;
  assign n5798 = n5797 ^ n5796 ;
  assign n5710 = n5564 ^ n5555 ;
  assign n5711 = ~n5561 & n5710 ;
  assign n5712 = n5711 ^ n5564 ;
  assign n5799 = n5798 ^ n5712 ;
  assign n5800 = n5799 ^ x29 ;
  assign n5709 = x82 & n2581 ;
  assign n5801 = n5800 ^ n5709 ;
  assign n5708 = x84 & n2422 ;
  assign n5802 = n5801 ^ n5708 ;
  assign n5707 = n1624 & n2423 ;
  assign n5803 = n5802 ^ n5707 ;
  assign n5805 = n5804 ^ n5803 ;
  assign n5809 = n5808 ^ n5805 ;
  assign n5810 = n5809 ^ x26 ;
  assign n5706 = x85 & n2018 ;
  assign n5811 = n5810 ^ n5706 ;
  assign n5705 = x87 & n2021 ;
  assign n5812 = n5811 ^ n5705 ;
  assign n5704 = n1982 & n2022 ;
  assign n5813 = n5812 ^ n5704 ;
  assign n5815 = n5814 ^ n5813 ;
  assign n5819 = n5818 ^ n5815 ;
  assign n5820 = n5819 ^ x23 ;
  assign n5703 = x88 & n1658 ;
  assign n5821 = n5820 ^ n5703 ;
  assign n5702 = x90 & n1661 ;
  assign n5822 = n5821 ^ n5702 ;
  assign n5701 = n1662 & n2386 ;
  assign n5823 = n5822 ^ n5701 ;
  assign n5825 = n5824 ^ n5823 ;
  assign n5829 = n5828 ^ n5825 ;
  assign n5830 = n5829 ^ x20 ;
  assign n5700 = x91 & n1327 ;
  assign n5831 = n5830 ^ n5700 ;
  assign n5699 = x93 & n1330 ;
  assign n5832 = n5831 ^ n5699 ;
  assign n5698 = n1331 & n2836 ;
  assign n5833 = n5832 ^ n5698 ;
  assign n5835 = n5834 ^ n5833 ;
  assign n5695 = n5595 ^ n5586 ;
  assign n5696 = ~n5592 & n5695 ;
  assign n5697 = n5696 ^ n5595 ;
  assign n5836 = n5835 ^ n5697 ;
  assign n5837 = n5836 ^ x17 ;
  assign n5694 = x94 & n1050 ;
  assign n5838 = n5837 ^ n5694 ;
  assign n5693 = x96 & n1053 ;
  assign n5839 = n5838 ^ n5693 ;
  assign n5692 = n1054 & n3323 ;
  assign n5840 = n5839 ^ n5692 ;
  assign n5842 = n5841 ^ n5840 ;
  assign n5846 = n5845 ^ n5842 ;
  assign n5847 = n5846 ^ x14 ;
  assign n5691 = x97 & n877 ;
  assign n5848 = n5847 ^ n5691 ;
  assign n5690 = x99 & n782 ;
  assign n5849 = n5848 ^ n5690 ;
  assign n5689 = n783 & n3843 ;
  assign n5850 = n5849 ^ n5689 ;
  assign n5852 = n5851 ^ n5850 ;
  assign n5686 = n5612 ^ n5603 ;
  assign n5687 = ~n5609 & n5686 ;
  assign n5688 = n5687 ^ n5612 ;
  assign n5853 = n5852 ^ n5688 ;
  assign n5854 = n5853 ^ x11 ;
  assign n5685 = x100 & n647 ;
  assign n5855 = n5854 ^ n5685 ;
  assign n5684 = x102 & ~n572 ;
  assign n5856 = n5855 ^ n5684 ;
  assign n5683 = ~n573 & n4410 ;
  assign n5857 = n5856 ^ n5683 ;
  assign n5859 = n5858 ^ n5857 ;
  assign n5680 = n5622 ^ n5613 ;
  assign n5681 = ~n5619 & n5680 ;
  assign n5682 = n5681 ^ n5622 ;
  assign n5860 = n5859 ^ n5682 ;
  assign n5861 = n5860 ^ x8 ;
  assign n5679 = x103 & n446 ;
  assign n5862 = n5861 ^ n5679 ;
  assign n5678 = x105 & n383 ;
  assign n5863 = n5862 ^ n5678 ;
  assign n5677 = n384 & ~n5023 ;
  assign n5864 = n5863 ^ n5677 ;
  assign n5866 = n5865 ^ n5864 ;
  assign n5674 = n5632 ^ n5623 ;
  assign n5675 = ~n5629 & n5674 ;
  assign n5676 = n5675 ^ n5632 ;
  assign n5867 = n5866 ^ n5676 ;
  assign n5868 = n5867 ^ x5 ;
  assign n5673 = x106 & n234 ;
  assign n5869 = n5868 ^ n5673 ;
  assign n5672 = x108 & n230 ;
  assign n5870 = n5869 ^ n5672 ;
  assign n5670 = n5006 ^ x108 ;
  assign n5671 = n231 & n5670 ;
  assign n5871 = n5870 ^ n5671 ;
  assign n5873 = n5872 ^ n5871 ;
  assign n5877 = n5876 ^ n5873 ;
  assign n5652 = x109 & n5430 ;
  assign n5654 = n5652 ^ n5431 ;
  assign n5655 = x110 & n5654 ;
  assign n5653 = ~x110 & ~n5652 ;
  assign n5656 = n5655 ^ n5653 ;
  assign n5658 = x111 ^ x1 ;
  assign n5657 = x111 ^ x2 ;
  assign n5659 = n5658 ^ n5657 ;
  assign n5660 = n5656 & n5659 ;
  assign n5661 = n5660 ^ n5658 ;
  assign n5878 = n5877 ^ n5661 ;
  assign n5665 = x2 & x109 ;
  assign n5666 = n5665 ^ x110 ;
  assign n5667 = ~x1 & n5666 ;
  assign n5662 = n5661 ^ n5432 ;
  assign n5668 = n5667 ^ n5662 ;
  assign n5669 = ~x0 & n5668 ;
  assign n5879 = n5878 ^ n5669 ;
  assign n5647 = n5645 ^ n5640 ;
  assign n5648 = ~n5642 & n5647 ;
  assign n5649 = n5648 ^ n5645 ;
  assign n5880 = n5879 ^ n5649 ;
  assign n6104 = n5877 ^ n5649 ;
  assign n6105 = ~n5879 & ~n6104 ;
  assign n6106 = n6105 ^ n5877 ;
  assign n6099 = x108 & n227 ;
  assign n6091 = n5860 ^ n5676 ;
  assign n6092 = ~n5866 & ~n6091 ;
  assign n6093 = n6092 ^ n5860 ;
  assign n6089 = x105 & n390 ;
  assign n6081 = n5853 ^ n5682 ;
  assign n6082 = ~n5859 & ~n6081 ;
  assign n6083 = n6082 ^ n5853 ;
  assign n6079 = x102 & n578 ;
  assign n6071 = n5846 ^ n5688 ;
  assign n6072 = ~n5852 & ~n6071 ;
  assign n6073 = n6072 ^ n5846 ;
  assign n6069 = x99 & n788 ;
  assign n6062 = x96 & n1058 ;
  assign n6054 = n5829 ^ n5697 ;
  assign n6055 = ~n5835 & ~n6054 ;
  assign n6056 = n6055 ^ n5829 ;
  assign n6052 = x93 & n1335 ;
  assign n6045 = x90 & n1666 ;
  assign n6038 = x87 & n2014 ;
  assign n6031 = x84 & n2429 ;
  assign n6023 = n5792 ^ n5712 ;
  assign n6024 = ~n5798 & ~n6023 ;
  assign n6025 = n6024 ^ n5792 ;
  assign n6021 = x81 & n2887 ;
  assign n6011 = x77 & n3375 ;
  assign n6010 = x79 & n3378 ;
  assign n6012 = n6011 ^ n6010 ;
  assign n6013 = n6012 ^ x35 ;
  assign n6009 = n1118 & n3379 ;
  assign n6014 = n6013 ^ n6009 ;
  assign n6008 = x78 & n3383 ;
  assign n6015 = n6014 ^ n6008 ;
  assign n6004 = x75 & n3924 ;
  assign n5994 = x71 & n4474 ;
  assign n5993 = x73 & n4471 ;
  assign n5995 = n5994 ^ n5993 ;
  assign n5996 = n5995 ^ x41 ;
  assign n5992 = n633 & n4472 ;
  assign n5997 = n5996 ^ n5992 ;
  assign n5991 = x72 & n4467 ;
  assign n5998 = n5997 ^ n5991 ;
  assign n5982 = n5760 ^ n5747 ;
  assign n5983 = ~n5752 & ~n5982 ;
  assign n5984 = n5983 ^ n5747 ;
  assign n5980 = x69 & n5102 ;
  assign n5972 = x48 ^ x47 ;
  assign n5973 = x64 & n5972 ;
  assign n5970 = x47 & ~n5742 ;
  assign n5971 = n5727 & n5970 ;
  assign n5974 = n5973 ^ n5971 ;
  assign n5963 = x47 ^ x45 ;
  assign n5964 = ~n5309 & n5963 ;
  assign n5965 = n5728 & n5964 ;
  assign n5966 = x65 & n5965 ;
  assign n5962 = x66 & n5736 ;
  assign n5967 = n5966 ^ n5962 ;
  assign n5968 = n5967 ^ x47 ;
  assign n5959 = ~n153 & ~n5728 ;
  assign n5960 = n5959 ^ n291 ;
  assign n5961 = n5309 & ~n5960 ;
  assign n5969 = n5968 ^ n5961 ;
  assign n5975 = n5974 ^ n5969 ;
  assign n5976 = n5975 ^ x44 ;
  assign n5956 = x68 & n5094 ;
  assign n5977 = n5976 ^ n5956 ;
  assign n5955 = x70 & n5097 ;
  assign n5978 = n5977 ^ n5955 ;
  assign n5954 = ~n436 & n5098 ;
  assign n5979 = n5978 ^ n5954 ;
  assign n5981 = n5980 ^ n5979 ;
  assign n5985 = n5984 ^ n5981 ;
  assign n5987 = n5985 ^ n5761 ;
  assign n5986 = n5985 ^ n5774 ;
  assign n5988 = n5987 ^ n5986 ;
  assign n5989 = ~n5766 & ~n5988 ;
  assign n5990 = n5989 ^ n5987 ;
  assign n5999 = n5998 ^ n5990 ;
  assign n6000 = n5999 ^ x38 ;
  assign n5953 = x74 & n3916 ;
  assign n6001 = n6000 ^ n5953 ;
  assign n5952 = x76 & n3919 ;
  assign n6002 = n6001 ^ n5952 ;
  assign n5951 = ~n853 & n3920 ;
  assign n6003 = n6002 ^ n5951 ;
  assign n6005 = n6004 ^ n6003 ;
  assign n5948 = n5784 ^ n5724 ;
  assign n5949 = n5776 & n5948 ;
  assign n5950 = n5949 ^ n5784 ;
  assign n6006 = n6005 ^ n5950 ;
  assign n5945 = n5785 ^ n5718 ;
  assign n5946 = ~n5791 & ~n5945 ;
  assign n5947 = n5946 ^ n5785 ;
  assign n6007 = n6006 ^ n5947 ;
  assign n6016 = n6015 ^ n6007 ;
  assign n6017 = n6016 ^ x32 ;
  assign n5944 = x80 & n2879 ;
  assign n6018 = n6017 ^ n5944 ;
  assign n5943 = x82 & n2882 ;
  assign n6019 = n6018 ^ n5943 ;
  assign n5942 = n1411 & n2883 ;
  assign n6020 = n6019 ^ n5942 ;
  assign n6022 = n6021 ^ n6020 ;
  assign n6026 = n6025 ^ n6022 ;
  assign n6027 = n6026 ^ x29 ;
  assign n5941 = x83 & n2581 ;
  assign n6028 = n6027 ^ n5941 ;
  assign n5940 = x85 & n2422 ;
  assign n6029 = n6028 ^ n5940 ;
  assign n5939 = n1743 & n2423 ;
  assign n6030 = n6029 ^ n5939 ;
  assign n6032 = n6031 ^ n6030 ;
  assign n5936 = n5808 ^ n5799 ;
  assign n5937 = n5805 & ~n5936 ;
  assign n5938 = n5937 ^ n5808 ;
  assign n6033 = n6032 ^ n5938 ;
  assign n6034 = n6033 ^ x26 ;
  assign n5935 = x86 & n2018 ;
  assign n6035 = n6034 ^ n5935 ;
  assign n5934 = x88 & n2021 ;
  assign n6036 = n6035 ^ n5934 ;
  assign n5933 = n2022 & n2119 ;
  assign n6037 = n6036 ^ n5933 ;
  assign n6039 = n6038 ^ n6037 ;
  assign n5930 = n5818 ^ n5809 ;
  assign n5931 = n5815 & ~n5930 ;
  assign n5932 = n5931 ^ n5818 ;
  assign n6040 = n6039 ^ n5932 ;
  assign n6041 = n6040 ^ x23 ;
  assign n5929 = x89 & n1658 ;
  assign n6042 = n6041 ^ n5929 ;
  assign n5928 = x91 & n1661 ;
  assign n6043 = n6042 ^ n5928 ;
  assign n5927 = n1662 & n2542 ;
  assign n6044 = n6043 ^ n5927 ;
  assign n6046 = n6045 ^ n6044 ;
  assign n5924 = n5828 ^ n5819 ;
  assign n5925 = n5825 & ~n5924 ;
  assign n5926 = n5925 ^ n5828 ;
  assign n6047 = n6046 ^ n5926 ;
  assign n6048 = n6047 ^ x20 ;
  assign n5923 = x92 & n1327 ;
  assign n6049 = n6048 ^ n5923 ;
  assign n5922 = x94 & n1330 ;
  assign n6050 = n6049 ^ n5922 ;
  assign n5921 = n1331 & n2997 ;
  assign n6051 = n6050 ^ n5921 ;
  assign n6053 = n6052 ^ n6051 ;
  assign n6057 = n6056 ^ n6053 ;
  assign n6058 = n6057 ^ x17 ;
  assign n5920 = x95 & n1050 ;
  assign n6059 = n6058 ^ n5920 ;
  assign n5919 = x97 & n1053 ;
  assign n6060 = n6059 ^ n5919 ;
  assign n5918 = n1054 & n3494 ;
  assign n6061 = n6060 ^ n5918 ;
  assign n6063 = n6062 ^ n6061 ;
  assign n5915 = n5845 ^ n5836 ;
  assign n5916 = n5842 & ~n5915 ;
  assign n5917 = n5916 ^ n5845 ;
  assign n6064 = n6063 ^ n5917 ;
  assign n6065 = n6064 ^ x14 ;
  assign n5914 = x98 & n877 ;
  assign n6066 = n6065 ^ n5914 ;
  assign n5913 = x100 & n782 ;
  assign n6067 = n6066 ^ n5913 ;
  assign n5912 = n783 & n4034 ;
  assign n6068 = n6067 ^ n5912 ;
  assign n6070 = n6069 ^ n6068 ;
  assign n6074 = n6073 ^ n6070 ;
  assign n6075 = n6074 ^ x11 ;
  assign n5911 = x101 & n647 ;
  assign n6076 = n6075 ^ n5911 ;
  assign n5910 = x103 & ~n572 ;
  assign n6077 = n6076 ^ n5910 ;
  assign n5909 = ~n573 & ~n4615 ;
  assign n6078 = n6077 ^ n5909 ;
  assign n6080 = n6079 ^ n6078 ;
  assign n6084 = n6083 ^ n6080 ;
  assign n6085 = n6084 ^ x8 ;
  assign n5908 = x104 & n446 ;
  assign n6086 = n6085 ^ n5908 ;
  assign n5907 = x106 & n383 ;
  assign n6087 = n6086 ^ n5907 ;
  assign n5906 = n384 & ~n5240 ;
  assign n6088 = n6087 ^ n5906 ;
  assign n6090 = n6089 ^ n6088 ;
  assign n6094 = n6093 ^ n6090 ;
  assign n6095 = n6094 ^ x5 ;
  assign n5905 = x107 & n234 ;
  assign n6096 = n6095 ^ n5905 ;
  assign n5904 = x109 & n230 ;
  assign n6097 = n6096 ^ n5904 ;
  assign n5902 = n5226 ^ x109 ;
  assign n5903 = n231 & n5902 ;
  assign n6098 = n6097 ^ n5903 ;
  assign n6100 = n6099 ^ n6098 ;
  assign n5899 = n5876 ^ n5867 ;
  assign n5900 = n5873 & ~n5899 ;
  assign n5901 = n5900 ^ n5876 ;
  assign n6101 = n6100 ^ n5901 ;
  assign n5884 = ~x111 & ~n5655 ;
  assign n5883 = x111 & ~n5653 ;
  assign n5885 = n5884 ^ n5883 ;
  assign n5887 = x112 ^ x1 ;
  assign n5886 = x112 ^ x2 ;
  assign n5888 = n5887 ^ n5886 ;
  assign n5889 = n5885 & n5888 ;
  assign n5890 = n5889 ^ n5887 ;
  assign n6102 = n6101 ^ n5890 ;
  assign n5894 = x2 & x110 ;
  assign n5895 = n5894 ^ x111 ;
  assign n5896 = ~x1 & n5895 ;
  assign n5891 = n5890 ^ n5657 ;
  assign n5897 = n5896 ^ n5891 ;
  assign n5898 = ~x0 & n5897 ;
  assign n6103 = n6102 ^ n5898 ;
  assign n6107 = n6106 ^ n6103 ;
  assign n6332 = n6094 ^ n5901 ;
  assign n6333 = n6100 & n6332 ;
  assign n6334 = n6333 ^ n6094 ;
  assign n6330 = x109 & n227 ;
  assign n6323 = x106 & n390 ;
  assign n6316 = x103 & n578 ;
  assign n6309 = x100 & n788 ;
  assign n6301 = n6057 ^ n5917 ;
  assign n6302 = ~n6063 & ~n6301 ;
  assign n6303 = n6302 ^ n6057 ;
  assign n6299 = x97 & n1058 ;
  assign n6292 = x94 & n1335 ;
  assign n6284 = n6040 ^ n5926 ;
  assign n6285 = n6046 & n6284 ;
  assign n6286 = n6285 ^ n6040 ;
  assign n6282 = x91 & n1666 ;
  assign n6274 = n6033 ^ n5932 ;
  assign n6275 = n6039 & n6274 ;
  assign n6276 = n6275 ^ n6033 ;
  assign n6272 = x88 & n2014 ;
  assign n6264 = n6026 ^ n5938 ;
  assign n6265 = n6032 & n6264 ;
  assign n6266 = n6265 ^ n6026 ;
  assign n6262 = x85 & n2429 ;
  assign n6255 = x82 & n2887 ;
  assign n6248 = x79 & n3383 ;
  assign n6241 = x76 & n3924 ;
  assign n6233 = n5998 ^ n5985 ;
  assign n6234 = n5990 & ~n6233 ;
  assign n6235 = n6234 ^ n5985 ;
  assign n6231 = x73 & n4467 ;
  assign n6224 = x70 & n5102 ;
  assign n6214 = x66 & n5965 ;
  assign n6213 = x68 & n5729 ;
  assign n6215 = n6214 ^ n6213 ;
  assign n6216 = n6215 ^ x47 ;
  assign n6212 = ~n340 & n5730 ;
  assign n6217 = n6216 ^ n6212 ;
  assign n6211 = x67 & n5736 ;
  assign n6218 = n6217 ^ n6211 ;
  assign n6207 = n5969 & ~n5973 ;
  assign n6208 = ~n5971 & n6207 ;
  assign n6209 = n6208 ^ n5969 ;
  assign n6204 = x65 ^ x48 ;
  assign n6205 = n5972 & ~n6204 ;
  assign n6200 = x47 & x48 ;
  assign n6201 = n6200 ^ x49 ;
  assign n6202 = ~x64 & n6201 ;
  assign n6196 = x49 ^ x47 ;
  assign n6203 = n6202 ^ n6196 ;
  assign n6206 = n6205 ^ n6203 ;
  assign n6210 = n6209 ^ n6206 ;
  assign n6219 = n6218 ^ n6210 ;
  assign n6220 = n6219 ^ x44 ;
  assign n6195 = x69 & n5094 ;
  assign n6221 = n6220 ^ n6195 ;
  assign n6194 = x71 & n5097 ;
  assign n6222 = n6221 ^ n6194 ;
  assign n6193 = ~n493 & n5098 ;
  assign n6223 = n6222 ^ n6193 ;
  assign n6225 = n6224 ^ n6223 ;
  assign n6190 = n5984 ^ n5975 ;
  assign n6191 = ~n5981 & ~n6190 ;
  assign n6192 = n6191 ^ n5984 ;
  assign n6226 = n6225 ^ n6192 ;
  assign n6227 = n6226 ^ x41 ;
  assign n6189 = x72 & n4474 ;
  assign n6228 = n6227 ^ n6189 ;
  assign n6188 = x74 & n4471 ;
  assign n6229 = n6228 ^ n6188 ;
  assign n6187 = n699 & n4472 ;
  assign n6230 = n6229 ^ n6187 ;
  assign n6232 = n6231 ^ n6230 ;
  assign n6236 = n6235 ^ n6232 ;
  assign n6237 = n6236 ^ x38 ;
  assign n6186 = x75 & n3916 ;
  assign n6238 = n6237 ^ n6186 ;
  assign n6185 = x77 & n3919 ;
  assign n6239 = n6238 ^ n6185 ;
  assign n6184 = ~n939 & n3920 ;
  assign n6240 = n6239 ^ n6184 ;
  assign n6242 = n6241 ^ n6240 ;
  assign n6181 = n5999 ^ n5950 ;
  assign n6182 = n6005 & n6181 ;
  assign n6183 = n6182 ^ n5999 ;
  assign n6243 = n6242 ^ n6183 ;
  assign n6244 = n6243 ^ x35 ;
  assign n6180 = x78 & n3375 ;
  assign n6245 = n6244 ^ n6180 ;
  assign n6179 = x80 & n3378 ;
  assign n6246 = n6245 ^ n6179 ;
  assign n6178 = n1206 & n3379 ;
  assign n6247 = n6246 ^ n6178 ;
  assign n6249 = n6248 ^ n6247 ;
  assign n6175 = n6015 ^ n5947 ;
  assign n6176 = n6007 & ~n6175 ;
  assign n6177 = n6176 ^ n6015 ;
  assign n6250 = n6249 ^ n6177 ;
  assign n6251 = n6250 ^ x32 ;
  assign n6174 = x81 & n2879 ;
  assign n6252 = n6251 ^ n6174 ;
  assign n6173 = x83 & n2882 ;
  assign n6253 = n6252 ^ n6173 ;
  assign n6172 = n1512 & n2883 ;
  assign n6254 = n6253 ^ n6172 ;
  assign n6256 = n6255 ^ n6254 ;
  assign n6169 = n6025 ^ n6016 ;
  assign n6170 = n6022 & n6169 ;
  assign n6171 = n6170 ^ n6025 ;
  assign n6257 = n6256 ^ n6171 ;
  assign n6258 = n6257 ^ x29 ;
  assign n6168 = x84 & n2581 ;
  assign n6259 = n6258 ^ n6168 ;
  assign n6167 = x86 & n2422 ;
  assign n6260 = n6259 ^ n6167 ;
  assign n6166 = n1857 & n2423 ;
  assign n6261 = n6260 ^ n6166 ;
  assign n6263 = n6262 ^ n6261 ;
  assign n6267 = n6266 ^ n6263 ;
  assign n6268 = n6267 ^ x26 ;
  assign n6165 = x87 & n2018 ;
  assign n6269 = n6268 ^ n6165 ;
  assign n6164 = x89 & n2021 ;
  assign n6270 = n6269 ^ n6164 ;
  assign n6163 = n2022 & n2249 ;
  assign n6271 = n6270 ^ n6163 ;
  assign n6273 = n6272 ^ n6271 ;
  assign n6277 = n6276 ^ n6273 ;
  assign n6278 = n6277 ^ x23 ;
  assign n6162 = x90 & n1658 ;
  assign n6279 = n6278 ^ n6162 ;
  assign n6161 = x92 & n1661 ;
  assign n6280 = n6279 ^ n6161 ;
  assign n6160 = n1662 & n2684 ;
  assign n6281 = n6280 ^ n6160 ;
  assign n6283 = n6282 ^ n6281 ;
  assign n6287 = n6286 ^ n6283 ;
  assign n6288 = n6287 ^ x20 ;
  assign n6159 = x93 & n1327 ;
  assign n6289 = n6288 ^ n6159 ;
  assign n6158 = x95 & n1330 ;
  assign n6290 = n6289 ^ n6158 ;
  assign n6157 = n1331 & n3159 ;
  assign n6291 = n6290 ^ n6157 ;
  assign n6293 = n6292 ^ n6291 ;
  assign n6154 = n6056 ^ n6047 ;
  assign n6155 = ~n6053 & ~n6154 ;
  assign n6156 = n6155 ^ n6056 ;
  assign n6294 = n6293 ^ n6156 ;
  assign n6295 = n6294 ^ x17 ;
  assign n6153 = x96 & n1050 ;
  assign n6296 = n6295 ^ n6153 ;
  assign n6152 = x98 & n1053 ;
  assign n6297 = n6296 ^ n6152 ;
  assign n6151 = n1054 & n3660 ;
  assign n6298 = n6297 ^ n6151 ;
  assign n6300 = n6299 ^ n6298 ;
  assign n6304 = n6303 ^ n6300 ;
  assign n6305 = n6304 ^ x14 ;
  assign n6150 = x99 & n877 ;
  assign n6306 = n6305 ^ n6150 ;
  assign n6149 = x101 & n782 ;
  assign n6307 = n6306 ^ n6149 ;
  assign n6148 = n783 & n4215 ;
  assign n6308 = n6307 ^ n6148 ;
  assign n6310 = n6309 ^ n6308 ;
  assign n6145 = n6073 ^ n6064 ;
  assign n6146 = n6070 & n6145 ;
  assign n6147 = n6146 ^ n6073 ;
  assign n6311 = n6310 ^ n6147 ;
  assign n6312 = n6311 ^ x11 ;
  assign n6144 = x102 & n647 ;
  assign n6313 = n6312 ^ n6144 ;
  assign n6143 = x104 & ~n572 ;
  assign n6314 = n6313 ^ n6143 ;
  assign n6142 = ~n573 & ~n4814 ;
  assign n6315 = n6314 ^ n6142 ;
  assign n6317 = n6316 ^ n6315 ;
  assign n6139 = n6083 ^ n6074 ;
  assign n6140 = ~n6080 & ~n6139 ;
  assign n6141 = n6140 ^ n6083 ;
  assign n6318 = n6317 ^ n6141 ;
  assign n6319 = n6318 ^ x8 ;
  assign n6138 = x105 & n446 ;
  assign n6320 = n6319 ^ n6138 ;
  assign n6137 = x107 & n383 ;
  assign n6321 = n6320 ^ n6137 ;
  assign n6136 = n384 & ~n5448 ;
  assign n6322 = n6321 ^ n6136 ;
  assign n6324 = n6323 ^ n6322 ;
  assign n6133 = n6093 ^ n6084 ;
  assign n6134 = n6090 & n6133 ;
  assign n6135 = n6134 ^ n6093 ;
  assign n6325 = n6324 ^ n6135 ;
  assign n6326 = n6325 ^ x5 ;
  assign n6132 = x108 & n234 ;
  assign n6327 = n6326 ^ n6132 ;
  assign n6131 = x110 & n230 ;
  assign n6328 = n6327 ^ n6131 ;
  assign n5650 = x110 ^ x109 ;
  assign n6129 = n5650 ^ n5430 ;
  assign n6130 = n231 & n6129 ;
  assign n6329 = n6328 ^ n6130 ;
  assign n6331 = n6330 ^ n6329 ;
  assign n6335 = n6334 ^ n6331 ;
  assign n6114 = x112 & ~n5884 ;
  assign n6113 = ~x112 & ~n5883 ;
  assign n6115 = n6114 ^ n6113 ;
  assign n6117 = x113 ^ x1 ;
  assign n6116 = x113 ^ x2 ;
  assign n6118 = n6117 ^ n6116 ;
  assign n6119 = n6115 & n6118 ;
  assign n6120 = n6119 ^ n6117 ;
  assign n6336 = n6335 ^ n6120 ;
  assign n6124 = x2 & x111 ;
  assign n6125 = n6124 ^ x112 ;
  assign n6126 = ~x1 & n6125 ;
  assign n6121 = n6120 ^ n5886 ;
  assign n6127 = n6126 ^ n6121 ;
  assign n6128 = ~x0 & n6127 ;
  assign n6337 = n6336 ^ n6128 ;
  assign n6108 = n6106 ^ n6101 ;
  assign n6109 = ~n6103 & ~n6108 ;
  assign n6110 = n6109 ^ n6106 ;
  assign n6338 = n6337 ^ n6110 ;
  assign n6575 = n6335 ^ n6110 ;
  assign n6576 = n6337 & ~n6575 ;
  assign n6577 = n6576 ^ n6335 ;
  assign n6570 = x110 & n227 ;
  assign n6562 = n6318 ^ n6135 ;
  assign n6563 = ~n6324 & n6562 ;
  assign n6564 = n6563 ^ n6318 ;
  assign n6560 = x107 & n390 ;
  assign n6552 = n6311 ^ n6141 ;
  assign n6553 = n6317 & ~n6552 ;
  assign n6554 = n6553 ^ n6311 ;
  assign n6550 = x104 & n578 ;
  assign n6542 = n6304 ^ n6147 ;
  assign n6543 = ~n6310 & n6542 ;
  assign n6544 = n6543 ^ n6304 ;
  assign n6540 = x101 & n788 ;
  assign n6533 = x98 & n1058 ;
  assign n6525 = n6287 ^ n6156 ;
  assign n6526 = ~n6293 & n6525 ;
  assign n6527 = n6526 ^ n6287 ;
  assign n6523 = x95 & n1335 ;
  assign n6516 = x92 & n1666 ;
  assign n6509 = x89 & n2014 ;
  assign n6502 = x86 & n2429 ;
  assign n6494 = n6250 ^ n6171 ;
  assign n6495 = n6256 & ~n6494 ;
  assign n6496 = n6495 ^ n6250 ;
  assign n6488 = x82 & n2879 ;
  assign n6487 = x84 & n2882 ;
  assign n6489 = n6488 ^ n6487 ;
  assign n6490 = n6489 ^ x32 ;
  assign n6486 = n1624 & n2883 ;
  assign n6491 = n6490 ^ n6486 ;
  assign n6485 = x83 & n2887 ;
  assign n6492 = n6491 ^ n6485 ;
  assign n6482 = x80 & n3383 ;
  assign n6474 = n6236 ^ n6183 ;
  assign n6475 = n6242 & n6474 ;
  assign n6476 = n6475 ^ n6236 ;
  assign n6472 = x77 & n3924 ;
  assign n6461 = x70 & n5094 ;
  assign n6460 = x72 & n5097 ;
  assign n6462 = n6461 ^ n6460 ;
  assign n6463 = n6462 ^ x44 ;
  assign n6459 = n556 & n5098 ;
  assign n6464 = n6463 ^ n6459 ;
  assign n6458 = x71 & n5102 ;
  assign n6465 = n6464 ^ n6458 ;
  assign n6455 = n6219 ^ n6192 ;
  assign n6456 = n6225 & ~n6455 ;
  assign n6445 = x67 & n5965 ;
  assign n6444 = x69 & n5729 ;
  assign n6446 = n6445 ^ n6444 ;
  assign n6447 = n6446 ^ x47 ;
  assign n6443 = ~n375 & n5730 ;
  assign n6448 = n6447 ^ n6443 ;
  assign n6442 = x68 & n5736 ;
  assign n6449 = n6448 ^ n6442 ;
  assign n6440 = x50 & ~n5973 ;
  assign n6441 = ~n6206 & n6440 ;
  assign n6450 = n6449 ^ n6441 ;
  assign n6425 = x64 & ~n6196 ;
  assign n6198 = x49 ^ x48 ;
  assign n6433 = ~n5972 & n6198 ;
  assign n6434 = x65 & n6433 ;
  assign n6427 = x50 ^ x49 ;
  assign n6428 = n5972 & ~n6427 ;
  assign n6429 = n6428 ^ n5972 ;
  assign n6430 = ~n150 & n6429 ;
  assign n6426 = x66 & n5972 ;
  assign n6431 = n6430 ^ n6426 ;
  assign n6432 = n6431 ^ x50 ;
  assign n6435 = n6434 ^ n6432 ;
  assign n6436 = n6435 ^ x47 ;
  assign n6437 = ~n6198 & n6436 ;
  assign n6438 = n6425 & n6437 ;
  assign n6439 = n6438 ^ n6435 ;
  assign n6451 = n6450 ^ n6439 ;
  assign n6422 = n6218 ^ n6209 ;
  assign n6423 = ~n6210 & n6422 ;
  assign n6424 = n6423 ^ n6218 ;
  assign n6452 = n6451 ^ n6424 ;
  assign n6453 = n6452 ^ n6219 ;
  assign n6457 = n6456 ^ n6453 ;
  assign n6466 = n6465 ^ n6457 ;
  assign n6412 = x73 & n4474 ;
  assign n6411 = x75 & n4471 ;
  assign n6413 = n6412 ^ n6411 ;
  assign n6414 = n6413 ^ x41 ;
  assign n6410 = ~n774 & n4472 ;
  assign n6415 = n6414 ^ n6410 ;
  assign n6409 = x74 & n4467 ;
  assign n6416 = n6415 ^ n6409 ;
  assign n6417 = n6416 ^ n6235 ;
  assign n6418 = n6417 ^ n6226 ;
  assign n6419 = n6418 ^ n6416 ;
  assign n6420 = n6232 & n6419 ;
  assign n6421 = n6420 ^ n6417 ;
  assign n6467 = n6466 ^ n6421 ;
  assign n6468 = n6467 ^ x38 ;
  assign n6408 = x76 & n3916 ;
  assign n6469 = n6468 ^ n6408 ;
  assign n6407 = x78 & n3919 ;
  assign n6470 = n6469 ^ n6407 ;
  assign n6406 = ~n1025 & n3920 ;
  assign n6471 = n6470 ^ n6406 ;
  assign n6473 = n6472 ^ n6471 ;
  assign n6477 = n6476 ^ n6473 ;
  assign n6478 = n6477 ^ x35 ;
  assign n6405 = x79 & n3375 ;
  assign n6479 = n6478 ^ n6405 ;
  assign n6404 = x81 & n3378 ;
  assign n6480 = n6479 ^ n6404 ;
  assign n6403 = n1305 & n3379 ;
  assign n6481 = n6480 ^ n6403 ;
  assign n6483 = n6482 ^ n6481 ;
  assign n6400 = n6243 ^ n6177 ;
  assign n6401 = n6249 & n6400 ;
  assign n6402 = n6401 ^ n6243 ;
  assign n6484 = n6483 ^ n6402 ;
  assign n6493 = n6492 ^ n6484 ;
  assign n6497 = n6496 ^ n6493 ;
  assign n6498 = n6497 ^ x29 ;
  assign n6399 = x85 & n2581 ;
  assign n6499 = n6498 ^ n6399 ;
  assign n6398 = x87 & n2422 ;
  assign n6500 = n6499 ^ n6398 ;
  assign n6397 = n1982 & n2423 ;
  assign n6501 = n6500 ^ n6397 ;
  assign n6503 = n6502 ^ n6501 ;
  assign n6394 = n6266 ^ n6257 ;
  assign n6395 = n6263 & ~n6394 ;
  assign n6396 = n6395 ^ n6266 ;
  assign n6504 = n6503 ^ n6396 ;
  assign n6505 = n6504 ^ x26 ;
  assign n6393 = x88 & n2018 ;
  assign n6506 = n6505 ^ n6393 ;
  assign n6392 = x90 & n2021 ;
  assign n6507 = n6506 ^ n6392 ;
  assign n6391 = n2022 & n2386 ;
  assign n6508 = n6507 ^ n6391 ;
  assign n6510 = n6509 ^ n6508 ;
  assign n6388 = n6276 ^ n6267 ;
  assign n6389 = n6273 & ~n6388 ;
  assign n6390 = n6389 ^ n6276 ;
  assign n6511 = n6510 ^ n6390 ;
  assign n6512 = n6511 ^ x23 ;
  assign n6387 = x91 & n1658 ;
  assign n6513 = n6512 ^ n6387 ;
  assign n6386 = x93 & n1661 ;
  assign n6514 = n6513 ^ n6386 ;
  assign n6385 = n1662 & n2836 ;
  assign n6515 = n6514 ^ n6385 ;
  assign n6517 = n6516 ^ n6515 ;
  assign n6382 = n6286 ^ n6277 ;
  assign n6383 = n6283 & ~n6382 ;
  assign n6384 = n6383 ^ n6286 ;
  assign n6518 = n6517 ^ n6384 ;
  assign n6519 = n6518 ^ x20 ;
  assign n6381 = x94 & n1327 ;
  assign n6520 = n6519 ^ n6381 ;
  assign n6380 = x96 & n1330 ;
  assign n6521 = n6520 ^ n6380 ;
  assign n6379 = n1331 & n3323 ;
  assign n6522 = n6521 ^ n6379 ;
  assign n6524 = n6523 ^ n6522 ;
  assign n6528 = n6527 ^ n6524 ;
  assign n6529 = n6528 ^ x17 ;
  assign n6378 = x97 & n1050 ;
  assign n6530 = n6529 ^ n6378 ;
  assign n6377 = x99 & n1053 ;
  assign n6531 = n6530 ^ n6377 ;
  assign n6376 = n1054 & n3843 ;
  assign n6532 = n6531 ^ n6376 ;
  assign n6534 = n6533 ^ n6532 ;
  assign n6373 = n6303 ^ n6294 ;
  assign n6374 = ~n6300 & ~n6373 ;
  assign n6375 = n6374 ^ n6303 ;
  assign n6535 = n6534 ^ n6375 ;
  assign n6536 = n6535 ^ x14 ;
  assign n6372 = x100 & n877 ;
  assign n6537 = n6536 ^ n6372 ;
  assign n6371 = x102 & n782 ;
  assign n6538 = n6537 ^ n6371 ;
  assign n6370 = n783 & n4410 ;
  assign n6539 = n6538 ^ n6370 ;
  assign n6541 = n6540 ^ n6539 ;
  assign n6545 = n6544 ^ n6541 ;
  assign n6546 = n6545 ^ x11 ;
  assign n6369 = x103 & n647 ;
  assign n6547 = n6546 ^ n6369 ;
  assign n6368 = x105 & ~n572 ;
  assign n6548 = n6547 ^ n6368 ;
  assign n6367 = ~n573 & ~n5023 ;
  assign n6549 = n6548 ^ n6367 ;
  assign n6551 = n6550 ^ n6549 ;
  assign n6555 = n6554 ^ n6551 ;
  assign n6556 = n6555 ^ x8 ;
  assign n6366 = x106 & n446 ;
  assign n6557 = n6556 ^ n6366 ;
  assign n6365 = x108 & n383 ;
  assign n6558 = n6557 ^ n6365 ;
  assign n6364 = n384 & n5670 ;
  assign n6559 = n6558 ^ n6364 ;
  assign n6561 = n6560 ^ n6559 ;
  assign n6565 = n6564 ^ n6561 ;
  assign n6566 = n6565 ^ x5 ;
  assign n6363 = x109 & n234 ;
  assign n6567 = n6566 ^ n6363 ;
  assign n6362 = x111 & n230 ;
  assign n6568 = n6567 ^ n6362 ;
  assign n6360 = n5656 ^ x111 ;
  assign n6361 = n231 & ~n6360 ;
  assign n6569 = n6568 ^ n6361 ;
  assign n6571 = n6570 ^ n6569 ;
  assign n6357 = n6334 ^ n6325 ;
  assign n6358 = ~n6331 & n6357 ;
  assign n6359 = n6358 ^ n6334 ;
  assign n6572 = n6571 ^ n6359 ;
  assign n6342 = ~x113 & ~n6114 ;
  assign n6341 = x113 & ~n6113 ;
  assign n6343 = n6342 ^ n6341 ;
  assign n6345 = x114 ^ x1 ;
  assign n6344 = x114 ^ x2 ;
  assign n6346 = n6345 ^ n6344 ;
  assign n6347 = n6343 & n6346 ;
  assign n6348 = n6347 ^ n6345 ;
  assign n6573 = n6572 ^ n6348 ;
  assign n6352 = x2 & x112 ;
  assign n6353 = n6352 ^ x113 ;
  assign n6354 = ~x1 & n6353 ;
  assign n6349 = n6348 ^ n6116 ;
  assign n6355 = n6354 ^ n6349 ;
  assign n6356 = ~x0 & n6355 ;
  assign n6574 = n6573 ^ n6356 ;
  assign n6578 = n6577 ^ n6574 ;
  assign n6811 = n6565 ^ n6359 ;
  assign n6812 = ~n6571 & ~n6811 ;
  assign n6813 = n6812 ^ n6565 ;
  assign n6809 = x111 & n227 ;
  assign n6802 = x108 & n390 ;
  assign n6795 = x105 & n578 ;
  assign n6788 = x102 & n788 ;
  assign n6780 = n6528 ^ n6375 ;
  assign n6781 = n6534 & ~n6780 ;
  assign n6782 = n6781 ^ n6528 ;
  assign n6778 = x99 & n1058 ;
  assign n6771 = x96 & n1335 ;
  assign n6763 = n6511 ^ n6384 ;
  assign n6764 = ~n6517 & ~n6763 ;
  assign n6765 = n6764 ^ n6511 ;
  assign n6761 = x93 & n1666 ;
  assign n6753 = n6504 ^ n6390 ;
  assign n6754 = ~n6510 & ~n6753 ;
  assign n6755 = n6754 ^ n6504 ;
  assign n6751 = x90 & n2014 ;
  assign n6743 = n6497 ^ n6396 ;
  assign n6744 = ~n6503 & ~n6743 ;
  assign n6745 = n6744 ^ n6497 ;
  assign n6741 = x87 & n2429 ;
  assign n6734 = x84 & n2887 ;
  assign n6732 = n1743 & n2883 ;
  assign n6728 = x83 & n2879 ;
  assign n6727 = x85 & n2882 ;
  assign n6729 = n6728 ^ n6727 ;
  assign n6730 = n6729 ^ x32 ;
  assign n6723 = n6477 ^ n6402 ;
  assign n6724 = ~n6483 & ~n6723 ;
  assign n6725 = n6724 ^ n6477 ;
  assign n6721 = x81 & n3383 ;
  assign n6713 = x75 & n4467 ;
  assign n6705 = n6465 ^ n6452 ;
  assign n6706 = n6457 & n6705 ;
  assign n6707 = n6706 ^ n6452 ;
  assign n6703 = x72 & n5102 ;
  assign n6692 = x68 & n5965 ;
  assign n6691 = x70 & n5729 ;
  assign n6693 = n6692 ^ n6691 ;
  assign n6694 = n6693 ^ x47 ;
  assign n6690 = ~n436 & n5730 ;
  assign n6695 = n6694 ^ n6690 ;
  assign n6689 = x69 & n5736 ;
  assign n6696 = n6695 ^ n6689 ;
  assign n6669 = n6452 ^ n6439 ;
  assign n6686 = n6441 ^ n6439 ;
  assign n6687 = n6669 & n6686 ;
  assign n6675 = x50 ^ x48 ;
  assign n6676 = ~n5972 & n6675 ;
  assign n6677 = n6427 & n6676 ;
  assign n6678 = x65 & n6677 ;
  assign n6674 = x67 & n6428 ;
  assign n6679 = n6678 ^ n6674 ;
  assign n6680 = n6679 ^ x50 ;
  assign n6673 = ~n291 & n6429 ;
  assign n6681 = n6680 ^ n6673 ;
  assign n6672 = x66 & n6433 ;
  assign n6682 = n6681 ^ n6672 ;
  assign n6670 = x51 ^ x50 ;
  assign n6671 = x64 & n6670 ;
  assign n6683 = n6682 ^ n6671 ;
  assign n6684 = n6683 ^ n6441 ;
  assign n6688 = n6687 ^ n6684 ;
  assign n6697 = n6696 ^ n6688 ;
  assign n6668 = n6424 & n6449 ;
  assign n6698 = n6697 ^ n6668 ;
  assign n6699 = n6698 ^ x44 ;
  assign n6667 = x71 & n5094 ;
  assign n6700 = n6699 ^ n6667 ;
  assign n6666 = x73 & n5097 ;
  assign n6701 = n6700 ^ n6666 ;
  assign n6665 = n633 & n5098 ;
  assign n6702 = n6701 ^ n6665 ;
  assign n6704 = n6703 ^ n6702 ;
  assign n6708 = n6707 ^ n6704 ;
  assign n6709 = n6708 ^ x41 ;
  assign n6664 = x74 & n4474 ;
  assign n6710 = n6709 ^ n6664 ;
  assign n6663 = x76 & n4471 ;
  assign n6711 = n6710 ^ n6663 ;
  assign n6662 = ~n853 & n4472 ;
  assign n6712 = n6711 ^ n6662 ;
  assign n6714 = n6713 ^ n6712 ;
  assign n6659 = n6466 ^ n6416 ;
  assign n6660 = ~n6421 & n6659 ;
  assign n6661 = n6660 ^ n6416 ;
  assign n6715 = n6714 ^ n6661 ;
  assign n6649 = x77 & n3916 ;
  assign n6648 = x79 & n3919 ;
  assign n6650 = n6649 ^ n6648 ;
  assign n6651 = n6650 ^ x38 ;
  assign n6647 = n1118 & n3920 ;
  assign n6652 = n6651 ^ n6647 ;
  assign n6646 = x78 & n3924 ;
  assign n6653 = n6652 ^ n6646 ;
  assign n6654 = n6653 ^ n6476 ;
  assign n6655 = n6654 ^ n6467 ;
  assign n6656 = n6655 ^ n6653 ;
  assign n6657 = n6473 & ~n6656 ;
  assign n6658 = n6657 ^ n6654 ;
  assign n6716 = n6715 ^ n6658 ;
  assign n6717 = n6716 ^ x35 ;
  assign n6645 = x80 & n3375 ;
  assign n6718 = n6717 ^ n6645 ;
  assign n6644 = x82 & n3378 ;
  assign n6719 = n6718 ^ n6644 ;
  assign n6643 = n1411 & n3379 ;
  assign n6720 = n6719 ^ n6643 ;
  assign n6722 = n6721 ^ n6720 ;
  assign n6726 = n6725 ^ n6722 ;
  assign n6731 = n6730 ^ n6726 ;
  assign n6733 = n6732 ^ n6731 ;
  assign n6735 = n6734 ^ n6733 ;
  assign n6640 = n6496 ^ n6492 ;
  assign n6641 = n6493 & n6640 ;
  assign n6642 = n6641 ^ n6496 ;
  assign n6736 = n6735 ^ n6642 ;
  assign n6737 = n6736 ^ x29 ;
  assign n6639 = x86 & n2581 ;
  assign n6738 = n6737 ^ n6639 ;
  assign n6638 = x88 & n2422 ;
  assign n6739 = n6738 ^ n6638 ;
  assign n6637 = n2119 & n2423 ;
  assign n6740 = n6739 ^ n6637 ;
  assign n6742 = n6741 ^ n6740 ;
  assign n6746 = n6745 ^ n6742 ;
  assign n6747 = n6746 ^ x26 ;
  assign n6636 = x89 & n2018 ;
  assign n6748 = n6747 ^ n6636 ;
  assign n6635 = x91 & n2021 ;
  assign n6749 = n6748 ^ n6635 ;
  assign n6634 = n2022 & n2542 ;
  assign n6750 = n6749 ^ n6634 ;
  assign n6752 = n6751 ^ n6750 ;
  assign n6756 = n6755 ^ n6752 ;
  assign n6757 = n6756 ^ x23 ;
  assign n6633 = x92 & n1658 ;
  assign n6758 = n6757 ^ n6633 ;
  assign n6632 = x94 & n1661 ;
  assign n6759 = n6758 ^ n6632 ;
  assign n6631 = n1662 & n2997 ;
  assign n6760 = n6759 ^ n6631 ;
  assign n6762 = n6761 ^ n6760 ;
  assign n6766 = n6765 ^ n6762 ;
  assign n6767 = n6766 ^ x20 ;
  assign n6630 = x95 & n1327 ;
  assign n6768 = n6767 ^ n6630 ;
  assign n6629 = x97 & n1330 ;
  assign n6769 = n6768 ^ n6629 ;
  assign n6628 = n1331 & n3494 ;
  assign n6770 = n6769 ^ n6628 ;
  assign n6772 = n6771 ^ n6770 ;
  assign n6625 = n6527 ^ n6518 ;
  assign n6626 = n6524 & n6625 ;
  assign n6627 = n6626 ^ n6527 ;
  assign n6773 = n6772 ^ n6627 ;
  assign n6774 = n6773 ^ x17 ;
  assign n6624 = x98 & n1050 ;
  assign n6775 = n6774 ^ n6624 ;
  assign n6623 = x100 & n1053 ;
  assign n6776 = n6775 ^ n6623 ;
  assign n6622 = n1054 & n4034 ;
  assign n6777 = n6776 ^ n6622 ;
  assign n6779 = n6778 ^ n6777 ;
  assign n6783 = n6782 ^ n6779 ;
  assign n6784 = n6783 ^ x14 ;
  assign n6621 = x101 & n877 ;
  assign n6785 = n6784 ^ n6621 ;
  assign n6620 = x103 & n782 ;
  assign n6786 = n6785 ^ n6620 ;
  assign n6619 = n783 & ~n4615 ;
  assign n6787 = n6786 ^ n6619 ;
  assign n6789 = n6788 ^ n6787 ;
  assign n6616 = n6544 ^ n6535 ;
  assign n6617 = n6541 & n6616 ;
  assign n6618 = n6617 ^ n6544 ;
  assign n6790 = n6789 ^ n6618 ;
  assign n6791 = n6790 ^ x11 ;
  assign n6615 = x104 & n647 ;
  assign n6792 = n6791 ^ n6615 ;
  assign n6614 = x106 & ~n572 ;
  assign n6793 = n6792 ^ n6614 ;
  assign n6613 = ~n573 & ~n5240 ;
  assign n6794 = n6793 ^ n6613 ;
  assign n6796 = n6795 ^ n6794 ;
  assign n6610 = n6554 ^ n6545 ;
  assign n6611 = ~n6551 & n6610 ;
  assign n6612 = n6611 ^ n6554 ;
  assign n6797 = n6796 ^ n6612 ;
  assign n6798 = n6797 ^ x8 ;
  assign n6609 = x107 & n446 ;
  assign n6799 = n6798 ^ n6609 ;
  assign n6608 = x109 & n383 ;
  assign n6800 = n6799 ^ n6608 ;
  assign n6607 = n384 & n5902 ;
  assign n6801 = n6800 ^ n6607 ;
  assign n6803 = n6802 ^ n6801 ;
  assign n6604 = n6564 ^ n6555 ;
  assign n6605 = ~n6561 & ~n6604 ;
  assign n6606 = n6605 ^ n6564 ;
  assign n6804 = n6803 ^ n6606 ;
  assign n6805 = n6804 ^ x5 ;
  assign n6603 = x110 & n234 ;
  assign n6806 = n6805 ^ n6603 ;
  assign n6602 = x112 & n230 ;
  assign n6807 = n6806 ^ n6602 ;
  assign n6600 = n5885 ^ x112 ;
  assign n6601 = n231 & ~n6600 ;
  assign n6808 = n6807 ^ n6601 ;
  assign n6810 = n6809 ^ n6808 ;
  assign n6814 = n6813 ^ n6810 ;
  assign n6585 = x114 & ~n6342 ;
  assign n6584 = ~x114 & ~n6341 ;
  assign n6586 = n6585 ^ n6584 ;
  assign n6588 = x115 ^ x1 ;
  assign n6587 = x115 ^ x2 ;
  assign n6589 = n6588 ^ n6587 ;
  assign n6590 = n6586 & n6589 ;
  assign n6591 = n6590 ^ n6588 ;
  assign n6815 = n6814 ^ n6591 ;
  assign n6595 = x2 & x113 ;
  assign n6596 = n6595 ^ x114 ;
  assign n6597 = ~x1 & n6596 ;
  assign n6592 = n6591 ^ n6344 ;
  assign n6598 = n6597 ^ n6592 ;
  assign n6599 = ~x0 & n6598 ;
  assign n6816 = n6815 ^ n6599 ;
  assign n6579 = n6577 ^ n6572 ;
  assign n6580 = n6574 & ~n6579 ;
  assign n6581 = n6580 ^ n6577 ;
  assign n6817 = n6816 ^ n6581 ;
  assign n7067 = n6814 ^ n6581 ;
  assign n7068 = n6816 & n7067 ;
  assign n7069 = n7068 ^ n6814 ;
  assign n7062 = x112 & n227 ;
  assign n7054 = n6797 ^ n6606 ;
  assign n7055 = n6803 & ~n7054 ;
  assign n7056 = n7055 ^ n6797 ;
  assign n7052 = x109 & n390 ;
  assign n7044 = n6790 ^ n6612 ;
  assign n7045 = n6796 & n7044 ;
  assign n7046 = n7045 ^ n6790 ;
  assign n7042 = x106 & n578 ;
  assign n7034 = n6783 ^ n6618 ;
  assign n7035 = ~n6789 & n7034 ;
  assign n7036 = n7035 ^ n6783 ;
  assign n7032 = x103 & n788 ;
  assign n7025 = x100 & n1058 ;
  assign n7017 = n6766 ^ n6627 ;
  assign n7018 = n6772 & ~n7017 ;
  assign n7019 = n7018 ^ n6766 ;
  assign n7015 = x97 & n1335 ;
  assign n7008 = x94 & n1666 ;
  assign n7001 = x91 & n2014 ;
  assign n6994 = x88 & n2429 ;
  assign n6986 = n6726 ^ n6642 ;
  assign n6987 = ~n6735 & ~n6986 ;
  assign n6988 = n6987 ^ n6726 ;
  assign n6980 = x84 & n2879 ;
  assign n6979 = x86 & n2882 ;
  assign n6981 = n6980 ^ n6979 ;
  assign n6982 = n6981 ^ x32 ;
  assign n6978 = n1857 & n2883 ;
  assign n6983 = n6982 ^ n6978 ;
  assign n6977 = x85 & n2887 ;
  assign n6984 = n6983 ^ n6977 ;
  assign n6974 = x82 & n3383 ;
  assign n6967 = x79 & n3924 ;
  assign n6959 = x73 & n5102 ;
  assign n6948 = x66 & n6677 ;
  assign n6947 = x68 & n6428 ;
  assign n6949 = n6948 ^ n6947 ;
  assign n6950 = n6949 ^ x50 ;
  assign n6946 = ~n340 & n6429 ;
  assign n6951 = n6950 ^ n6946 ;
  assign n6945 = x67 & n6433 ;
  assign n6952 = n6951 ^ n6945 ;
  assign n6939 = x50 & x51 ;
  assign n6940 = n6939 ^ x52 ;
  assign n6941 = ~x64 & n6940 ;
  assign n6935 = x52 ^ x50 ;
  assign n6942 = n6941 ^ n6935 ;
  assign n6933 = x65 ^ x51 ;
  assign n6934 = n6670 & ~n6933 ;
  assign n6943 = n6942 ^ n6934 ;
  assign n6910 = n6441 & n6683 ;
  assign n6911 = n6439 & n6910 ;
  assign n6912 = n6911 ^ n6683 ;
  assign n6932 = n6682 & ~n6912 ;
  assign n6944 = n6943 ^ n6932 ;
  assign n6953 = n6952 ^ n6944 ;
  assign n6924 = n6696 ^ n6668 ;
  assign n6925 = n6924 ^ n6683 ;
  assign n6926 = n6688 & n6925 ;
  assign n6916 = x69 & n5965 ;
  assign n6915 = x71 & n5729 ;
  assign n6917 = n6916 ^ n6915 ;
  assign n6918 = n6917 ^ x47 ;
  assign n6914 = ~n493 & n5730 ;
  assign n6919 = n6918 ^ n6914 ;
  assign n6913 = x70 & n5736 ;
  assign n6920 = n6919 ^ n6913 ;
  assign n6922 = n6920 ^ n6668 ;
  assign n6923 = n6922 ^ n6912 ;
  assign n6927 = n6926 ^ n6923 ;
  assign n6921 = n6920 ^ n6912 ;
  assign n6928 = n6927 ^ n6921 ;
  assign n6929 = ~n6696 & ~n6926 ;
  assign n6930 = n6928 & n6929 ;
  assign n6931 = n6930 ^ n6927 ;
  assign n6954 = n6953 ^ n6931 ;
  assign n6955 = n6954 ^ x44 ;
  assign n6909 = x72 & n5094 ;
  assign n6956 = n6955 ^ n6909 ;
  assign n6908 = x74 & n5097 ;
  assign n6957 = n6956 ^ n6908 ;
  assign n6907 = n699 & n5098 ;
  assign n6958 = n6957 ^ n6907 ;
  assign n6960 = n6959 ^ n6958 ;
  assign n6904 = n6707 ^ n6698 ;
  assign n6905 = ~n6704 & n6904 ;
  assign n6906 = n6905 ^ n6707 ;
  assign n6961 = n6960 ^ n6906 ;
  assign n6894 = x75 & n4474 ;
  assign n6893 = x77 & n4471 ;
  assign n6895 = n6894 ^ n6893 ;
  assign n6896 = n6895 ^ x41 ;
  assign n6892 = ~n939 & n4472 ;
  assign n6897 = n6896 ^ n6892 ;
  assign n6891 = x76 & n4467 ;
  assign n6898 = n6897 ^ n6891 ;
  assign n6899 = n6898 ^ n6708 ;
  assign n6900 = n6899 ^ n6661 ;
  assign n6901 = n6900 ^ n6898 ;
  assign n6902 = n6714 & n6901 ;
  assign n6903 = n6902 ^ n6899 ;
  assign n6962 = n6961 ^ n6903 ;
  assign n6963 = n6962 ^ x38 ;
  assign n6890 = x78 & n3916 ;
  assign n6964 = n6963 ^ n6890 ;
  assign n6889 = x80 & n3919 ;
  assign n6965 = n6964 ^ n6889 ;
  assign n6888 = n1206 & n3920 ;
  assign n6966 = n6965 ^ n6888 ;
  assign n6968 = n6967 ^ n6966 ;
  assign n6885 = n6715 ^ n6653 ;
  assign n6886 = n6658 & n6885 ;
  assign n6887 = n6886 ^ n6653 ;
  assign n6969 = n6968 ^ n6887 ;
  assign n6970 = n6969 ^ x35 ;
  assign n6884 = x81 & n3375 ;
  assign n6971 = n6970 ^ n6884 ;
  assign n6883 = x83 & n3378 ;
  assign n6972 = n6971 ^ n6883 ;
  assign n6882 = n1512 & n3379 ;
  assign n6973 = n6972 ^ n6882 ;
  assign n6975 = n6974 ^ n6973 ;
  assign n6879 = n6725 ^ n6716 ;
  assign n6880 = ~n6722 & ~n6879 ;
  assign n6881 = n6880 ^ n6725 ;
  assign n6976 = n6975 ^ n6881 ;
  assign n6985 = n6984 ^ n6976 ;
  assign n6989 = n6988 ^ n6985 ;
  assign n6990 = n6989 ^ x29 ;
  assign n6878 = x87 & n2581 ;
  assign n6991 = n6990 ^ n6878 ;
  assign n6877 = x89 & n2422 ;
  assign n6992 = n6991 ^ n6877 ;
  assign n6876 = n2249 & n2423 ;
  assign n6993 = n6992 ^ n6876 ;
  assign n6995 = n6994 ^ n6993 ;
  assign n6873 = n6745 ^ n6736 ;
  assign n6874 = n6742 & n6873 ;
  assign n6875 = n6874 ^ n6745 ;
  assign n6996 = n6995 ^ n6875 ;
  assign n6997 = n6996 ^ x26 ;
  assign n6872 = x90 & n2018 ;
  assign n6998 = n6997 ^ n6872 ;
  assign n6871 = x92 & n2021 ;
  assign n6999 = n6998 ^ n6871 ;
  assign n6870 = n2022 & n2684 ;
  assign n7000 = n6999 ^ n6870 ;
  assign n7002 = n7001 ^ n7000 ;
  assign n6867 = n6755 ^ n6746 ;
  assign n6868 = ~n6752 & ~n6867 ;
  assign n6869 = n6868 ^ n6755 ;
  assign n7003 = n7002 ^ n6869 ;
  assign n7004 = n7003 ^ x23 ;
  assign n6866 = x93 & n1658 ;
  assign n7005 = n7004 ^ n6866 ;
  assign n6865 = x95 & n1661 ;
  assign n7006 = n7005 ^ n6865 ;
  assign n6864 = n1662 & n3159 ;
  assign n7007 = n7006 ^ n6864 ;
  assign n7009 = n7008 ^ n7007 ;
  assign n6861 = n6765 ^ n6756 ;
  assign n6862 = n6762 & n6861 ;
  assign n6863 = n6862 ^ n6765 ;
  assign n7010 = n7009 ^ n6863 ;
  assign n7011 = n7010 ^ x20 ;
  assign n6860 = x96 & n1327 ;
  assign n7012 = n7011 ^ n6860 ;
  assign n6859 = x98 & n1330 ;
  assign n7013 = n7012 ^ n6859 ;
  assign n6858 = n1331 & n3660 ;
  assign n7014 = n7013 ^ n6858 ;
  assign n7016 = n7015 ^ n7014 ;
  assign n7020 = n7019 ^ n7016 ;
  assign n7021 = n7020 ^ x17 ;
  assign n6857 = x99 & n1050 ;
  assign n7022 = n7021 ^ n6857 ;
  assign n6856 = x101 & n1053 ;
  assign n7023 = n7022 ^ n6856 ;
  assign n6855 = n1054 & n4215 ;
  assign n7024 = n7023 ^ n6855 ;
  assign n7026 = n7025 ^ n7024 ;
  assign n6852 = n6782 ^ n6773 ;
  assign n6853 = n6779 & ~n6852 ;
  assign n6854 = n6853 ^ n6782 ;
  assign n7027 = n7026 ^ n6854 ;
  assign n7028 = n7027 ^ x14 ;
  assign n6851 = x102 & n877 ;
  assign n7029 = n7028 ^ n6851 ;
  assign n6850 = x104 & n782 ;
  assign n7030 = n7029 ^ n6850 ;
  assign n6849 = n783 & ~n4814 ;
  assign n7031 = n7030 ^ n6849 ;
  assign n7033 = n7032 ^ n7031 ;
  assign n7037 = n7036 ^ n7033 ;
  assign n7038 = n7037 ^ x11 ;
  assign n6848 = x105 & n647 ;
  assign n7039 = n7038 ^ n6848 ;
  assign n6847 = x107 & ~n572 ;
  assign n7040 = n7039 ^ n6847 ;
  assign n6846 = ~n573 & ~n5448 ;
  assign n7041 = n7040 ^ n6846 ;
  assign n7043 = n7042 ^ n7041 ;
  assign n7047 = n7046 ^ n7043 ;
  assign n7048 = n7047 ^ x8 ;
  assign n6845 = x108 & n446 ;
  assign n7049 = n7048 ^ n6845 ;
  assign n6844 = x110 & n383 ;
  assign n7050 = n7049 ^ n6844 ;
  assign n6843 = n384 & n6129 ;
  assign n7051 = n7050 ^ n6843 ;
  assign n7053 = n7052 ^ n7051 ;
  assign n7057 = n7056 ^ n7053 ;
  assign n7058 = n7057 ^ x5 ;
  assign n6842 = x111 & n234 ;
  assign n7059 = n7058 ^ n6842 ;
  assign n6841 = x113 & n230 ;
  assign n7060 = n7059 ^ n6841 ;
  assign n6839 = n6115 ^ x113 ;
  assign n6840 = n231 & ~n6839 ;
  assign n7061 = n7060 ^ n6840 ;
  assign n7063 = n7062 ^ n7061 ;
  assign n6836 = n6813 ^ n6804 ;
  assign n6837 = n6810 & n6836 ;
  assign n6838 = n6837 ^ n6813 ;
  assign n7064 = n7063 ^ n6838 ;
  assign n6821 = ~x115 & ~n6585 ;
  assign n6820 = x115 & ~n6584 ;
  assign n6822 = n6821 ^ n6820 ;
  assign n6824 = x116 ^ x1 ;
  assign n6823 = x116 ^ x2 ;
  assign n6825 = n6824 ^ n6823 ;
  assign n6826 = n6822 & n6825 ;
  assign n6827 = n6826 ^ n6824 ;
  assign n7065 = n7064 ^ n6827 ;
  assign n6831 = x2 & x114 ;
  assign n6832 = n6831 ^ x115 ;
  assign n6833 = ~n255 & n6832 ;
  assign n6828 = n6827 ^ n6587 ;
  assign n6834 = n6833 ^ n6828 ;
  assign n6835 = ~x0 & n6834 ;
  assign n7066 = n7065 ^ n6835 ;
  assign n7070 = n7069 ^ n7066 ;
  assign n7315 = n7057 ^ n6838 ;
  assign n7316 = n7063 & ~n7315 ;
  assign n7317 = n7316 ^ n7057 ;
  assign n7313 = x113 & n227 ;
  assign n7306 = x110 & n390 ;
  assign n7299 = x107 & n578 ;
  assign n7292 = x104 & n788 ;
  assign n7284 = n7020 ^ n6854 ;
  assign n7285 = ~n7026 & ~n7284 ;
  assign n7286 = n7285 ^ n7020 ;
  assign n7282 = x101 & n1058 ;
  assign n7275 = x98 & n1335 ;
  assign n7267 = n7003 ^ n6863 ;
  assign n7268 = n7009 & ~n7267 ;
  assign n7269 = n7268 ^ n7003 ;
  assign n7265 = x95 & n1666 ;
  assign n7257 = n6996 ^ n6869 ;
  assign n7258 = ~n7002 & n7257 ;
  assign n7259 = n7258 ^ n6996 ;
  assign n7255 = x92 & n2014 ;
  assign n7247 = n6989 ^ n6875 ;
  assign n7248 = n6995 & ~n7247 ;
  assign n7249 = n7248 ^ n6989 ;
  assign n7245 = x89 & n2429 ;
  assign n7238 = x86 & n2887 ;
  assign n7230 = n6969 ^ n6881 ;
  assign n7231 = n6975 & ~n7230 ;
  assign n7232 = n7231 ^ n6969 ;
  assign n7228 = x83 & n3383 ;
  assign n7218 = x79 & n3916 ;
  assign n7217 = x81 & n3919 ;
  assign n7219 = n7218 ^ n7217 ;
  assign n7220 = n7219 ^ x38 ;
  assign n7216 = n1305 & n3920 ;
  assign n7221 = n7220 ^ n7216 ;
  assign n7215 = x80 & n3924 ;
  assign n7222 = n7221 ^ n7215 ;
  assign n7211 = x77 & n4467 ;
  assign n7204 = x74 & n5102 ;
  assign n7197 = x71 & n5736 ;
  assign n7190 = x68 & n6433 ;
  assign n7183 = x53 & ~n6671 ;
  assign n7184 = ~n6943 & n7183 ;
  assign n6937 = x52 ^ x51 ;
  assign n7179 = ~n6670 & n6937 ;
  assign n7180 = x65 & n7179 ;
  assign n7168 = x53 ^ x52 ;
  assign n7174 = n6670 & ~n7168 ;
  assign n7175 = n7174 ^ n6670 ;
  assign n7176 = ~n150 & n7175 ;
  assign n7173 = x66 & n6670 ;
  assign n7177 = n7176 ^ n7173 ;
  assign n7178 = n7177 ^ x53 ;
  assign n7181 = n7180 ^ n7178 ;
  assign n7169 = x53 ^ x51 ;
  assign n7170 = ~n6670 & n7169 ;
  assign n7171 = n7168 & n7170 ;
  assign n7172 = x64 & n7171 ;
  assign n7182 = n7181 ^ n7172 ;
  assign n7185 = n7184 ^ n7182 ;
  assign n7186 = n7185 ^ x50 ;
  assign n7167 = x67 & n6677 ;
  assign n7187 = n7186 ^ n7167 ;
  assign n7166 = x69 & n6428 ;
  assign n7188 = n7187 ^ n7166 ;
  assign n7165 = ~n375 & n6429 ;
  assign n7189 = n7188 ^ n7165 ;
  assign n7191 = n7190 ^ n7189 ;
  assign n7162 = n6952 ^ n6943 ;
  assign n7163 = ~n6944 & n7162 ;
  assign n7164 = n7163 ^ n6952 ;
  assign n7192 = n7191 ^ n7164 ;
  assign n7193 = n7192 ^ x47 ;
  assign n7161 = x70 & n5965 ;
  assign n7194 = n7193 ^ n7161 ;
  assign n7160 = x72 & n5729 ;
  assign n7195 = n7194 ^ n7160 ;
  assign n7159 = n556 & n5730 ;
  assign n7196 = n7195 ^ n7159 ;
  assign n7198 = n7197 ^ n7196 ;
  assign n7156 = n6953 ^ n6920 ;
  assign n7157 = n6931 & n7156 ;
  assign n7158 = n7157 ^ n6920 ;
  assign n7199 = n7198 ^ n7158 ;
  assign n7200 = n7199 ^ x44 ;
  assign n7155 = x73 & n5094 ;
  assign n7201 = n7200 ^ n7155 ;
  assign n7154 = x75 & n5097 ;
  assign n7202 = n7201 ^ n7154 ;
  assign n7153 = ~n774 & n5098 ;
  assign n7203 = n7202 ^ n7153 ;
  assign n7205 = n7204 ^ n7203 ;
  assign n7150 = n6954 ^ n6906 ;
  assign n7151 = n6960 & n7150 ;
  assign n7152 = n7151 ^ n6954 ;
  assign n7206 = n7205 ^ n7152 ;
  assign n7207 = n7206 ^ x41 ;
  assign n7149 = x76 & n4474 ;
  assign n7208 = n7207 ^ n7149 ;
  assign n7148 = x78 & n4471 ;
  assign n7209 = n7208 ^ n7148 ;
  assign n7147 = ~n1025 & n4472 ;
  assign n7210 = n7209 ^ n7147 ;
  assign n7212 = n7211 ^ n7210 ;
  assign n7144 = n6961 ^ n6898 ;
  assign n7145 = n6903 & n7144 ;
  assign n7146 = n7145 ^ n6898 ;
  assign n7213 = n7212 ^ n7146 ;
  assign n7141 = n6962 ^ n6887 ;
  assign n7142 = n6968 & n7141 ;
  assign n7143 = n7142 ^ n6962 ;
  assign n7214 = n7213 ^ n7143 ;
  assign n7223 = n7222 ^ n7214 ;
  assign n7224 = n7223 ^ x35 ;
  assign n7140 = x82 & n3375 ;
  assign n7225 = n7224 ^ n7140 ;
  assign n7139 = x84 & n3378 ;
  assign n7226 = n7225 ^ n7139 ;
  assign n7138 = n1624 & n3379 ;
  assign n7227 = n7226 ^ n7138 ;
  assign n7229 = n7228 ^ n7227 ;
  assign n7233 = n7232 ^ n7229 ;
  assign n7234 = n7233 ^ x32 ;
  assign n7137 = x85 & n2879 ;
  assign n7235 = n7234 ^ n7137 ;
  assign n7136 = x87 & n2882 ;
  assign n7236 = n7235 ^ n7136 ;
  assign n7135 = n1982 & n2883 ;
  assign n7237 = n7236 ^ n7135 ;
  assign n7239 = n7238 ^ n7237 ;
  assign n7132 = n6988 ^ n6984 ;
  assign n7133 = n6985 & ~n7132 ;
  assign n7134 = n7133 ^ n6988 ;
  assign n7240 = n7239 ^ n7134 ;
  assign n7241 = n7240 ^ x29 ;
  assign n7131 = x88 & n2581 ;
  assign n7242 = n7241 ^ n7131 ;
  assign n7130 = x90 & n2422 ;
  assign n7243 = n7242 ^ n7130 ;
  assign n7129 = n2386 & n2423 ;
  assign n7244 = n7243 ^ n7129 ;
  assign n7246 = n7245 ^ n7244 ;
  assign n7250 = n7249 ^ n7246 ;
  assign n7251 = n7250 ^ x26 ;
  assign n7128 = x91 & n2018 ;
  assign n7252 = n7251 ^ n7128 ;
  assign n7127 = x93 & n2021 ;
  assign n7253 = n7252 ^ n7127 ;
  assign n7126 = n2022 & n2836 ;
  assign n7254 = n7253 ^ n7126 ;
  assign n7256 = n7255 ^ n7254 ;
  assign n7260 = n7259 ^ n7256 ;
  assign n7261 = n7260 ^ x23 ;
  assign n7125 = x94 & n1658 ;
  assign n7262 = n7261 ^ n7125 ;
  assign n7124 = x96 & n1661 ;
  assign n7263 = n7262 ^ n7124 ;
  assign n7123 = n1662 & n3323 ;
  assign n7264 = n7263 ^ n7123 ;
  assign n7266 = n7265 ^ n7264 ;
  assign n7270 = n7269 ^ n7266 ;
  assign n7271 = n7270 ^ x20 ;
  assign n7122 = x97 & n1327 ;
  assign n7272 = n7271 ^ n7122 ;
  assign n7121 = x99 & n1330 ;
  assign n7273 = n7272 ^ n7121 ;
  assign n7120 = n1331 & n3843 ;
  assign n7274 = n7273 ^ n7120 ;
  assign n7276 = n7275 ^ n7274 ;
  assign n7117 = n7019 ^ n7010 ;
  assign n7118 = n7016 & ~n7117 ;
  assign n7119 = n7118 ^ n7019 ;
  assign n7277 = n7276 ^ n7119 ;
  assign n7278 = n7277 ^ x17 ;
  assign n7116 = x100 & n1050 ;
  assign n7279 = n7278 ^ n7116 ;
  assign n7115 = x102 & n1053 ;
  assign n7280 = n7279 ^ n7115 ;
  assign n7114 = n1054 & n4410 ;
  assign n7281 = n7280 ^ n7114 ;
  assign n7283 = n7282 ^ n7281 ;
  assign n7287 = n7286 ^ n7283 ;
  assign n7288 = n7287 ^ x14 ;
  assign n7113 = x103 & n877 ;
  assign n7289 = n7288 ^ n7113 ;
  assign n7112 = x105 & n782 ;
  assign n7290 = n7289 ^ n7112 ;
  assign n7111 = n783 & ~n5023 ;
  assign n7291 = n7290 ^ n7111 ;
  assign n7293 = n7292 ^ n7291 ;
  assign n7108 = n7036 ^ n7027 ;
  assign n7109 = n7033 & n7108 ;
  assign n7110 = n7109 ^ n7036 ;
  assign n7294 = n7293 ^ n7110 ;
  assign n7295 = n7294 ^ x11 ;
  assign n7107 = x106 & n647 ;
  assign n7296 = n7295 ^ n7107 ;
  assign n7106 = x108 & ~n572 ;
  assign n7297 = n7296 ^ n7106 ;
  assign n7105 = ~n573 & n5670 ;
  assign n7298 = n7297 ^ n7105 ;
  assign n7300 = n7299 ^ n7298 ;
  assign n7102 = n7046 ^ n7037 ;
  assign n7103 = ~n7043 & n7102 ;
  assign n7104 = n7103 ^ n7046 ;
  assign n7301 = n7300 ^ n7104 ;
  assign n7302 = n7301 ^ x8 ;
  assign n7101 = x109 & n446 ;
  assign n7303 = n7302 ^ n7101 ;
  assign n7100 = x111 & n383 ;
  assign n7304 = n7303 ^ n7100 ;
  assign n7099 = n384 & ~n6360 ;
  assign n7305 = n7304 ^ n7099 ;
  assign n7307 = n7306 ^ n7305 ;
  assign n7096 = n7056 ^ n7047 ;
  assign n7097 = ~n7053 & n7096 ;
  assign n7098 = n7097 ^ n7056 ;
  assign n7308 = n7307 ^ n7098 ;
  assign n7309 = n7308 ^ x5 ;
  assign n7095 = x112 & n234 ;
  assign n7310 = n7309 ^ n7095 ;
  assign n7094 = x114 & n230 ;
  assign n7311 = n7310 ^ n7094 ;
  assign n7092 = n6343 ^ x114 ;
  assign n7093 = n231 & ~n7092 ;
  assign n7312 = n7311 ^ n7093 ;
  assign n7314 = n7313 ^ n7312 ;
  assign n7318 = n7317 ^ n7314 ;
  assign n7077 = x116 & ~n6821 ;
  assign n7076 = ~x116 & ~n6820 ;
  assign n7078 = n7077 ^ n7076 ;
  assign n7080 = x117 ^ x1 ;
  assign n7079 = x117 ^ x2 ;
  assign n7081 = n7080 ^ n7079 ;
  assign n7082 = n7078 & n7081 ;
  assign n7083 = n7082 ^ n7080 ;
  assign n7319 = n7318 ^ n7083 ;
  assign n7087 = x2 & x115 ;
  assign n7088 = n7087 ^ x116 ;
  assign n7089 = ~n255 & n7088 ;
  assign n7084 = n7083 ^ n6823 ;
  assign n7090 = n7089 ^ n7084 ;
  assign n7091 = ~x0 & n7090 ;
  assign n7320 = n7319 ^ n7091 ;
  assign n7071 = n7069 ^ n7064 ;
  assign n7072 = n7066 & ~n7071 ;
  assign n7073 = n7072 ^ n7069 ;
  assign n7321 = n7320 ^ n7073 ;
  assign n7565 = n7318 ^ n7073 ;
  assign n7566 = n7320 & n7565 ;
  assign n7567 = n7566 ^ n7318 ;
  assign n7560 = x114 & n227 ;
  assign n7552 = n7301 ^ n7098 ;
  assign n7553 = n7307 & n7552 ;
  assign n7554 = n7553 ^ n7301 ;
  assign n7550 = x111 & n390 ;
  assign n7542 = n7294 ^ n7104 ;
  assign n7543 = n7300 & n7542 ;
  assign n7544 = n7543 ^ n7294 ;
  assign n7536 = x107 & n647 ;
  assign n7535 = x109 & ~n572 ;
  assign n7537 = n7536 ^ n7535 ;
  assign n7538 = n7537 ^ x11 ;
  assign n7534 = ~n573 & n5902 ;
  assign n7539 = n7538 ^ n7534 ;
  assign n7533 = x108 & n578 ;
  assign n7540 = n7539 ^ n7533 ;
  assign n7529 = n7287 ^ n7110 ;
  assign n7530 = ~n7293 & n7529 ;
  assign n7531 = n7530 ^ n7287 ;
  assign n7527 = x105 & n788 ;
  assign n7520 = x102 & n1058 ;
  assign n7512 = n7270 ^ n7119 ;
  assign n7513 = n7276 & n7512 ;
  assign n7514 = n7513 ^ n7270 ;
  assign n7510 = x99 & n1335 ;
  assign n7503 = x96 & n1666 ;
  assign n7496 = x93 & n2014 ;
  assign n7489 = x90 & n2429 ;
  assign n7481 = n7233 ^ n7134 ;
  assign n7482 = n7239 & ~n7481 ;
  assign n7483 = n7482 ^ n7233 ;
  assign n7479 = x87 & n2887 ;
  assign n7472 = x84 & n3383 ;
  assign n7465 = x81 & n3924 ;
  assign n7457 = x75 & n5102 ;
  assign n7450 = x72 & n5736 ;
  assign n7442 = n7185 ^ n7164 ;
  assign n7443 = n7191 & n7442 ;
  assign n7444 = n7443 ^ n7185 ;
  assign n7440 = x69 & n6433 ;
  assign n7429 = x65 & n7171 ;
  assign n7428 = x67 & n7174 ;
  assign n7430 = n7429 ^ n7428 ;
  assign n7431 = n7430 ^ x53 ;
  assign n7427 = ~n291 & n7175 ;
  assign n7432 = n7431 ^ n7427 ;
  assign n7426 = x66 & n7179 ;
  assign n7433 = n7432 ^ n7426 ;
  assign n7424 = x54 ^ x53 ;
  assign n7425 = x64 & n7424 ;
  assign n7434 = n7433 ^ n7425 ;
  assign n7423 = n7182 & n7184 ;
  assign n7435 = n7434 ^ n7423 ;
  assign n7436 = n7435 ^ x50 ;
  assign n7422 = x68 & n6677 ;
  assign n7437 = n7436 ^ n7422 ;
  assign n7421 = x70 & n6428 ;
  assign n7438 = n7437 ^ n7421 ;
  assign n7420 = ~n436 & n6429 ;
  assign n7439 = n7438 ^ n7420 ;
  assign n7441 = n7440 ^ n7439 ;
  assign n7445 = n7444 ^ n7441 ;
  assign n7446 = n7445 ^ x47 ;
  assign n7419 = x71 & n5965 ;
  assign n7447 = n7446 ^ n7419 ;
  assign n7418 = x73 & n5729 ;
  assign n7448 = n7447 ^ n7418 ;
  assign n7417 = n633 & n5730 ;
  assign n7449 = n7448 ^ n7417 ;
  assign n7451 = n7450 ^ n7449 ;
  assign n7414 = n7192 ^ n7158 ;
  assign n7415 = n7198 & n7414 ;
  assign n7416 = n7415 ^ n7192 ;
  assign n7452 = n7451 ^ n7416 ;
  assign n7453 = n7452 ^ x44 ;
  assign n7413 = x74 & n5094 ;
  assign n7454 = n7453 ^ n7413 ;
  assign n7412 = x76 & n5097 ;
  assign n7455 = n7454 ^ n7412 ;
  assign n7411 = ~n853 & n5098 ;
  assign n7456 = n7455 ^ n7411 ;
  assign n7458 = n7457 ^ n7456 ;
  assign n7408 = n7199 ^ n7152 ;
  assign n7409 = n7205 & n7408 ;
  assign n7410 = n7409 ^ n7199 ;
  assign n7459 = n7458 ^ n7410 ;
  assign n7398 = x77 & n4474 ;
  assign n7397 = x79 & n4471 ;
  assign n7399 = n7398 ^ n7397 ;
  assign n7400 = n7399 ^ x41 ;
  assign n7396 = n1118 & n4472 ;
  assign n7401 = n7400 ^ n7396 ;
  assign n7395 = x78 & n4467 ;
  assign n7402 = n7401 ^ n7395 ;
  assign n7403 = n7402 ^ n7206 ;
  assign n7404 = n7403 ^ n7146 ;
  assign n7405 = n7404 ^ n7402 ;
  assign n7406 = n7212 & n7405 ;
  assign n7407 = n7406 ^ n7403 ;
  assign n7460 = n7459 ^ n7407 ;
  assign n7461 = n7460 ^ x38 ;
  assign n7394 = x80 & n3916 ;
  assign n7462 = n7461 ^ n7394 ;
  assign n7393 = x82 & n3919 ;
  assign n7463 = n7462 ^ n7393 ;
  assign n7392 = n1411 & n3920 ;
  assign n7464 = n7463 ^ n7392 ;
  assign n7466 = n7465 ^ n7464 ;
  assign n7389 = n7222 ^ n7143 ;
  assign n7390 = ~n7214 & n7389 ;
  assign n7391 = n7390 ^ n7222 ;
  assign n7467 = n7466 ^ n7391 ;
  assign n7468 = n7467 ^ x35 ;
  assign n7388 = x83 & n3375 ;
  assign n7469 = n7468 ^ n7388 ;
  assign n7387 = x85 & n3378 ;
  assign n7470 = n7469 ^ n7387 ;
  assign n7386 = n1743 & n3379 ;
  assign n7471 = n7470 ^ n7386 ;
  assign n7473 = n7472 ^ n7471 ;
  assign n7383 = n7232 ^ n7223 ;
  assign n7384 = ~n7229 & n7383 ;
  assign n7385 = n7384 ^ n7232 ;
  assign n7474 = n7473 ^ n7385 ;
  assign n7475 = n7474 ^ x32 ;
  assign n7382 = x86 & n2879 ;
  assign n7476 = n7475 ^ n7382 ;
  assign n7381 = x88 & n2882 ;
  assign n7477 = n7476 ^ n7381 ;
  assign n7380 = n2119 & n2883 ;
  assign n7478 = n7477 ^ n7380 ;
  assign n7480 = n7479 ^ n7478 ;
  assign n7484 = n7483 ^ n7480 ;
  assign n7485 = n7484 ^ x29 ;
  assign n7379 = x89 & n2581 ;
  assign n7486 = n7485 ^ n7379 ;
  assign n7378 = x91 & n2422 ;
  assign n7487 = n7486 ^ n7378 ;
  assign n7377 = n2423 & n2542 ;
  assign n7488 = n7487 ^ n7377 ;
  assign n7490 = n7489 ^ n7488 ;
  assign n7374 = n7249 ^ n7240 ;
  assign n7375 = n7246 & ~n7374 ;
  assign n7376 = n7375 ^ n7249 ;
  assign n7491 = n7490 ^ n7376 ;
  assign n7492 = n7491 ^ x26 ;
  assign n7373 = x92 & n2018 ;
  assign n7493 = n7492 ^ n7373 ;
  assign n7372 = x94 & n2021 ;
  assign n7494 = n7493 ^ n7372 ;
  assign n7371 = n2022 & n2997 ;
  assign n7495 = n7494 ^ n7371 ;
  assign n7497 = n7496 ^ n7495 ;
  assign n7368 = n7259 ^ n7250 ;
  assign n7369 = n7256 & n7368 ;
  assign n7370 = n7369 ^ n7259 ;
  assign n7498 = n7497 ^ n7370 ;
  assign n7499 = n7498 ^ x23 ;
  assign n7367 = x95 & n1658 ;
  assign n7500 = n7499 ^ n7367 ;
  assign n7366 = x97 & n1661 ;
  assign n7501 = n7500 ^ n7366 ;
  assign n7365 = n1662 & n3494 ;
  assign n7502 = n7501 ^ n7365 ;
  assign n7504 = n7503 ^ n7502 ;
  assign n7362 = n7269 ^ n7260 ;
  assign n7363 = ~n7266 & n7362 ;
  assign n7364 = n7363 ^ n7269 ;
  assign n7505 = n7504 ^ n7364 ;
  assign n7506 = n7505 ^ x20 ;
  assign n7361 = x98 & n1327 ;
  assign n7507 = n7506 ^ n7361 ;
  assign n7360 = x100 & n1330 ;
  assign n7508 = n7507 ^ n7360 ;
  assign n7359 = n1331 & n4034 ;
  assign n7509 = n7508 ^ n7359 ;
  assign n7511 = n7510 ^ n7509 ;
  assign n7515 = n7514 ^ n7511 ;
  assign n7516 = n7515 ^ x17 ;
  assign n7358 = x101 & n1050 ;
  assign n7517 = n7516 ^ n7358 ;
  assign n7357 = x103 & n1053 ;
  assign n7518 = n7517 ^ n7357 ;
  assign n7356 = n1054 & ~n4615 ;
  assign n7519 = n7518 ^ n7356 ;
  assign n7521 = n7520 ^ n7519 ;
  assign n7353 = n7286 ^ n7277 ;
  assign n7354 = ~n7283 & ~n7353 ;
  assign n7355 = n7354 ^ n7286 ;
  assign n7522 = n7521 ^ n7355 ;
  assign n7523 = n7522 ^ x14 ;
  assign n7352 = x104 & n877 ;
  assign n7524 = n7523 ^ n7352 ;
  assign n7351 = x106 & n782 ;
  assign n7525 = n7524 ^ n7351 ;
  assign n7350 = n783 & ~n5240 ;
  assign n7526 = n7525 ^ n7350 ;
  assign n7528 = n7527 ^ n7526 ;
  assign n7532 = n7531 ^ n7528 ;
  assign n7541 = n7540 ^ n7532 ;
  assign n7545 = n7544 ^ n7541 ;
  assign n7546 = n7545 ^ x8 ;
  assign n7349 = x110 & n446 ;
  assign n7547 = n7546 ^ n7349 ;
  assign n7348 = x112 & n383 ;
  assign n7548 = n7547 ^ n7348 ;
  assign n7347 = n384 & ~n6600 ;
  assign n7549 = n7548 ^ n7347 ;
  assign n7551 = n7550 ^ n7549 ;
  assign n7555 = n7554 ^ n7551 ;
  assign n7556 = n7555 ^ x5 ;
  assign n7346 = x113 & n234 ;
  assign n7557 = n7556 ^ n7346 ;
  assign n7345 = x115 & n230 ;
  assign n7558 = n7557 ^ n7345 ;
  assign n7343 = n6586 ^ x115 ;
  assign n7344 = n231 & ~n7343 ;
  assign n7559 = n7558 ^ n7344 ;
  assign n7561 = n7560 ^ n7559 ;
  assign n7340 = n7317 ^ n7308 ;
  assign n7341 = ~n7314 & n7340 ;
  assign n7342 = n7341 ^ n7317 ;
  assign n7562 = n7561 ^ n7342 ;
  assign n7325 = ~x117 & ~n7077 ;
  assign n7324 = x117 & ~n7076 ;
  assign n7326 = n7325 ^ n7324 ;
  assign n7328 = x118 ^ x1 ;
  assign n7327 = x118 ^ x2 ;
  assign n7329 = n7328 ^ n7327 ;
  assign n7330 = n7326 & n7329 ;
  assign n7331 = n7330 ^ n7328 ;
  assign n7563 = n7562 ^ n7331 ;
  assign n7335 = x2 & x116 ;
  assign n7336 = n7335 ^ x117 ;
  assign n7337 = ~x1 & n7336 ;
  assign n7332 = n7331 ^ n7079 ;
  assign n7338 = n7337 ^ n7332 ;
  assign n7339 = ~x0 & n7338 ;
  assign n7564 = n7563 ^ n7339 ;
  assign n7568 = n7567 ^ n7564 ;
  assign n7818 = n7555 ^ n7342 ;
  assign n7819 = ~n7561 & ~n7818 ;
  assign n7820 = n7819 ^ n7555 ;
  assign n7816 = x115 & n227 ;
  assign n7809 = x112 & n390 ;
  assign n7802 = x109 & n578 ;
  assign n7795 = x106 & n788 ;
  assign n7787 = n7515 ^ n7355 ;
  assign n7788 = ~n7521 & n7787 ;
  assign n7789 = n7788 ^ n7515 ;
  assign n7785 = x103 & n1058 ;
  assign n7778 = x100 & n1335 ;
  assign n7770 = n7498 ^ n7364 ;
  assign n7771 = ~n7504 & ~n7770 ;
  assign n7772 = n7771 ^ n7498 ;
  assign n7768 = x97 & n1666 ;
  assign n7760 = n7491 ^ n7370 ;
  assign n7761 = n7497 & ~n7760 ;
  assign n7762 = n7761 ^ n7491 ;
  assign n7758 = x94 & n2014 ;
  assign n7750 = n7484 ^ n7376 ;
  assign n7751 = n7490 & n7750 ;
  assign n7752 = n7751 ^ n7484 ;
  assign n7748 = x91 & n2429 ;
  assign n7741 = x88 & n2887 ;
  assign n7733 = n7467 ^ n7385 ;
  assign n7734 = n7473 & n7733 ;
  assign n7735 = n7734 ^ n7467 ;
  assign n7731 = x85 & n3383 ;
  assign n7724 = x82 & n3924 ;
  assign n7717 = x79 & n4467 ;
  assign n7708 = n7445 ^ n7416 ;
  assign n7709 = n7451 & n7708 ;
  assign n7710 = n7709 ^ n7445 ;
  assign n7706 = x73 & n5736 ;
  assign n7699 = x70 & n6433 ;
  assign n7691 = ~n7425 & n7433 ;
  assign n7692 = ~n7423 & n7691 ;
  assign n7693 = n7692 ^ n7433 ;
  assign n7685 = x66 & n7171 ;
  assign n7684 = x68 & n7174 ;
  assign n7686 = n7685 ^ n7684 ;
  assign n7687 = n7686 ^ x53 ;
  assign n7683 = ~n340 & n7175 ;
  assign n7688 = n7687 ^ n7683 ;
  assign n7682 = x67 & n7179 ;
  assign n7689 = n7688 ^ n7682 ;
  assign n7679 = x65 ^ x54 ;
  assign n7680 = n7424 & ~n7679 ;
  assign n7675 = x53 & x54 ;
  assign n7676 = n7675 ^ x55 ;
  assign n7677 = ~x64 & n7676 ;
  assign n7671 = x55 ^ x53 ;
  assign n7678 = n7677 ^ n7671 ;
  assign n7681 = n7680 ^ n7678 ;
  assign n7690 = n7689 ^ n7681 ;
  assign n7694 = n7693 ^ n7690 ;
  assign n7695 = n7694 ^ x50 ;
  assign n7670 = x69 & n6677 ;
  assign n7696 = n7695 ^ n7670 ;
  assign n7669 = x71 & n6428 ;
  assign n7697 = n7696 ^ n7669 ;
  assign n7668 = ~n493 & n6429 ;
  assign n7698 = n7697 ^ n7668 ;
  assign n7700 = n7699 ^ n7698 ;
  assign n7665 = n7444 ^ n7435 ;
  assign n7666 = ~n7441 & n7665 ;
  assign n7667 = n7666 ^ n7444 ;
  assign n7701 = n7700 ^ n7667 ;
  assign n7702 = n7701 ^ x47 ;
  assign n7664 = x72 & n5965 ;
  assign n7703 = n7702 ^ n7664 ;
  assign n7663 = x74 & n5729 ;
  assign n7704 = n7703 ^ n7663 ;
  assign n7662 = n699 & n5730 ;
  assign n7705 = n7704 ^ n7662 ;
  assign n7707 = n7706 ^ n7705 ;
  assign n7711 = n7710 ^ n7707 ;
  assign n7652 = x75 & n5094 ;
  assign n7651 = x77 & n5097 ;
  assign n7653 = n7652 ^ n7651 ;
  assign n7654 = n7653 ^ x44 ;
  assign n7650 = ~n939 & n5098 ;
  assign n7655 = n7654 ^ n7650 ;
  assign n7649 = x76 & n5102 ;
  assign n7656 = n7655 ^ n7649 ;
  assign n7657 = n7656 ^ n7452 ;
  assign n7658 = n7657 ^ n7410 ;
  assign n7659 = n7658 ^ n7656 ;
  assign n7660 = n7458 & n7659 ;
  assign n7661 = n7660 ^ n7657 ;
  assign n7712 = n7711 ^ n7661 ;
  assign n7713 = n7712 ^ x41 ;
  assign n7648 = x78 & n4474 ;
  assign n7714 = n7713 ^ n7648 ;
  assign n7647 = x80 & n4471 ;
  assign n7715 = n7714 ^ n7647 ;
  assign n7646 = n1206 & n4472 ;
  assign n7716 = n7715 ^ n7646 ;
  assign n7718 = n7717 ^ n7716 ;
  assign n7643 = n7459 ^ n7402 ;
  assign n7644 = n7407 & n7643 ;
  assign n7645 = n7644 ^ n7402 ;
  assign n7719 = n7718 ^ n7645 ;
  assign n7720 = n7719 ^ x38 ;
  assign n7642 = x81 & n3916 ;
  assign n7721 = n7720 ^ n7642 ;
  assign n7641 = x83 & n3919 ;
  assign n7722 = n7721 ^ n7641 ;
  assign n7640 = n1512 & n3920 ;
  assign n7723 = n7722 ^ n7640 ;
  assign n7725 = n7724 ^ n7723 ;
  assign n7637 = n7460 ^ n7391 ;
  assign n7638 = n7466 & n7637 ;
  assign n7639 = n7638 ^ n7460 ;
  assign n7726 = n7725 ^ n7639 ;
  assign n7727 = n7726 ^ x35 ;
  assign n7636 = x84 & n3375 ;
  assign n7728 = n7727 ^ n7636 ;
  assign n7635 = x86 & n3378 ;
  assign n7729 = n7728 ^ n7635 ;
  assign n7634 = n1857 & n3379 ;
  assign n7730 = n7729 ^ n7634 ;
  assign n7732 = n7731 ^ n7730 ;
  assign n7736 = n7735 ^ n7732 ;
  assign n7737 = n7736 ^ x32 ;
  assign n7633 = x87 & n2879 ;
  assign n7738 = n7737 ^ n7633 ;
  assign n7632 = x89 & n2882 ;
  assign n7739 = n7738 ^ n7632 ;
  assign n7631 = n2249 & n2883 ;
  assign n7740 = n7739 ^ n7631 ;
  assign n7742 = n7741 ^ n7740 ;
  assign n7628 = n7483 ^ n7474 ;
  assign n7629 = ~n7480 & n7628 ;
  assign n7630 = n7629 ^ n7483 ;
  assign n7743 = n7742 ^ n7630 ;
  assign n7744 = n7743 ^ x29 ;
  assign n7627 = x90 & n2581 ;
  assign n7745 = n7744 ^ n7627 ;
  assign n7626 = x92 & n2422 ;
  assign n7746 = n7745 ^ n7626 ;
  assign n7625 = n2423 & n2684 ;
  assign n7747 = n7746 ^ n7625 ;
  assign n7749 = n7748 ^ n7747 ;
  assign n7753 = n7752 ^ n7749 ;
  assign n7754 = n7753 ^ x26 ;
  assign n7624 = x93 & n2018 ;
  assign n7755 = n7754 ^ n7624 ;
  assign n7623 = x95 & n2021 ;
  assign n7756 = n7755 ^ n7623 ;
  assign n7622 = n2022 & n3159 ;
  assign n7757 = n7756 ^ n7622 ;
  assign n7759 = n7758 ^ n7757 ;
  assign n7763 = n7762 ^ n7759 ;
  assign n7764 = n7763 ^ x23 ;
  assign n7621 = x96 & n1658 ;
  assign n7765 = n7764 ^ n7621 ;
  assign n7620 = x98 & n1661 ;
  assign n7766 = n7765 ^ n7620 ;
  assign n7619 = n1662 & n3660 ;
  assign n7767 = n7766 ^ n7619 ;
  assign n7769 = n7768 ^ n7767 ;
  assign n7773 = n7772 ^ n7769 ;
  assign n7774 = n7773 ^ x20 ;
  assign n7618 = x99 & n1327 ;
  assign n7775 = n7774 ^ n7618 ;
  assign n7617 = x101 & n1330 ;
  assign n7776 = n7775 ^ n7617 ;
  assign n7616 = n1331 & n4215 ;
  assign n7777 = n7776 ^ n7616 ;
  assign n7779 = n7778 ^ n7777 ;
  assign n7613 = n7514 ^ n7505 ;
  assign n7614 = n7511 & ~n7613 ;
  assign n7615 = n7614 ^ n7514 ;
  assign n7780 = n7779 ^ n7615 ;
  assign n7781 = n7780 ^ x17 ;
  assign n7612 = x102 & n1050 ;
  assign n7782 = n7781 ^ n7612 ;
  assign n7611 = x104 & n1053 ;
  assign n7783 = n7782 ^ n7611 ;
  assign n7610 = n1054 & ~n4814 ;
  assign n7784 = n7783 ^ n7610 ;
  assign n7786 = n7785 ^ n7784 ;
  assign n7790 = n7789 ^ n7786 ;
  assign n7791 = n7790 ^ x14 ;
  assign n7609 = x105 & n877 ;
  assign n7792 = n7791 ^ n7609 ;
  assign n7608 = x107 & n782 ;
  assign n7793 = n7792 ^ n7608 ;
  assign n7607 = n783 & ~n5448 ;
  assign n7794 = n7793 ^ n7607 ;
  assign n7796 = n7795 ^ n7794 ;
  assign n7604 = n7531 ^ n7522 ;
  assign n7605 = ~n7528 & ~n7604 ;
  assign n7606 = n7605 ^ n7531 ;
  assign n7797 = n7796 ^ n7606 ;
  assign n7798 = n7797 ^ x11 ;
  assign n7603 = x108 & n647 ;
  assign n7799 = n7798 ^ n7603 ;
  assign n7602 = x110 & ~n572 ;
  assign n7800 = n7799 ^ n7602 ;
  assign n7601 = ~n573 & n6129 ;
  assign n7801 = n7800 ^ n7601 ;
  assign n7803 = n7802 ^ n7801 ;
  assign n7598 = n7544 ^ n7540 ;
  assign n7599 = n7541 & n7598 ;
  assign n7600 = n7599 ^ n7544 ;
  assign n7804 = n7803 ^ n7600 ;
  assign n7805 = n7804 ^ x8 ;
  assign n7597 = x111 & n446 ;
  assign n7806 = n7805 ^ n7597 ;
  assign n7596 = x113 & n383 ;
  assign n7807 = n7806 ^ n7596 ;
  assign n7595 = n384 & ~n6839 ;
  assign n7808 = n7807 ^ n7595 ;
  assign n7810 = n7809 ^ n7808 ;
  assign n7592 = n7554 ^ n7545 ;
  assign n7593 = n7551 & ~n7592 ;
  assign n7594 = n7593 ^ n7554 ;
  assign n7811 = n7810 ^ n7594 ;
  assign n7812 = n7811 ^ x5 ;
  assign n7591 = x114 & n234 ;
  assign n7813 = n7812 ^ n7591 ;
  assign n7590 = x116 & n230 ;
  assign n7814 = n7813 ^ n7590 ;
  assign n7588 = n6822 ^ x116 ;
  assign n7589 = n231 & ~n7588 ;
  assign n7815 = n7814 ^ n7589 ;
  assign n7817 = n7816 ^ n7815 ;
  assign n7821 = n7820 ^ n7817 ;
  assign n7572 = x118 ^ x117 ;
  assign n7574 = n7326 & n7572 ;
  assign n7576 = x119 ^ x1 ;
  assign n7575 = x119 ^ x2 ;
  assign n7577 = n7576 ^ n7575 ;
  assign n7578 = ~n7574 & n7577 ;
  assign n7579 = n7578 ^ n7576 ;
  assign n7822 = n7821 ^ n7579 ;
  assign n7583 = x2 & x117 ;
  assign n7584 = n7583 ^ x118 ;
  assign n7585 = ~x1 & n7584 ;
  assign n7580 = n7579 ^ n7327 ;
  assign n7586 = n7585 ^ n7580 ;
  assign n7587 = ~x0 & n7586 ;
  assign n7823 = n7822 ^ n7587 ;
  assign n7569 = n7567 ^ n7562 ;
  assign n7570 = n7564 & ~n7569 ;
  assign n7571 = n7570 ^ n7567 ;
  assign n7824 = n7823 ^ n7571 ;
  assign n8093 = n7821 ^ n7571 ;
  assign n8094 = n7823 & n8093 ;
  assign n8095 = n8094 ^ n7821 ;
  assign n8088 = x116 & n227 ;
  assign n8080 = n7804 ^ n7594 ;
  assign n8081 = ~n7810 & ~n8080 ;
  assign n8082 = n8081 ^ n7804 ;
  assign n8078 = x113 & n390 ;
  assign n8070 = n7797 ^ n7600 ;
  assign n8071 = ~n7803 & ~n8070 ;
  assign n8072 = n8071 ^ n7797 ;
  assign n8068 = x110 & n578 ;
  assign n8060 = n7790 ^ n7606 ;
  assign n8061 = n7796 & ~n8060 ;
  assign n8062 = n8061 ^ n7790 ;
  assign n8058 = x107 & n788 ;
  assign n8051 = x104 & n1058 ;
  assign n8043 = n7773 ^ n7615 ;
  assign n8044 = ~n7779 & ~n8043 ;
  assign n8045 = n8044 ^ n7773 ;
  assign n8041 = x101 & n1335 ;
  assign n8034 = x98 & n1666 ;
  assign n8027 = x95 & n2014 ;
  assign n8020 = x92 & n2429 ;
  assign n8012 = n7736 ^ n7630 ;
  assign n8013 = n7742 & n8012 ;
  assign n8014 = n8013 ^ n7736 ;
  assign n8010 = x89 & n2887 ;
  assign n8003 = x86 & n3383 ;
  assign n7995 = n7719 ^ n7639 ;
  assign n7996 = n7725 & n7995 ;
  assign n7997 = n7996 ^ n7719 ;
  assign n7993 = x83 & n3924 ;
  assign n7984 = x77 & n5102 ;
  assign n7977 = x74 & n5736 ;
  assign n7969 = n7694 ^ n7667 ;
  assign n7970 = n7700 & n7969 ;
  assign n7971 = n7970 ^ n7694 ;
  assign n7967 = x71 & n6433 ;
  assign n7956 = x67 & n7171 ;
  assign n7955 = x69 & n7174 ;
  assign n7957 = n7956 ^ n7955 ;
  assign n7958 = n7957 ^ x53 ;
  assign n7954 = ~n375 & n7175 ;
  assign n7959 = n7958 ^ n7954 ;
  assign n7953 = x68 & n7179 ;
  assign n7960 = n7959 ^ n7953 ;
  assign n7949 = x56 & ~n7425 ;
  assign n7950 = ~n7681 & n7949 ;
  assign n7951 = n7950 ^ x56 ;
  assign n7946 = x66 & n7424 ;
  assign n7933 = x56 ^ x55 ;
  assign n7938 = n7424 & ~n7933 ;
  assign n7939 = n7938 ^ n7424 ;
  assign n7942 = x65 & n7939 ;
  assign n7673 = x55 ^ x54 ;
  assign n7934 = ~n7424 & ~n7673 ;
  assign n7935 = n7933 & n7934 ;
  assign n7943 = n7942 ^ n7935 ;
  assign n7944 = ~x64 & n7943 ;
  assign n7945 = n7944 ^ n7935 ;
  assign n7947 = n7946 ^ n7945 ;
  assign n7931 = ~n7424 & n7673 ;
  assign n7932 = x65 & n7931 ;
  assign n7948 = n7947 ^ n7932 ;
  assign n7952 = n7951 ^ n7948 ;
  assign n7961 = n7960 ^ n7952 ;
  assign n7928 = n7693 ^ n7689 ;
  assign n7929 = ~n7690 & n7928 ;
  assign n7930 = n7929 ^ n7693 ;
  assign n7962 = n7961 ^ n7930 ;
  assign n7963 = n7962 ^ x50 ;
  assign n7927 = x70 & n6677 ;
  assign n7964 = n7963 ^ n7927 ;
  assign n7926 = x72 & n6428 ;
  assign n7965 = n7964 ^ n7926 ;
  assign n7925 = n556 & n6429 ;
  assign n7966 = n7965 ^ n7925 ;
  assign n7968 = n7967 ^ n7966 ;
  assign n7972 = n7971 ^ n7968 ;
  assign n7973 = n7972 ^ x47 ;
  assign n7924 = x73 & n5965 ;
  assign n7974 = n7973 ^ n7924 ;
  assign n7923 = x75 & n5729 ;
  assign n7975 = n7974 ^ n7923 ;
  assign n7922 = ~n774 & n5730 ;
  assign n7976 = n7975 ^ n7922 ;
  assign n7978 = n7977 ^ n7976 ;
  assign n7919 = n7710 ^ n7701 ;
  assign n7920 = ~n7707 & n7919 ;
  assign n7921 = n7920 ^ n7710 ;
  assign n7979 = n7978 ^ n7921 ;
  assign n7980 = n7979 ^ x44 ;
  assign n7918 = x76 & n5094 ;
  assign n7981 = n7980 ^ n7918 ;
  assign n7917 = x78 & n5097 ;
  assign n7982 = n7981 ^ n7917 ;
  assign n7916 = ~n1025 & n5098 ;
  assign n7983 = n7982 ^ n7916 ;
  assign n7985 = n7984 ^ n7983 ;
  assign n7911 = x79 & n4474 ;
  assign n7910 = x81 & n4471 ;
  assign n7912 = n7911 ^ n7910 ;
  assign n7913 = n7912 ^ x41 ;
  assign n7909 = n1305 & n4472 ;
  assign n7914 = n7913 ^ n7909 ;
  assign n7908 = x80 & n4467 ;
  assign n7915 = n7914 ^ n7908 ;
  assign n7986 = n7985 ^ n7915 ;
  assign n7905 = n7711 ^ n7656 ;
  assign n7906 = n7661 & n7905 ;
  assign n7907 = n7906 ^ n7656 ;
  assign n7987 = n7986 ^ n7907 ;
  assign n7902 = n7712 ^ n7645 ;
  assign n7903 = n7718 & n7902 ;
  assign n7904 = n7903 ^ n7712 ;
  assign n7988 = n7987 ^ n7904 ;
  assign n7989 = n7988 ^ x38 ;
  assign n7901 = x82 & n3916 ;
  assign n7990 = n7989 ^ n7901 ;
  assign n7900 = x84 & n3919 ;
  assign n7991 = n7990 ^ n7900 ;
  assign n7899 = n1624 & n3920 ;
  assign n7992 = n7991 ^ n7899 ;
  assign n7994 = n7993 ^ n7992 ;
  assign n7998 = n7997 ^ n7994 ;
  assign n7999 = n7998 ^ x35 ;
  assign n7898 = x85 & n3375 ;
  assign n8000 = n7999 ^ n7898 ;
  assign n7897 = x87 & n3378 ;
  assign n8001 = n8000 ^ n7897 ;
  assign n7896 = n1982 & n3379 ;
  assign n8002 = n8001 ^ n7896 ;
  assign n8004 = n8003 ^ n8002 ;
  assign n7893 = n7735 ^ n7726 ;
  assign n7894 = ~n7732 & n7893 ;
  assign n7895 = n7894 ^ n7735 ;
  assign n8005 = n8004 ^ n7895 ;
  assign n8006 = n8005 ^ x32 ;
  assign n7892 = x88 & n2879 ;
  assign n8007 = n8006 ^ n7892 ;
  assign n7891 = x90 & n2882 ;
  assign n8008 = n8007 ^ n7891 ;
  assign n7890 = n2386 & n2883 ;
  assign n8009 = n8008 ^ n7890 ;
  assign n8011 = n8010 ^ n8009 ;
  assign n8015 = n8014 ^ n8011 ;
  assign n8016 = n8015 ^ x29 ;
  assign n7889 = x91 & n2581 ;
  assign n8017 = n8016 ^ n7889 ;
  assign n7888 = x93 & n2422 ;
  assign n8018 = n8017 ^ n7888 ;
  assign n7887 = n2423 & n2836 ;
  assign n8019 = n8018 ^ n7887 ;
  assign n8021 = n8020 ^ n8019 ;
  assign n7884 = n7752 ^ n7743 ;
  assign n7885 = ~n7749 & n7884 ;
  assign n7886 = n7885 ^ n7752 ;
  assign n8022 = n8021 ^ n7886 ;
  assign n8023 = n8022 ^ x26 ;
  assign n7883 = x94 & n2018 ;
  assign n8024 = n8023 ^ n7883 ;
  assign n7882 = x96 & n2021 ;
  assign n8025 = n8024 ^ n7882 ;
  assign n7881 = n2022 & n3323 ;
  assign n8026 = n8025 ^ n7881 ;
  assign n8028 = n8027 ^ n8026 ;
  assign n7878 = n7762 ^ n7753 ;
  assign n7879 = ~n7759 & n7878 ;
  assign n7880 = n7879 ^ n7762 ;
  assign n8029 = n8028 ^ n7880 ;
  assign n8030 = n8029 ^ x23 ;
  assign n7877 = x97 & n1658 ;
  assign n8031 = n8030 ^ n7877 ;
  assign n7876 = x99 & n1661 ;
  assign n8032 = n8031 ^ n7876 ;
  assign n7875 = n1662 & n3843 ;
  assign n8033 = n8032 ^ n7875 ;
  assign n8035 = n8034 ^ n8033 ;
  assign n7872 = n7772 ^ n7763 ;
  assign n7873 = ~n7769 & ~n7872 ;
  assign n7874 = n7873 ^ n7772 ;
  assign n8036 = n8035 ^ n7874 ;
  assign n8037 = n8036 ^ x20 ;
  assign n7871 = x100 & n1327 ;
  assign n8038 = n8037 ^ n7871 ;
  assign n7870 = x102 & n1330 ;
  assign n8039 = n8038 ^ n7870 ;
  assign n7869 = n1331 & n4410 ;
  assign n8040 = n8039 ^ n7869 ;
  assign n8042 = n8041 ^ n8040 ;
  assign n8046 = n8045 ^ n8042 ;
  assign n8047 = n8046 ^ x17 ;
  assign n7868 = x103 & n1050 ;
  assign n8048 = n8047 ^ n7868 ;
  assign n7867 = x105 & n1053 ;
  assign n8049 = n8048 ^ n7867 ;
  assign n7866 = n1054 & ~n5023 ;
  assign n8050 = n8049 ^ n7866 ;
  assign n8052 = n8051 ^ n8050 ;
  assign n7863 = n7789 ^ n7780 ;
  assign n7864 = n7786 & n7863 ;
  assign n7865 = n7864 ^ n7789 ;
  assign n8053 = n8052 ^ n7865 ;
  assign n8054 = n8053 ^ x14 ;
  assign n7862 = x106 & n877 ;
  assign n8055 = n8054 ^ n7862 ;
  assign n7861 = x108 & n782 ;
  assign n8056 = n8055 ^ n7861 ;
  assign n7860 = n783 & n5670 ;
  assign n8057 = n8056 ^ n7860 ;
  assign n8059 = n8058 ^ n8057 ;
  assign n8063 = n8062 ^ n8059 ;
  assign n8064 = n8063 ^ x11 ;
  assign n7859 = x109 & n647 ;
  assign n8065 = n8064 ^ n7859 ;
  assign n7858 = x111 & ~n572 ;
  assign n8066 = n8065 ^ n7858 ;
  assign n7857 = ~n573 & ~n6360 ;
  assign n8067 = n8066 ^ n7857 ;
  assign n8069 = n8068 ^ n8067 ;
  assign n8073 = n8072 ^ n8069 ;
  assign n8074 = n8073 ^ x8 ;
  assign n7856 = x112 & n446 ;
  assign n8075 = n8074 ^ n7856 ;
  assign n7855 = x114 & n383 ;
  assign n8076 = n8075 ^ n7855 ;
  assign n7854 = n384 & ~n7092 ;
  assign n8077 = n8076 ^ n7854 ;
  assign n8079 = n8078 ^ n8077 ;
  assign n8083 = n8082 ^ n8079 ;
  assign n8084 = n8083 ^ x5 ;
  assign n7853 = x115 & n234 ;
  assign n8085 = n8084 ^ n7853 ;
  assign n7852 = x117 & n230 ;
  assign n8086 = n8085 ^ n7852 ;
  assign n7850 = n7078 ^ x117 ;
  assign n7851 = n231 & ~n7850 ;
  assign n8087 = n8086 ^ n7851 ;
  assign n8089 = n8088 ^ n8087 ;
  assign n7847 = n7820 ^ n7811 ;
  assign n7848 = n7817 & n7847 ;
  assign n7849 = n7848 ^ n7820 ;
  assign n8090 = n8089 ^ n7849 ;
  assign n7825 = x119 ^ x118 ;
  assign n7831 = ~x119 & n7326 ;
  assign n7832 = n7831 ^ n7324 ;
  assign n7833 = n7825 & ~n7832 ;
  assign n7835 = x120 ^ x1 ;
  assign n7834 = x120 ^ x2 ;
  assign n7836 = n7835 ^ n7834 ;
  assign n7837 = ~n7833 & n7836 ;
  assign n7838 = n7837 ^ n7835 ;
  assign n8091 = n8090 ^ n7838 ;
  assign n7842 = x2 & x118 ;
  assign n7843 = n7842 ^ x119 ;
  assign n7844 = ~x1 & n7843 ;
  assign n7839 = n7838 ^ n7575 ;
  assign n7845 = n7844 ^ n7839 ;
  assign n7846 = ~x0 & n7845 ;
  assign n8092 = n8091 ^ n7846 ;
  assign n8096 = n8095 ^ n8092 ;
  assign n8362 = n8083 ^ n7849 ;
  assign n8363 = ~n8089 & n8362 ;
  assign n8364 = n8363 ^ n8083 ;
  assign n8360 = x117 & n227 ;
  assign n8353 = x114 & n390 ;
  assign n8346 = x111 & n578 ;
  assign n8339 = x108 & n788 ;
  assign n8331 = n8046 ^ n7865 ;
  assign n8332 = n8052 & ~n8331 ;
  assign n8333 = n8332 ^ n8046 ;
  assign n8329 = x105 & n1058 ;
  assign n8322 = x102 & n1335 ;
  assign n8314 = n8029 ^ n7874 ;
  assign n8315 = n8035 & ~n8314 ;
  assign n8316 = n8315 ^ n8029 ;
  assign n8312 = x99 & n1666 ;
  assign n8304 = n8022 ^ n7880 ;
  assign n8305 = n8028 & n8304 ;
  assign n8306 = n8305 ^ n8022 ;
  assign n8302 = x96 & n2014 ;
  assign n8294 = n8015 ^ n7886 ;
  assign n8295 = n8021 & n8294 ;
  assign n8296 = n8295 ^ n8015 ;
  assign n8292 = x93 & n2429 ;
  assign n8285 = x90 & n2887 ;
  assign n8277 = n7998 ^ n7895 ;
  assign n8278 = n8004 & n8277 ;
  assign n8279 = n8278 ^ n7998 ;
  assign n8275 = x87 & n3383 ;
  assign n8268 = x84 & n3924 ;
  assign n8260 = n7915 ^ n7904 ;
  assign n8261 = n7987 & n8260 ;
  assign n8262 = n8261 ^ n7915 ;
  assign n8258 = x81 & n4467 ;
  assign n8249 = n7972 ^ n7921 ;
  assign n8250 = n7978 & n8249 ;
  assign n8251 = n8250 ^ n7972 ;
  assign n8247 = x75 & n5736 ;
  assign n8234 = x65 & n7935 ;
  assign n8233 = x66 & n7931 ;
  assign n8235 = n8234 ^ n8233 ;
  assign n8236 = n8235 ^ x56 ;
  assign n8230 = ~n153 & ~n7933 ;
  assign n8231 = n8230 ^ n291 ;
  assign n8232 = n7424 & ~n8231 ;
  assign n8237 = n8236 ^ n8232 ;
  assign n8223 = x57 ^ x56 ;
  assign n8224 = x64 & n8223 ;
  assign n8238 = n8237 ^ n8224 ;
  assign n8225 = ~n7948 & n7950 ;
  assign n8226 = ~n8224 & ~n8225 ;
  assign n8227 = n8226 ^ n8225 ;
  assign n8239 = n8238 ^ n8227 ;
  assign n8240 = n8239 ^ n8226 ;
  assign n8220 = n7960 ^ n7930 ;
  assign n8221 = n7961 & n8220 ;
  assign n8213 = x68 & n7171 ;
  assign n8212 = x70 & n7174 ;
  assign n8214 = n8213 ^ n8212 ;
  assign n8215 = n8214 ^ x53 ;
  assign n8211 = ~n436 & n7175 ;
  assign n8216 = n8215 ^ n8211 ;
  assign n8210 = x69 & n7179 ;
  assign n8217 = n8216 ^ n8210 ;
  assign n8218 = n8217 ^ n7960 ;
  assign n8222 = n8221 ^ n8218 ;
  assign n8241 = n8240 ^ n8222 ;
  assign n8200 = x71 & n6677 ;
  assign n8199 = x73 & n6428 ;
  assign n8201 = n8200 ^ n8199 ;
  assign n8202 = n8201 ^ x50 ;
  assign n8198 = n633 & n6429 ;
  assign n8203 = n8202 ^ n8198 ;
  assign n8197 = x72 & n6433 ;
  assign n8204 = n8203 ^ n8197 ;
  assign n8205 = n8204 ^ n7971 ;
  assign n8206 = n8205 ^ n7962 ;
  assign n8207 = n8206 ^ n8204 ;
  assign n8208 = ~n7968 & n8207 ;
  assign n8209 = n8208 ^ n8205 ;
  assign n8242 = n8241 ^ n8209 ;
  assign n8243 = n8242 ^ x47 ;
  assign n8196 = x74 & n5965 ;
  assign n8244 = n8243 ^ n8196 ;
  assign n8195 = x76 & n5729 ;
  assign n8245 = n8244 ^ n8195 ;
  assign n8194 = ~n853 & n5730 ;
  assign n8246 = n8245 ^ n8194 ;
  assign n8248 = n8247 ^ n8246 ;
  assign n8252 = n8251 ^ n8248 ;
  assign n8184 = x77 & n5094 ;
  assign n8183 = x79 & n5097 ;
  assign n8185 = n8184 ^ n8183 ;
  assign n8186 = n8185 ^ x44 ;
  assign n8182 = n1118 & n5098 ;
  assign n8187 = n8186 ^ n8182 ;
  assign n8181 = x78 & n5102 ;
  assign n8188 = n8187 ^ n8181 ;
  assign n8189 = n8188 ^ n7979 ;
  assign n8190 = n8189 ^ n7907 ;
  assign n8191 = n8190 ^ n8188 ;
  assign n8192 = n7985 & n8191 ;
  assign n8193 = n8192 ^ n8189 ;
  assign n8253 = n8252 ^ n8193 ;
  assign n8254 = n8253 ^ x41 ;
  assign n8180 = x80 & n4474 ;
  assign n8255 = n8254 ^ n8180 ;
  assign n8179 = x82 & n4471 ;
  assign n8256 = n8255 ^ n8179 ;
  assign n8178 = n1411 & n4472 ;
  assign n8257 = n8256 ^ n8178 ;
  assign n8259 = n8258 ^ n8257 ;
  assign n8263 = n8262 ^ n8259 ;
  assign n8264 = n8263 ^ x38 ;
  assign n8177 = x83 & n3916 ;
  assign n8265 = n8264 ^ n8177 ;
  assign n8176 = x85 & n3919 ;
  assign n8266 = n8265 ^ n8176 ;
  assign n8175 = n1743 & n3920 ;
  assign n8267 = n8266 ^ n8175 ;
  assign n8269 = n8268 ^ n8267 ;
  assign n8172 = n7997 ^ n7988 ;
  assign n8173 = ~n7994 & n8172 ;
  assign n8174 = n8173 ^ n7997 ;
  assign n8270 = n8269 ^ n8174 ;
  assign n8271 = n8270 ^ x35 ;
  assign n8171 = x86 & n3375 ;
  assign n8272 = n8271 ^ n8171 ;
  assign n8170 = x88 & n3378 ;
  assign n8273 = n8272 ^ n8170 ;
  assign n8169 = n2119 & n3379 ;
  assign n8274 = n8273 ^ n8169 ;
  assign n8276 = n8275 ^ n8274 ;
  assign n8280 = n8279 ^ n8276 ;
  assign n8281 = n8280 ^ x32 ;
  assign n8168 = x89 & n2879 ;
  assign n8282 = n8281 ^ n8168 ;
  assign n8167 = x91 & n2882 ;
  assign n8283 = n8282 ^ n8167 ;
  assign n8166 = n2542 & n2883 ;
  assign n8284 = n8283 ^ n8166 ;
  assign n8286 = n8285 ^ n8284 ;
  assign n8163 = n8014 ^ n8005 ;
  assign n8164 = ~n8011 & n8163 ;
  assign n8165 = n8164 ^ n8014 ;
  assign n8287 = n8286 ^ n8165 ;
  assign n8288 = n8287 ^ x29 ;
  assign n8162 = x92 & n2581 ;
  assign n8289 = n8288 ^ n8162 ;
  assign n8161 = x94 & n2422 ;
  assign n8290 = n8289 ^ n8161 ;
  assign n8160 = n2423 & n2997 ;
  assign n8291 = n8290 ^ n8160 ;
  assign n8293 = n8292 ^ n8291 ;
  assign n8297 = n8296 ^ n8293 ;
  assign n8298 = n8297 ^ x26 ;
  assign n8159 = x95 & n2018 ;
  assign n8299 = n8298 ^ n8159 ;
  assign n8158 = x97 & n2021 ;
  assign n8300 = n8299 ^ n8158 ;
  assign n8157 = n2022 & n3494 ;
  assign n8301 = n8300 ^ n8157 ;
  assign n8303 = n8302 ^ n8301 ;
  assign n8307 = n8306 ^ n8303 ;
  assign n8308 = n8307 ^ x23 ;
  assign n8156 = x98 & n1658 ;
  assign n8309 = n8308 ^ n8156 ;
  assign n8155 = x100 & n1661 ;
  assign n8310 = n8309 ^ n8155 ;
  assign n8154 = n1662 & n4034 ;
  assign n8311 = n8310 ^ n8154 ;
  assign n8313 = n8312 ^ n8311 ;
  assign n8317 = n8316 ^ n8313 ;
  assign n8318 = n8317 ^ x20 ;
  assign n8153 = x101 & n1327 ;
  assign n8319 = n8318 ^ n8153 ;
  assign n8152 = x103 & n1330 ;
  assign n8320 = n8319 ^ n8152 ;
  assign n8151 = n1331 & ~n4615 ;
  assign n8321 = n8320 ^ n8151 ;
  assign n8323 = n8322 ^ n8321 ;
  assign n8148 = n8045 ^ n8036 ;
  assign n8149 = n8042 & n8148 ;
  assign n8150 = n8149 ^ n8045 ;
  assign n8324 = n8323 ^ n8150 ;
  assign n8325 = n8324 ^ x17 ;
  assign n8147 = x104 & n1050 ;
  assign n8326 = n8325 ^ n8147 ;
  assign n8146 = x106 & n1053 ;
  assign n8327 = n8326 ^ n8146 ;
  assign n8145 = n1054 & ~n5240 ;
  assign n8328 = n8327 ^ n8145 ;
  assign n8330 = n8329 ^ n8328 ;
  assign n8334 = n8333 ^ n8330 ;
  assign n8335 = n8334 ^ x14 ;
  assign n8144 = x107 & n877 ;
  assign n8336 = n8335 ^ n8144 ;
  assign n8143 = x109 & n782 ;
  assign n8337 = n8336 ^ n8143 ;
  assign n8142 = n783 & n5902 ;
  assign n8338 = n8337 ^ n8142 ;
  assign n8340 = n8339 ^ n8338 ;
  assign n8139 = n8062 ^ n8053 ;
  assign n8140 = n8059 & ~n8139 ;
  assign n8141 = n8140 ^ n8062 ;
  assign n8341 = n8340 ^ n8141 ;
  assign n8342 = n8341 ^ x11 ;
  assign n8138 = x110 & n647 ;
  assign n8343 = n8342 ^ n8138 ;
  assign n8137 = x112 & ~n572 ;
  assign n8344 = n8343 ^ n8137 ;
  assign n8136 = ~n573 & ~n6600 ;
  assign n8345 = n8344 ^ n8136 ;
  assign n8347 = n8346 ^ n8345 ;
  assign n8133 = n8072 ^ n8063 ;
  assign n8134 = n8069 & n8133 ;
  assign n8135 = n8134 ^ n8072 ;
  assign n8348 = n8347 ^ n8135 ;
  assign n8349 = n8348 ^ x8 ;
  assign n8132 = x113 & n446 ;
  assign n8350 = n8349 ^ n8132 ;
  assign n8131 = x115 & n383 ;
  assign n8351 = n8350 ^ n8131 ;
  assign n8130 = n384 & ~n7343 ;
  assign n8352 = n8351 ^ n8130 ;
  assign n8354 = n8353 ^ n8352 ;
  assign n8127 = n8082 ^ n8073 ;
  assign n8128 = ~n8079 & ~n8127 ;
  assign n8129 = n8128 ^ n8082 ;
  assign n8355 = n8354 ^ n8129 ;
  assign n8356 = n8355 ^ x5 ;
  assign n8126 = x116 & n234 ;
  assign n8357 = n8356 ^ n8126 ;
  assign n8125 = x118 & n230 ;
  assign n8358 = n8357 ^ n8125 ;
  assign n8122 = n7326 ^ x117 ;
  assign n8123 = n8122 ^ n7572 ;
  assign n8124 = n231 & ~n8123 ;
  assign n8359 = n8358 ^ n8124 ;
  assign n8361 = n8360 ^ n8359 ;
  assign n8365 = n8364 ^ n8361 ;
  assign n8102 = x120 ^ x117 ;
  assign n8100 = x120 ^ x119 ;
  assign n8103 = n7825 & n8100 ;
  assign n8104 = n7326 & n8103 ;
  assign n8105 = n8102 & n8104 ;
  assign n8106 = n8105 ^ n8103 ;
  assign n8107 = n8106 ^ x119 ;
  assign n8108 = n8107 ^ x120 ;
  assign n8110 = x121 ^ x1 ;
  assign n8109 = x121 ^ x2 ;
  assign n8111 = n8110 ^ n8109 ;
  assign n8112 = ~n8108 & n8111 ;
  assign n8113 = n8112 ^ n8110 ;
  assign n8366 = n8365 ^ n8113 ;
  assign n8117 = x2 & x119 ;
  assign n8118 = n8117 ^ x120 ;
  assign n8119 = ~x1 & n8118 ;
  assign n8114 = n8113 ^ n7834 ;
  assign n8120 = n8119 ^ n8114 ;
  assign n8121 = ~x0 & n8120 ;
  assign n8367 = n8366 ^ n8121 ;
  assign n8097 = n8095 ^ n8090 ;
  assign n8098 = ~n8092 & n8097 ;
  assign n8099 = n8098 ^ n8095 ;
  assign n8368 = n8367 ^ n8099 ;
  assign n8635 = n8365 ^ n8099 ;
  assign n8636 = n8367 & n8635 ;
  assign n8637 = n8636 ^ n8365 ;
  assign n8629 = n8348 ^ n8129 ;
  assign n8630 = n8354 & ~n8629 ;
  assign n8631 = n8630 ^ n8348 ;
  assign n8627 = x115 & n390 ;
  assign n8619 = n8341 ^ n8135 ;
  assign n8620 = ~n8347 & n8619 ;
  assign n8621 = n8620 ^ n8341 ;
  assign n8617 = x112 & n578 ;
  assign n8609 = n8334 ^ n8141 ;
  assign n8610 = ~n8340 & ~n8609 ;
  assign n8611 = n8610 ^ n8334 ;
  assign n8607 = x109 & n788 ;
  assign n8600 = x106 & n1058 ;
  assign n8592 = n8317 ^ n8150 ;
  assign n8593 = n8323 & ~n8592 ;
  assign n8594 = n8593 ^ n8317 ;
  assign n8590 = x103 & n1335 ;
  assign n8583 = x100 & n1666 ;
  assign n8576 = x97 & n2014 ;
  assign n8565 = x93 & n2581 ;
  assign n8564 = x95 & n2422 ;
  assign n8566 = n8565 ^ n8564 ;
  assign n8567 = n8566 ^ x29 ;
  assign n8563 = n2423 & n3159 ;
  assign n8568 = n8567 ^ n8563 ;
  assign n8562 = x94 & n2429 ;
  assign n8569 = n8568 ^ n8562 ;
  assign n8558 = n8280 ^ n8165 ;
  assign n8559 = n8286 & n8558 ;
  assign n8560 = n8559 ^ n8280 ;
  assign n8556 = x91 & n2887 ;
  assign n8549 = x88 & n3383 ;
  assign n8541 = n8263 ^ n8174 ;
  assign n8542 = n8269 & n8541 ;
  assign n8543 = n8542 ^ n8263 ;
  assign n8539 = x85 & n3924 ;
  assign n8532 = x82 & n4467 ;
  assign n8525 = x79 & n5102 ;
  assign n8518 = x76 & n5736 ;
  assign n8511 = x73 & n6433 ;
  assign n8504 = x70 & n7179 ;
  assign n8494 = x66 & n7935 ;
  assign n8493 = x68 & n7938 ;
  assign n8495 = n8494 ^ n8493 ;
  assign n8496 = n8495 ^ x56 ;
  assign n8492 = ~n340 & n7939 ;
  assign n8497 = n8496 ^ n8492 ;
  assign n8491 = x67 & n7931 ;
  assign n8498 = n8497 ^ n8491 ;
  assign n8489 = ~n8226 & n8237 ;
  assign n8486 = x65 ^ x57 ;
  assign n8487 = n8223 & ~n8486 ;
  assign n8482 = x56 & x57 ;
  assign n8483 = n8482 ^ x58 ;
  assign n8484 = ~x64 & n8483 ;
  assign n8478 = x58 ^ x56 ;
  assign n8485 = n8484 ^ n8478 ;
  assign n8488 = n8487 ^ n8485 ;
  assign n8490 = n8489 ^ n8488 ;
  assign n8499 = n8498 ^ n8490 ;
  assign n8500 = n8499 ^ x53 ;
  assign n8477 = x69 & n7171 ;
  assign n8501 = n8500 ^ n8477 ;
  assign n8476 = x71 & n7174 ;
  assign n8502 = n8501 ^ n8476 ;
  assign n8475 = ~n493 & n7175 ;
  assign n8503 = n8502 ^ n8475 ;
  assign n8505 = n8504 ^ n8503 ;
  assign n8472 = n8240 ^ n8217 ;
  assign n8473 = n8222 & n8472 ;
  assign n8474 = n8473 ^ n8217 ;
  assign n8506 = n8505 ^ n8474 ;
  assign n8507 = n8506 ^ x50 ;
  assign n8471 = x72 & n6677 ;
  assign n8508 = n8507 ^ n8471 ;
  assign n8470 = x74 & n6428 ;
  assign n8509 = n8508 ^ n8470 ;
  assign n8469 = n699 & n6429 ;
  assign n8510 = n8509 ^ n8469 ;
  assign n8512 = n8511 ^ n8510 ;
  assign n8466 = n8241 ^ n8204 ;
  assign n8467 = n8209 & n8466 ;
  assign n8468 = n8467 ^ n8204 ;
  assign n8513 = n8512 ^ n8468 ;
  assign n8514 = n8513 ^ x47 ;
  assign n8465 = x75 & n5965 ;
  assign n8515 = n8514 ^ n8465 ;
  assign n8464 = x77 & n5729 ;
  assign n8516 = n8515 ^ n8464 ;
  assign n8463 = ~n939 & n5730 ;
  assign n8517 = n8516 ^ n8463 ;
  assign n8519 = n8518 ^ n8517 ;
  assign n8460 = n8251 ^ n8242 ;
  assign n8461 = ~n8248 & n8460 ;
  assign n8462 = n8461 ^ n8251 ;
  assign n8520 = n8519 ^ n8462 ;
  assign n8521 = n8520 ^ x44 ;
  assign n8459 = x78 & n5094 ;
  assign n8522 = n8521 ^ n8459 ;
  assign n8458 = x80 & n5097 ;
  assign n8523 = n8522 ^ n8458 ;
  assign n8457 = n1206 & n5098 ;
  assign n8524 = n8523 ^ n8457 ;
  assign n8526 = n8525 ^ n8524 ;
  assign n8454 = n8252 ^ n8188 ;
  assign n8455 = n8193 & n8454 ;
  assign n8456 = n8455 ^ n8188 ;
  assign n8527 = n8526 ^ n8456 ;
  assign n8528 = n8527 ^ x41 ;
  assign n8453 = x81 & n4474 ;
  assign n8529 = n8528 ^ n8453 ;
  assign n8452 = x83 & n4471 ;
  assign n8530 = n8529 ^ n8452 ;
  assign n8451 = n1512 & n4472 ;
  assign n8531 = n8530 ^ n8451 ;
  assign n8533 = n8532 ^ n8531 ;
  assign n8448 = n8262 ^ n8253 ;
  assign n8449 = ~n8259 & n8448 ;
  assign n8450 = n8449 ^ n8262 ;
  assign n8534 = n8533 ^ n8450 ;
  assign n8535 = n8534 ^ x38 ;
  assign n8447 = x84 & n3916 ;
  assign n8536 = n8535 ^ n8447 ;
  assign n8446 = x86 & n3919 ;
  assign n8537 = n8536 ^ n8446 ;
  assign n8445 = n1857 & n3920 ;
  assign n8538 = n8537 ^ n8445 ;
  assign n8540 = n8539 ^ n8538 ;
  assign n8544 = n8543 ^ n8540 ;
  assign n8545 = n8544 ^ x35 ;
  assign n8444 = x87 & n3375 ;
  assign n8546 = n8545 ^ n8444 ;
  assign n8443 = x89 & n3378 ;
  assign n8547 = n8546 ^ n8443 ;
  assign n8442 = n2249 & n3379 ;
  assign n8548 = n8547 ^ n8442 ;
  assign n8550 = n8549 ^ n8548 ;
  assign n8439 = n8279 ^ n8270 ;
  assign n8440 = ~n8276 & n8439 ;
  assign n8441 = n8440 ^ n8279 ;
  assign n8551 = n8550 ^ n8441 ;
  assign n8552 = n8551 ^ x32 ;
  assign n8438 = x90 & n2879 ;
  assign n8553 = n8552 ^ n8438 ;
  assign n8437 = x92 & n2882 ;
  assign n8554 = n8553 ^ n8437 ;
  assign n8436 = n2684 & n2883 ;
  assign n8555 = n8554 ^ n8436 ;
  assign n8557 = n8556 ^ n8555 ;
  assign n8561 = n8560 ^ n8557 ;
  assign n8570 = n8569 ^ n8561 ;
  assign n8433 = n8296 ^ n8287 ;
  assign n8434 = ~n8293 & n8433 ;
  assign n8435 = n8434 ^ n8296 ;
  assign n8571 = n8570 ^ n8435 ;
  assign n8572 = n8571 ^ x26 ;
  assign n8432 = x96 & n2018 ;
  assign n8573 = n8572 ^ n8432 ;
  assign n8431 = x98 & n2021 ;
  assign n8574 = n8573 ^ n8431 ;
  assign n8430 = n2022 & n3660 ;
  assign n8575 = n8574 ^ n8430 ;
  assign n8577 = n8576 ^ n8575 ;
  assign n8427 = n8306 ^ n8297 ;
  assign n8428 = ~n8303 & n8427 ;
  assign n8429 = n8428 ^ n8306 ;
  assign n8578 = n8577 ^ n8429 ;
  assign n8579 = n8578 ^ x23 ;
  assign n8426 = x99 & n1658 ;
  assign n8580 = n8579 ^ n8426 ;
  assign n8425 = x101 & n1661 ;
  assign n8581 = n8580 ^ n8425 ;
  assign n8424 = n1662 & n4215 ;
  assign n8582 = n8581 ^ n8424 ;
  assign n8584 = n8583 ^ n8582 ;
  assign n8421 = n8316 ^ n8307 ;
  assign n8422 = ~n8313 & n8421 ;
  assign n8423 = n8422 ^ n8316 ;
  assign n8585 = n8584 ^ n8423 ;
  assign n8586 = n8585 ^ x20 ;
  assign n8420 = x102 & n1327 ;
  assign n8587 = n8586 ^ n8420 ;
  assign n8419 = x104 & n1330 ;
  assign n8588 = n8587 ^ n8419 ;
  assign n8418 = n1331 & ~n4814 ;
  assign n8589 = n8588 ^ n8418 ;
  assign n8591 = n8590 ^ n8589 ;
  assign n8595 = n8594 ^ n8591 ;
  assign n8596 = n8595 ^ x17 ;
  assign n8417 = x105 & n1050 ;
  assign n8597 = n8596 ^ n8417 ;
  assign n8416 = x107 & n1053 ;
  assign n8598 = n8597 ^ n8416 ;
  assign n8415 = n1054 & ~n5448 ;
  assign n8599 = n8598 ^ n8415 ;
  assign n8601 = n8600 ^ n8599 ;
  assign n8412 = n8333 ^ n8324 ;
  assign n8413 = n8330 & ~n8412 ;
  assign n8414 = n8413 ^ n8333 ;
  assign n8602 = n8601 ^ n8414 ;
  assign n8603 = n8602 ^ x14 ;
  assign n8411 = x108 & n877 ;
  assign n8604 = n8603 ^ n8411 ;
  assign n8410 = x110 & n782 ;
  assign n8605 = n8604 ^ n8410 ;
  assign n8409 = n783 & n6129 ;
  assign n8606 = n8605 ^ n8409 ;
  assign n8608 = n8607 ^ n8606 ;
  assign n8612 = n8611 ^ n8608 ;
  assign n8613 = n8612 ^ x11 ;
  assign n8408 = x111 & n647 ;
  assign n8614 = n8613 ^ n8408 ;
  assign n8407 = x113 & ~n572 ;
  assign n8615 = n8614 ^ n8407 ;
  assign n8406 = ~n573 & ~n6839 ;
  assign n8616 = n8615 ^ n8406 ;
  assign n8618 = n8617 ^ n8616 ;
  assign n8622 = n8621 ^ n8618 ;
  assign n8623 = n8622 ^ x8 ;
  assign n8405 = x114 & n446 ;
  assign n8624 = n8623 ^ n8405 ;
  assign n8404 = x116 & n383 ;
  assign n8625 = n8624 ^ n8404 ;
  assign n8403 = n384 & ~n7588 ;
  assign n8626 = n8625 ^ n8403 ;
  assign n8628 = n8627 ^ n8626 ;
  assign n8632 = n8631 ^ n8628 ;
  assign n8397 = x117 & n234 ;
  assign n8396 = x119 & n230 ;
  assign n8398 = n8397 ^ n8396 ;
  assign n8399 = n8398 ^ x5 ;
  assign n8394 = n7574 ^ x119 ;
  assign n8395 = n231 & n8394 ;
  assign n8400 = n8399 ^ n8395 ;
  assign n8393 = x118 & n227 ;
  assign n8401 = n8400 ^ n8393 ;
  assign n8387 = x2 & x120 ;
  assign n8388 = n8387 ^ x121 ;
  assign n8389 = ~x1 & n8388 ;
  assign n8372 = x120 & n8107 ;
  assign n8374 = n8372 ^ n8108 ;
  assign n8375 = x121 & n8374 ;
  assign n8373 = ~x121 & ~n8372 ;
  assign n8376 = n8375 ^ n8373 ;
  assign n8378 = x122 ^ x1 ;
  assign n8377 = x122 ^ x2 ;
  assign n8379 = n8378 ^ n8377 ;
  assign n8380 = n8376 & n8379 ;
  assign n8381 = n8380 ^ n8378 ;
  assign n8384 = n8381 ^ n8109 ;
  assign n8390 = n8389 ^ n8384 ;
  assign n8391 = ~x0 & n8390 ;
  assign n8392 = n8391 ^ n8381 ;
  assign n8402 = n8401 ^ n8392 ;
  assign n8633 = n8632 ^ n8402 ;
  assign n8369 = n8364 ^ n8355 ;
  assign n8370 = n8361 & n8369 ;
  assign n8371 = n8370 ^ n8364 ;
  assign n8634 = n8633 ^ n8371 ;
  assign n8638 = n8637 ^ n8634 ;
  assign n8918 = x119 & n227 ;
  assign n8908 = x2 & x121 ;
  assign n8909 = n8908 ^ x122 ;
  assign n8910 = ~x1 & n8909 ;
  assign n8896 = ~x122 & ~n8375 ;
  assign n8895 = x122 & ~n8373 ;
  assign n8897 = n8896 ^ n8895 ;
  assign n8899 = x123 ^ x1 ;
  assign n8898 = x123 ^ x2 ;
  assign n8900 = n8899 ^ n8898 ;
  assign n8901 = n8897 & n8900 ;
  assign n8902 = n8901 ^ n8899 ;
  assign n8905 = n8902 ^ n8377 ;
  assign n8911 = n8910 ^ n8905 ;
  assign n8912 = ~x0 & n8911 ;
  assign n8913 = n8912 ^ n8902 ;
  assign n8914 = n8913 ^ x5 ;
  assign n8894 = x118 & n234 ;
  assign n8915 = n8914 ^ n8894 ;
  assign n8893 = x120 & n230 ;
  assign n8916 = n8915 ^ n8893 ;
  assign n8891 = n7833 ^ x120 ;
  assign n8892 = n231 & n8891 ;
  assign n8917 = n8916 ^ n8892 ;
  assign n8919 = n8918 ^ n8917 ;
  assign n8888 = x116 & n390 ;
  assign n8881 = x113 & n578 ;
  assign n8874 = x110 & n788 ;
  assign n8866 = n8595 ^ n8414 ;
  assign n8867 = n8601 & n8866 ;
  assign n8868 = n8867 ^ n8595 ;
  assign n8864 = x107 & n1058 ;
  assign n8857 = x104 & n1335 ;
  assign n8849 = n8578 ^ n8423 ;
  assign n8850 = n8584 & n8849 ;
  assign n8851 = n8850 ^ n8578 ;
  assign n8847 = x101 & n1666 ;
  assign n8839 = n8571 ^ n8429 ;
  assign n8840 = n8577 & n8839 ;
  assign n8841 = n8840 ^ n8571 ;
  assign n8837 = x98 & n2014 ;
  assign n8830 = x95 & n2429 ;
  assign n8828 = n2423 & n3323 ;
  assign n8824 = x94 & n2581 ;
  assign n8823 = x96 & n2422 ;
  assign n8825 = n8824 ^ n8823 ;
  assign n8826 = n8825 ^ x29 ;
  assign n8820 = x92 & n2887 ;
  assign n8812 = n8544 ^ n8441 ;
  assign n8813 = n8550 & n8812 ;
  assign n8814 = n8813 ^ n8544 ;
  assign n8810 = x89 & n3383 ;
  assign n8803 = x86 & n3924 ;
  assign n8795 = n8527 ^ n8450 ;
  assign n8796 = n8533 & n8795 ;
  assign n8797 = n8796 ^ n8527 ;
  assign n8793 = x83 & n4467 ;
  assign n8786 = x80 & n5102 ;
  assign n8777 = x71 & n7179 ;
  assign n8767 = x67 & n7935 ;
  assign n8766 = x69 & n7938 ;
  assign n8768 = n8767 ^ n8766 ;
  assign n8769 = n8768 ^ x56 ;
  assign n8765 = ~n375 & n7939 ;
  assign n8770 = n8769 ^ n8765 ;
  assign n8764 = x68 & n7931 ;
  assign n8771 = n8770 ^ n8764 ;
  assign n8755 = x59 & ~n8224 ;
  assign n8756 = ~n8488 & n8755 ;
  assign n8757 = n8756 ^ x59 ;
  assign n8752 = x66 & n8223 ;
  assign n8739 = x59 ^ x58 ;
  assign n8744 = n8223 & ~n8739 ;
  assign n8745 = n8744 ^ n8223 ;
  assign n8748 = x65 & n8745 ;
  assign n8480 = x58 ^ x57 ;
  assign n8740 = ~n8223 & ~n8480 ;
  assign n8741 = n8739 & n8740 ;
  assign n8749 = n8748 ^ n8741 ;
  assign n8750 = ~x64 & n8749 ;
  assign n8751 = n8750 ^ n8741 ;
  assign n8753 = n8752 ^ n8751 ;
  assign n8737 = ~n8223 & n8480 ;
  assign n8738 = x65 & n8737 ;
  assign n8754 = n8753 ^ n8738 ;
  assign n8758 = n8757 ^ n8754 ;
  assign n8759 = n8758 ^ n8498 ;
  assign n8760 = n8759 ^ n8488 ;
  assign n8761 = n8760 ^ n8758 ;
  assign n8762 = ~n8490 & n8761 ;
  assign n8763 = n8762 ^ n8759 ;
  assign n8772 = n8771 ^ n8763 ;
  assign n8773 = n8772 ^ x53 ;
  assign n8736 = x70 & n7171 ;
  assign n8774 = n8773 ^ n8736 ;
  assign n8735 = x72 & n7174 ;
  assign n8775 = n8774 ^ n8735 ;
  assign n8734 = n556 & n7175 ;
  assign n8776 = n8775 ^ n8734 ;
  assign n8778 = n8777 ^ n8776 ;
  assign n8731 = n8499 ^ n8474 ;
  assign n8732 = n8505 & n8731 ;
  assign n8733 = n8732 ^ n8499 ;
  assign n8779 = n8778 ^ n8733 ;
  assign n8721 = x73 & n6677 ;
  assign n8720 = x75 & n6428 ;
  assign n8722 = n8721 ^ n8720 ;
  assign n8723 = n8722 ^ x50 ;
  assign n8719 = ~n774 & n6429 ;
  assign n8724 = n8723 ^ n8719 ;
  assign n8718 = x74 & n6433 ;
  assign n8725 = n8724 ^ n8718 ;
  assign n8726 = n8725 ^ n8506 ;
  assign n8727 = n8726 ^ n8468 ;
  assign n8728 = n8727 ^ n8725 ;
  assign n8729 = n8512 & n8728 ;
  assign n8730 = n8729 ^ n8726 ;
  assign n8780 = n8779 ^ n8730 ;
  assign n8715 = n8513 ^ n8462 ;
  assign n8716 = n8519 & n8715 ;
  assign n8708 = x76 & n5965 ;
  assign n8707 = x78 & n5729 ;
  assign n8709 = n8708 ^ n8707 ;
  assign n8710 = n8709 ^ x47 ;
  assign n8706 = ~n1025 & n5730 ;
  assign n8711 = n8710 ^ n8706 ;
  assign n8705 = x77 & n5736 ;
  assign n8712 = n8711 ^ n8705 ;
  assign n8713 = n8712 ^ n8513 ;
  assign n8717 = n8716 ^ n8713 ;
  assign n8781 = n8780 ^ n8717 ;
  assign n8782 = n8781 ^ x44 ;
  assign n8704 = x79 & n5094 ;
  assign n8783 = n8782 ^ n8704 ;
  assign n8703 = x81 & n5097 ;
  assign n8784 = n8783 ^ n8703 ;
  assign n8702 = n1305 & n5098 ;
  assign n8785 = n8784 ^ n8702 ;
  assign n8787 = n8786 ^ n8785 ;
  assign n8699 = n8520 ^ n8456 ;
  assign n8700 = n8526 & n8699 ;
  assign n8701 = n8700 ^ n8520 ;
  assign n8788 = n8787 ^ n8701 ;
  assign n8789 = n8788 ^ x41 ;
  assign n8698 = x82 & n4474 ;
  assign n8790 = n8789 ^ n8698 ;
  assign n8697 = x84 & n4471 ;
  assign n8791 = n8790 ^ n8697 ;
  assign n8696 = n1624 & n4472 ;
  assign n8792 = n8791 ^ n8696 ;
  assign n8794 = n8793 ^ n8792 ;
  assign n8798 = n8797 ^ n8794 ;
  assign n8799 = n8798 ^ x38 ;
  assign n8695 = x85 & n3916 ;
  assign n8800 = n8799 ^ n8695 ;
  assign n8694 = x87 & n3919 ;
  assign n8801 = n8800 ^ n8694 ;
  assign n8693 = n1982 & n3920 ;
  assign n8802 = n8801 ^ n8693 ;
  assign n8804 = n8803 ^ n8802 ;
  assign n8690 = n8543 ^ n8534 ;
  assign n8691 = ~n8540 & n8690 ;
  assign n8692 = n8691 ^ n8543 ;
  assign n8805 = n8804 ^ n8692 ;
  assign n8806 = n8805 ^ x35 ;
  assign n8689 = x88 & n3375 ;
  assign n8807 = n8806 ^ n8689 ;
  assign n8688 = x90 & n3378 ;
  assign n8808 = n8807 ^ n8688 ;
  assign n8687 = n2386 & n3379 ;
  assign n8809 = n8808 ^ n8687 ;
  assign n8811 = n8810 ^ n8809 ;
  assign n8815 = n8814 ^ n8811 ;
  assign n8816 = n8815 ^ x32 ;
  assign n8686 = x91 & n2879 ;
  assign n8817 = n8816 ^ n8686 ;
  assign n8685 = x93 & n2882 ;
  assign n8818 = n8817 ^ n8685 ;
  assign n8684 = n2836 & n2883 ;
  assign n8819 = n8818 ^ n8684 ;
  assign n8821 = n8820 ^ n8819 ;
  assign n8681 = n8560 ^ n8551 ;
  assign n8682 = ~n8557 & n8681 ;
  assign n8683 = n8682 ^ n8560 ;
  assign n8822 = n8821 ^ n8683 ;
  assign n8827 = n8826 ^ n8822 ;
  assign n8829 = n8828 ^ n8827 ;
  assign n8831 = n8830 ^ n8829 ;
  assign n8678 = n8569 ^ n8435 ;
  assign n8679 = n8570 & n8678 ;
  assign n8680 = n8679 ^ n8569 ;
  assign n8832 = n8831 ^ n8680 ;
  assign n8833 = n8832 ^ x26 ;
  assign n8677 = x97 & n2018 ;
  assign n8834 = n8833 ^ n8677 ;
  assign n8676 = x99 & n2021 ;
  assign n8835 = n8834 ^ n8676 ;
  assign n8675 = n2022 & n3843 ;
  assign n8836 = n8835 ^ n8675 ;
  assign n8838 = n8837 ^ n8836 ;
  assign n8842 = n8841 ^ n8838 ;
  assign n8843 = n8842 ^ x23 ;
  assign n8674 = x100 & n1658 ;
  assign n8844 = n8843 ^ n8674 ;
  assign n8673 = x102 & n1661 ;
  assign n8845 = n8844 ^ n8673 ;
  assign n8672 = n1662 & n4410 ;
  assign n8846 = n8845 ^ n8672 ;
  assign n8848 = n8847 ^ n8846 ;
  assign n8852 = n8851 ^ n8848 ;
  assign n8853 = n8852 ^ x20 ;
  assign n8671 = x103 & n1327 ;
  assign n8854 = n8853 ^ n8671 ;
  assign n8670 = x105 & n1330 ;
  assign n8855 = n8854 ^ n8670 ;
  assign n8669 = n1331 & ~n5023 ;
  assign n8856 = n8855 ^ n8669 ;
  assign n8858 = n8857 ^ n8856 ;
  assign n8666 = n8594 ^ n8585 ;
  assign n8667 = ~n8591 & n8666 ;
  assign n8668 = n8667 ^ n8594 ;
  assign n8859 = n8858 ^ n8668 ;
  assign n8860 = n8859 ^ x17 ;
  assign n8665 = x106 & n1050 ;
  assign n8861 = n8860 ^ n8665 ;
  assign n8664 = x108 & n1053 ;
  assign n8862 = n8861 ^ n8664 ;
  assign n8663 = n1054 & n5670 ;
  assign n8863 = n8862 ^ n8663 ;
  assign n8865 = n8864 ^ n8863 ;
  assign n8869 = n8868 ^ n8865 ;
  assign n8870 = n8869 ^ x14 ;
  assign n8662 = x109 & n877 ;
  assign n8871 = n8870 ^ n8662 ;
  assign n8661 = x111 & n782 ;
  assign n8872 = n8871 ^ n8661 ;
  assign n8660 = n783 & ~n6360 ;
  assign n8873 = n8872 ^ n8660 ;
  assign n8875 = n8874 ^ n8873 ;
  assign n8657 = n8611 ^ n8602 ;
  assign n8658 = ~n8608 & ~n8657 ;
  assign n8659 = n8658 ^ n8611 ;
  assign n8876 = n8875 ^ n8659 ;
  assign n8877 = n8876 ^ x11 ;
  assign n8656 = x112 & n647 ;
  assign n8878 = n8877 ^ n8656 ;
  assign n8655 = x114 & ~n572 ;
  assign n8879 = n8878 ^ n8655 ;
  assign n8654 = ~n573 & ~n7092 ;
  assign n8880 = n8879 ^ n8654 ;
  assign n8882 = n8881 ^ n8880 ;
  assign n8651 = n8621 ^ n8612 ;
  assign n8652 = n8618 & n8651 ;
  assign n8653 = n8652 ^ n8621 ;
  assign n8883 = n8882 ^ n8653 ;
  assign n8884 = n8883 ^ x8 ;
  assign n8650 = x115 & n446 ;
  assign n8885 = n8884 ^ n8650 ;
  assign n8649 = x117 & n383 ;
  assign n8886 = n8885 ^ n8649 ;
  assign n8648 = n384 & ~n7850 ;
  assign n8887 = n8886 ^ n8648 ;
  assign n8889 = n8888 ^ n8887 ;
  assign n8645 = n8631 ^ n8622 ;
  assign n8646 = ~n8628 & n8645 ;
  assign n8647 = n8646 ^ n8631 ;
  assign n8890 = n8889 ^ n8647 ;
  assign n8920 = n8919 ^ n8890 ;
  assign n8639 = n8637 ^ n8632 ;
  assign n8642 = n8639 ^ n8392 ;
  assign n8643 = n8642 ^ n8371 ;
  assign n8644 = ~n8402 & ~n8643 ;
  assign n8921 = n8920 ^ n8644 ;
  assign n8640 = n8632 ^ n8371 ;
  assign n8641 = ~n8639 & n8640 ;
  assign n8922 = n8921 ^ n8641 ;
  assign n9209 = n8883 ^ n8647 ;
  assign n9210 = n8889 & n9209 ;
  assign n9211 = n9210 ^ n8883 ;
  assign n9207 = x117 & n390 ;
  assign n9199 = n8876 ^ n8653 ;
  assign n9200 = ~n8882 & n9199 ;
  assign n9201 = n9200 ^ n8876 ;
  assign n9197 = x114 & n578 ;
  assign n9189 = n8869 ^ n8659 ;
  assign n9190 = n8875 & ~n9189 ;
  assign n9191 = n9190 ^ n8869 ;
  assign n9187 = x111 & n788 ;
  assign n9180 = x108 & n1058 ;
  assign n9172 = n8852 ^ n8668 ;
  assign n9173 = n8858 & n9172 ;
  assign n9174 = n9173 ^ n8852 ;
  assign n9170 = x105 & n1335 ;
  assign n9163 = x102 & n1666 ;
  assign n9156 = x99 & n2014 ;
  assign n9148 = n8822 ^ n8680 ;
  assign n9149 = n8831 & n9148 ;
  assign n9150 = n9149 ^ n8822 ;
  assign n9142 = x95 & n2581 ;
  assign n9141 = x97 & n2422 ;
  assign n9143 = n9142 ^ n9141 ;
  assign n9144 = n9143 ^ x29 ;
  assign n9140 = n2423 & n3494 ;
  assign n9145 = n9144 ^ n9140 ;
  assign n9139 = x96 & n2429 ;
  assign n9146 = n9145 ^ n9139 ;
  assign n9135 = n8815 ^ n8683 ;
  assign n9136 = n8821 & n9135 ;
  assign n9137 = n9136 ^ n8815 ;
  assign n9133 = x93 & n2887 ;
  assign n9126 = x90 & n3383 ;
  assign n9118 = n8798 ^ n8692 ;
  assign n9119 = n8804 & n9118 ;
  assign n9120 = n9119 ^ n8798 ;
  assign n9116 = x87 & n3924 ;
  assign n9109 = x84 & n4467 ;
  assign n9102 = x81 & n5102 ;
  assign n9095 = x78 & n5736 ;
  assign n9088 = x75 & n6433 ;
  assign n9080 = n8772 ^ n8733 ;
  assign n9081 = n8778 & n9080 ;
  assign n9082 = n9081 ^ n8772 ;
  assign n9078 = x72 & n7179 ;
  assign n9070 = n8771 ^ n8758 ;
  assign n9071 = n8763 & n9070 ;
  assign n9072 = n9071 ^ n8758 ;
  assign n9068 = x69 & n7931 ;
  assign n9058 = x65 & n8741 ;
  assign n9057 = x66 & n8737 ;
  assign n9059 = n9058 ^ n9057 ;
  assign n9060 = n9059 ^ x59 ;
  assign n9054 = ~n153 & ~n8739 ;
  assign n9055 = n9054 ^ n291 ;
  assign n9056 = n8223 & ~n9055 ;
  assign n9061 = n9060 ^ n9056 ;
  assign n9046 = x60 ^ x59 ;
  assign n9047 = x64 & n9046 ;
  assign n9048 = ~n8754 & n8756 ;
  assign n9050 = ~n9047 & ~n9048 ;
  assign n9062 = n9061 ^ n9050 ;
  assign n9049 = n9048 ^ n9047 ;
  assign n9051 = n9050 ^ n9049 ;
  assign n9063 = n9062 ^ n9051 ;
  assign n9064 = n9063 ^ x56 ;
  assign n9045 = x68 & n7935 ;
  assign n9065 = n9064 ^ n9045 ;
  assign n9044 = x70 & n7938 ;
  assign n9066 = n9065 ^ n9044 ;
  assign n9043 = ~n436 & n7939 ;
  assign n9067 = n9066 ^ n9043 ;
  assign n9069 = n9068 ^ n9067 ;
  assign n9073 = n9072 ^ n9069 ;
  assign n9074 = n9073 ^ x53 ;
  assign n9042 = x71 & n7171 ;
  assign n9075 = n9074 ^ n9042 ;
  assign n9041 = x73 & n7174 ;
  assign n9076 = n9075 ^ n9041 ;
  assign n9040 = n633 & n7175 ;
  assign n9077 = n9076 ^ n9040 ;
  assign n9079 = n9078 ^ n9077 ;
  assign n9083 = n9082 ^ n9079 ;
  assign n9084 = n9083 ^ x50 ;
  assign n9039 = x74 & n6677 ;
  assign n9085 = n9084 ^ n9039 ;
  assign n9038 = x76 & n6428 ;
  assign n9086 = n9085 ^ n9038 ;
  assign n9037 = ~n853 & n6429 ;
  assign n9087 = n9086 ^ n9037 ;
  assign n9089 = n9088 ^ n9087 ;
  assign n9034 = n8779 ^ n8725 ;
  assign n9035 = n8730 & n9034 ;
  assign n9036 = n9035 ^ n8725 ;
  assign n9090 = n9089 ^ n9036 ;
  assign n9091 = n9090 ^ x47 ;
  assign n9033 = x77 & n5965 ;
  assign n9092 = n9091 ^ n9033 ;
  assign n9032 = x79 & n5729 ;
  assign n9093 = n9092 ^ n9032 ;
  assign n9031 = n1118 & n5730 ;
  assign n9094 = n9093 ^ n9031 ;
  assign n9096 = n9095 ^ n9094 ;
  assign n9028 = n8780 ^ n8712 ;
  assign n9029 = n8717 & n9028 ;
  assign n9030 = n9029 ^ n8712 ;
  assign n9097 = n9096 ^ n9030 ;
  assign n9098 = n9097 ^ x44 ;
  assign n9027 = x80 & n5094 ;
  assign n9099 = n9098 ^ n9027 ;
  assign n9026 = x82 & n5097 ;
  assign n9100 = n9099 ^ n9026 ;
  assign n9025 = n1411 & n5098 ;
  assign n9101 = n9100 ^ n9025 ;
  assign n9103 = n9102 ^ n9101 ;
  assign n9022 = n8781 ^ n8701 ;
  assign n9023 = n8787 & n9022 ;
  assign n9024 = n9023 ^ n8781 ;
  assign n9104 = n9103 ^ n9024 ;
  assign n9105 = n9104 ^ x41 ;
  assign n9021 = x83 & n4474 ;
  assign n9106 = n9105 ^ n9021 ;
  assign n9020 = x85 & n4471 ;
  assign n9107 = n9106 ^ n9020 ;
  assign n9019 = n1743 & n4472 ;
  assign n9108 = n9107 ^ n9019 ;
  assign n9110 = n9109 ^ n9108 ;
  assign n9016 = n8797 ^ n8788 ;
  assign n9017 = ~n8794 & n9016 ;
  assign n9018 = n9017 ^ n8797 ;
  assign n9111 = n9110 ^ n9018 ;
  assign n9112 = n9111 ^ x38 ;
  assign n9015 = x86 & n3916 ;
  assign n9113 = n9112 ^ n9015 ;
  assign n9014 = x88 & n3919 ;
  assign n9114 = n9113 ^ n9014 ;
  assign n9013 = n2119 & n3920 ;
  assign n9115 = n9114 ^ n9013 ;
  assign n9117 = n9116 ^ n9115 ;
  assign n9121 = n9120 ^ n9117 ;
  assign n9122 = n9121 ^ x35 ;
  assign n9012 = x89 & n3375 ;
  assign n9123 = n9122 ^ n9012 ;
  assign n9011 = x91 & n3378 ;
  assign n9124 = n9123 ^ n9011 ;
  assign n9010 = n2542 & n3379 ;
  assign n9125 = n9124 ^ n9010 ;
  assign n9127 = n9126 ^ n9125 ;
  assign n9007 = n8814 ^ n8805 ;
  assign n9008 = ~n8811 & n9007 ;
  assign n9009 = n9008 ^ n8814 ;
  assign n9128 = n9127 ^ n9009 ;
  assign n9129 = n9128 ^ x32 ;
  assign n9006 = x92 & n2879 ;
  assign n9130 = n9129 ^ n9006 ;
  assign n9005 = x94 & n2882 ;
  assign n9131 = n9130 ^ n9005 ;
  assign n9004 = n2883 & n2997 ;
  assign n9132 = n9131 ^ n9004 ;
  assign n9134 = n9133 ^ n9132 ;
  assign n9138 = n9137 ^ n9134 ;
  assign n9147 = n9146 ^ n9138 ;
  assign n9151 = n9150 ^ n9147 ;
  assign n9152 = n9151 ^ x26 ;
  assign n9003 = x98 & n2018 ;
  assign n9153 = n9152 ^ n9003 ;
  assign n9002 = x100 & n2021 ;
  assign n9154 = n9153 ^ n9002 ;
  assign n9001 = n2022 & n4034 ;
  assign n9155 = n9154 ^ n9001 ;
  assign n9157 = n9156 ^ n9155 ;
  assign n8998 = n8841 ^ n8832 ;
  assign n8999 = ~n8838 & n8998 ;
  assign n9000 = n8999 ^ n8841 ;
  assign n9158 = n9157 ^ n9000 ;
  assign n9159 = n9158 ^ x23 ;
  assign n8997 = x101 & n1658 ;
  assign n9160 = n9159 ^ n8997 ;
  assign n8996 = x103 & n1661 ;
  assign n9161 = n9160 ^ n8996 ;
  assign n8995 = n1662 & ~n4615 ;
  assign n9162 = n9161 ^ n8995 ;
  assign n9164 = n9163 ^ n9162 ;
  assign n8992 = n8851 ^ n8842 ;
  assign n8993 = ~n8848 & n8992 ;
  assign n8994 = n8993 ^ n8851 ;
  assign n9165 = n9164 ^ n8994 ;
  assign n9166 = n9165 ^ x20 ;
  assign n8991 = x104 & n1327 ;
  assign n9167 = n9166 ^ n8991 ;
  assign n8990 = x106 & n1330 ;
  assign n9168 = n9167 ^ n8990 ;
  assign n8989 = n1331 & ~n5240 ;
  assign n9169 = n9168 ^ n8989 ;
  assign n9171 = n9170 ^ n9169 ;
  assign n9175 = n9174 ^ n9171 ;
  assign n9176 = n9175 ^ x17 ;
  assign n8988 = x107 & n1050 ;
  assign n9177 = n9176 ^ n8988 ;
  assign n8987 = x109 & n1053 ;
  assign n9178 = n9177 ^ n8987 ;
  assign n8986 = n1054 & n5902 ;
  assign n9179 = n9178 ^ n8986 ;
  assign n9181 = n9180 ^ n9179 ;
  assign n8983 = n8868 ^ n8859 ;
  assign n8984 = ~n8865 & n8983 ;
  assign n8985 = n8984 ^ n8868 ;
  assign n9182 = n9181 ^ n8985 ;
  assign n9183 = n9182 ^ x14 ;
  assign n8982 = x110 & n877 ;
  assign n9184 = n9183 ^ n8982 ;
  assign n8981 = x112 & n782 ;
  assign n9185 = n9184 ^ n8981 ;
  assign n8980 = n783 & ~n6600 ;
  assign n9186 = n9185 ^ n8980 ;
  assign n9188 = n9187 ^ n9186 ;
  assign n9192 = n9191 ^ n9188 ;
  assign n9193 = n9192 ^ x11 ;
  assign n8979 = x113 & n647 ;
  assign n9194 = n9193 ^ n8979 ;
  assign n8978 = x115 & ~n572 ;
  assign n9195 = n9194 ^ n8978 ;
  assign n8977 = ~n573 & ~n7343 ;
  assign n9196 = n9195 ^ n8977 ;
  assign n9198 = n9197 ^ n9196 ;
  assign n9202 = n9201 ^ n9198 ;
  assign n9203 = n9202 ^ x8 ;
  assign n8976 = x116 & n446 ;
  assign n9204 = n9203 ^ n8976 ;
  assign n8975 = x118 & n383 ;
  assign n9205 = n9204 ^ n8975 ;
  assign n8974 = n384 & ~n8123 ;
  assign n9206 = n9205 ^ n8974 ;
  assign n9208 = n9207 ^ n9206 ;
  assign n9212 = n9211 ^ n9208 ;
  assign n8971 = n8913 ^ n8890 ;
  assign n8972 = n8919 & n8971 ;
  assign n8973 = n8972 ^ n8913 ;
  assign n9213 = n9212 ^ n8973 ;
  assign n8965 = x119 & n234 ;
  assign n8964 = x121 & n230 ;
  assign n8966 = n8965 ^ n8964 ;
  assign n8967 = n8966 ^ x5 ;
  assign n8962 = n8108 ^ x121 ;
  assign n8963 = n231 & n8962 ;
  assign n8968 = n8967 ^ n8963 ;
  assign n8961 = x120 & n227 ;
  assign n8969 = n8968 ^ n8961 ;
  assign n8955 = x2 & x122 ;
  assign n8956 = n8955 ^ x123 ;
  assign n8957 = ~x1 & n8956 ;
  assign n8944 = x123 ^ x122 ;
  assign n8945 = n8897 & n8944 ;
  assign n8947 = x124 ^ x1 ;
  assign n8946 = x124 ^ x2 ;
  assign n8948 = n8947 ^ n8946 ;
  assign n8949 = ~n8945 & n8948 ;
  assign n8950 = n8949 ^ n8947 ;
  assign n8952 = n8950 ^ n8898 ;
  assign n8958 = n8957 ^ n8952 ;
  assign n8959 = ~x0 & n8958 ;
  assign n8960 = n8959 ^ n8950 ;
  assign n8970 = n8969 ^ n8960 ;
  assign n9214 = n9213 ^ n8970 ;
  assign n8923 = n8392 & n8401 ;
  assign n8924 = n8632 & n8923 ;
  assign n8925 = ~n8371 & n8924 ;
  assign n8926 = n8637 & ~n8925 ;
  assign n8928 = n8923 ^ n8402 ;
  assign n8929 = ~n8632 & ~n8928 ;
  assign n8936 = ~n8920 & n8929 ;
  assign n8937 = n8371 & n8936 ;
  assign n8930 = n8371 & ~n8929 ;
  assign n8931 = n8924 ^ n8632 ;
  assign n8932 = n8931 ^ n8402 ;
  assign n8933 = n8930 & n8932 ;
  assign n8934 = n8933 ^ n8929 ;
  assign n8927 = n8920 ^ n8634 ;
  assign n8935 = n8934 ^ n8927 ;
  assign n8938 = n8937 ^ n8935 ;
  assign n8939 = n8926 & ~n8938 ;
  assign n8940 = n8939 ^ n8925 ;
  assign n8941 = n8920 & ~n8934 ;
  assign n8942 = ~n8940 & n8941 ;
  assign n8943 = n8942 ^ n8940 ;
  assign n9215 = n9214 ^ n8943 ;
  assign n9508 = x115 & n578 ;
  assign n9501 = x112 & n788 ;
  assign n9493 = n9175 ^ n8985 ;
  assign n9494 = n9181 & n9493 ;
  assign n9495 = n9494 ^ n9175 ;
  assign n9491 = x109 & n1058 ;
  assign n9484 = x106 & n1335 ;
  assign n9476 = n9158 ^ n8994 ;
  assign n9477 = n9164 & n9476 ;
  assign n9478 = n9477 ^ n9158 ;
  assign n9474 = x103 & n1666 ;
  assign n9466 = n9151 ^ n9000 ;
  assign n9467 = n9157 & n9466 ;
  assign n9468 = n9467 ^ n9151 ;
  assign n9464 = x100 & n2014 ;
  assign n9457 = x97 & n2429 ;
  assign n9455 = n2423 & n3660 ;
  assign n9451 = x96 & n2581 ;
  assign n9450 = x98 & n2422 ;
  assign n9452 = n9451 ^ n9450 ;
  assign n9453 = n9452 ^ x29 ;
  assign n9447 = x94 & n2887 ;
  assign n9439 = n9121 ^ n9009 ;
  assign n9440 = n9127 & n9439 ;
  assign n9441 = n9440 ^ n9121 ;
  assign n9437 = x91 & n3383 ;
  assign n9430 = x88 & n3924 ;
  assign n9422 = n9104 ^ n9018 ;
  assign n9423 = n9110 & n9422 ;
  assign n9424 = n9423 ^ n9104 ;
  assign n9420 = x85 & n4467 ;
  assign n9413 = x82 & n5102 ;
  assign n9406 = x79 & n5736 ;
  assign n9398 = x73 & n7179 ;
  assign n9387 = x69 & n7935 ;
  assign n9386 = x71 & n7938 ;
  assign n9388 = n9387 ^ n9386 ;
  assign n9389 = n9388 ^ x56 ;
  assign n9385 = ~n493 & n7939 ;
  assign n9390 = n9389 ^ n9385 ;
  assign n9384 = x70 & n7931 ;
  assign n9391 = n9390 ^ n9384 ;
  assign n9381 = ~n9050 & n9061 ;
  assign n9378 = x65 ^ x60 ;
  assign n9379 = n9046 & ~n9378 ;
  assign n9374 = x59 & x60 ;
  assign n9375 = n9374 ^ x61 ;
  assign n9376 = ~x64 & n9375 ;
  assign n9370 = x61 ^ x59 ;
  assign n9377 = n9376 ^ n9370 ;
  assign n9380 = n9379 ^ n9377 ;
  assign n9382 = n9381 ^ n9380 ;
  assign n9366 = ~n340 & n8745 ;
  assign n9365 = x67 & n8737 ;
  assign n9367 = n9366 ^ n9365 ;
  assign n9363 = x66 & n8741 ;
  assign n9362 = x68 & n8744 ;
  assign n9364 = n9363 ^ n9362 ;
  assign n9368 = n9367 ^ n9364 ;
  assign n9369 = n9368 ^ x59 ;
  assign n9383 = n9382 ^ n9369 ;
  assign n9392 = n9391 ^ n9383 ;
  assign n9359 = n9072 ^ n9063 ;
  assign n9360 = ~n9069 & n9359 ;
  assign n9361 = n9360 ^ n9072 ;
  assign n9393 = n9392 ^ n9361 ;
  assign n9394 = n9393 ^ x53 ;
  assign n9358 = x72 & n7171 ;
  assign n9395 = n9394 ^ n9358 ;
  assign n9357 = x74 & n7174 ;
  assign n9396 = n9395 ^ n9357 ;
  assign n9356 = n699 & n7175 ;
  assign n9397 = n9396 ^ n9356 ;
  assign n9399 = n9398 ^ n9397 ;
  assign n9353 = n9082 ^ n9073 ;
  assign n9354 = ~n9079 & n9353 ;
  assign n9355 = n9354 ^ n9082 ;
  assign n9400 = n9399 ^ n9355 ;
  assign n9343 = x75 & n6677 ;
  assign n9342 = x77 & n6428 ;
  assign n9344 = n9343 ^ n9342 ;
  assign n9345 = n9344 ^ x50 ;
  assign n9341 = ~n939 & n6429 ;
  assign n9346 = n9345 ^ n9341 ;
  assign n9340 = x76 & n6433 ;
  assign n9347 = n9346 ^ n9340 ;
  assign n9348 = n9347 ^ n9083 ;
  assign n9349 = n9348 ^ n9036 ;
  assign n9350 = n9349 ^ n9347 ;
  assign n9351 = n9089 & n9350 ;
  assign n9352 = n9351 ^ n9348 ;
  assign n9401 = n9400 ^ n9352 ;
  assign n9402 = n9401 ^ x47 ;
  assign n9339 = x78 & n5965 ;
  assign n9403 = n9402 ^ n9339 ;
  assign n9338 = x80 & n5729 ;
  assign n9404 = n9403 ^ n9338 ;
  assign n9337 = n1206 & n5730 ;
  assign n9405 = n9404 ^ n9337 ;
  assign n9407 = n9406 ^ n9405 ;
  assign n9334 = n9090 ^ n9030 ;
  assign n9335 = n9096 & n9334 ;
  assign n9336 = n9335 ^ n9090 ;
  assign n9408 = n9407 ^ n9336 ;
  assign n9409 = n9408 ^ x44 ;
  assign n9333 = x81 & n5094 ;
  assign n9410 = n9409 ^ n9333 ;
  assign n9332 = x83 & n5097 ;
  assign n9411 = n9410 ^ n9332 ;
  assign n9331 = n1512 & n5098 ;
  assign n9412 = n9411 ^ n9331 ;
  assign n9414 = n9413 ^ n9412 ;
  assign n9328 = n9097 ^ n9024 ;
  assign n9329 = n9103 & n9328 ;
  assign n9330 = n9329 ^ n9097 ;
  assign n9415 = n9414 ^ n9330 ;
  assign n9416 = n9415 ^ x41 ;
  assign n9327 = x84 & n4474 ;
  assign n9417 = n9416 ^ n9327 ;
  assign n9326 = x86 & n4471 ;
  assign n9418 = n9417 ^ n9326 ;
  assign n9325 = n1857 & n4472 ;
  assign n9419 = n9418 ^ n9325 ;
  assign n9421 = n9420 ^ n9419 ;
  assign n9425 = n9424 ^ n9421 ;
  assign n9426 = n9425 ^ x38 ;
  assign n9324 = x87 & n3916 ;
  assign n9427 = n9426 ^ n9324 ;
  assign n9323 = x89 & n3919 ;
  assign n9428 = n9427 ^ n9323 ;
  assign n9322 = n2249 & n3920 ;
  assign n9429 = n9428 ^ n9322 ;
  assign n9431 = n9430 ^ n9429 ;
  assign n9319 = n9120 ^ n9111 ;
  assign n9320 = ~n9117 & n9319 ;
  assign n9321 = n9320 ^ n9120 ;
  assign n9432 = n9431 ^ n9321 ;
  assign n9433 = n9432 ^ x35 ;
  assign n9318 = x90 & n3375 ;
  assign n9434 = n9433 ^ n9318 ;
  assign n9317 = x92 & n3378 ;
  assign n9435 = n9434 ^ n9317 ;
  assign n9316 = n2684 & n3379 ;
  assign n9436 = n9435 ^ n9316 ;
  assign n9438 = n9437 ^ n9436 ;
  assign n9442 = n9441 ^ n9438 ;
  assign n9443 = n9442 ^ x32 ;
  assign n9315 = x93 & n2879 ;
  assign n9444 = n9443 ^ n9315 ;
  assign n9314 = x95 & n2882 ;
  assign n9445 = n9444 ^ n9314 ;
  assign n9313 = n2883 & n3159 ;
  assign n9446 = n9445 ^ n9313 ;
  assign n9448 = n9447 ^ n9446 ;
  assign n9310 = n9137 ^ n9128 ;
  assign n9311 = ~n9134 & n9310 ;
  assign n9312 = n9311 ^ n9137 ;
  assign n9449 = n9448 ^ n9312 ;
  assign n9454 = n9453 ^ n9449 ;
  assign n9456 = n9455 ^ n9454 ;
  assign n9458 = n9457 ^ n9456 ;
  assign n9307 = n9150 ^ n9146 ;
  assign n9308 = ~n9147 & n9307 ;
  assign n9309 = n9308 ^ n9150 ;
  assign n9459 = n9458 ^ n9309 ;
  assign n9460 = n9459 ^ x26 ;
  assign n9306 = x99 & n2018 ;
  assign n9461 = n9460 ^ n9306 ;
  assign n9305 = x101 & n2021 ;
  assign n9462 = n9461 ^ n9305 ;
  assign n9304 = n2022 & n4215 ;
  assign n9463 = n9462 ^ n9304 ;
  assign n9465 = n9464 ^ n9463 ;
  assign n9469 = n9468 ^ n9465 ;
  assign n9470 = n9469 ^ x23 ;
  assign n9303 = x102 & n1658 ;
  assign n9471 = n9470 ^ n9303 ;
  assign n9302 = x104 & n1661 ;
  assign n9472 = n9471 ^ n9302 ;
  assign n9301 = n1662 & ~n4814 ;
  assign n9473 = n9472 ^ n9301 ;
  assign n9475 = n9474 ^ n9473 ;
  assign n9479 = n9478 ^ n9475 ;
  assign n9480 = n9479 ^ x20 ;
  assign n9300 = x105 & n1327 ;
  assign n9481 = n9480 ^ n9300 ;
  assign n9299 = x107 & n1330 ;
  assign n9482 = n9481 ^ n9299 ;
  assign n9298 = n1331 & ~n5448 ;
  assign n9483 = n9482 ^ n9298 ;
  assign n9485 = n9484 ^ n9483 ;
  assign n9295 = n9174 ^ n9165 ;
  assign n9296 = ~n9171 & n9295 ;
  assign n9297 = n9296 ^ n9174 ;
  assign n9486 = n9485 ^ n9297 ;
  assign n9487 = n9486 ^ x17 ;
  assign n9294 = x108 & n1050 ;
  assign n9488 = n9487 ^ n9294 ;
  assign n9293 = x110 & n1053 ;
  assign n9489 = n9488 ^ n9293 ;
  assign n9292 = n1054 & n6129 ;
  assign n9490 = n9489 ^ n9292 ;
  assign n9492 = n9491 ^ n9490 ;
  assign n9496 = n9495 ^ n9492 ;
  assign n9497 = n9496 ^ x14 ;
  assign n9291 = x111 & n877 ;
  assign n9498 = n9497 ^ n9291 ;
  assign n9290 = x113 & n782 ;
  assign n9499 = n9498 ^ n9290 ;
  assign n9289 = n783 & ~n6839 ;
  assign n9500 = n9499 ^ n9289 ;
  assign n9502 = n9501 ^ n9500 ;
  assign n9286 = n9191 ^ n9182 ;
  assign n9287 = ~n9188 & n9286 ;
  assign n9288 = n9287 ^ n9191 ;
  assign n9503 = n9502 ^ n9288 ;
  assign n9504 = n9503 ^ x11 ;
  assign n9285 = x114 & n647 ;
  assign n9505 = n9504 ^ n9285 ;
  assign n9284 = x116 & ~n572 ;
  assign n9506 = n9505 ^ n9284 ;
  assign n9283 = ~n573 & ~n7588 ;
  assign n9507 = n9506 ^ n9283 ;
  assign n9509 = n9508 ^ n9507 ;
  assign n9280 = n9201 ^ n9192 ;
  assign n9281 = ~n9198 & ~n9280 ;
  assign n9282 = n9281 ^ n9201 ;
  assign n9510 = n9509 ^ n9282 ;
  assign n9273 = x2 & x123 ;
  assign n9274 = n9273 ^ x124 ;
  assign n9275 = ~x1 & n9274 ;
  assign n9256 = ~x124 & n8896 ;
  assign n9257 = ~x123 & x124 ;
  assign n9258 = n8895 & n9257 ;
  assign n9259 = n9258 ^ x123 ;
  assign n9260 = n9256 & n9259 ;
  assign n9261 = n9260 ^ n9259 ;
  assign n9262 = n9261 ^ x124 ;
  assign n9263 = x125 ^ x1 ;
  assign n9264 = n9263 ^ x2 ;
  assign n9265 = n9264 ^ x125 ;
  assign n9266 = ~n9262 & n9265 ;
  assign n9267 = n9266 ^ n9263 ;
  assign n9270 = n9267 ^ n8946 ;
  assign n9276 = n9275 ^ n9270 ;
  assign n9277 = ~x0 & n9276 ;
  assign n9278 = n9277 ^ n9267 ;
  assign n9250 = x120 & n234 ;
  assign n9249 = x122 & n230 ;
  assign n9251 = n9250 ^ n9249 ;
  assign n9252 = n9251 ^ x5 ;
  assign n9247 = n8376 ^ x122 ;
  assign n9248 = n231 & ~n9247 ;
  assign n9253 = n9252 ^ n9248 ;
  assign n9246 = x121 & n227 ;
  assign n9254 = n9253 ^ n9246 ;
  assign n9241 = x117 & n446 ;
  assign n9240 = x119 & n383 ;
  assign n9242 = n9241 ^ n9240 ;
  assign n9243 = n9242 ^ x8 ;
  assign n9239 = n384 & n8394 ;
  assign n9244 = n9243 ^ n9239 ;
  assign n9238 = x118 & n390 ;
  assign n9245 = n9244 ^ n9238 ;
  assign n9255 = n9254 ^ n9245 ;
  assign n9279 = n9278 ^ n9255 ;
  assign n9511 = n9510 ^ n9279 ;
  assign n9235 = n9211 ^ n9202 ;
  assign n9236 = n9208 & ~n9235 ;
  assign n9237 = n9236 ^ n9211 ;
  assign n9512 = n9511 ^ n9237 ;
  assign n9217 = n8960 & n8969 ;
  assign n9216 = ~n8973 & n9212 ;
  assign n9220 = n9216 ^ n9213 ;
  assign n9221 = n9217 & n9220 ;
  assign n9218 = n9217 ^ n8970 ;
  assign n9219 = n9216 & ~n9218 ;
  assign n9222 = n9221 ^ n9219 ;
  assign n9223 = n9218 ^ n9212 ;
  assign n9224 = n9218 ^ n8973 ;
  assign n9225 = ~n9223 & ~n9224 ;
  assign n9226 = n9225 ^ n9212 ;
  assign n9227 = ~n9217 & n9226 ;
  assign n9228 = n9227 ^ n8943 ;
  assign n9229 = n9228 ^ n9227 ;
  assign n9230 = n9227 ^ n9214 ;
  assign n9231 = n9230 ^ n9227 ;
  assign n9232 = n9229 & ~n9231 ;
  assign n9233 = n9232 ^ n9227 ;
  assign n9234 = ~n9222 & ~n9233 ;
  assign n9513 = n9512 ^ n9234 ;
  assign n9812 = n9222 ^ n9214 ;
  assign n9813 = n9812 ^ n9227 ;
  assign n9811 = ~n9219 & ~n9512 ;
  assign n9814 = n9813 ^ n9811 ;
  assign n9815 = ~n8943 & ~n9814 ;
  assign n9816 = n9512 ^ n9220 ;
  assign n9817 = n9816 ^ n9217 ;
  assign n9818 = n9815 & ~n9817 ;
  assign n9819 = n9818 ^ n9814 ;
  assign n9820 = ~n9226 & ~n9512 ;
  assign n9821 = n9819 & n9820 ;
  assign n9822 = n9821 ^ n9819 ;
  assign n9514 = n9510 ^ n9245 ;
  assign n9515 = n9514 ^ n9254 ;
  assign n9516 = n9515 ^ n9237 ;
  assign n9800 = x119 & n390 ;
  assign n9797 = x120 & n383 ;
  assign n9795 = x118 & n446 ;
  assign n9789 = x121 & n234 ;
  assign n9788 = x123 & n230 ;
  assign n9790 = n9789 ^ n9788 ;
  assign n9791 = n9790 ^ x5 ;
  assign n9786 = n8897 ^ x123 ;
  assign n9787 = n231 & ~n9786 ;
  assign n9792 = n9791 ^ n9787 ;
  assign n9785 = x122 & n227 ;
  assign n9793 = n9792 ^ n9785 ;
  assign n9794 = n9793 ^ x8 ;
  assign n9796 = n9795 ^ n9794 ;
  assign n9798 = n9797 ^ n9796 ;
  assign n9784 = n384 & n8891 ;
  assign n9799 = n9798 ^ n9784 ;
  assign n9801 = n9800 ^ n9799 ;
  assign n9780 = n9503 ^ n9282 ;
  assign n9781 = n9509 & ~n9780 ;
  assign n9782 = n9781 ^ n9503 ;
  assign n9778 = x116 & n578 ;
  assign n9770 = n9496 ^ n9288 ;
  assign n9771 = n9502 & n9770 ;
  assign n9772 = n9771 ^ n9496 ;
  assign n9768 = x113 & n788 ;
  assign n9761 = x110 & n1058 ;
  assign n9753 = n9479 ^ n9297 ;
  assign n9754 = n9485 & n9753 ;
  assign n9755 = n9754 ^ n9479 ;
  assign n9751 = x107 & n1335 ;
  assign n9744 = x104 & n1666 ;
  assign n9737 = x101 & n2014 ;
  assign n9729 = n9449 ^ n9309 ;
  assign n9730 = n9458 & n9729 ;
  assign n9731 = n9730 ^ n9449 ;
  assign n9723 = x97 & n2581 ;
  assign n9722 = x99 & n2422 ;
  assign n9724 = n9723 ^ n9722 ;
  assign n9725 = n9724 ^ x29 ;
  assign n9721 = n2423 & n3843 ;
  assign n9726 = n9725 ^ n9721 ;
  assign n9720 = x98 & n2429 ;
  assign n9727 = n9726 ^ n9720 ;
  assign n9716 = n9442 ^ n9312 ;
  assign n9717 = n9448 & n9716 ;
  assign n9718 = n9717 ^ n9442 ;
  assign n9714 = x95 & n2887 ;
  assign n9707 = x92 & n3383 ;
  assign n9699 = n9425 ^ n9321 ;
  assign n9700 = n9431 & n9699 ;
  assign n9701 = n9700 ^ n9425 ;
  assign n9697 = x89 & n3924 ;
  assign n9690 = x86 & n4467 ;
  assign n9683 = x83 & n5102 ;
  assign n9675 = n9401 ^ n9336 ;
  assign n9676 = n9407 & n9675 ;
  assign n9677 = n9676 ^ n9401 ;
  assign n9668 = n9391 ^ n9361 ;
  assign n9669 = n9392 & n9668 ;
  assign n9670 = n9669 ^ n9391 ;
  assign n9666 = x71 & n7931 ;
  assign n9659 = n9380 ^ n9369 ;
  assign n9660 = ~n9382 & n9659 ;
  assign n9654 = ~n375 & n8745 ;
  assign n9653 = x68 & n8737 ;
  assign n9655 = n9654 ^ n9653 ;
  assign n9651 = x67 & n8741 ;
  assign n9650 = x69 & n8744 ;
  assign n9652 = n9651 ^ n9650 ;
  assign n9656 = n9655 ^ n9652 ;
  assign n9646 = x62 & ~n9047 ;
  assign n9647 = ~n9380 & n9646 ;
  assign n9648 = n9647 ^ x62 ;
  assign n9643 = x66 & n9046 ;
  assign n9630 = x62 ^ x61 ;
  assign n9635 = n9046 & ~n9630 ;
  assign n9636 = n9635 ^ n9046 ;
  assign n9639 = x65 & n9636 ;
  assign n9372 = x61 ^ x60 ;
  assign n9631 = ~n9046 & ~n9372 ;
  assign n9632 = n9630 & n9631 ;
  assign n9640 = n9639 ^ n9632 ;
  assign n9641 = ~x64 & n9640 ;
  assign n9642 = n9641 ^ n9632 ;
  assign n9644 = n9643 ^ n9642 ;
  assign n9628 = ~n9046 & n9372 ;
  assign n9629 = x65 & n9628 ;
  assign n9645 = n9644 ^ n9629 ;
  assign n9649 = n9648 ^ n9645 ;
  assign n9657 = n9656 ^ n9649 ;
  assign n9658 = n9657 ^ n9368 ;
  assign n9661 = n9660 ^ n9658 ;
  assign n9662 = n9661 ^ x56 ;
  assign n9627 = x70 & n7935 ;
  assign n9663 = n9662 ^ n9627 ;
  assign n9626 = x72 & n7938 ;
  assign n9664 = n9663 ^ n9626 ;
  assign n9625 = n556 & n7939 ;
  assign n9665 = n9664 ^ n9625 ;
  assign n9667 = n9666 ^ n9665 ;
  assign n9671 = n9670 ^ n9667 ;
  assign n9622 = n9393 ^ n9355 ;
  assign n9623 = n9399 & n9622 ;
  assign n9615 = x73 & n7171 ;
  assign n9614 = x75 & n7174 ;
  assign n9616 = n9615 ^ n9614 ;
  assign n9617 = n9616 ^ x53 ;
  assign n9613 = ~n774 & n7175 ;
  assign n9618 = n9617 ^ n9613 ;
  assign n9612 = x74 & n7179 ;
  assign n9619 = n9618 ^ n9612 ;
  assign n9620 = n9619 ^ n9393 ;
  assign n9624 = n9623 ^ n9620 ;
  assign n9672 = n9671 ^ n9624 ;
  assign n9606 = x79 & n5965 ;
  assign n9605 = x81 & n5729 ;
  assign n9607 = n9606 ^ n9605 ;
  assign n9608 = n9607 ^ x47 ;
  assign n9604 = n1305 & n5730 ;
  assign n9609 = n9608 ^ n9604 ;
  assign n9603 = x80 & n5736 ;
  assign n9610 = n9609 ^ n9603 ;
  assign n9598 = x76 & n6677 ;
  assign n9597 = x78 & n6428 ;
  assign n9599 = n9598 ^ n9597 ;
  assign n9600 = n9599 ^ x50 ;
  assign n9596 = ~n1025 & n6429 ;
  assign n9601 = n9600 ^ n9596 ;
  assign n9595 = x77 & n6433 ;
  assign n9602 = n9601 ^ n9595 ;
  assign n9611 = n9610 ^ n9602 ;
  assign n9673 = n9672 ^ n9611 ;
  assign n9592 = n9400 ^ n9347 ;
  assign n9593 = n9352 & n9592 ;
  assign n9594 = n9593 ^ n9347 ;
  assign n9674 = n9673 ^ n9594 ;
  assign n9678 = n9677 ^ n9674 ;
  assign n9679 = n9678 ^ x44 ;
  assign n9591 = x82 & n5094 ;
  assign n9680 = n9679 ^ n9591 ;
  assign n9590 = x84 & n5097 ;
  assign n9681 = n9680 ^ n9590 ;
  assign n9589 = n1624 & n5098 ;
  assign n9682 = n9681 ^ n9589 ;
  assign n9684 = n9683 ^ n9682 ;
  assign n9586 = n9408 ^ n9330 ;
  assign n9587 = n9414 & n9586 ;
  assign n9588 = n9587 ^ n9408 ;
  assign n9685 = n9684 ^ n9588 ;
  assign n9686 = n9685 ^ x41 ;
  assign n9585 = x85 & n4474 ;
  assign n9687 = n9686 ^ n9585 ;
  assign n9584 = x87 & n4471 ;
  assign n9688 = n9687 ^ n9584 ;
  assign n9583 = n1982 & n4472 ;
  assign n9689 = n9688 ^ n9583 ;
  assign n9691 = n9690 ^ n9689 ;
  assign n9580 = n9424 ^ n9415 ;
  assign n9581 = ~n9421 & n9580 ;
  assign n9582 = n9581 ^ n9424 ;
  assign n9692 = n9691 ^ n9582 ;
  assign n9693 = n9692 ^ x38 ;
  assign n9579 = x88 & n3916 ;
  assign n9694 = n9693 ^ n9579 ;
  assign n9578 = x90 & n3919 ;
  assign n9695 = n9694 ^ n9578 ;
  assign n9577 = n2386 & n3920 ;
  assign n9696 = n9695 ^ n9577 ;
  assign n9698 = n9697 ^ n9696 ;
  assign n9702 = n9701 ^ n9698 ;
  assign n9703 = n9702 ^ x35 ;
  assign n9576 = x91 & n3375 ;
  assign n9704 = n9703 ^ n9576 ;
  assign n9575 = x93 & n3378 ;
  assign n9705 = n9704 ^ n9575 ;
  assign n9574 = n2836 & n3379 ;
  assign n9706 = n9705 ^ n9574 ;
  assign n9708 = n9707 ^ n9706 ;
  assign n9571 = n9441 ^ n9432 ;
  assign n9572 = ~n9438 & n9571 ;
  assign n9573 = n9572 ^ n9441 ;
  assign n9709 = n9708 ^ n9573 ;
  assign n9710 = n9709 ^ x32 ;
  assign n9570 = x94 & n2879 ;
  assign n9711 = n9710 ^ n9570 ;
  assign n9569 = x96 & n2882 ;
  assign n9712 = n9711 ^ n9569 ;
  assign n9568 = n2883 & n3323 ;
  assign n9713 = n9712 ^ n9568 ;
  assign n9715 = n9714 ^ n9713 ;
  assign n9719 = n9718 ^ n9715 ;
  assign n9728 = n9727 ^ n9719 ;
  assign n9732 = n9731 ^ n9728 ;
  assign n9733 = n9732 ^ x26 ;
  assign n9567 = x100 & n2018 ;
  assign n9734 = n9733 ^ n9567 ;
  assign n9566 = x102 & n2021 ;
  assign n9735 = n9734 ^ n9566 ;
  assign n9565 = n2022 & n4410 ;
  assign n9736 = n9735 ^ n9565 ;
  assign n9738 = n9737 ^ n9736 ;
  assign n9562 = n9468 ^ n9459 ;
  assign n9563 = ~n9465 & n9562 ;
  assign n9564 = n9563 ^ n9468 ;
  assign n9739 = n9738 ^ n9564 ;
  assign n9740 = n9739 ^ x23 ;
  assign n9561 = x103 & n1658 ;
  assign n9741 = n9740 ^ n9561 ;
  assign n9560 = x105 & n1661 ;
  assign n9742 = n9741 ^ n9560 ;
  assign n9559 = n1662 & ~n5023 ;
  assign n9743 = n9742 ^ n9559 ;
  assign n9745 = n9744 ^ n9743 ;
  assign n9556 = n9478 ^ n9469 ;
  assign n9557 = ~n9475 & n9556 ;
  assign n9558 = n9557 ^ n9478 ;
  assign n9746 = n9745 ^ n9558 ;
  assign n9747 = n9746 ^ x20 ;
  assign n9555 = x106 & n1327 ;
  assign n9748 = n9747 ^ n9555 ;
  assign n9554 = x108 & n1330 ;
  assign n9749 = n9748 ^ n9554 ;
  assign n9553 = n1331 & n5670 ;
  assign n9750 = n9749 ^ n9553 ;
  assign n9752 = n9751 ^ n9750 ;
  assign n9756 = n9755 ^ n9752 ;
  assign n9757 = n9756 ^ x17 ;
  assign n9552 = x109 & n1050 ;
  assign n9758 = n9757 ^ n9552 ;
  assign n9551 = x111 & n1053 ;
  assign n9759 = n9758 ^ n9551 ;
  assign n9550 = n1054 & ~n6360 ;
  assign n9760 = n9759 ^ n9550 ;
  assign n9762 = n9761 ^ n9760 ;
  assign n9547 = n9495 ^ n9486 ;
  assign n9548 = ~n9492 & n9547 ;
  assign n9549 = n9548 ^ n9495 ;
  assign n9763 = n9762 ^ n9549 ;
  assign n9764 = n9763 ^ x14 ;
  assign n9546 = x112 & n877 ;
  assign n9765 = n9764 ^ n9546 ;
  assign n9545 = x114 & n782 ;
  assign n9766 = n9765 ^ n9545 ;
  assign n9544 = n783 & ~n7092 ;
  assign n9767 = n9766 ^ n9544 ;
  assign n9769 = n9768 ^ n9767 ;
  assign n9773 = n9772 ^ n9769 ;
  assign n9774 = n9773 ^ x11 ;
  assign n9543 = x115 & n647 ;
  assign n9775 = n9774 ^ n9543 ;
  assign n9542 = x117 & ~n572 ;
  assign n9776 = n9775 ^ n9542 ;
  assign n9541 = ~n573 & ~n7850 ;
  assign n9777 = n9776 ^ n9541 ;
  assign n9779 = n9778 ^ n9777 ;
  assign n9783 = n9782 ^ n9779 ;
  assign n9802 = n9801 ^ n9783 ;
  assign n9522 = ~x124 & x125 ;
  assign n9525 = ~n9261 & n9522 ;
  assign n9520 = x125 ^ x124 ;
  assign n9523 = n9522 ^ n9520 ;
  assign n9524 = n9259 & n9523 ;
  assign n9526 = n9525 ^ n9524 ;
  assign n9528 = x126 ^ x1 ;
  assign n9527 = x126 ^ x2 ;
  assign n9529 = n9528 ^ n9527 ;
  assign n9530 = ~n9526 & n9529 ;
  assign n9531 = n9530 ^ n9528 ;
  assign n9803 = n9802 ^ n9531 ;
  assign n9536 = x2 & x124 ;
  assign n9537 = n9536 ^ x125 ;
  assign n9538 = ~n255 & n9537 ;
  assign n9532 = x125 ^ x2 ;
  assign n9533 = n9532 ^ n9531 ;
  assign n9539 = n9538 ^ n9533 ;
  assign n9540 = ~x0 & n9539 ;
  assign n9804 = n9803 ^ n9540 ;
  assign n9517 = n9245 ^ n9237 ;
  assign n9518 = ~n9514 & ~n9517 ;
  assign n9519 = n9518 ^ n9510 ;
  assign n9805 = n9804 ^ n9519 ;
  assign n9806 = n9805 ^ n9278 ;
  assign n9807 = n9806 ^ n9254 ;
  assign n9808 = n9807 ^ n9805 ;
  assign n9809 = n9516 & n9808 ;
  assign n9810 = n9809 ^ n9806 ;
  assign n9823 = n9822 ^ n9810 ;
  assign n10118 = n9822 ^ n9805 ;
  assign n10119 = ~n9810 & n10118 ;
  assign n10120 = n10119 ^ n9805 ;
  assign n10114 = n9802 ^ n9519 ;
  assign n10115 = n9804 & ~n10114 ;
  assign n10116 = n10115 ^ n9802 ;
  assign n10109 = x120 & n390 ;
  assign n10106 = x121 & n383 ;
  assign n10104 = x119 & n446 ;
  assign n10098 = x122 & n234 ;
  assign n10097 = x124 & n230 ;
  assign n10099 = n10098 ^ n10097 ;
  assign n10100 = n10099 ^ x5 ;
  assign n10095 = n8945 ^ x124 ;
  assign n10096 = n231 & n10095 ;
  assign n10101 = n10100 ^ n10096 ;
  assign n10094 = x123 & n227 ;
  assign n10102 = n10101 ^ n10094 ;
  assign n10103 = n10102 ^ x8 ;
  assign n10105 = n10104 ^ n10103 ;
  assign n10107 = n10106 ^ n10105 ;
  assign n10093 = n384 & n8962 ;
  assign n10108 = n10107 ^ n10093 ;
  assign n10110 = n10109 ^ n10108 ;
  assign n10090 = x117 & n578 ;
  assign n10083 = x114 & n788 ;
  assign n10075 = n9756 ^ n9549 ;
  assign n10076 = n9762 & n10075 ;
  assign n10077 = n10076 ^ n9756 ;
  assign n10073 = x111 & n1058 ;
  assign n10066 = x108 & n1335 ;
  assign n10058 = n9739 ^ n9558 ;
  assign n10059 = n9745 & n10058 ;
  assign n10060 = n10059 ^ n9739 ;
  assign n10056 = x105 & n1666 ;
  assign n10048 = n9732 ^ n9564 ;
  assign n10049 = n9738 & n10048 ;
  assign n10050 = n10049 ^ n9732 ;
  assign n10046 = x102 & n2014 ;
  assign n10039 = x99 & n2429 ;
  assign n10032 = x96 & n2887 ;
  assign n10024 = n9702 ^ n9573 ;
  assign n10025 = n9708 & n10024 ;
  assign n10026 = n10025 ^ n9702 ;
  assign n10022 = x93 & n3383 ;
  assign n10015 = x90 & n3924 ;
  assign n10007 = n9685 ^ n9582 ;
  assign n10008 = n9691 & n10007 ;
  assign n10009 = n10008 ^ n9685 ;
  assign n10005 = x87 & n4467 ;
  assign n9998 = x84 & n5102 ;
  assign n9991 = x81 & n5736 ;
  assign n9981 = x77 & n6677 ;
  assign n9980 = x79 & n6428 ;
  assign n9982 = n9981 ^ n9980 ;
  assign n9983 = n9982 ^ x50 ;
  assign n9979 = n1118 & n6429 ;
  assign n9984 = n9983 ^ n9979 ;
  assign n9978 = x78 & n6433 ;
  assign n9985 = n9984 ^ n9978 ;
  assign n9974 = x75 & n7179 ;
  assign n9966 = x69 & n8737 ;
  assign n9956 = x65 & n9632 ;
  assign n9955 = x66 & n9628 ;
  assign n9957 = n9956 ^ n9955 ;
  assign n9952 = ~n153 & n9630 ;
  assign n9953 = n9952 ^ x67 ;
  assign n9954 = n9046 & n9953 ;
  assign n9958 = n9957 ^ n9954 ;
  assign n9959 = n9958 ^ x62 ;
  assign n9948 = x63 ^ x62 ;
  assign n9949 = x64 & n9948 ;
  assign n9960 = n9959 ^ n9949 ;
  assign n9947 = ~n9645 & n9647 ;
  assign n9961 = n9960 ^ n9947 ;
  assign n9962 = n9961 ^ x59 ;
  assign n9946 = x68 & n8741 ;
  assign n9963 = n9962 ^ n9946 ;
  assign n9945 = x70 & n8744 ;
  assign n9964 = n9963 ^ n9945 ;
  assign n9944 = ~n436 & n8745 ;
  assign n9965 = n9964 ^ n9944 ;
  assign n9967 = n9966 ^ n9965 ;
  assign n9934 = n9380 & n9381 ;
  assign n9935 = n9934 ^ n9382 ;
  assign n9936 = n9369 & ~n9658 ;
  assign n9937 = n9935 & n9936 ;
  assign n9938 = n9934 ^ n9649 ;
  assign n9939 = n9656 ^ x59 ;
  assign n9940 = n9939 ^ n9649 ;
  assign n9941 = n9938 & n9940 ;
  assign n9942 = n9941 ^ n9649 ;
  assign n9943 = ~n9937 & ~n9942 ;
  assign n9968 = n9967 ^ n9943 ;
  assign n9924 = x71 & n7935 ;
  assign n9923 = x73 & n7938 ;
  assign n9925 = n9924 ^ n9923 ;
  assign n9926 = n9925 ^ x56 ;
  assign n9922 = n633 & n7939 ;
  assign n9927 = n9926 ^ n9922 ;
  assign n9921 = x72 & n7931 ;
  assign n9928 = n9927 ^ n9921 ;
  assign n9929 = n9928 ^ n9670 ;
  assign n9930 = n9929 ^ n9661 ;
  assign n9931 = n9930 ^ n9928 ;
  assign n9932 = ~n9667 & n9931 ;
  assign n9933 = n9932 ^ n9929 ;
  assign n9969 = n9968 ^ n9933 ;
  assign n9970 = n9969 ^ x53 ;
  assign n9920 = x74 & n7171 ;
  assign n9971 = n9970 ^ n9920 ;
  assign n9919 = x76 & n7174 ;
  assign n9972 = n9971 ^ n9919 ;
  assign n9918 = ~n853 & n7175 ;
  assign n9973 = n9972 ^ n9918 ;
  assign n9975 = n9974 ^ n9973 ;
  assign n9915 = n9671 ^ n9619 ;
  assign n9916 = n9624 & n9915 ;
  assign n9917 = n9916 ^ n9619 ;
  assign n9976 = n9975 ^ n9917 ;
  assign n9911 = n9672 ^ n9602 ;
  assign n9912 = n9602 ^ n9594 ;
  assign n9913 = n9911 & ~n9912 ;
  assign n9914 = n9913 ^ n9672 ;
  assign n9977 = n9976 ^ n9914 ;
  assign n9986 = n9985 ^ n9977 ;
  assign n9987 = n9986 ^ x47 ;
  assign n9910 = x80 & n5965 ;
  assign n9988 = n9987 ^ n9910 ;
  assign n9909 = x82 & n5729 ;
  assign n9989 = n9988 ^ n9909 ;
  assign n9908 = n1411 & n5730 ;
  assign n9990 = n9989 ^ n9908 ;
  assign n9992 = n9991 ^ n9990 ;
  assign n9905 = n9677 ^ n9610 ;
  assign n9906 = ~n9674 & n9905 ;
  assign n9907 = n9906 ^ n9677 ;
  assign n9993 = n9992 ^ n9907 ;
  assign n9994 = n9993 ^ x44 ;
  assign n9904 = x83 & n5094 ;
  assign n9995 = n9994 ^ n9904 ;
  assign n9903 = x85 & n5097 ;
  assign n9996 = n9995 ^ n9903 ;
  assign n9902 = n1743 & n5098 ;
  assign n9997 = n9996 ^ n9902 ;
  assign n9999 = n9998 ^ n9997 ;
  assign n9899 = n9678 ^ n9588 ;
  assign n9900 = n9684 & n9899 ;
  assign n9901 = n9900 ^ n9678 ;
  assign n10000 = n9999 ^ n9901 ;
  assign n10001 = n10000 ^ x41 ;
  assign n9898 = x86 & n4474 ;
  assign n10002 = n10001 ^ n9898 ;
  assign n9897 = x88 & n4471 ;
  assign n10003 = n10002 ^ n9897 ;
  assign n9896 = n2119 & n4472 ;
  assign n10004 = n10003 ^ n9896 ;
  assign n10006 = n10005 ^ n10004 ;
  assign n10010 = n10009 ^ n10006 ;
  assign n10011 = n10010 ^ x38 ;
  assign n9895 = x89 & n3916 ;
  assign n10012 = n10011 ^ n9895 ;
  assign n9894 = x91 & n3919 ;
  assign n10013 = n10012 ^ n9894 ;
  assign n9893 = n2542 & n3920 ;
  assign n10014 = n10013 ^ n9893 ;
  assign n10016 = n10015 ^ n10014 ;
  assign n9890 = n9701 ^ n9692 ;
  assign n9891 = ~n9698 & n9890 ;
  assign n9892 = n9891 ^ n9701 ;
  assign n10017 = n10016 ^ n9892 ;
  assign n10018 = n10017 ^ x35 ;
  assign n9889 = x92 & n3375 ;
  assign n10019 = n10018 ^ n9889 ;
  assign n9888 = x94 & n3378 ;
  assign n10020 = n10019 ^ n9888 ;
  assign n9887 = n2997 & n3379 ;
  assign n10021 = n10020 ^ n9887 ;
  assign n10023 = n10022 ^ n10021 ;
  assign n10027 = n10026 ^ n10023 ;
  assign n10028 = n10027 ^ x32 ;
  assign n9886 = x95 & n2879 ;
  assign n10029 = n10028 ^ n9886 ;
  assign n9885 = x97 & n2882 ;
  assign n10030 = n10029 ^ n9885 ;
  assign n9884 = n2883 & n3494 ;
  assign n10031 = n10030 ^ n9884 ;
  assign n10033 = n10032 ^ n10031 ;
  assign n9881 = n9718 ^ n9709 ;
  assign n9882 = ~n9715 & n9881 ;
  assign n9883 = n9882 ^ n9718 ;
  assign n10034 = n10033 ^ n9883 ;
  assign n10035 = n10034 ^ x29 ;
  assign n9880 = x98 & n2581 ;
  assign n10036 = n10035 ^ n9880 ;
  assign n9879 = x100 & n2422 ;
  assign n10037 = n10036 ^ n9879 ;
  assign n9878 = n2423 & n4034 ;
  assign n10038 = n10037 ^ n9878 ;
  assign n10040 = n10039 ^ n10038 ;
  assign n9875 = n9731 ^ n9727 ;
  assign n9876 = ~n9728 & n9875 ;
  assign n9877 = n9876 ^ n9731 ;
  assign n10041 = n10040 ^ n9877 ;
  assign n10042 = n10041 ^ x26 ;
  assign n9874 = x101 & n2018 ;
  assign n10043 = n10042 ^ n9874 ;
  assign n9873 = x103 & n2021 ;
  assign n10044 = n10043 ^ n9873 ;
  assign n9872 = n2022 & ~n4615 ;
  assign n10045 = n10044 ^ n9872 ;
  assign n10047 = n10046 ^ n10045 ;
  assign n10051 = n10050 ^ n10047 ;
  assign n10052 = n10051 ^ x23 ;
  assign n9871 = x104 & n1658 ;
  assign n10053 = n10052 ^ n9871 ;
  assign n9870 = x106 & n1661 ;
  assign n10054 = n10053 ^ n9870 ;
  assign n9869 = n1662 & ~n5240 ;
  assign n10055 = n10054 ^ n9869 ;
  assign n10057 = n10056 ^ n10055 ;
  assign n10061 = n10060 ^ n10057 ;
  assign n10062 = n10061 ^ x20 ;
  assign n9868 = x107 & n1327 ;
  assign n10063 = n10062 ^ n9868 ;
  assign n9867 = x109 & n1330 ;
  assign n10064 = n10063 ^ n9867 ;
  assign n9866 = n1331 & n5902 ;
  assign n10065 = n10064 ^ n9866 ;
  assign n10067 = n10066 ^ n10065 ;
  assign n9863 = n9755 ^ n9746 ;
  assign n9864 = ~n9752 & n9863 ;
  assign n9865 = n9864 ^ n9755 ;
  assign n10068 = n10067 ^ n9865 ;
  assign n10069 = n10068 ^ x17 ;
  assign n9862 = x110 & n1050 ;
  assign n10070 = n10069 ^ n9862 ;
  assign n9861 = x112 & n1053 ;
  assign n10071 = n10070 ^ n9861 ;
  assign n9860 = n1054 & ~n6600 ;
  assign n10072 = n10071 ^ n9860 ;
  assign n10074 = n10073 ^ n10072 ;
  assign n10078 = n10077 ^ n10074 ;
  assign n10079 = n10078 ^ x14 ;
  assign n9859 = x113 & n877 ;
  assign n10080 = n10079 ^ n9859 ;
  assign n9858 = x115 & n782 ;
  assign n10081 = n10080 ^ n9858 ;
  assign n9857 = n783 & ~n7343 ;
  assign n10082 = n10081 ^ n9857 ;
  assign n10084 = n10083 ^ n10082 ;
  assign n9854 = n9772 ^ n9763 ;
  assign n9855 = ~n9769 & n9854 ;
  assign n9856 = n9855 ^ n9772 ;
  assign n10085 = n10084 ^ n9856 ;
  assign n10086 = n10085 ^ x11 ;
  assign n9853 = x116 & n647 ;
  assign n10087 = n10086 ^ n9853 ;
  assign n9852 = x118 & ~n572 ;
  assign n10088 = n10087 ^ n9852 ;
  assign n9851 = ~n573 & ~n8123 ;
  assign n10089 = n10088 ^ n9851 ;
  assign n10091 = n10090 ^ n10089 ;
  assign n9848 = n9782 ^ n9773 ;
  assign n9849 = ~n9779 & n9848 ;
  assign n9850 = n9849 ^ n9782 ;
  assign n10092 = n10091 ^ n9850 ;
  assign n10111 = n10110 ^ n10092 ;
  assign n9842 = x2 & x125 ;
  assign n9843 = n9842 ^ x126 ;
  assign n9844 = ~x1 & n9843 ;
  assign n9828 = x125 & ~x126 ;
  assign n9831 = ~n9525 & n9828 ;
  assign n9827 = x126 ^ x125 ;
  assign n9829 = n9828 ^ n9827 ;
  assign n9830 = ~n9524 & n9829 ;
  assign n9832 = n9831 ^ n9830 ;
  assign n9834 = x127 ^ x1 ;
  assign n9833 = x127 ^ x2 ;
  assign n9835 = n9834 ^ n9833 ;
  assign n9836 = ~n9832 & n9835 ;
  assign n9837 = n9836 ^ n9834 ;
  assign n9839 = n9837 ^ n9527 ;
  assign n9845 = n9844 ^ n9839 ;
  assign n9846 = ~x0 & n9845 ;
  assign n9847 = n9846 ^ n9837 ;
  assign n10112 = n10111 ^ n9847 ;
  assign n9824 = n9793 ^ n9783 ;
  assign n9825 = n9801 & n9824 ;
  assign n9826 = n9825 ^ n9793 ;
  assign n10113 = n10112 ^ n9826 ;
  assign n10117 = n10116 ^ n10113 ;
  assign n10121 = n10120 ^ n10117 ;
  assign n10414 = x121 & n390 ;
  assign n10411 = x122 & n383 ;
  assign n10409 = x120 & n446 ;
  assign n10403 = x123 & n234 ;
  assign n10402 = x125 & n230 ;
  assign n10404 = n10403 ^ n10402 ;
  assign n10405 = n10404 ^ x5 ;
  assign n10400 = n9520 ^ n9261 ;
  assign n10401 = n231 & n10400 ;
  assign n10406 = n10405 ^ n10401 ;
  assign n10399 = x124 & n227 ;
  assign n10407 = n10406 ^ n10399 ;
  assign n10408 = n10407 ^ x8 ;
  assign n10410 = n10409 ^ n10408 ;
  assign n10412 = n10411 ^ n10410 ;
  assign n10398 = n384 & ~n9247 ;
  assign n10413 = n10412 ^ n10398 ;
  assign n10415 = n10414 ^ n10413 ;
  assign n10394 = n10085 ^ n9850 ;
  assign n10395 = ~n10091 & ~n10394 ;
  assign n10396 = n10395 ^ n10085 ;
  assign n10392 = x118 & n578 ;
  assign n10384 = n10078 ^ n9856 ;
  assign n10385 = ~n10084 & ~n10384 ;
  assign n10386 = n10385 ^ n10078 ;
  assign n10382 = x115 & n788 ;
  assign n10375 = x112 & n1058 ;
  assign n10367 = n10061 ^ n9865 ;
  assign n10368 = ~n10067 & ~n10367 ;
  assign n10369 = n10368 ^ n10061 ;
  assign n10365 = x109 & n1335 ;
  assign n10358 = x106 & n1666 ;
  assign n10351 = x103 & n2014 ;
  assign n10343 = n10034 ^ n9877 ;
  assign n10344 = ~n10040 & ~n10343 ;
  assign n10345 = n10344 ^ n10034 ;
  assign n10341 = x100 & n2429 ;
  assign n10333 = n10027 ^ n9883 ;
  assign n10334 = ~n10033 & ~n10333 ;
  assign n10335 = n10334 ^ n10027 ;
  assign n10331 = x97 & n2887 ;
  assign n10324 = x94 & n3383 ;
  assign n10316 = n10010 ^ n9892 ;
  assign n10317 = ~n10016 & ~n10316 ;
  assign n10318 = n10317 ^ n10010 ;
  assign n10314 = x91 & n3924 ;
  assign n10307 = x88 & n4467 ;
  assign n10300 = x85 & n5102 ;
  assign n10292 = n9986 ^ n9907 ;
  assign n10293 = ~n9992 & ~n10292 ;
  assign n10294 = n10293 ^ n9986 ;
  assign n10290 = x82 & n5736 ;
  assign n10283 = x79 & n6433 ;
  assign n10275 = x73 & n7931 ;
  assign n10267 = n9961 ^ n9943 ;
  assign n10268 = n9967 & ~n10267 ;
  assign n10269 = n10268 ^ n9961 ;
  assign n10265 = x70 & n8737 ;
  assign n10256 = ~x63 & x64 ;
  assign n330 = x65 ^ x64 ;
  assign n10257 = n10256 ^ n330 ;
  assign n10258 = ~n9948 & n10257 ;
  assign n10246 = x66 & n9632 ;
  assign n10245 = x68 & n9635 ;
  assign n10247 = n10246 ^ n10245 ;
  assign n10248 = n10247 ^ x62 ;
  assign n10244 = ~n340 & n9636 ;
  assign n10249 = n10248 ^ n10244 ;
  assign n10243 = x67 & n9628 ;
  assign n10250 = n10249 ^ n10243 ;
  assign n10251 = n10250 ^ x65 ;
  assign n10259 = n10258 ^ n10251 ;
  assign n10236 = x62 & n9949 ;
  assign n10235 = n9958 ^ n9949 ;
  assign n10237 = n10236 ^ n10235 ;
  assign n10238 = n10237 ^ n9947 ;
  assign n10239 = n9949 ^ n9947 ;
  assign n10240 = ~n10236 & ~n10239 ;
  assign n10241 = ~n10238 & n10240 ;
  assign n10242 = n10241 ^ n10237 ;
  assign n10260 = n10259 ^ n10242 ;
  assign n10261 = n10260 ^ x59 ;
  assign n10234 = x69 & n8741 ;
  assign n10262 = n10261 ^ n10234 ;
  assign n10233 = x71 & n8744 ;
  assign n10263 = n10262 ^ n10233 ;
  assign n10232 = ~n493 & n8745 ;
  assign n10264 = n10263 ^ n10232 ;
  assign n10266 = n10265 ^ n10264 ;
  assign n10270 = n10269 ^ n10266 ;
  assign n10271 = n10270 ^ x56 ;
  assign n10231 = x72 & n7935 ;
  assign n10272 = n10271 ^ n10231 ;
  assign n10230 = x74 & n7938 ;
  assign n10273 = n10272 ^ n10230 ;
  assign n10229 = n699 & n7939 ;
  assign n10274 = n10273 ^ n10229 ;
  assign n10276 = n10275 ^ n10274 ;
  assign n10226 = n9968 ^ n9928 ;
  assign n10227 = n9933 & ~n10226 ;
  assign n10228 = n10227 ^ n9928 ;
  assign n10277 = n10276 ^ n10228 ;
  assign n10216 = x75 & n7171 ;
  assign n10215 = x77 & n7174 ;
  assign n10217 = n10216 ^ n10215 ;
  assign n10218 = n10217 ^ x53 ;
  assign n10214 = ~n939 & n7175 ;
  assign n10219 = n10218 ^ n10214 ;
  assign n10213 = x76 & n7179 ;
  assign n10220 = n10219 ^ n10213 ;
  assign n10221 = n10220 ^ n9969 ;
  assign n10222 = n10221 ^ n9917 ;
  assign n10223 = n10222 ^ n10220 ;
  assign n10224 = ~n9975 & ~n10223 ;
  assign n10225 = n10224 ^ n10221 ;
  assign n10278 = n10277 ^ n10225 ;
  assign n10279 = n10278 ^ x50 ;
  assign n10212 = x78 & n6677 ;
  assign n10280 = n10279 ^ n10212 ;
  assign n10211 = x80 & n6428 ;
  assign n10281 = n10280 ^ n10211 ;
  assign n10210 = n1206 & n6429 ;
  assign n10282 = n10281 ^ n10210 ;
  assign n10284 = n10283 ^ n10282 ;
  assign n10207 = n9985 ^ n9914 ;
  assign n10208 = n9977 & n10207 ;
  assign n10209 = n10208 ^ n9985 ;
  assign n10285 = n10284 ^ n10209 ;
  assign n10286 = n10285 ^ x47 ;
  assign n10206 = x81 & n5965 ;
  assign n10287 = n10286 ^ n10206 ;
  assign n10205 = x83 & n5729 ;
  assign n10288 = n10287 ^ n10205 ;
  assign n10204 = n1512 & n5730 ;
  assign n10289 = n10288 ^ n10204 ;
  assign n10291 = n10290 ^ n10289 ;
  assign n10295 = n10294 ^ n10291 ;
  assign n10296 = n10295 ^ x44 ;
  assign n10203 = x84 & n5094 ;
  assign n10297 = n10296 ^ n10203 ;
  assign n10202 = x86 & n5097 ;
  assign n10298 = n10297 ^ n10202 ;
  assign n10201 = n1857 & n5098 ;
  assign n10299 = n10298 ^ n10201 ;
  assign n10301 = n10300 ^ n10299 ;
  assign n10198 = n9993 ^ n9901 ;
  assign n10199 = ~n9999 & ~n10198 ;
  assign n10200 = n10199 ^ n9993 ;
  assign n10302 = n10301 ^ n10200 ;
  assign n10303 = n10302 ^ x41 ;
  assign n10197 = x87 & n4474 ;
  assign n10304 = n10303 ^ n10197 ;
  assign n10196 = x89 & n4471 ;
  assign n10305 = n10304 ^ n10196 ;
  assign n10195 = n2249 & n4472 ;
  assign n10306 = n10305 ^ n10195 ;
  assign n10308 = n10307 ^ n10306 ;
  assign n10192 = n10009 ^ n10000 ;
  assign n10193 = n10006 & ~n10192 ;
  assign n10194 = n10193 ^ n10009 ;
  assign n10309 = n10308 ^ n10194 ;
  assign n10310 = n10309 ^ x38 ;
  assign n10191 = x90 & n3916 ;
  assign n10311 = n10310 ^ n10191 ;
  assign n10190 = x92 & n3919 ;
  assign n10312 = n10311 ^ n10190 ;
  assign n10189 = n2684 & n3920 ;
  assign n10313 = n10312 ^ n10189 ;
  assign n10315 = n10314 ^ n10313 ;
  assign n10319 = n10318 ^ n10315 ;
  assign n10320 = n10319 ^ x35 ;
  assign n10188 = x93 & n3375 ;
  assign n10321 = n10320 ^ n10188 ;
  assign n10187 = x95 & n3378 ;
  assign n10322 = n10321 ^ n10187 ;
  assign n10186 = n3159 & n3379 ;
  assign n10323 = n10322 ^ n10186 ;
  assign n10325 = n10324 ^ n10323 ;
  assign n10183 = n10026 ^ n10017 ;
  assign n10184 = n10023 & ~n10183 ;
  assign n10185 = n10184 ^ n10026 ;
  assign n10326 = n10325 ^ n10185 ;
  assign n10327 = n10326 ^ x32 ;
  assign n10182 = x96 & n2879 ;
  assign n10328 = n10327 ^ n10182 ;
  assign n10181 = x98 & n2882 ;
  assign n10329 = n10328 ^ n10181 ;
  assign n10180 = n2883 & n3660 ;
  assign n10330 = n10329 ^ n10180 ;
  assign n10332 = n10331 ^ n10330 ;
  assign n10336 = n10335 ^ n10332 ;
  assign n10337 = n10336 ^ x29 ;
  assign n10179 = x99 & n2581 ;
  assign n10338 = n10337 ^ n10179 ;
  assign n10178 = x101 & n2422 ;
  assign n10339 = n10338 ^ n10178 ;
  assign n10177 = n2423 & n4215 ;
  assign n10340 = n10339 ^ n10177 ;
  assign n10342 = n10341 ^ n10340 ;
  assign n10346 = n10345 ^ n10342 ;
  assign n10347 = n10346 ^ x26 ;
  assign n10176 = x102 & n2018 ;
  assign n10348 = n10347 ^ n10176 ;
  assign n10175 = x104 & n2021 ;
  assign n10349 = n10348 ^ n10175 ;
  assign n10174 = n2022 & ~n4814 ;
  assign n10350 = n10349 ^ n10174 ;
  assign n10352 = n10351 ^ n10350 ;
  assign n10171 = n10050 ^ n10041 ;
  assign n10172 = n10047 & ~n10171 ;
  assign n10173 = n10172 ^ n10050 ;
  assign n10353 = n10352 ^ n10173 ;
  assign n10354 = n10353 ^ x23 ;
  assign n10170 = x105 & n1658 ;
  assign n10355 = n10354 ^ n10170 ;
  assign n10169 = x107 & n1661 ;
  assign n10356 = n10355 ^ n10169 ;
  assign n10168 = n1662 & ~n5448 ;
  assign n10357 = n10356 ^ n10168 ;
  assign n10359 = n10358 ^ n10357 ;
  assign n10165 = n10060 ^ n10051 ;
  assign n10166 = n10057 & ~n10165 ;
  assign n10167 = n10166 ^ n10060 ;
  assign n10360 = n10359 ^ n10167 ;
  assign n10361 = n10360 ^ x20 ;
  assign n10164 = x108 & n1327 ;
  assign n10362 = n10361 ^ n10164 ;
  assign n10163 = x110 & n1330 ;
  assign n10363 = n10362 ^ n10163 ;
  assign n10162 = n1331 & n6129 ;
  assign n10364 = n10363 ^ n10162 ;
  assign n10366 = n10365 ^ n10364 ;
  assign n10370 = n10369 ^ n10366 ;
  assign n10371 = n10370 ^ x17 ;
  assign n10161 = x111 & n1050 ;
  assign n10372 = n10371 ^ n10161 ;
  assign n10160 = x113 & n1053 ;
  assign n10373 = n10372 ^ n10160 ;
  assign n10159 = n1054 & ~n6839 ;
  assign n10374 = n10373 ^ n10159 ;
  assign n10376 = n10375 ^ n10374 ;
  assign n10156 = n10077 ^ n10068 ;
  assign n10157 = n10074 & ~n10156 ;
  assign n10158 = n10157 ^ n10077 ;
  assign n10377 = n10376 ^ n10158 ;
  assign n10378 = n10377 ^ x14 ;
  assign n10155 = x114 & n877 ;
  assign n10379 = n10378 ^ n10155 ;
  assign n10154 = x116 & n782 ;
  assign n10380 = n10379 ^ n10154 ;
  assign n10153 = n783 & ~n7588 ;
  assign n10381 = n10380 ^ n10153 ;
  assign n10383 = n10382 ^ n10381 ;
  assign n10387 = n10386 ^ n10383 ;
  assign n10388 = n10387 ^ x11 ;
  assign n10152 = x117 & n647 ;
  assign n10389 = n10388 ^ n10152 ;
  assign n10151 = x119 & ~n572 ;
  assign n10390 = n10389 ^ n10151 ;
  assign n10150 = ~n573 & n8394 ;
  assign n10391 = n10390 ^ n10150 ;
  assign n10393 = n10392 ^ n10391 ;
  assign n10397 = n10396 ^ n10393 ;
  assign n10416 = n10415 ^ n10397 ;
  assign n10128 = x2 & ~x127 ;
  assign n10135 = ~x126 & x127 ;
  assign n10138 = ~n9831 & n10135 ;
  assign n10130 = x127 ^ x126 ;
  assign n10136 = n10135 ^ n10130 ;
  assign n10137 = ~n9830 & n10136 ;
  assign n10139 = n10138 ^ n10137 ;
  assign n10140 = n10129 & ~n10139 ;
  assign n10141 = n10140 ^ x1 ;
  assign n10132 = ~x2 & ~n10130 ;
  assign n10133 = n10132 ^ x126 ;
  assign n10134 = n10129 & ~n10133 ;
  assign n10142 = n10141 ^ n10134 ;
  assign n10143 = ~x0 & n10142 ;
  assign n10144 = n10143 ^ n10141 ;
  assign n10145 = n10128 & ~n10144 ;
  assign n10147 = ~x1 & x126 ;
  assign n10148 = n10145 & n10147 ;
  assign n10146 = n10145 ^ n10144 ;
  assign n10149 = n10148 ^ n10146 ;
  assign n10417 = n10416 ^ n10149 ;
  assign n10125 = n10102 ^ n10092 ;
  assign n10126 = n10110 & ~n10125 ;
  assign n10127 = n10126 ^ n10102 ;
  assign n10418 = n10417 ^ n10127 ;
  assign n10419 = n10418 ^ n9847 ;
  assign n10420 = n10419 ^ n10418 ;
  assign n10421 = n10420 ^ n9826 ;
  assign n10422 = ~n10112 & n10421 ;
  assign n10423 = n10422 ^ n10419 ;
  assign n10122 = n10120 ^ n10116 ;
  assign n10123 = n10117 & ~n10122 ;
  assign n10124 = n10123 ^ n10120 ;
  assign n10424 = n10423 ^ n10124 ;
  assign n10708 = n10418 ^ n10124 ;
  assign n10709 = n10423 & ~n10708 ;
  assign n10710 = n10709 ^ n10418 ;
  assign n10699 = x125 & n227 ;
  assign n10692 = x119 & n578 ;
  assign n10689 = x120 & ~n572 ;
  assign n10687 = x118 & n647 ;
  assign n10681 = x121 & n446 ;
  assign n10680 = x123 & n383 ;
  assign n10682 = n10681 ^ n10680 ;
  assign n10683 = n10682 ^ x8 ;
  assign n10679 = n384 & ~n9786 ;
  assign n10684 = n10683 ^ n10679 ;
  assign n10678 = x122 & n390 ;
  assign n10685 = n10684 ^ n10678 ;
  assign n10686 = n10685 ^ x11 ;
  assign n10688 = n10687 ^ n10686 ;
  assign n10690 = n10689 ^ n10688 ;
  assign n10677 = ~n573 & n8891 ;
  assign n10691 = n10690 ^ n10677 ;
  assign n10693 = n10692 ^ n10691 ;
  assign n10674 = x116 & n788 ;
  assign n10666 = n10370 ^ n10158 ;
  assign n10667 = n10376 & n10666 ;
  assign n10668 = n10667 ^ n10370 ;
  assign n10664 = x113 & n1058 ;
  assign n10657 = x110 & n1335 ;
  assign n10649 = n10353 ^ n10167 ;
  assign n10650 = ~n10359 & ~n10649 ;
  assign n10651 = n10650 ^ n10353 ;
  assign n10647 = x107 & n1666 ;
  assign n10639 = n10346 ^ n10173 ;
  assign n10640 = ~n10352 & ~n10639 ;
  assign n10641 = n10640 ^ n10346 ;
  assign n10637 = x104 & n2014 ;
  assign n10630 = x101 & n2429 ;
  assign n10623 = x98 & n2887 ;
  assign n10615 = n10319 ^ n10185 ;
  assign n10616 = ~n10325 & ~n10615 ;
  assign n10617 = n10616 ^ n10319 ;
  assign n10613 = x95 & n3383 ;
  assign n10606 = x92 & n3924 ;
  assign n10598 = n10302 ^ n10194 ;
  assign n10599 = n10308 & n10598 ;
  assign n10600 = n10599 ^ n10302 ;
  assign n10596 = x89 & n4467 ;
  assign n10589 = x86 & n5102 ;
  assign n10582 = x83 & n5736 ;
  assign n10575 = x80 & n6433 ;
  assign n10566 = x71 & n8737 ;
  assign n10556 = x67 & n9632 ;
  assign n10555 = x69 & n9635 ;
  assign n10557 = n10556 ^ n10555 ;
  assign n10558 = n10557 ^ x62 ;
  assign n10554 = ~n375 & n9636 ;
  assign n10559 = n10558 ^ n10554 ;
  assign n10553 = x68 & n9628 ;
  assign n10560 = n10559 ^ n10553 ;
  assign n10549 = x63 & x65 ;
  assign n10550 = n10549 ^ x66 ;
  assign n10551 = ~n9948 & n10550 ;
  assign n10540 = n10250 ^ n10242 ;
  assign n10541 = n10259 & ~n10540 ;
  assign n10542 = n10541 ^ n10250 ;
  assign n10543 = n10542 ^ x66 ;
  assign n10552 = n10551 ^ n10543 ;
  assign n10561 = n10560 ^ n10552 ;
  assign n10562 = n10561 ^ x59 ;
  assign n10539 = x70 & n8741 ;
  assign n10563 = n10562 ^ n10539 ;
  assign n10538 = x72 & n8744 ;
  assign n10564 = n10563 ^ n10538 ;
  assign n10537 = n556 & n8745 ;
  assign n10565 = n10564 ^ n10537 ;
  assign n10567 = n10566 ^ n10565 ;
  assign n10534 = n10269 ^ n10260 ;
  assign n10535 = n10266 & ~n10534 ;
  assign n10536 = n10535 ^ n10269 ;
  assign n10568 = n10567 ^ n10536 ;
  assign n10524 = x73 & n7935 ;
  assign n10523 = x75 & n7938 ;
  assign n10525 = n10524 ^ n10523 ;
  assign n10526 = n10525 ^ x56 ;
  assign n10522 = ~n774 & n7939 ;
  assign n10527 = n10526 ^ n10522 ;
  assign n10521 = x74 & n7931 ;
  assign n10528 = n10527 ^ n10521 ;
  assign n10529 = n10528 ^ n10270 ;
  assign n10530 = n10529 ^ n10228 ;
  assign n10531 = n10530 ^ n10528 ;
  assign n10532 = ~n10276 & ~n10531 ;
  assign n10533 = n10532 ^ n10529 ;
  assign n10569 = n10568 ^ n10533 ;
  assign n10511 = x76 & n7171 ;
  assign n10510 = x78 & n7174 ;
  assign n10512 = n10511 ^ n10510 ;
  assign n10513 = n10512 ^ x53 ;
  assign n10509 = ~n1025 & n7175 ;
  assign n10514 = n10513 ^ n10509 ;
  assign n10508 = x77 & n7179 ;
  assign n10515 = n10514 ^ n10508 ;
  assign n10517 = n10515 ^ n10220 ;
  assign n10516 = n10515 ^ n10277 ;
  assign n10518 = n10517 ^ n10516 ;
  assign n10519 = ~n10225 & ~n10518 ;
  assign n10520 = n10519 ^ n10517 ;
  assign n10570 = n10569 ^ n10520 ;
  assign n10571 = n10570 ^ x50 ;
  assign n10507 = x79 & n6677 ;
  assign n10572 = n10571 ^ n10507 ;
  assign n10506 = x81 & n6428 ;
  assign n10573 = n10572 ^ n10506 ;
  assign n10505 = n1305 & n6429 ;
  assign n10574 = n10573 ^ n10505 ;
  assign n10576 = n10575 ^ n10574 ;
  assign n10502 = n10278 ^ n10209 ;
  assign n10503 = n10284 & n10502 ;
  assign n10504 = n10503 ^ n10278 ;
  assign n10577 = n10576 ^ n10504 ;
  assign n10578 = n10577 ^ x47 ;
  assign n10501 = x82 & n5965 ;
  assign n10579 = n10578 ^ n10501 ;
  assign n10500 = x84 & n5729 ;
  assign n10580 = n10579 ^ n10500 ;
  assign n10499 = n1624 & n5730 ;
  assign n10581 = n10580 ^ n10499 ;
  assign n10583 = n10582 ^ n10581 ;
  assign n10496 = n10294 ^ n10285 ;
  assign n10497 = ~n10291 & ~n10496 ;
  assign n10498 = n10497 ^ n10294 ;
  assign n10584 = n10583 ^ n10498 ;
  assign n10585 = n10584 ^ x44 ;
  assign n10495 = x85 & n5094 ;
  assign n10586 = n10585 ^ n10495 ;
  assign n10494 = x87 & n5097 ;
  assign n10587 = n10586 ^ n10494 ;
  assign n10493 = n1982 & n5098 ;
  assign n10588 = n10587 ^ n10493 ;
  assign n10590 = n10589 ^ n10588 ;
  assign n10490 = n10295 ^ n10200 ;
  assign n10491 = ~n10301 & n10490 ;
  assign n10492 = n10491 ^ n10295 ;
  assign n10591 = n10590 ^ n10492 ;
  assign n10592 = n10591 ^ x41 ;
  assign n10489 = x88 & n4474 ;
  assign n10593 = n10592 ^ n10489 ;
  assign n10488 = x90 & n4471 ;
  assign n10594 = n10593 ^ n10488 ;
  assign n10487 = n2386 & n4472 ;
  assign n10595 = n10594 ^ n10487 ;
  assign n10597 = n10596 ^ n10595 ;
  assign n10601 = n10600 ^ n10597 ;
  assign n10602 = n10601 ^ x38 ;
  assign n10486 = x91 & n3916 ;
  assign n10603 = n10602 ^ n10486 ;
  assign n10485 = x93 & n3919 ;
  assign n10604 = n10603 ^ n10485 ;
  assign n10484 = n2836 & n3920 ;
  assign n10605 = n10604 ^ n10484 ;
  assign n10607 = n10606 ^ n10605 ;
  assign n10481 = n10318 ^ n10309 ;
  assign n10482 = ~n10315 & ~n10481 ;
  assign n10483 = n10482 ^ n10318 ;
  assign n10608 = n10607 ^ n10483 ;
  assign n10609 = n10608 ^ x35 ;
  assign n10480 = x94 & n3375 ;
  assign n10610 = n10609 ^ n10480 ;
  assign n10479 = x96 & n3378 ;
  assign n10611 = n10610 ^ n10479 ;
  assign n10478 = n3323 & n3379 ;
  assign n10612 = n10611 ^ n10478 ;
  assign n10614 = n10613 ^ n10612 ;
  assign n10618 = n10617 ^ n10614 ;
  assign n10619 = n10618 ^ x32 ;
  assign n10477 = x97 & n2879 ;
  assign n10620 = n10619 ^ n10477 ;
  assign n10476 = x99 & n2882 ;
  assign n10621 = n10620 ^ n10476 ;
  assign n10475 = n2883 & n3843 ;
  assign n10622 = n10621 ^ n10475 ;
  assign n10624 = n10623 ^ n10622 ;
  assign n10472 = n10335 ^ n10326 ;
  assign n10473 = n10332 & n10472 ;
  assign n10474 = n10473 ^ n10335 ;
  assign n10625 = n10624 ^ n10474 ;
  assign n10626 = n10625 ^ x29 ;
  assign n10471 = x100 & n2581 ;
  assign n10627 = n10626 ^ n10471 ;
  assign n10470 = x102 & n2422 ;
  assign n10628 = n10627 ^ n10470 ;
  assign n10469 = n2423 & n4410 ;
  assign n10629 = n10628 ^ n10469 ;
  assign n10631 = n10630 ^ n10629 ;
  assign n10466 = n10345 ^ n10336 ;
  assign n10467 = ~n10342 & ~n10466 ;
  assign n10468 = n10467 ^ n10345 ;
  assign n10632 = n10631 ^ n10468 ;
  assign n10633 = n10632 ^ x26 ;
  assign n10465 = x103 & n2018 ;
  assign n10634 = n10633 ^ n10465 ;
  assign n10464 = x105 & n2021 ;
  assign n10635 = n10634 ^ n10464 ;
  assign n10463 = n2022 & ~n5023 ;
  assign n10636 = n10635 ^ n10463 ;
  assign n10638 = n10637 ^ n10636 ;
  assign n10642 = n10641 ^ n10638 ;
  assign n10643 = n10642 ^ x23 ;
  assign n10462 = x106 & n1658 ;
  assign n10644 = n10643 ^ n10462 ;
  assign n10461 = x108 & n1661 ;
  assign n10645 = n10644 ^ n10461 ;
  assign n10460 = n1662 & n5670 ;
  assign n10646 = n10645 ^ n10460 ;
  assign n10648 = n10647 ^ n10646 ;
  assign n10652 = n10651 ^ n10648 ;
  assign n10653 = n10652 ^ x20 ;
  assign n10459 = x109 & n1327 ;
  assign n10654 = n10653 ^ n10459 ;
  assign n10458 = x111 & n1330 ;
  assign n10655 = n10654 ^ n10458 ;
  assign n10457 = n1331 & ~n6360 ;
  assign n10656 = n10655 ^ n10457 ;
  assign n10658 = n10657 ^ n10656 ;
  assign n10454 = n10369 ^ n10360 ;
  assign n10455 = n10366 & n10454 ;
  assign n10456 = n10455 ^ n10369 ;
  assign n10659 = n10658 ^ n10456 ;
  assign n10660 = n10659 ^ x17 ;
  assign n10453 = x112 & n1050 ;
  assign n10661 = n10660 ^ n10453 ;
  assign n10452 = x114 & n1053 ;
  assign n10662 = n10661 ^ n10452 ;
  assign n10451 = n1054 & ~n7092 ;
  assign n10663 = n10662 ^ n10451 ;
  assign n10665 = n10664 ^ n10663 ;
  assign n10669 = n10668 ^ n10665 ;
  assign n10670 = n10669 ^ x14 ;
  assign n10450 = x115 & n877 ;
  assign n10671 = n10670 ^ n10450 ;
  assign n10449 = x117 & n782 ;
  assign n10672 = n10671 ^ n10449 ;
  assign n10448 = n783 & ~n7850 ;
  assign n10673 = n10672 ^ n10448 ;
  assign n10675 = n10674 ^ n10673 ;
  assign n10445 = n10386 ^ n10377 ;
  assign n10446 = ~n10383 & ~n10445 ;
  assign n10447 = n10446 ^ n10386 ;
  assign n10676 = n10675 ^ n10447 ;
  assign n10694 = n10693 ^ n10676 ;
  assign n10695 = n10694 ^ x5 ;
  assign n10444 = x124 & n234 ;
  assign n10696 = n10695 ^ n10444 ;
  assign n10443 = x126 & n230 ;
  assign n10697 = n10696 ^ n10443 ;
  assign n10441 = n9526 ^ x126 ;
  assign n10442 = n231 & n10441 ;
  assign n10698 = n10697 ^ n10442 ;
  assign n10700 = n10699 ^ n10698 ;
  assign n10438 = n10396 ^ n10387 ;
  assign n10439 = n10393 & n10438 ;
  assign n10440 = n10439 ^ n10396 ;
  assign n10701 = n10700 ^ n10440 ;
  assign n10425 = x127 & n10129 ;
  assign n10426 = n10138 ^ x2 ;
  assign n10429 = x0 & ~n10426 ;
  assign n10430 = n10429 ^ x2 ;
  assign n10431 = n10425 & n10430 ;
  assign n10432 = n10431 ^ x2 ;
  assign n10433 = n10432 ^ n10407 ;
  assign n10434 = n10433 ^ n10397 ;
  assign n10435 = n10434 ^ n10432 ;
  assign n10436 = n10415 & n10435 ;
  assign n10437 = n10436 ^ n10433 ;
  assign n10702 = n10701 ^ n10437 ;
  assign n10703 = n10702 ^ n10149 ;
  assign n10704 = n10703 ^ n10702 ;
  assign n10705 = n10704 ^ n10127 ;
  assign n10706 = n10417 & n10705 ;
  assign n10707 = n10706 ^ n10703 ;
  assign n10711 = n10710 ^ n10707 ;
  assign n10975 = x125 & n234 ;
  assign n10974 = x127 & n230 ;
  assign n10976 = n10975 ^ n10974 ;
  assign n10977 = n10976 ^ x5 ;
  assign n10972 = n9832 ^ x127 ;
  assign n10973 = n231 & n10972 ;
  assign n10978 = n10977 ^ n10973 ;
  assign n10971 = x126 & n227 ;
  assign n10979 = n10978 ^ n10971 ;
  assign n10960 = x122 & n446 ;
  assign n10959 = x124 & n383 ;
  assign n10961 = n10960 ^ n10959 ;
  assign n10962 = n10961 ^ x8 ;
  assign n10958 = n384 & n10095 ;
  assign n10963 = n10962 ^ n10958 ;
  assign n10957 = x123 & n390 ;
  assign n10964 = n10963 ^ n10957 ;
  assign n10948 = n10669 ^ n10447 ;
  assign n10949 = n10675 & ~n10948 ;
  assign n10950 = n10949 ^ n10669 ;
  assign n10946 = x120 & n578 ;
  assign n10939 = x117 & n788 ;
  assign n10931 = n10652 ^ n10456 ;
  assign n10932 = ~n10658 & n10931 ;
  assign n10933 = n10932 ^ n10652 ;
  assign n10929 = x114 & n1058 ;
  assign n10922 = x111 & n1335 ;
  assign n10915 = x108 & n1666 ;
  assign n10907 = n10625 ^ n10468 ;
  assign n10908 = n10631 & ~n10907 ;
  assign n10909 = n10908 ^ n10625 ;
  assign n10905 = x105 & n2014 ;
  assign n10897 = n10618 ^ n10474 ;
  assign n10898 = ~n10624 & n10897 ;
  assign n10899 = n10898 ^ n10618 ;
  assign n10895 = x102 & n2429 ;
  assign n10888 = x99 & n2887 ;
  assign n10880 = n10601 ^ n10483 ;
  assign n10881 = ~n10607 & n10880 ;
  assign n10882 = n10881 ^ n10601 ;
  assign n10878 = x96 & n3383 ;
  assign n10871 = x93 & n3924 ;
  assign n10864 = x90 & n4467 ;
  assign n10856 = n10577 ^ n10498 ;
  assign n10857 = ~n10583 & n10856 ;
  assign n10858 = n10857 ^ n10577 ;
  assign n10854 = x87 & n5102 ;
  assign n10846 = n10570 ^ n10504 ;
  assign n10847 = ~n10576 & ~n10846 ;
  assign n10848 = n10847 ^ n10570 ;
  assign n10844 = x84 & n5736 ;
  assign n10837 = x81 & n6433 ;
  assign n10830 = x78 & n7179 ;
  assign n10822 = n10561 ^ n10536 ;
  assign n10823 = n10567 & n10822 ;
  assign n10824 = n10823 ^ n10561 ;
  assign n10820 = x75 & n7931 ;
  assign n10812 = n10560 ^ n10542 ;
  assign n10813 = n10552 & n10812 ;
  assign n10814 = n10813 ^ n10542 ;
  assign n10805 = x71 & n8741 ;
  assign n10804 = x73 & n8744 ;
  assign n10806 = n10805 ^ n10804 ;
  assign n10807 = n10806 ^ x59 ;
  assign n10803 = n633 & n8745 ;
  assign n10808 = n10807 ^ n10803 ;
  assign n10802 = x72 & n8737 ;
  assign n10809 = n10808 ^ n10802 ;
  assign n10798 = ~n436 & n9636 ;
  assign n10797 = x69 & n9628 ;
  assign n10799 = n10798 ^ n10797 ;
  assign n10795 = x68 & n9632 ;
  assign n10794 = x70 & n9635 ;
  assign n10796 = n10795 ^ n10794 ;
  assign n10800 = n10799 ^ n10796 ;
  assign n10792 = x63 & x67 ;
  assign n10793 = n10792 ^ x2 ;
  assign n10801 = n10800 ^ n10793 ;
  assign n10810 = n10809 ^ n10801 ;
  assign n10789 = x63 & x66 ;
  assign n10790 = n10789 ^ x67 ;
  assign n10791 = x62 & ~n10790 ;
  assign n10811 = n10810 ^ n10791 ;
  assign n10815 = n10814 ^ n10811 ;
  assign n10816 = n10815 ^ x56 ;
  assign n10786 = x74 & n7935 ;
  assign n10817 = n10816 ^ n10786 ;
  assign n10785 = x76 & n7938 ;
  assign n10818 = n10817 ^ n10785 ;
  assign n10784 = ~n853 & n7939 ;
  assign n10819 = n10818 ^ n10784 ;
  assign n10821 = n10820 ^ n10819 ;
  assign n10825 = n10824 ^ n10821 ;
  assign n10826 = n10825 ^ x53 ;
  assign n10783 = x77 & n7171 ;
  assign n10827 = n10826 ^ n10783 ;
  assign n10782 = x79 & n7174 ;
  assign n10828 = n10827 ^ n10782 ;
  assign n10781 = n1118 & n7175 ;
  assign n10829 = n10828 ^ n10781 ;
  assign n10831 = n10830 ^ n10829 ;
  assign n10778 = n10568 ^ n10528 ;
  assign n10779 = ~n10533 & n10778 ;
  assign n10780 = n10779 ^ n10528 ;
  assign n10832 = n10831 ^ n10780 ;
  assign n10833 = n10832 ^ x50 ;
  assign n10777 = x80 & n6677 ;
  assign n10834 = n10833 ^ n10777 ;
  assign n10776 = x82 & n6428 ;
  assign n10835 = n10834 ^ n10776 ;
  assign n10775 = n1411 & n6429 ;
  assign n10836 = n10835 ^ n10775 ;
  assign n10838 = n10837 ^ n10836 ;
  assign n10772 = n10569 ^ n10515 ;
  assign n10773 = n10520 & ~n10772 ;
  assign n10774 = n10773 ^ n10515 ;
  assign n10839 = n10838 ^ n10774 ;
  assign n10840 = n10839 ^ x47 ;
  assign n10771 = x83 & n5965 ;
  assign n10841 = n10840 ^ n10771 ;
  assign n10770 = x85 & n5729 ;
  assign n10842 = n10841 ^ n10770 ;
  assign n10769 = n1743 & n5730 ;
  assign n10843 = n10842 ^ n10769 ;
  assign n10845 = n10844 ^ n10843 ;
  assign n10849 = n10848 ^ n10845 ;
  assign n10850 = n10849 ^ x44 ;
  assign n10768 = x86 & n5094 ;
  assign n10851 = n10850 ^ n10768 ;
  assign n10767 = x88 & n5097 ;
  assign n10852 = n10851 ^ n10767 ;
  assign n10766 = n2119 & n5098 ;
  assign n10853 = n10852 ^ n10766 ;
  assign n10855 = n10854 ^ n10853 ;
  assign n10859 = n10858 ^ n10855 ;
  assign n10860 = n10859 ^ x41 ;
  assign n10765 = x89 & n4474 ;
  assign n10861 = n10860 ^ n10765 ;
  assign n10764 = x91 & n4471 ;
  assign n10862 = n10861 ^ n10764 ;
  assign n10763 = n2542 & n4472 ;
  assign n10863 = n10862 ^ n10763 ;
  assign n10865 = n10864 ^ n10863 ;
  assign n10760 = n10584 ^ n10492 ;
  assign n10761 = n10590 & ~n10760 ;
  assign n10762 = n10761 ^ n10584 ;
  assign n10866 = n10865 ^ n10762 ;
  assign n10867 = n10866 ^ x38 ;
  assign n10759 = x92 & n3916 ;
  assign n10868 = n10867 ^ n10759 ;
  assign n10758 = x94 & n3919 ;
  assign n10869 = n10868 ^ n10758 ;
  assign n10757 = n2997 & n3920 ;
  assign n10870 = n10869 ^ n10757 ;
  assign n10872 = n10871 ^ n10870 ;
  assign n10754 = n10600 ^ n10591 ;
  assign n10755 = n10597 & ~n10754 ;
  assign n10756 = n10755 ^ n10600 ;
  assign n10873 = n10872 ^ n10756 ;
  assign n10874 = n10873 ^ x35 ;
  assign n10753 = x95 & n3375 ;
  assign n10875 = n10874 ^ n10753 ;
  assign n10752 = x97 & n3378 ;
  assign n10876 = n10875 ^ n10752 ;
  assign n10751 = n3379 & n3494 ;
  assign n10877 = n10876 ^ n10751 ;
  assign n10879 = n10878 ^ n10877 ;
  assign n10883 = n10882 ^ n10879 ;
  assign n10884 = n10883 ^ x32 ;
  assign n10750 = x98 & n2879 ;
  assign n10885 = n10884 ^ n10750 ;
  assign n10749 = x100 & n2882 ;
  assign n10886 = n10885 ^ n10749 ;
  assign n10748 = n2883 & n4034 ;
  assign n10887 = n10886 ^ n10748 ;
  assign n10889 = n10888 ^ n10887 ;
  assign n10745 = n10617 ^ n10608 ;
  assign n10746 = ~n10614 & ~n10745 ;
  assign n10747 = n10746 ^ n10617 ;
  assign n10890 = n10889 ^ n10747 ;
  assign n10891 = n10890 ^ x29 ;
  assign n10744 = x101 & n2581 ;
  assign n10892 = n10891 ^ n10744 ;
  assign n10743 = x103 & n2422 ;
  assign n10893 = n10892 ^ n10743 ;
  assign n10742 = n2423 & ~n4615 ;
  assign n10894 = n10893 ^ n10742 ;
  assign n10896 = n10895 ^ n10894 ;
  assign n10900 = n10899 ^ n10896 ;
  assign n10901 = n10900 ^ x26 ;
  assign n10741 = x104 & n2018 ;
  assign n10902 = n10901 ^ n10741 ;
  assign n10740 = x106 & n2021 ;
  assign n10903 = n10902 ^ n10740 ;
  assign n10739 = n2022 & ~n5240 ;
  assign n10904 = n10903 ^ n10739 ;
  assign n10906 = n10905 ^ n10904 ;
  assign n10910 = n10909 ^ n10906 ;
  assign n10911 = n10910 ^ x23 ;
  assign n10738 = x107 & n1658 ;
  assign n10912 = n10911 ^ n10738 ;
  assign n10737 = x109 & n1661 ;
  assign n10913 = n10912 ^ n10737 ;
  assign n10736 = n1662 & n5902 ;
  assign n10914 = n10913 ^ n10736 ;
  assign n10916 = n10915 ^ n10914 ;
  assign n10733 = n10641 ^ n10632 ;
  assign n10734 = n10638 & n10733 ;
  assign n10735 = n10734 ^ n10641 ;
  assign n10917 = n10916 ^ n10735 ;
  assign n10918 = n10917 ^ x20 ;
  assign n10732 = x110 & n1327 ;
  assign n10919 = n10918 ^ n10732 ;
  assign n10731 = x112 & n1330 ;
  assign n10920 = n10919 ^ n10731 ;
  assign n10730 = n1331 & ~n6600 ;
  assign n10921 = n10920 ^ n10730 ;
  assign n10923 = n10922 ^ n10921 ;
  assign n10727 = n10651 ^ n10642 ;
  assign n10728 = ~n10648 & ~n10727 ;
  assign n10729 = n10728 ^ n10651 ;
  assign n10924 = n10923 ^ n10729 ;
  assign n10925 = n10924 ^ x17 ;
  assign n10726 = x113 & n1050 ;
  assign n10926 = n10925 ^ n10726 ;
  assign n10725 = x115 & n1053 ;
  assign n10927 = n10926 ^ n10725 ;
  assign n10724 = n1054 & ~n7343 ;
  assign n10928 = n10927 ^ n10724 ;
  assign n10930 = n10929 ^ n10928 ;
  assign n10934 = n10933 ^ n10930 ;
  assign n10935 = n10934 ^ x14 ;
  assign n10723 = x116 & n877 ;
  assign n10936 = n10935 ^ n10723 ;
  assign n10722 = x118 & n782 ;
  assign n10937 = n10936 ^ n10722 ;
  assign n10721 = n783 & ~n8123 ;
  assign n10938 = n10937 ^ n10721 ;
  assign n10940 = n10939 ^ n10938 ;
  assign n10718 = n10668 ^ n10659 ;
  assign n10719 = ~n10665 & n10718 ;
  assign n10720 = n10719 ^ n10668 ;
  assign n10941 = n10940 ^ n10720 ;
  assign n10942 = n10941 ^ x11 ;
  assign n10717 = x119 & n647 ;
  assign n10943 = n10942 ^ n10717 ;
  assign n10716 = x121 & ~n572 ;
  assign n10944 = n10943 ^ n10716 ;
  assign n10715 = ~n573 & n8962 ;
  assign n10945 = n10944 ^ n10715 ;
  assign n10947 = n10946 ^ n10945 ;
  assign n10951 = n10950 ^ n10947 ;
  assign n10952 = n10951 ^ n10685 ;
  assign n10953 = n10952 ^ n10676 ;
  assign n10954 = n10953 ^ n10951 ;
  assign n10955 = n10693 & ~n10954 ;
  assign n10956 = n10955 ^ n10952 ;
  assign n10965 = n10964 ^ n10956 ;
  assign n10966 = n10965 ^ n10694 ;
  assign n10967 = n10966 ^ n10965 ;
  assign n10968 = n10967 ^ n10440 ;
  assign n10969 = ~n10700 & n10968 ;
  assign n10970 = n10969 ^ n10966 ;
  assign n10980 = n10979 ^ n10970 ;
  assign n10982 = n10980 ^ n10701 ;
  assign n10981 = n10980 ^ n10432 ;
  assign n10983 = n10982 ^ n10981 ;
  assign n10984 = n10437 & n10983 ;
  assign n10985 = n10984 ^ n10981 ;
  assign n10712 = n10710 ^ n10702 ;
  assign n10713 = ~n10707 & n10712 ;
  assign n10714 = n10713 ^ n10710 ;
  assign n10986 = n10985 ^ n10714 ;
  assign n11253 = n10980 ^ n10714 ;
  assign n11254 = ~n10985 & ~n11253 ;
  assign n11255 = n11254 ^ n10980 ;
  assign n11249 = n10979 ^ n10965 ;
  assign n11250 = ~n10970 & n11249 ;
  assign n11251 = n11250 ^ n10965 ;
  assign n11245 = n10964 ^ n10951 ;
  assign n11246 = n10956 & n11245 ;
  assign n11247 = n11246 ^ n10951 ;
  assign n11243 = x127 & n227 ;
  assign n11237 = x124 & n390 ;
  assign n11229 = n10934 ^ n10720 ;
  assign n11230 = n10940 & n11229 ;
  assign n11231 = n11230 ^ n10934 ;
  assign n11227 = x121 & n578 ;
  assign n11220 = x118 & n788 ;
  assign n11212 = n10917 ^ n10729 ;
  assign n11213 = n10923 & ~n11212 ;
  assign n11214 = n11213 ^ n10917 ;
  assign n11210 = x115 & n1058 ;
  assign n11202 = n10910 ^ n10735 ;
  assign n11203 = ~n10916 & n11202 ;
  assign n11204 = n11203 ^ n10910 ;
  assign n11200 = x112 & n1335 ;
  assign n11193 = x109 & n1666 ;
  assign n11186 = x106 & n2014 ;
  assign n11178 = n10883 ^ n10747 ;
  assign n11179 = ~n10889 & n11178 ;
  assign n11180 = n11179 ^ n10883 ;
  assign n11176 = x103 & n2429 ;
  assign n11169 = x100 & n2887 ;
  assign n11161 = n10866 ^ n10756 ;
  assign n11162 = n10872 & n11161 ;
  assign n11163 = n11162 ^ n10866 ;
  assign n11159 = x97 & n3383 ;
  assign n11152 = x94 & n3924 ;
  assign n11145 = x91 & n4467 ;
  assign n11138 = x88 & n5102 ;
  assign n11131 = x85 & n5736 ;
  assign n11119 = x78 & n7171 ;
  assign n11118 = x80 & n7174 ;
  assign n11120 = n11119 ^ n11118 ;
  assign n11121 = n11120 ^ x53 ;
  assign n11117 = n1206 & n7175 ;
  assign n11122 = n11121 ^ n11117 ;
  assign n11116 = x79 & n7179 ;
  assign n11123 = n11122 ^ n11116 ;
  assign n11109 = x75 & n7935 ;
  assign n11108 = x77 & n7938 ;
  assign n11110 = n11109 ^ n11108 ;
  assign n11111 = n11110 ^ x56 ;
  assign n11107 = ~n939 & n7939 ;
  assign n11112 = n11111 ^ n11107 ;
  assign n11106 = x76 & n7931 ;
  assign n11113 = n11112 ^ n11106 ;
  assign n11100 = x63 & x68 ;
  assign n11101 = n11100 ^ x2 ;
  assign n11097 = ~n493 & n9636 ;
  assign n11096 = x70 & n9628 ;
  assign n11098 = n11097 ^ n11096 ;
  assign n11094 = x69 & n9632 ;
  assign n11093 = x71 & n9635 ;
  assign n11095 = n11094 ^ n11093 ;
  assign n11099 = n11098 ^ n11095 ;
  assign n11102 = n11101 ^ n11099 ;
  assign n11087 = x62 ^ x2 ;
  assign n11088 = n11087 ^ n10800 ;
  assign n11089 = n10800 ^ n10792 ;
  assign n11090 = n11089 ^ n10791 ;
  assign n11091 = n11088 & ~n11090 ;
  assign n11092 = n11091 ^ x2 ;
  assign n11103 = n11102 ^ n11092 ;
  assign n11085 = n10792 ^ x68 ;
  assign n11086 = x62 & ~n11085 ;
  assign n11104 = n11103 ^ n11086 ;
  assign n11080 = x72 & n8741 ;
  assign n11079 = x74 & n8744 ;
  assign n11081 = n11080 ^ n11079 ;
  assign n11082 = n11081 ^ x59 ;
  assign n11078 = n699 & n8745 ;
  assign n11083 = n11082 ^ n11078 ;
  assign n11077 = x73 & n8737 ;
  assign n11084 = n11083 ^ n11077 ;
  assign n11105 = n11104 ^ n11084 ;
  assign n11114 = n11113 ^ n11105 ;
  assign n11074 = n10814 ^ n10809 ;
  assign n11075 = ~n10811 & n11074 ;
  assign n11076 = n11075 ^ n10814 ;
  assign n11115 = n11114 ^ n11076 ;
  assign n11124 = n11123 ^ n11115 ;
  assign n11071 = n10824 ^ n10815 ;
  assign n11072 = ~n10821 & n11071 ;
  assign n11073 = n11072 ^ n10824 ;
  assign n11125 = n11124 ^ n11073 ;
  assign n11061 = x81 & n6677 ;
  assign n11060 = x83 & n6428 ;
  assign n11062 = n11061 ^ n11060 ;
  assign n11063 = n11062 ^ x50 ;
  assign n11059 = n1512 & n6429 ;
  assign n11064 = n11063 ^ n11059 ;
  assign n11058 = x82 & n6433 ;
  assign n11065 = n11064 ^ n11058 ;
  assign n11066 = n11065 ^ n10825 ;
  assign n11067 = n11066 ^ n10780 ;
  assign n11068 = n11067 ^ n11065 ;
  assign n11069 = n10831 & n11068 ;
  assign n11070 = n11069 ^ n11066 ;
  assign n11126 = n11125 ^ n11070 ;
  assign n11127 = n11126 ^ x47 ;
  assign n11057 = x84 & n5965 ;
  assign n11128 = n11127 ^ n11057 ;
  assign n11056 = x86 & n5729 ;
  assign n11129 = n11128 ^ n11056 ;
  assign n11055 = n1857 & n5730 ;
  assign n11130 = n11129 ^ n11055 ;
  assign n11132 = n11131 ^ n11130 ;
  assign n11052 = n10832 ^ n10774 ;
  assign n11053 = n10838 & n11052 ;
  assign n11054 = n11053 ^ n10832 ;
  assign n11133 = n11132 ^ n11054 ;
  assign n11134 = n11133 ^ x44 ;
  assign n11051 = x87 & n5094 ;
  assign n11135 = n11134 ^ n11051 ;
  assign n11050 = x89 & n5097 ;
  assign n11136 = n11135 ^ n11050 ;
  assign n11049 = n2249 & n5098 ;
  assign n11137 = n11136 ^ n11049 ;
  assign n11139 = n11138 ^ n11137 ;
  assign n11046 = n10848 ^ n10839 ;
  assign n11047 = ~n10845 & ~n11046 ;
  assign n11048 = n11047 ^ n10848 ;
  assign n11140 = n11139 ^ n11048 ;
  assign n11141 = n11140 ^ x41 ;
  assign n11045 = x90 & n4474 ;
  assign n11142 = n11141 ^ n11045 ;
  assign n11044 = x92 & n4471 ;
  assign n11143 = n11142 ^ n11044 ;
  assign n11043 = n2684 & n4472 ;
  assign n11144 = n11143 ^ n11043 ;
  assign n11146 = n11145 ^ n11144 ;
  assign n11040 = n10858 ^ n10849 ;
  assign n11041 = n10855 & n11040 ;
  assign n11042 = n11041 ^ n10858 ;
  assign n11147 = n11146 ^ n11042 ;
  assign n11148 = n11147 ^ x38 ;
  assign n11039 = x93 & n3916 ;
  assign n11149 = n11148 ^ n11039 ;
  assign n11038 = x95 & n3919 ;
  assign n11150 = n11149 ^ n11038 ;
  assign n11037 = n3159 & n3920 ;
  assign n11151 = n11150 ^ n11037 ;
  assign n11153 = n11152 ^ n11151 ;
  assign n11034 = n10859 ^ n10762 ;
  assign n11035 = n10865 & n11034 ;
  assign n11036 = n11035 ^ n10859 ;
  assign n11154 = n11153 ^ n11036 ;
  assign n11155 = n11154 ^ x35 ;
  assign n11033 = x96 & n3375 ;
  assign n11156 = n11155 ^ n11033 ;
  assign n11032 = x98 & n3378 ;
  assign n11157 = n11156 ^ n11032 ;
  assign n11031 = n3379 & n3660 ;
  assign n11158 = n11157 ^ n11031 ;
  assign n11160 = n11159 ^ n11158 ;
  assign n11164 = n11163 ^ n11160 ;
  assign n11165 = n11164 ^ x32 ;
  assign n11030 = x99 & n2879 ;
  assign n11166 = n11165 ^ n11030 ;
  assign n11029 = x101 & n2882 ;
  assign n11167 = n11166 ^ n11029 ;
  assign n11028 = n2883 & n4215 ;
  assign n11168 = n11167 ^ n11028 ;
  assign n11170 = n11169 ^ n11168 ;
  assign n11025 = n10882 ^ n10873 ;
  assign n11026 = ~n10879 & ~n11025 ;
  assign n11027 = n11026 ^ n10882 ;
  assign n11171 = n11170 ^ n11027 ;
  assign n11172 = n11171 ^ x29 ;
  assign n11024 = x102 & n2581 ;
  assign n11173 = n11172 ^ n11024 ;
  assign n11023 = x104 & n2422 ;
  assign n11174 = n11173 ^ n11023 ;
  assign n11022 = n2423 & ~n4814 ;
  assign n11175 = n11174 ^ n11022 ;
  assign n11177 = n11176 ^ n11175 ;
  assign n11181 = n11180 ^ n11177 ;
  assign n11182 = n11181 ^ x26 ;
  assign n11021 = x105 & n2018 ;
  assign n11183 = n11182 ^ n11021 ;
  assign n11020 = x107 & n2021 ;
  assign n11184 = n11183 ^ n11020 ;
  assign n11019 = n2022 & ~n5448 ;
  assign n11185 = n11184 ^ n11019 ;
  assign n11187 = n11186 ^ n11185 ;
  assign n11016 = n10899 ^ n10890 ;
  assign n11017 = ~n10896 & ~n11016 ;
  assign n11018 = n11017 ^ n10899 ;
  assign n11188 = n11187 ^ n11018 ;
  assign n11189 = n11188 ^ x23 ;
  assign n11015 = x108 & n1658 ;
  assign n11190 = n11189 ^ n11015 ;
  assign n11014 = x110 & n1661 ;
  assign n11191 = n11190 ^ n11014 ;
  assign n11013 = n1662 & n6129 ;
  assign n11192 = n11191 ^ n11013 ;
  assign n11194 = n11193 ^ n11192 ;
  assign n11010 = n10909 ^ n10900 ;
  assign n11011 = n10906 & ~n11010 ;
  assign n11012 = n11011 ^ n10909 ;
  assign n11195 = n11194 ^ n11012 ;
  assign n11196 = n11195 ^ x20 ;
  assign n11009 = x111 & n1327 ;
  assign n11197 = n11196 ^ n11009 ;
  assign n11008 = x113 & n1330 ;
  assign n11198 = n11197 ^ n11008 ;
  assign n11007 = n1331 & ~n6839 ;
  assign n11199 = n11198 ^ n11007 ;
  assign n11201 = n11200 ^ n11199 ;
  assign n11205 = n11204 ^ n11201 ;
  assign n11206 = n11205 ^ x17 ;
  assign n11006 = x114 & n1050 ;
  assign n11207 = n11206 ^ n11006 ;
  assign n11005 = x116 & n1053 ;
  assign n11208 = n11207 ^ n11005 ;
  assign n11004 = n1054 & ~n7588 ;
  assign n11209 = n11208 ^ n11004 ;
  assign n11211 = n11210 ^ n11209 ;
  assign n11215 = n11214 ^ n11211 ;
  assign n11216 = n11215 ^ x14 ;
  assign n11003 = x117 & n877 ;
  assign n11217 = n11216 ^ n11003 ;
  assign n11002 = x119 & n782 ;
  assign n11218 = n11217 ^ n11002 ;
  assign n11001 = n783 & n8394 ;
  assign n11219 = n11218 ^ n11001 ;
  assign n11221 = n11220 ^ n11219 ;
  assign n10998 = n10933 ^ n10924 ;
  assign n10999 = n10930 & n10998 ;
  assign n11000 = n10999 ^ n10933 ;
  assign n11222 = n11221 ^ n11000 ;
  assign n11223 = n11222 ^ x11 ;
  assign n10997 = x120 & n647 ;
  assign n11224 = n11223 ^ n10997 ;
  assign n10996 = x122 & ~n572 ;
  assign n11225 = n11224 ^ n10996 ;
  assign n10995 = ~n573 & ~n9247 ;
  assign n11226 = n11225 ^ n10995 ;
  assign n11228 = n11227 ^ n11226 ;
  assign n11232 = n11231 ^ n11228 ;
  assign n11233 = n11232 ^ x8 ;
  assign n10994 = x123 & n446 ;
  assign n11234 = n11233 ^ n10994 ;
  assign n10993 = x125 & n383 ;
  assign n11235 = n11234 ^ n10993 ;
  assign n10992 = n384 & n10400 ;
  assign n11236 = n11235 ^ n10992 ;
  assign n11238 = n11237 ^ n11236 ;
  assign n10989 = n10950 ^ n10941 ;
  assign n10990 = ~n10947 & n10989 ;
  assign n10991 = n10990 ^ n10950 ;
  assign n11239 = n11238 ^ n10991 ;
  assign n11240 = n11239 ^ x5 ;
  assign n10988 = x126 & n234 ;
  assign n11241 = n11240 ^ n10988 ;
  assign n10987 = n231 & n10139 ;
  assign n11242 = n11241 ^ n10987 ;
  assign n11244 = n11243 ^ n11242 ;
  assign n11248 = n11247 ^ n11244 ;
  assign n11252 = n11251 ^ n11248 ;
  assign n11256 = n11255 ^ n11252 ;
  assign n11525 = n11232 ^ n10991 ;
  assign n11526 = ~n11238 & ~n11525 ;
  assign n11527 = n11526 ^ n11232 ;
  assign n11521 = x125 & n390 ;
  assign n11513 = n11215 ^ n11000 ;
  assign n11514 = n11221 & ~n11513 ;
  assign n11515 = n11514 ^ n11215 ;
  assign n11511 = x122 & n578 ;
  assign n11504 = x119 & n788 ;
  assign n11497 = x116 & n1058 ;
  assign n11489 = n11188 ^ n11012 ;
  assign n11490 = ~n11194 & ~n11489 ;
  assign n11491 = n11490 ^ n11188 ;
  assign n11487 = x113 & n1335 ;
  assign n11479 = n11181 ^ n11018 ;
  assign n11480 = n11187 & ~n11479 ;
  assign n11481 = n11480 ^ n11181 ;
  assign n11477 = x110 & n1666 ;
  assign n11470 = x107 & n2014 ;
  assign n11462 = n11164 ^ n11027 ;
  assign n11463 = n11170 & ~n11462 ;
  assign n11464 = n11463 ^ n11164 ;
  assign n11460 = x104 & n2429 ;
  assign n11453 = x101 & n2887 ;
  assign n11446 = x98 & n3383 ;
  assign n11438 = n11140 ^ n11042 ;
  assign n11439 = ~n11146 & n11438 ;
  assign n11440 = n11439 ^ n11140 ;
  assign n11436 = x95 & n3924 ;
  assign n11428 = n11133 ^ n11048 ;
  assign n11429 = n11139 & ~n11428 ;
  assign n11430 = n11429 ^ n11133 ;
  assign n11426 = x92 & n4467 ;
  assign n11418 = n11126 ^ n11054 ;
  assign n11419 = n11132 & n11418 ;
  assign n11420 = n11419 ^ n11126 ;
  assign n11416 = x89 & n5102 ;
  assign n11406 = x85 & n5965 ;
  assign n11405 = x87 & n5729 ;
  assign n11407 = n11406 ^ n11405 ;
  assign n11408 = n11407 ^ x47 ;
  assign n11404 = n1982 & n5730 ;
  assign n11409 = n11408 ^ n11404 ;
  assign n11403 = x86 & n5736 ;
  assign n11410 = n11409 ^ n11403 ;
  assign n11394 = n11123 ^ n11073 ;
  assign n11395 = n11124 & n11394 ;
  assign n11396 = n11395 ^ n11123 ;
  assign n11388 = x82 & n6677 ;
  assign n11387 = x84 & n6428 ;
  assign n11389 = n11388 ^ n11387 ;
  assign n11390 = n11389 ^ x50 ;
  assign n11386 = n1624 & n6429 ;
  assign n11391 = n11390 ^ n11386 ;
  assign n11385 = x83 & n6433 ;
  assign n11392 = n11391 ^ n11385 ;
  assign n11382 = x80 & n7179 ;
  assign n11380 = n1305 & n7175 ;
  assign n11376 = x79 & n7171 ;
  assign n11375 = x81 & n7174 ;
  assign n11377 = n11376 ^ n11375 ;
  assign n11378 = n11377 ^ x53 ;
  assign n11370 = n11100 ^ x69 ;
  assign n11371 = x62 & ~n11370 ;
  assign n11368 = x63 & x69 ;
  assign n11364 = n556 & n9636 ;
  assign n11363 = x71 & n9628 ;
  assign n11365 = n11364 ^ n11363 ;
  assign n11361 = x70 & n9632 ;
  assign n11360 = x72 & n9635 ;
  assign n11362 = n11361 ^ n11360 ;
  assign n11366 = n11365 ^ n11362 ;
  assign n11367 = n11366 ^ x2 ;
  assign n11369 = n11368 ^ n11367 ;
  assign n11372 = n11371 ^ n11369 ;
  assign n11355 = n11099 ^ n11087 ;
  assign n11356 = n11100 ^ n11099 ;
  assign n11357 = n11356 ^ n11086 ;
  assign n11358 = n11355 & ~n11357 ;
  assign n11349 = x73 & n8741 ;
  assign n11348 = x75 & n8744 ;
  assign n11350 = n11349 ^ n11348 ;
  assign n11351 = n11350 ^ x59 ;
  assign n11347 = ~n774 & n8745 ;
  assign n11352 = n11351 ^ n11347 ;
  assign n11346 = x74 & n8737 ;
  assign n11353 = n11352 ^ n11346 ;
  assign n11354 = n11353 ^ x2 ;
  assign n11359 = n11358 ^ n11354 ;
  assign n11373 = n11372 ^ n11359 ;
  assign n11343 = ~n1025 & n7939 ;
  assign n11341 = x76 & n7935 ;
  assign n11337 = n11092 ^ n11084 ;
  assign n11338 = ~n11104 & n11337 ;
  assign n11339 = n11338 ^ n11084 ;
  assign n11335 = x78 & n7938 ;
  assign n11336 = n11335 ^ x56 ;
  assign n11340 = n11339 ^ n11336 ;
  assign n11342 = n11341 ^ n11340 ;
  assign n11344 = n11343 ^ n11342 ;
  assign n11334 = x77 & n7931 ;
  assign n11345 = n11344 ^ n11334 ;
  assign n11374 = n11373 ^ n11345 ;
  assign n11379 = n11378 ^ n11374 ;
  assign n11381 = n11380 ^ n11379 ;
  assign n11383 = n11382 ^ n11381 ;
  assign n11331 = n11113 ^ n11076 ;
  assign n11332 = n11114 & n11331 ;
  assign n11333 = n11332 ^ n11113 ;
  assign n11384 = n11383 ^ n11333 ;
  assign n11393 = n11392 ^ n11384 ;
  assign n11397 = n11396 ^ n11393 ;
  assign n11399 = n11397 ^ n11065 ;
  assign n11398 = n11397 ^ n11125 ;
  assign n11400 = n11399 ^ n11398 ;
  assign n11401 = n11070 & n11400 ;
  assign n11402 = n11401 ^ n11399 ;
  assign n11411 = n11410 ^ n11402 ;
  assign n11412 = n11411 ^ x44 ;
  assign n11330 = x88 & n5094 ;
  assign n11413 = n11412 ^ n11330 ;
  assign n11329 = x90 & n5097 ;
  assign n11414 = n11413 ^ n11329 ;
  assign n11328 = n2386 & n5098 ;
  assign n11415 = n11414 ^ n11328 ;
  assign n11417 = n11416 ^ n11415 ;
  assign n11421 = n11420 ^ n11417 ;
  assign n11422 = n11421 ^ x41 ;
  assign n11327 = x91 & n4474 ;
  assign n11423 = n11422 ^ n11327 ;
  assign n11326 = x93 & n4471 ;
  assign n11424 = n11423 ^ n11326 ;
  assign n11325 = n2836 & n4472 ;
  assign n11425 = n11424 ^ n11325 ;
  assign n11427 = n11426 ^ n11425 ;
  assign n11431 = n11430 ^ n11427 ;
  assign n11432 = n11431 ^ x38 ;
  assign n11324 = x94 & n3916 ;
  assign n11433 = n11432 ^ n11324 ;
  assign n11323 = x96 & n3919 ;
  assign n11434 = n11433 ^ n11323 ;
  assign n11322 = n3323 & n3920 ;
  assign n11435 = n11434 ^ n11322 ;
  assign n11437 = n11436 ^ n11435 ;
  assign n11441 = n11440 ^ n11437 ;
  assign n11442 = n11441 ^ x35 ;
  assign n11321 = x97 & n3375 ;
  assign n11443 = n11442 ^ n11321 ;
  assign n11320 = x99 & n3378 ;
  assign n11444 = n11443 ^ n11320 ;
  assign n11319 = n3379 & n3843 ;
  assign n11445 = n11444 ^ n11319 ;
  assign n11447 = n11446 ^ n11445 ;
  assign n11316 = n11147 ^ n11036 ;
  assign n11317 = n11153 & n11316 ;
  assign n11318 = n11317 ^ n11147 ;
  assign n11448 = n11447 ^ n11318 ;
  assign n11449 = n11448 ^ x32 ;
  assign n11315 = x100 & n2879 ;
  assign n11450 = n11449 ^ n11315 ;
  assign n11314 = x102 & n2882 ;
  assign n11451 = n11450 ^ n11314 ;
  assign n11313 = n2883 & n4410 ;
  assign n11452 = n11451 ^ n11313 ;
  assign n11454 = n11453 ^ n11452 ;
  assign n11310 = n11163 ^ n11154 ;
  assign n11311 = ~n11160 & n11310 ;
  assign n11312 = n11311 ^ n11163 ;
  assign n11455 = n11454 ^ n11312 ;
  assign n11456 = n11455 ^ x29 ;
  assign n11309 = x103 & n2581 ;
  assign n11457 = n11456 ^ n11309 ;
  assign n11308 = x105 & n2422 ;
  assign n11458 = n11457 ^ n11308 ;
  assign n11307 = n2423 & ~n5023 ;
  assign n11459 = n11458 ^ n11307 ;
  assign n11461 = n11460 ^ n11459 ;
  assign n11465 = n11464 ^ n11461 ;
  assign n11466 = n11465 ^ x26 ;
  assign n11306 = x106 & n2018 ;
  assign n11467 = n11466 ^ n11306 ;
  assign n11305 = x108 & n2021 ;
  assign n11468 = n11467 ^ n11305 ;
  assign n11304 = n2022 & n5670 ;
  assign n11469 = n11468 ^ n11304 ;
  assign n11471 = n11470 ^ n11469 ;
  assign n11301 = n11180 ^ n11171 ;
  assign n11302 = n11177 & n11301 ;
  assign n11303 = n11302 ^ n11180 ;
  assign n11472 = n11471 ^ n11303 ;
  assign n11473 = n11472 ^ x23 ;
  assign n11300 = x109 & n1658 ;
  assign n11474 = n11473 ^ n11300 ;
  assign n11299 = x111 & n1661 ;
  assign n11475 = n11474 ^ n11299 ;
  assign n11298 = n1662 & ~n6360 ;
  assign n11476 = n11475 ^ n11298 ;
  assign n11478 = n11477 ^ n11476 ;
  assign n11482 = n11481 ^ n11478 ;
  assign n11483 = n11482 ^ x20 ;
  assign n11297 = x112 & n1327 ;
  assign n11484 = n11483 ^ n11297 ;
  assign n11296 = x114 & n1330 ;
  assign n11485 = n11484 ^ n11296 ;
  assign n11295 = n1331 & ~n7092 ;
  assign n11486 = n11485 ^ n11295 ;
  assign n11488 = n11487 ^ n11486 ;
  assign n11492 = n11491 ^ n11488 ;
  assign n11493 = n11492 ^ x17 ;
  assign n11294 = x115 & n1050 ;
  assign n11494 = n11493 ^ n11294 ;
  assign n11293 = x117 & n1053 ;
  assign n11495 = n11494 ^ n11293 ;
  assign n11292 = n1054 & ~n7850 ;
  assign n11496 = n11495 ^ n11292 ;
  assign n11498 = n11497 ^ n11496 ;
  assign n11289 = n11204 ^ n11195 ;
  assign n11290 = n11201 & n11289 ;
  assign n11291 = n11290 ^ n11204 ;
  assign n11499 = n11498 ^ n11291 ;
  assign n11500 = n11499 ^ x14 ;
  assign n11288 = x118 & n877 ;
  assign n11501 = n11500 ^ n11288 ;
  assign n11287 = x120 & n782 ;
  assign n11502 = n11501 ^ n11287 ;
  assign n11286 = n783 & n8891 ;
  assign n11503 = n11502 ^ n11286 ;
  assign n11505 = n11504 ^ n11503 ;
  assign n11283 = n11214 ^ n11205 ;
  assign n11284 = ~n11211 & n11283 ;
  assign n11285 = n11284 ^ n11214 ;
  assign n11506 = n11505 ^ n11285 ;
  assign n11507 = n11506 ^ x11 ;
  assign n11282 = x121 & n647 ;
  assign n11508 = n11507 ^ n11282 ;
  assign n11281 = x123 & ~n572 ;
  assign n11509 = n11508 ^ n11281 ;
  assign n11280 = ~n573 & ~n9786 ;
  assign n11510 = n11509 ^ n11280 ;
  assign n11512 = n11511 ^ n11510 ;
  assign n11516 = n11515 ^ n11512 ;
  assign n11517 = n11516 ^ x8 ;
  assign n11279 = x124 & n446 ;
  assign n11518 = n11517 ^ n11279 ;
  assign n11278 = x126 & n383 ;
  assign n11519 = n11518 ^ n11278 ;
  assign n11277 = n384 & n10441 ;
  assign n11520 = n11519 ^ n11277 ;
  assign n11522 = n11521 ^ n11520 ;
  assign n11274 = n11231 ^ n11222 ;
  assign n11275 = n11228 & ~n11274 ;
  assign n11276 = n11275 ^ n11231 ;
  assign n11523 = n11522 ^ n11276 ;
  assign n11263 = x127 & n233 ;
  assign n11264 = n11263 ^ n229 ;
  assign n11265 = n10138 ^ x127 ;
  assign n11270 = n198 & n11265 ;
  assign n11271 = n11270 ^ n11263 ;
  assign n11272 = n11264 & ~n11271 ;
  assign n11273 = n11272 ^ x4 ;
  assign n11524 = n11523 ^ n11273 ;
  assign n11528 = n11527 ^ n11524 ;
  assign n11260 = n11247 ^ n11239 ;
  assign n11261 = n11244 & ~n11260 ;
  assign n11262 = n11261 ^ n11247 ;
  assign n11529 = n11528 ^ n11262 ;
  assign n11257 = n11255 ^ n11251 ;
  assign n11258 = n11252 & ~n11257 ;
  assign n11259 = n11258 ^ n11255 ;
  assign n11530 = n11529 ^ n11259 ;
  assign n11804 = ~n11262 & ~n11523 ;
  assign n11805 = n11259 & ~n11528 ;
  assign n11806 = n11804 & n11805 ;
  assign n11531 = n11527 ^ n11273 ;
  assign n11789 = n11516 ^ n11276 ;
  assign n11790 = n11522 & n11789 ;
  assign n11791 = n11790 ^ n11516 ;
  assign n11787 = x126 & n390 ;
  assign n11780 = x123 & n578 ;
  assign n11772 = n11499 ^ n11285 ;
  assign n11773 = n11505 & n11772 ;
  assign n11774 = n11773 ^ n11499 ;
  assign n11770 = x120 & n788 ;
  assign n11762 = n11492 ^ n11291 ;
  assign n11763 = ~n11498 & n11762 ;
  assign n11764 = n11763 ^ n11492 ;
  assign n11760 = x117 & n1058 ;
  assign n11753 = x114 & n1335 ;
  assign n11746 = x111 & n1666 ;
  assign n11738 = n11465 ^ n11303 ;
  assign n11739 = ~n11471 & n11738 ;
  assign n11740 = n11739 ^ n11465 ;
  assign n11736 = x108 & n2014 ;
  assign n11729 = x105 & n2429 ;
  assign n11721 = n11448 ^ n11312 ;
  assign n11722 = ~n11454 & ~n11721 ;
  assign n11723 = n11722 ^ n11448 ;
  assign n11719 = x102 & n2887 ;
  assign n11712 = x99 & n3383 ;
  assign n11705 = x96 & n3924 ;
  assign n11698 = x93 & n4467 ;
  assign n11691 = x90 & n5102 ;
  assign n11681 = x86 & n5965 ;
  assign n11680 = x88 & n5729 ;
  assign n11682 = n11681 ^ n11680 ;
  assign n11683 = n11682 ^ x47 ;
  assign n11679 = n2119 & n5730 ;
  assign n11684 = n11683 ^ n11679 ;
  assign n11678 = x87 & n5736 ;
  assign n11685 = n11684 ^ n11678 ;
  assign n11670 = x84 & n6433 ;
  assign n11662 = n11374 ^ n11333 ;
  assign n11663 = n11383 & n11662 ;
  assign n11664 = n11663 ^ n11374 ;
  assign n11656 = x80 & n7171 ;
  assign n11655 = x82 & n7174 ;
  assign n11657 = n11656 ^ n11655 ;
  assign n11658 = n11657 ^ x53 ;
  assign n11654 = n1411 & n7175 ;
  assign n11659 = n11658 ^ n11654 ;
  assign n11653 = x81 & n7179 ;
  assign n11660 = n11659 ^ n11653 ;
  assign n11649 = x75 & n8737 ;
  assign n11639 = x71 & n9632 ;
  assign n11638 = x73 & n9635 ;
  assign n11640 = n11639 ^ n11638 ;
  assign n11641 = n11640 ^ x62 ;
  assign n11637 = n633 & n9636 ;
  assign n11642 = n11641 ^ n11637 ;
  assign n11636 = x72 & n9628 ;
  assign n11643 = n11642 ^ n11636 ;
  assign n11630 = n11366 ^ n11087 ;
  assign n11631 = n11371 ^ n11368 ;
  assign n11632 = n11631 ^ n11366 ;
  assign n11633 = n11630 & ~n11632 ;
  assign n11634 = n11633 ^ x2 ;
  assign n11626 = n11368 ^ x70 ;
  assign n11627 = ~n9948 & n11626 ;
  assign n11628 = n11627 ^ x70 ;
  assign n11625 = x5 ^ x2 ;
  assign n11629 = n11628 ^ n11625 ;
  assign n11635 = n11634 ^ n11629 ;
  assign n11644 = n11643 ^ n11635 ;
  assign n11645 = n11644 ^ x59 ;
  assign n11624 = x74 & n8741 ;
  assign n11646 = n11645 ^ n11624 ;
  assign n11623 = x76 & n8744 ;
  assign n11647 = n11646 ^ n11623 ;
  assign n11622 = ~n853 & n8745 ;
  assign n11648 = n11647 ^ n11622 ;
  assign n11650 = n11649 ^ n11648 ;
  assign n11619 = n11372 ^ n11353 ;
  assign n11620 = n11359 & n11619 ;
  assign n11621 = n11620 ^ n11353 ;
  assign n11651 = n11650 ^ n11621 ;
  assign n11609 = x77 & n7935 ;
  assign n11608 = x79 & n7938 ;
  assign n11610 = n11609 ^ n11608 ;
  assign n11611 = n11610 ^ x56 ;
  assign n11607 = n1118 & n7939 ;
  assign n11612 = n11611 ^ n11607 ;
  assign n11606 = x78 & n7931 ;
  assign n11613 = n11612 ^ n11606 ;
  assign n11614 = n11613 ^ n11373 ;
  assign n11615 = n11614 ^ n11339 ;
  assign n11616 = n11615 ^ n11613 ;
  assign n11617 = ~n11345 & n11616 ;
  assign n11618 = n11617 ^ n11614 ;
  assign n11652 = n11651 ^ n11618 ;
  assign n11661 = n11660 ^ n11652 ;
  assign n11665 = n11664 ^ n11661 ;
  assign n11666 = n11665 ^ x50 ;
  assign n11605 = x83 & n6677 ;
  assign n11667 = n11666 ^ n11605 ;
  assign n11604 = x85 & n6428 ;
  assign n11668 = n11667 ^ n11604 ;
  assign n11603 = n1743 & n6429 ;
  assign n11669 = n11668 ^ n11603 ;
  assign n11671 = n11670 ^ n11669 ;
  assign n11600 = n11396 ^ n11392 ;
  assign n11601 = ~n11393 & n11600 ;
  assign n11602 = n11601 ^ n11396 ;
  assign n11672 = n11671 ^ n11602 ;
  assign n11674 = n11672 ^ n11397 ;
  assign n11673 = n11672 ^ n11410 ;
  assign n11675 = n11674 ^ n11673 ;
  assign n11676 = n11402 & n11675 ;
  assign n11677 = n11676 ^ n11674 ;
  assign n11686 = n11685 ^ n11677 ;
  assign n11687 = n11686 ^ x44 ;
  assign n11599 = x89 & n5094 ;
  assign n11688 = n11687 ^ n11599 ;
  assign n11598 = x91 & n5097 ;
  assign n11689 = n11688 ^ n11598 ;
  assign n11597 = n2542 & n5098 ;
  assign n11690 = n11689 ^ n11597 ;
  assign n11692 = n11691 ^ n11690 ;
  assign n11594 = n11420 ^ n11411 ;
  assign n11595 = ~n11417 & n11594 ;
  assign n11596 = n11595 ^ n11420 ;
  assign n11693 = n11692 ^ n11596 ;
  assign n11694 = n11693 ^ x41 ;
  assign n11593 = x92 & n4474 ;
  assign n11695 = n11694 ^ n11593 ;
  assign n11592 = x94 & n4471 ;
  assign n11696 = n11695 ^ n11592 ;
  assign n11591 = n2997 & n4472 ;
  assign n11697 = n11696 ^ n11591 ;
  assign n11699 = n11698 ^ n11697 ;
  assign n11588 = n11430 ^ n11421 ;
  assign n11589 = ~n11427 & n11588 ;
  assign n11590 = n11589 ^ n11430 ;
  assign n11700 = n11699 ^ n11590 ;
  assign n11701 = n11700 ^ x38 ;
  assign n11587 = x95 & n3916 ;
  assign n11702 = n11701 ^ n11587 ;
  assign n11586 = x97 & n3919 ;
  assign n11703 = n11702 ^ n11586 ;
  assign n11585 = n3494 & n3920 ;
  assign n11704 = n11703 ^ n11585 ;
  assign n11706 = n11705 ^ n11704 ;
  assign n11582 = n11440 ^ n11431 ;
  assign n11583 = ~n11437 & ~n11582 ;
  assign n11584 = n11583 ^ n11440 ;
  assign n11707 = n11706 ^ n11584 ;
  assign n11708 = n11707 ^ x35 ;
  assign n11581 = x98 & n3375 ;
  assign n11709 = n11708 ^ n11581 ;
  assign n11580 = x100 & n3378 ;
  assign n11710 = n11709 ^ n11580 ;
  assign n11579 = n3379 & n4034 ;
  assign n11711 = n11710 ^ n11579 ;
  assign n11713 = n11712 ^ n11711 ;
  assign n11576 = n11441 ^ n11318 ;
  assign n11577 = ~n11447 & ~n11576 ;
  assign n11578 = n11577 ^ n11441 ;
  assign n11714 = n11713 ^ n11578 ;
  assign n11715 = n11714 ^ x32 ;
  assign n11575 = x101 & n2879 ;
  assign n11716 = n11715 ^ n11575 ;
  assign n11574 = x103 & n2882 ;
  assign n11717 = n11716 ^ n11574 ;
  assign n11573 = n2883 & ~n4615 ;
  assign n11718 = n11717 ^ n11573 ;
  assign n11720 = n11719 ^ n11718 ;
  assign n11724 = n11723 ^ n11720 ;
  assign n11725 = n11724 ^ x29 ;
  assign n11572 = x104 & n2581 ;
  assign n11726 = n11725 ^ n11572 ;
  assign n11571 = x106 & n2422 ;
  assign n11727 = n11726 ^ n11571 ;
  assign n11570 = n2423 & ~n5240 ;
  assign n11728 = n11727 ^ n11570 ;
  assign n11730 = n11729 ^ n11728 ;
  assign n11567 = n11464 ^ n11455 ;
  assign n11568 = n11461 & ~n11567 ;
  assign n11569 = n11568 ^ n11464 ;
  assign n11731 = n11730 ^ n11569 ;
  assign n11732 = n11731 ^ x26 ;
  assign n11566 = x107 & n2018 ;
  assign n11733 = n11732 ^ n11566 ;
  assign n11565 = x109 & n2021 ;
  assign n11734 = n11733 ^ n11565 ;
  assign n11564 = n2022 & n5902 ;
  assign n11735 = n11734 ^ n11564 ;
  assign n11737 = n11736 ^ n11735 ;
  assign n11741 = n11740 ^ n11737 ;
  assign n11742 = n11741 ^ x23 ;
  assign n11563 = x110 & n1658 ;
  assign n11743 = n11742 ^ n11563 ;
  assign n11562 = x112 & n1661 ;
  assign n11744 = n11743 ^ n11562 ;
  assign n11561 = n1662 & ~n6600 ;
  assign n11745 = n11744 ^ n11561 ;
  assign n11747 = n11746 ^ n11745 ;
  assign n11558 = n11481 ^ n11472 ;
  assign n11559 = ~n11478 & n11558 ;
  assign n11560 = n11559 ^ n11481 ;
  assign n11748 = n11747 ^ n11560 ;
  assign n11749 = n11748 ^ x20 ;
  assign n11557 = x113 & n1327 ;
  assign n11750 = n11749 ^ n11557 ;
  assign n11556 = x115 & n1330 ;
  assign n11751 = n11750 ^ n11556 ;
  assign n11555 = n1331 & ~n7343 ;
  assign n11752 = n11751 ^ n11555 ;
  assign n11754 = n11753 ^ n11752 ;
  assign n11552 = n11491 ^ n11482 ;
  assign n11553 = ~n11488 & ~n11552 ;
  assign n11554 = n11553 ^ n11491 ;
  assign n11755 = n11754 ^ n11554 ;
  assign n11756 = n11755 ^ x17 ;
  assign n11551 = x116 & n1050 ;
  assign n11757 = n11756 ^ n11551 ;
  assign n11550 = x118 & n1053 ;
  assign n11758 = n11757 ^ n11550 ;
  assign n11549 = n1054 & ~n8123 ;
  assign n11759 = n11758 ^ n11549 ;
  assign n11761 = n11760 ^ n11759 ;
  assign n11765 = n11764 ^ n11761 ;
  assign n11766 = n11765 ^ x14 ;
  assign n11548 = x119 & n877 ;
  assign n11767 = n11766 ^ n11548 ;
  assign n11547 = x121 & n782 ;
  assign n11768 = n11767 ^ n11547 ;
  assign n11546 = n783 & n8962 ;
  assign n11769 = n11768 ^ n11546 ;
  assign n11771 = n11770 ^ n11769 ;
  assign n11775 = n11774 ^ n11771 ;
  assign n11776 = n11775 ^ x11 ;
  assign n11545 = x122 & n647 ;
  assign n11777 = n11776 ^ n11545 ;
  assign n11544 = x124 & ~n572 ;
  assign n11778 = n11777 ^ n11544 ;
  assign n11543 = ~n573 & n10095 ;
  assign n11779 = n11778 ^ n11543 ;
  assign n11781 = n11780 ^ n11779 ;
  assign n11540 = n11515 ^ n11506 ;
  assign n11541 = ~n11512 & n11540 ;
  assign n11542 = n11541 ^ n11515 ;
  assign n11782 = n11781 ^ n11542 ;
  assign n11783 = n11782 ^ x8 ;
  assign n11539 = x125 & n446 ;
  assign n11784 = n11783 ^ n11539 ;
  assign n11538 = x127 & n383 ;
  assign n11785 = n11784 ^ n11538 ;
  assign n11537 = n384 & n10972 ;
  assign n11786 = n11785 ^ n11537 ;
  assign n11788 = n11787 ^ n11786 ;
  assign n11792 = n11791 ^ n11788 ;
  assign n11533 = n11527 ^ n11523 ;
  assign n11793 = n11792 ^ n11533 ;
  assign n11532 = n11262 ^ n11259 ;
  assign n11534 = n11533 ^ n11273 ;
  assign n11535 = n11534 ^ n11262 ;
  assign n11536 = n11532 & ~n11535 ;
  assign n11794 = n11793 ^ n11536 ;
  assign n11795 = n11794 ^ n11792 ;
  assign n11796 = n11795 ^ n11536 ;
  assign n11797 = n11796 ^ n11795 ;
  assign n11798 = n11795 ^ n11259 ;
  assign n11799 = n11798 ^ n11795 ;
  assign n11800 = n11797 & ~n11799 ;
  assign n11801 = n11800 ^ n11795 ;
  assign n11802 = ~n11531 & n11801 ;
  assign n11803 = n11802 ^ n11794 ;
  assign n11807 = n11806 ^ n11803 ;
  assign n12062 = n11273 & ~n11527 ;
  assign n12063 = n12062 ^ n11531 ;
  assign n12064 = n11804 ^ n11259 ;
  assign n12065 = n12064 ^ n11804 ;
  assign n12066 = n11523 ^ n11262 ;
  assign n12067 = n12066 ^ n11804 ;
  assign n12068 = ~n12065 & n12067 ;
  assign n12069 = n12068 ^ n11804 ;
  assign n12070 = ~n11792 & ~n12069 ;
  assign n12071 = n12070 ^ n12064 ;
  assign n12072 = ~n12063 & n12071 ;
  assign n12073 = n12062 ^ n11792 ;
  assign n12074 = n12062 ^ n11523 ;
  assign n12075 = n12074 ^ n11532 ;
  assign n12076 = n12075 ^ n12074 ;
  assign n12077 = n12062 ^ n11262 ;
  assign n12078 = n12077 ^ n12074 ;
  assign n12079 = n12076 & n12078 ;
  assign n12080 = n12079 ^ n12074 ;
  assign n12081 = n12073 & ~n12080 ;
  assign n12082 = n12081 ^ n11792 ;
  assign n12083 = ~n12072 & ~n12082 ;
  assign n12057 = n11775 ^ n11542 ;
  assign n12058 = n11781 & n12057 ;
  assign n12059 = n12058 ^ n11775 ;
  assign n12055 = x127 & n390 ;
  assign n12049 = x124 & n578 ;
  assign n12038 = x120 & n877 ;
  assign n12037 = x122 & n782 ;
  assign n12039 = n12038 ^ n12037 ;
  assign n12040 = n12039 ^ x14 ;
  assign n12036 = n783 & ~n9247 ;
  assign n12041 = n12040 ^ n12036 ;
  assign n12035 = x121 & n788 ;
  assign n12042 = n12041 ^ n12035 ;
  assign n12031 = n11748 ^ n11554 ;
  assign n12032 = n11754 & ~n12031 ;
  assign n12033 = n12032 ^ n11748 ;
  assign n12029 = x118 & n1058 ;
  assign n12021 = n11741 ^ n11560 ;
  assign n12022 = n11747 & n12021 ;
  assign n12023 = n12022 ^ n11741 ;
  assign n12019 = x115 & n1335 ;
  assign n12012 = x112 & n1666 ;
  assign n12004 = n11724 ^ n11569 ;
  assign n12005 = ~n11730 & ~n12004 ;
  assign n12006 = n12005 ^ n11724 ;
  assign n12002 = x109 & n2014 ;
  assign n11995 = x106 & n2429 ;
  assign n11988 = x103 & n2887 ;
  assign n11980 = n11700 ^ n11584 ;
  assign n11981 = n11706 & ~n11980 ;
  assign n11982 = n11981 ^ n11700 ;
  assign n11978 = x100 & n3383 ;
  assign n11970 = n11693 ^ n11590 ;
  assign n11971 = n11699 & n11970 ;
  assign n11972 = n11971 ^ n11693 ;
  assign n11968 = x97 & n3924 ;
  assign n11960 = n11686 ^ n11596 ;
  assign n11961 = n11692 & n11960 ;
  assign n11962 = n11961 ^ n11686 ;
  assign n11958 = x94 & n4467 ;
  assign n11950 = n11685 ^ n11672 ;
  assign n11951 = n11677 & n11950 ;
  assign n11952 = n11951 ^ n11672 ;
  assign n11944 = x90 & n5094 ;
  assign n11943 = x92 & n5097 ;
  assign n11945 = n11944 ^ n11943 ;
  assign n11946 = n11945 ^ x44 ;
  assign n11942 = n2684 & n5098 ;
  assign n11947 = n11946 ^ n11942 ;
  assign n11941 = x91 & n5102 ;
  assign n11948 = n11947 ^ n11941 ;
  assign n11937 = n11665 ^ n11602 ;
  assign n11938 = n11671 & n11937 ;
  assign n11939 = n11938 ^ n11665 ;
  assign n11931 = x87 & n5965 ;
  assign n11930 = x89 & n5729 ;
  assign n11932 = n11931 ^ n11930 ;
  assign n11933 = n11932 ^ x47 ;
  assign n11929 = n2249 & n5730 ;
  assign n11934 = n11933 ^ n11929 ;
  assign n11928 = x88 & n5736 ;
  assign n11935 = n11934 ^ n11928 ;
  assign n11921 = x84 & n6677 ;
  assign n11920 = x86 & n6428 ;
  assign n11922 = n11921 ^ n11920 ;
  assign n11923 = n11922 ^ x50 ;
  assign n11919 = n1857 & n6429 ;
  assign n11924 = n11923 ^ n11919 ;
  assign n11918 = x85 & n6433 ;
  assign n11925 = n11924 ^ n11918 ;
  assign n11911 = x81 & n7171 ;
  assign n11910 = x83 & n7174 ;
  assign n11912 = n11911 ^ n11910 ;
  assign n11913 = n11912 ^ x53 ;
  assign n11909 = n1512 & n7175 ;
  assign n11914 = n11913 ^ n11909 ;
  assign n11908 = x82 & n7179 ;
  assign n11915 = n11914 ^ n11908 ;
  assign n11905 = x79 & n7931 ;
  assign n11894 = x75 & n8741 ;
  assign n11893 = x77 & n8744 ;
  assign n11895 = n11894 ^ n11893 ;
  assign n11896 = n11895 ^ x59 ;
  assign n11892 = ~n939 & n8745 ;
  assign n11897 = n11896 ^ n11892 ;
  assign n11891 = x76 & n8737 ;
  assign n11898 = n11897 ^ n11891 ;
  assign n11885 = x72 & n9632 ;
  assign n11884 = x74 & n9635 ;
  assign n11886 = n11885 ^ n11884 ;
  assign n11887 = n11886 ^ x62 ;
  assign n11883 = n699 & n9636 ;
  assign n11888 = n11887 ^ n11883 ;
  assign n11882 = x73 & n9628 ;
  assign n11889 = n11888 ^ n11882 ;
  assign n11877 = n11628 ^ x5 ;
  assign n11878 = n11625 & n11877 ;
  assign n11879 = n11878 ^ x2 ;
  assign n11874 = x62 & ~x63 ;
  assign n11875 = n11874 ^ x62 ;
  assign n11876 = x70 & n11875 ;
  assign n11880 = n11879 ^ n11876 ;
  assign n11873 = x71 & n9948 ;
  assign n11881 = n11880 ^ n11873 ;
  assign n11890 = n11889 ^ n11881 ;
  assign n11899 = n11898 ^ n11890 ;
  assign n11870 = n11643 ^ n11634 ;
  assign n11871 = ~n11635 & n11870 ;
  assign n11872 = n11871 ^ n11643 ;
  assign n11900 = n11899 ^ n11872 ;
  assign n11901 = n11900 ^ x56 ;
  assign n11869 = x78 & n7935 ;
  assign n11902 = n11901 ^ n11869 ;
  assign n11868 = x80 & n7938 ;
  assign n11903 = n11902 ^ n11868 ;
  assign n11867 = n1206 & n7939 ;
  assign n11904 = n11903 ^ n11867 ;
  assign n11906 = n11905 ^ n11904 ;
  assign n11864 = n11644 ^ n11621 ;
  assign n11865 = n11650 & n11864 ;
  assign n11866 = n11865 ^ n11644 ;
  assign n11907 = n11906 ^ n11866 ;
  assign n11916 = n11915 ^ n11907 ;
  assign n11861 = n11651 ^ n11613 ;
  assign n11862 = n11618 & n11861 ;
  assign n11863 = n11862 ^ n11613 ;
  assign n11917 = n11916 ^ n11863 ;
  assign n11926 = n11925 ^ n11917 ;
  assign n11858 = n11664 ^ n11660 ;
  assign n11859 = ~n11661 & n11858 ;
  assign n11860 = n11859 ^ n11664 ;
  assign n11927 = n11926 ^ n11860 ;
  assign n11936 = n11935 ^ n11927 ;
  assign n11940 = n11939 ^ n11936 ;
  assign n11949 = n11948 ^ n11940 ;
  assign n11953 = n11952 ^ n11949 ;
  assign n11954 = n11953 ^ x41 ;
  assign n11857 = x93 & n4474 ;
  assign n11955 = n11954 ^ n11857 ;
  assign n11856 = x95 & n4471 ;
  assign n11956 = n11955 ^ n11856 ;
  assign n11855 = n3159 & n4472 ;
  assign n11957 = n11956 ^ n11855 ;
  assign n11959 = n11958 ^ n11957 ;
  assign n11963 = n11962 ^ n11959 ;
  assign n11964 = n11963 ^ x38 ;
  assign n11854 = x96 & n3916 ;
  assign n11965 = n11964 ^ n11854 ;
  assign n11853 = x98 & n3919 ;
  assign n11966 = n11965 ^ n11853 ;
  assign n11852 = n3660 & n3920 ;
  assign n11967 = n11966 ^ n11852 ;
  assign n11969 = n11968 ^ n11967 ;
  assign n11973 = n11972 ^ n11969 ;
  assign n11974 = n11973 ^ x35 ;
  assign n11851 = x99 & n3375 ;
  assign n11975 = n11974 ^ n11851 ;
  assign n11850 = x101 & n3378 ;
  assign n11976 = n11975 ^ n11850 ;
  assign n11849 = n3379 & n4215 ;
  assign n11977 = n11976 ^ n11849 ;
  assign n11979 = n11978 ^ n11977 ;
  assign n11983 = n11982 ^ n11979 ;
  assign n11984 = n11983 ^ x32 ;
  assign n11848 = x102 & n2879 ;
  assign n11985 = n11984 ^ n11848 ;
  assign n11847 = x104 & n2882 ;
  assign n11986 = n11985 ^ n11847 ;
  assign n11846 = n2883 & ~n4814 ;
  assign n11987 = n11986 ^ n11846 ;
  assign n11989 = n11988 ^ n11987 ;
  assign n11843 = n11707 ^ n11578 ;
  assign n11844 = ~n11713 & n11843 ;
  assign n11845 = n11844 ^ n11707 ;
  assign n11990 = n11989 ^ n11845 ;
  assign n11991 = n11990 ^ x29 ;
  assign n11842 = x105 & n2581 ;
  assign n11992 = n11991 ^ n11842 ;
  assign n11841 = x107 & n2422 ;
  assign n11993 = n11992 ^ n11841 ;
  assign n11840 = n2423 & ~n5448 ;
  assign n11994 = n11993 ^ n11840 ;
  assign n11996 = n11995 ^ n11994 ;
  assign n11837 = n11723 ^ n11714 ;
  assign n11838 = ~n11720 & ~n11837 ;
  assign n11839 = n11838 ^ n11723 ;
  assign n11997 = n11996 ^ n11839 ;
  assign n11998 = n11997 ^ x26 ;
  assign n11836 = x108 & n2018 ;
  assign n11999 = n11998 ^ n11836 ;
  assign n11835 = x110 & n2021 ;
  assign n12000 = n11999 ^ n11835 ;
  assign n11834 = n2022 & n6129 ;
  assign n12001 = n12000 ^ n11834 ;
  assign n12003 = n12002 ^ n12001 ;
  assign n12007 = n12006 ^ n12003 ;
  assign n12008 = n12007 ^ x23 ;
  assign n11833 = x111 & n1658 ;
  assign n12009 = n12008 ^ n11833 ;
  assign n11832 = x113 & n1661 ;
  assign n12010 = n12009 ^ n11832 ;
  assign n11831 = n1662 & ~n6839 ;
  assign n12011 = n12010 ^ n11831 ;
  assign n12013 = n12012 ^ n12011 ;
  assign n11828 = n11740 ^ n11731 ;
  assign n11829 = n11737 & n11828 ;
  assign n11830 = n11829 ^ n11740 ;
  assign n12014 = n12013 ^ n11830 ;
  assign n12015 = n12014 ^ x20 ;
  assign n11827 = x114 & n1327 ;
  assign n12016 = n12015 ^ n11827 ;
  assign n11826 = x116 & n1330 ;
  assign n12017 = n12016 ^ n11826 ;
  assign n11825 = n1331 & ~n7588 ;
  assign n12018 = n12017 ^ n11825 ;
  assign n12020 = n12019 ^ n12018 ;
  assign n12024 = n12023 ^ n12020 ;
  assign n12025 = n12024 ^ x17 ;
  assign n11824 = x117 & n1050 ;
  assign n12026 = n12025 ^ n11824 ;
  assign n11823 = x119 & n1053 ;
  assign n12027 = n12026 ^ n11823 ;
  assign n11822 = n1054 & n8394 ;
  assign n12028 = n12027 ^ n11822 ;
  assign n12030 = n12029 ^ n12028 ;
  assign n12034 = n12033 ^ n12030 ;
  assign n12043 = n12042 ^ n12034 ;
  assign n11819 = n11764 ^ n11755 ;
  assign n11820 = n11761 & n11819 ;
  assign n11821 = n11820 ^ n11764 ;
  assign n12044 = n12043 ^ n11821 ;
  assign n12045 = n12044 ^ x11 ;
  assign n11818 = x123 & n647 ;
  assign n12046 = n12045 ^ n11818 ;
  assign n11817 = x125 & ~n572 ;
  assign n12047 = n12046 ^ n11817 ;
  assign n11816 = ~n573 & n10400 ;
  assign n12048 = n12047 ^ n11816 ;
  assign n12050 = n12049 ^ n12048 ;
  assign n11813 = n11774 ^ n11765 ;
  assign n11814 = ~n11771 & n11813 ;
  assign n11815 = n11814 ^ n11774 ;
  assign n12051 = n12050 ^ n11815 ;
  assign n12052 = n12051 ^ x8 ;
  assign n11812 = x126 & n446 ;
  assign n12053 = n12052 ^ n11812 ;
  assign n11811 = n384 & n10139 ;
  assign n12054 = n12053 ^ n11811 ;
  assign n12056 = n12055 ^ n12054 ;
  assign n12060 = n12059 ^ n12056 ;
  assign n11808 = n11791 ^ n11782 ;
  assign n11809 = ~n11788 & n11808 ;
  assign n11810 = n11809 ^ n11791 ;
  assign n12061 = n12060 ^ n11810 ;
  assign n12084 = n12083 ^ n12061 ;
  assign n12348 = n12044 ^ n11815 ;
  assign n12349 = ~n12050 & ~n12348 ;
  assign n12350 = n12349 ^ n12044 ;
  assign n12343 = n12042 ^ n11821 ;
  assign n12344 = n12043 & ~n12343 ;
  assign n12345 = n12344 ^ n12042 ;
  assign n12341 = x125 & n578 ;
  assign n12334 = x122 & n788 ;
  assign n12327 = x119 & n1058 ;
  assign n12319 = n12007 ^ n11830 ;
  assign n12320 = ~n12013 & n12319 ;
  assign n12321 = n12320 ^ n12007 ;
  assign n12317 = x116 & n1335 ;
  assign n12310 = x113 & n1666 ;
  assign n12302 = n11990 ^ n11839 ;
  assign n12303 = ~n11996 & n12302 ;
  assign n12304 = n12303 ^ n11990 ;
  assign n12300 = x110 & n2014 ;
  assign n12293 = x107 & n2429 ;
  assign n12286 = x104 & n2887 ;
  assign n12279 = x101 & n3383 ;
  assign n12272 = x98 & n3924 ;
  assign n12261 = x94 & n4474 ;
  assign n12260 = x96 & n4471 ;
  assign n12262 = n12261 ^ n12260 ;
  assign n12263 = n12262 ^ x41 ;
  assign n12259 = n3323 & n4472 ;
  assign n12264 = n12263 ^ n12259 ;
  assign n12258 = x95 & n4467 ;
  assign n12265 = n12264 ^ n12258 ;
  assign n12251 = x91 & n5094 ;
  assign n12250 = x93 & n5097 ;
  assign n12252 = n12251 ^ n12250 ;
  assign n12253 = n12252 ^ x44 ;
  assign n12249 = n2836 & n5098 ;
  assign n12254 = n12253 ^ n12249 ;
  assign n12248 = x92 & n5102 ;
  assign n12255 = n12254 ^ n12248 ;
  assign n12240 = x85 & n6677 ;
  assign n12239 = x87 & n6428 ;
  assign n12241 = n12240 ^ n12239 ;
  assign n12242 = n12241 ^ x50 ;
  assign n12238 = n1982 & n6429 ;
  assign n12243 = n12242 ^ n12238 ;
  assign n12237 = x86 & n6433 ;
  assign n12244 = n12243 ^ n12237 ;
  assign n12230 = x82 & n7171 ;
  assign n12229 = x84 & n7174 ;
  assign n12231 = n12230 ^ n12229 ;
  assign n12232 = n12231 ^ x53 ;
  assign n12228 = n1624 & n7175 ;
  assign n12233 = n12232 ^ n12228 ;
  assign n12227 = x83 & n7179 ;
  assign n12234 = n12233 ^ n12227 ;
  assign n12223 = n11898 ^ n11872 ;
  assign n12224 = n11899 & n12223 ;
  assign n12225 = n12224 ^ n11898 ;
  assign n12217 = x79 & n7935 ;
  assign n12216 = x81 & n7938 ;
  assign n12218 = n12217 ^ n12216 ;
  assign n12219 = n12218 ^ x56 ;
  assign n12215 = n1305 & n7939 ;
  assign n12220 = n12219 ^ n12215 ;
  assign n12214 = x80 & n7931 ;
  assign n12221 = n12220 ^ n12214 ;
  assign n12201 = ~x72 & n9948 ;
  assign n12202 = n12201 ^ n11876 ;
  assign n12203 = x71 & n12202 ;
  assign n12204 = n12203 ^ n11876 ;
  assign n12205 = n9948 ^ x71 ;
  assign n12206 = n11874 ^ x63 ;
  assign n12207 = n12206 ^ n12202 ;
  assign n12208 = n12205 & n12207 ;
  assign n12432 = ~n12204 & ~n12208 ;
  assign n12198 = n11889 ^ n11879 ;
  assign n12199 = ~n11881 & ~n12198 ;
  assign n12200 = n12199 ^ n11889 ;
  assign n12212 = ~n12432 ^ n12200 ;
  assign n12195 = ~n1025 & n8745 ;
  assign n12193 = x76 & n8741 ;
  assign n12187 = x73 & n9632 ;
  assign n12186 = x75 & n9635 ;
  assign n12188 = n12187 ^ n12186 ;
  assign n12189 = n12188 ^ x62 ;
  assign n12185 = ~n774 & n9636 ;
  assign n12190 = n12189 ^ n12185 ;
  assign n12184 = x74 & n9628 ;
  assign n12191 = n12190 ^ n12184 ;
  assign n12182 = x78 & n8744 ;
  assign n12183 = n12182 ^ x59 ;
  assign n12192 = n12191 ^ n12183 ;
  assign n12194 = n12193 ^ n12192 ;
  assign n12196 = n12195 ^ n12194 ;
  assign n12181 = x77 & n8737 ;
  assign n12197 = n12196 ^ n12181 ;
  assign n12213 = n12212 ^ n12197 ;
  assign n12222 = n12221 ^ n12213 ;
  assign n12226 = n12225 ^ n12222 ;
  assign n12235 = n12234 ^ n12226 ;
  assign n12178 = n11900 ^ n11866 ;
  assign n12179 = n11906 & n12178 ;
  assign n12180 = n12179 ^ n11900 ;
  assign n12236 = n12235 ^ n12180 ;
  assign n12245 = n12244 ^ n12236 ;
  assign n12175 = n11915 ^ n11863 ;
  assign n12176 = n11916 & n12175 ;
  assign n12177 = n12176 ^ n11915 ;
  assign n12246 = n12245 ^ n12177 ;
  assign n12172 = n2386 & n5730 ;
  assign n12170 = x88 & n5965 ;
  assign n12166 = n11925 ^ n11860 ;
  assign n12167 = n11926 & n12166 ;
  assign n12168 = n12167 ^ n11925 ;
  assign n12164 = x90 & n5729 ;
  assign n12165 = n12164 ^ x47 ;
  assign n12169 = n12168 ^ n12165 ;
  assign n12171 = n12170 ^ n12169 ;
  assign n12173 = n12172 ^ n12171 ;
  assign n12163 = x89 & n5736 ;
  assign n12174 = n12173 ^ n12163 ;
  assign n12247 = n12246 ^ n12174 ;
  assign n12256 = n12255 ^ n12247 ;
  assign n12160 = n11939 ^ n11935 ;
  assign n12161 = ~n11936 & n12160 ;
  assign n12162 = n12161 ^ n11939 ;
  assign n12257 = n12256 ^ n12162 ;
  assign n12266 = n12265 ^ n12257 ;
  assign n12157 = n11952 ^ n11948 ;
  assign n12158 = ~n11949 & n12157 ;
  assign n12159 = n12158 ^ n11952 ;
  assign n12267 = n12266 ^ n12159 ;
  assign n12268 = n12267 ^ x38 ;
  assign n12156 = x97 & n3916 ;
  assign n12269 = n12268 ^ n12156 ;
  assign n12155 = x99 & n3919 ;
  assign n12270 = n12269 ^ n12155 ;
  assign n12154 = n3843 & n3920 ;
  assign n12271 = n12270 ^ n12154 ;
  assign n12273 = n12272 ^ n12271 ;
  assign n12151 = n11962 ^ n11953 ;
  assign n12152 = ~n11959 & n12151 ;
  assign n12153 = n12152 ^ n11962 ;
  assign n12274 = n12273 ^ n12153 ;
  assign n12275 = n12274 ^ x35 ;
  assign n12150 = x100 & n3375 ;
  assign n12276 = n12275 ^ n12150 ;
  assign n12149 = x102 & n3378 ;
  assign n12277 = n12276 ^ n12149 ;
  assign n12148 = n3379 & n4410 ;
  assign n12278 = n12277 ^ n12148 ;
  assign n12280 = n12279 ^ n12278 ;
  assign n12145 = n11972 ^ n11963 ;
  assign n12146 = ~n11969 & n12145 ;
  assign n12147 = n12146 ^ n11972 ;
  assign n12281 = n12280 ^ n12147 ;
  assign n12282 = n12281 ^ x32 ;
  assign n12144 = x103 & n2879 ;
  assign n12283 = n12282 ^ n12144 ;
  assign n12143 = x105 & n2882 ;
  assign n12284 = n12283 ^ n12143 ;
  assign n12142 = n2883 & ~n5023 ;
  assign n12285 = n12284 ^ n12142 ;
  assign n12287 = n12286 ^ n12285 ;
  assign n12139 = n11982 ^ n11973 ;
  assign n12140 = ~n11979 & n12139 ;
  assign n12141 = n12140 ^ n11982 ;
  assign n12288 = n12287 ^ n12141 ;
  assign n12289 = n12288 ^ x29 ;
  assign n12138 = x106 & n2581 ;
  assign n12290 = n12289 ^ n12138 ;
  assign n12137 = x108 & n2422 ;
  assign n12291 = n12290 ^ n12137 ;
  assign n12136 = n2423 & n5670 ;
  assign n12292 = n12291 ^ n12136 ;
  assign n12294 = n12293 ^ n12292 ;
  assign n12133 = n11983 ^ n11845 ;
  assign n12134 = n11989 & ~n12133 ;
  assign n12135 = n12134 ^ n11983 ;
  assign n12295 = n12294 ^ n12135 ;
  assign n12296 = n12295 ^ x26 ;
  assign n12132 = x109 & n2018 ;
  assign n12297 = n12296 ^ n12132 ;
  assign n12131 = x111 & n2021 ;
  assign n12298 = n12297 ^ n12131 ;
  assign n12130 = n2022 & ~n6360 ;
  assign n12299 = n12298 ^ n12130 ;
  assign n12301 = n12300 ^ n12299 ;
  assign n12305 = n12304 ^ n12301 ;
  assign n12306 = n12305 ^ x23 ;
  assign n12129 = x112 & n1658 ;
  assign n12307 = n12306 ^ n12129 ;
  assign n12128 = x114 & n1661 ;
  assign n12308 = n12307 ^ n12128 ;
  assign n12127 = n1662 & ~n7092 ;
  assign n12309 = n12308 ^ n12127 ;
  assign n12311 = n12310 ^ n12309 ;
  assign n12124 = n12006 ^ n11997 ;
  assign n12125 = ~n12003 & ~n12124 ;
  assign n12126 = n12125 ^ n12006 ;
  assign n12312 = n12311 ^ n12126 ;
  assign n12313 = n12312 ^ x20 ;
  assign n12123 = x115 & n1327 ;
  assign n12314 = n12313 ^ n12123 ;
  assign n12122 = x117 & n1330 ;
  assign n12315 = n12314 ^ n12122 ;
  assign n12121 = n1331 & ~n7850 ;
  assign n12316 = n12315 ^ n12121 ;
  assign n12318 = n12317 ^ n12316 ;
  assign n12322 = n12321 ^ n12318 ;
  assign n12323 = n12322 ^ x17 ;
  assign n12120 = x118 & n1050 ;
  assign n12324 = n12323 ^ n12120 ;
  assign n12119 = x120 & n1053 ;
  assign n12325 = n12324 ^ n12119 ;
  assign n12118 = n1054 & n8891 ;
  assign n12326 = n12325 ^ n12118 ;
  assign n12328 = n12327 ^ n12326 ;
  assign n12115 = n12023 ^ n12014 ;
  assign n12116 = ~n12020 & n12115 ;
  assign n12117 = n12116 ^ n12023 ;
  assign n12329 = n12328 ^ n12117 ;
  assign n12330 = n12329 ^ x14 ;
  assign n12114 = x121 & n877 ;
  assign n12331 = n12330 ^ n12114 ;
  assign n12113 = x123 & n782 ;
  assign n12332 = n12331 ^ n12113 ;
  assign n12112 = n783 & ~n9786 ;
  assign n12333 = n12332 ^ n12112 ;
  assign n12335 = n12334 ^ n12333 ;
  assign n12109 = n12033 ^ n12024 ;
  assign n12110 = ~n12030 & n12109 ;
  assign n12111 = n12110 ^ n12033 ;
  assign n12336 = n12335 ^ n12111 ;
  assign n12337 = n12336 ^ x11 ;
  assign n12108 = x124 & n647 ;
  assign n12338 = n12337 ^ n12108 ;
  assign n12107 = x126 & ~n572 ;
  assign n12339 = n12338 ^ n12107 ;
  assign n12106 = ~n573 & n10441 ;
  assign n12340 = n12339 ^ n12106 ;
  assign n12342 = n12341 ^ n12340 ;
  assign n12346 = n12345 ^ n12342 ;
  assign n12093 = ~x7 & x127 ;
  assign n12094 = n12093 ^ x8 ;
  assign n12095 = ~n10138 & ~n12094 ;
  assign n12096 = n12095 ^ x8 ;
  assign n12097 = n329 & ~n12096 ;
  assign n12098 = n328 ^ x8 ;
  assign n12101 = x127 & n382 ;
  assign n12102 = ~n12098 & n12101 ;
  assign n12103 = n12102 ^ n12098 ;
  assign n12104 = n12103 ^ n328 ;
  assign n12105 = ~n12097 & n12104 ;
  assign n12347 = n12346 ^ n12105 ;
  assign n12351 = n12350 ^ n12347 ;
  assign n12088 = n12059 ^ n12051 ;
  assign n12089 = n12056 & ~n12088 ;
  assign n12090 = n12089 ^ n12059 ;
  assign n12352 = n12351 ^ n12090 ;
  assign n12085 = n12083 ^ n11810 ;
  assign n12086 = n12061 & ~n12085 ;
  assign n12087 = n12086 ^ n12083 ;
  assign n12353 = n12352 ^ n12087 ;
  assign n12354 = n12350 ^ n12346 ;
  assign n12355 = ~n12347 & ~n12354 ;
  assign n12599 = n12355 ^ n12347 ;
  assign n12591 = x125 & n647 ;
  assign n12590 = x127 & ~n572 ;
  assign n12592 = n12591 ^ n12590 ;
  assign n12593 = n12592 ^ x11 ;
  assign n12589 = ~n573 & n10972 ;
  assign n12594 = n12593 ^ n12589 ;
  assign n12588 = x126 & n578 ;
  assign n12595 = n12594 ^ n12588 ;
  assign n12584 = n12329 ^ n12111 ;
  assign n12585 = n12335 & n12584 ;
  assign n12586 = n12585 ^ n12329 ;
  assign n12582 = x123 & n788 ;
  assign n12574 = n12322 ^ n12117 ;
  assign n12575 = n12328 & n12574 ;
  assign n12576 = n12575 ^ n12322 ;
  assign n12572 = x120 & n1058 ;
  assign n12565 = x117 & n1335 ;
  assign n12557 = n12305 ^ n12126 ;
  assign n12558 = n12311 & ~n12557 ;
  assign n12559 = n12558 ^ n12305 ;
  assign n12555 = x114 & n1666 ;
  assign n12548 = x111 & n2014 ;
  assign n12541 = x108 & n2429 ;
  assign n12533 = n12281 ^ n12141 ;
  assign n12534 = ~n12287 & ~n12533 ;
  assign n12535 = n12534 ^ n12281 ;
  assign n12531 = x105 & n2887 ;
  assign n12523 = n12274 ^ n12147 ;
  assign n12524 = ~n12280 & ~n12523 ;
  assign n12525 = n12524 ^ n12274 ;
  assign n12521 = x102 & n3383 ;
  assign n12513 = n12267 ^ n12153 ;
  assign n12514 = ~n12273 & ~n12513 ;
  assign n12515 = n12514 ^ n12267 ;
  assign n12511 = x99 & n3924 ;
  assign n12503 = n12265 ^ n12159 ;
  assign n12504 = ~n12266 & n12503 ;
  assign n12505 = n12504 ^ n12265 ;
  assign n12497 = x95 & n4474 ;
  assign n12496 = x97 & n4471 ;
  assign n12498 = n12497 ^ n12496 ;
  assign n12499 = n12498 ^ x41 ;
  assign n12495 = n3494 & n4472 ;
  assign n12500 = n12499 ^ n12495 ;
  assign n12494 = x96 & n4467 ;
  assign n12501 = n12500 ^ n12494 ;
  assign n12488 = x92 & n5094 ;
  assign n12487 = x94 & n5097 ;
  assign n12489 = n12488 ^ n12487 ;
  assign n12490 = n12489 ^ x44 ;
  assign n12486 = n2997 & n5098 ;
  assign n12491 = n12490 ^ n12486 ;
  assign n12485 = x93 & n5102 ;
  assign n12492 = n12491 ^ n12485 ;
  assign n12482 = n12247 ^ n12162 ;
  assign n12483 = ~n12256 & ~n12482 ;
  assign n12473 = x89 & n5965 ;
  assign n12472 = x91 & n5729 ;
  assign n12474 = n12473 ^ n12472 ;
  assign n12475 = n12474 ^ x47 ;
  assign n12471 = n2542 & n5730 ;
  assign n12476 = n12475 ^ n12471 ;
  assign n12470 = x90 & n5736 ;
  assign n12477 = n12476 ^ n12470 ;
  assign n12466 = n12244 ^ n12177 ;
  assign n12467 = ~n12245 & n12466 ;
  assign n12468 = n12467 ^ n12244 ;
  assign n12460 = x86 & n6677 ;
  assign n12459 = x88 & n6428 ;
  assign n12461 = n12460 ^ n12459 ;
  assign n12462 = n12461 ^ x50 ;
  assign n12458 = n2119 & n6429 ;
  assign n12463 = n12462 ^ n12458 ;
  assign n12457 = x87 & n6433 ;
  assign n12464 = n12463 ^ n12457 ;
  assign n12453 = n12234 ^ n12180 ;
  assign n12454 = ~n12235 & n12453 ;
  assign n12455 = n12454 ^ n12234 ;
  assign n12451 = x84 & n7179 ;
  assign n12444 = x81 & n7931 ;
  assign n12442 = n1411 & n7939 ;
  assign n12438 = x80 & n7935 ;
  assign n12437 = x82 & n7938 ;
  assign n12439 = n12438 ^ n12437 ;
  assign n12440 = n12439 ^ x56 ;
  assign n12433 = ~n12200 & n12432 ;
  assign n12434 = n12433 ^ n12208 ;
  assign n12425 = x74 & n9632 ;
  assign n12424 = x76 & n9635 ;
  assign n12426 = n12425 ^ n12424 ;
  assign n12427 = n12426 ^ x62 ;
  assign n12423 = ~n853 & n9636 ;
  assign n12428 = n12427 ^ n12423 ;
  assign n12422 = x75 & n9628 ;
  assign n12429 = n12428 ^ n12422 ;
  assign n12430 = n12429 ^ x8 ;
  assign n12418 = x73 ^ x71 ;
  assign n12419 = ~n11875 & n12418 ;
  assign n12420 = n12419 ^ n416 ;
  assign n12421 = n12206 & n12420 ;
  assign n12431 = n12430 ^ n12421 ;
  assign n12435 = n12434 ^ n12431 ;
  assign n12408 = x77 & n8741 ;
  assign n12407 = x79 & n8744 ;
  assign n12409 = n12408 ^ n12407 ;
  assign n12410 = n12409 ^ x59 ;
  assign n12406 = n1118 & n8745 ;
  assign n12411 = n12410 ^ n12406 ;
  assign n12405 = x78 & n8737 ;
  assign n12412 = n12411 ^ n12405 ;
  assign n12413 = n12412 ^ n12212 ;
  assign n12414 = n12413 ^ n12191 ;
  assign n12415 = n12414 ^ n12412 ;
  assign n12416 = ~n12197 & ~n12415 ;
  assign n12417 = n12416 ^ n12413 ;
  assign n12436 = n12435 ^ n12417 ;
  assign n12441 = n12440 ^ n12436 ;
  assign n12443 = n12442 ^ n12441 ;
  assign n12445 = n12444 ^ n12443 ;
  assign n12402 = n12225 ^ n12221 ;
  assign n12403 = n12222 & n12402 ;
  assign n12404 = n12403 ^ n12225 ;
  assign n12446 = n12445 ^ n12404 ;
  assign n12447 = n12446 ^ x53 ;
  assign n12401 = x83 & n7171 ;
  assign n12448 = n12447 ^ n12401 ;
  assign n12400 = x85 & n7174 ;
  assign n12449 = n12448 ^ n12400 ;
  assign n12399 = n1743 & n7175 ;
  assign n12450 = n12449 ^ n12399 ;
  assign n12452 = n12451 ^ n12450 ;
  assign n12456 = n12455 ^ n12452 ;
  assign n12465 = n12464 ^ n12456 ;
  assign n12469 = n12468 ^ n12465 ;
  assign n12478 = n12477 ^ n12469 ;
  assign n12396 = n12246 ^ n12168 ;
  assign n12397 = ~n12174 & ~n12396 ;
  assign n12398 = n12397 ^ n12246 ;
  assign n12479 = n12478 ^ n12398 ;
  assign n12480 = n12479 ^ n12247 ;
  assign n12484 = n12483 ^ n12480 ;
  assign n12493 = n12492 ^ n12484 ;
  assign n12502 = n12501 ^ n12493 ;
  assign n12506 = n12505 ^ n12502 ;
  assign n12507 = n12506 ^ x38 ;
  assign n12395 = x98 & n3916 ;
  assign n12508 = n12507 ^ n12395 ;
  assign n12394 = x100 & n3919 ;
  assign n12509 = n12508 ^ n12394 ;
  assign n12393 = n3920 & n4034 ;
  assign n12510 = n12509 ^ n12393 ;
  assign n12512 = n12511 ^ n12510 ;
  assign n12516 = n12515 ^ n12512 ;
  assign n12517 = n12516 ^ x35 ;
  assign n12392 = x101 & n3375 ;
  assign n12518 = n12517 ^ n12392 ;
  assign n12391 = x103 & n3378 ;
  assign n12519 = n12518 ^ n12391 ;
  assign n12390 = n3379 & ~n4615 ;
  assign n12520 = n12519 ^ n12390 ;
  assign n12522 = n12521 ^ n12520 ;
  assign n12526 = n12525 ^ n12522 ;
  assign n12527 = n12526 ^ x32 ;
  assign n12389 = x104 & n2879 ;
  assign n12528 = n12527 ^ n12389 ;
  assign n12388 = x106 & n2882 ;
  assign n12529 = n12528 ^ n12388 ;
  assign n12387 = n2883 & ~n5240 ;
  assign n12530 = n12529 ^ n12387 ;
  assign n12532 = n12531 ^ n12530 ;
  assign n12536 = n12535 ^ n12532 ;
  assign n12537 = n12536 ^ x29 ;
  assign n12386 = x107 & n2581 ;
  assign n12538 = n12537 ^ n12386 ;
  assign n12385 = x109 & n2422 ;
  assign n12539 = n12538 ^ n12385 ;
  assign n12384 = n2423 & n5902 ;
  assign n12540 = n12539 ^ n12384 ;
  assign n12542 = n12541 ^ n12540 ;
  assign n12381 = n12288 ^ n12135 ;
  assign n12382 = ~n12294 & ~n12381 ;
  assign n12383 = n12382 ^ n12288 ;
  assign n12543 = n12542 ^ n12383 ;
  assign n12544 = n12543 ^ x26 ;
  assign n12380 = x110 & n2018 ;
  assign n12545 = n12544 ^ n12380 ;
  assign n12379 = x112 & n2021 ;
  assign n12546 = n12545 ^ n12379 ;
  assign n12378 = n2022 & ~n6600 ;
  assign n12547 = n12546 ^ n12378 ;
  assign n12549 = n12548 ^ n12547 ;
  assign n12375 = n12304 ^ n12295 ;
  assign n12376 = n12301 & n12375 ;
  assign n12377 = n12376 ^ n12304 ;
  assign n12550 = n12549 ^ n12377 ;
  assign n12551 = n12550 ^ x23 ;
  assign n12374 = x113 & n1658 ;
  assign n12552 = n12551 ^ n12374 ;
  assign n12373 = x115 & n1661 ;
  assign n12553 = n12552 ^ n12373 ;
  assign n12372 = n1662 & ~n7343 ;
  assign n12554 = n12553 ^ n12372 ;
  assign n12556 = n12555 ^ n12554 ;
  assign n12560 = n12559 ^ n12556 ;
  assign n12561 = n12560 ^ x20 ;
  assign n12371 = x116 & n1327 ;
  assign n12562 = n12561 ^ n12371 ;
  assign n12370 = x118 & n1330 ;
  assign n12563 = n12562 ^ n12370 ;
  assign n12369 = n1331 & ~n8123 ;
  assign n12564 = n12563 ^ n12369 ;
  assign n12566 = n12565 ^ n12564 ;
  assign n12366 = n12321 ^ n12312 ;
  assign n12367 = n12318 & n12366 ;
  assign n12368 = n12367 ^ n12321 ;
  assign n12567 = n12566 ^ n12368 ;
  assign n12568 = n12567 ^ x17 ;
  assign n12365 = x119 & n1050 ;
  assign n12569 = n12568 ^ n12365 ;
  assign n12364 = x121 & n1053 ;
  assign n12570 = n12569 ^ n12364 ;
  assign n12363 = n1054 & n8962 ;
  assign n12571 = n12570 ^ n12363 ;
  assign n12573 = n12572 ^ n12571 ;
  assign n12577 = n12576 ^ n12573 ;
  assign n12578 = n12577 ^ x14 ;
  assign n12362 = x122 & n877 ;
  assign n12579 = n12578 ^ n12362 ;
  assign n12361 = x124 & n782 ;
  assign n12580 = n12579 ^ n12361 ;
  assign n12360 = n783 & n10095 ;
  assign n12581 = n12580 ^ n12360 ;
  assign n12583 = n12582 ^ n12581 ;
  assign n12587 = n12586 ^ n12583 ;
  assign n12596 = n12595 ^ n12587 ;
  assign n12357 = n12345 ^ n12336 ;
  assign n12358 = ~n12342 & n12357 ;
  assign n12359 = n12358 ^ n12345 ;
  assign n12597 = n12596 ^ n12359 ;
  assign n12600 = n12599 ^ n12597 ;
  assign n12356 = n12355 ^ n12350 ;
  assign n12598 = n12597 ^ n12356 ;
  assign n12601 = n12600 ^ n12598 ;
  assign n12602 = n12601 ^ n12090 ;
  assign n12603 = n12090 ^ n12087 ;
  assign n12604 = ~n12602 & n12603 ;
  assign n12605 = n12604 ^ n12600 ;
  assign n12853 = n12597 ^ n12346 ;
  assign n12854 = n12354 & ~n12853 ;
  assign n12855 = n12597 ^ n12105 ;
  assign n12856 = n12854 & ~n12855 ;
  assign n12857 = n12856 ^ n12597 ;
  assign n12871 = n12857 ^ n12356 ;
  assign n12872 = n12871 ^ n12087 ;
  assign n12873 = n12872 ^ n12090 ;
  assign n12858 = n12857 ^ n12087 ;
  assign n12859 = n12858 ^ n12087 ;
  assign n12860 = n12859 ^ n12090 ;
  assign n12850 = n12356 ^ n12090 ;
  assign n12849 = n12597 ^ n12090 ;
  assign n12851 = n12850 ^ n12849 ;
  assign n12852 = ~n12090 & ~n12851 ;
  assign n12861 = n12860 ^ n12852 ;
  assign n12862 = n12850 ^ n12603 ;
  assign n12863 = ~n12851 & n12862 ;
  assign n12864 = n12863 ^ n12603 ;
  assign n12865 = n12860 & ~n12864 ;
  assign n12866 = n12861 & n12865 ;
  assign n12867 = n12866 ^ n12863 ;
  assign n12868 = n12867 ^ n12858 ;
  assign n12869 = n12868 ^ n12603 ;
  assign n12870 = n12869 ^ n12356 ;
  assign n12874 = n12873 ^ n12870 ;
  assign n12845 = n12595 ^ n12359 ;
  assign n12846 = ~n12596 & n12845 ;
  assign n12847 = n12846 ^ n12595 ;
  assign n12842 = x127 & n578 ;
  assign n12836 = x124 & n788 ;
  assign n12828 = n12560 ^ n12368 ;
  assign n12829 = n12566 & ~n12828 ;
  assign n12830 = n12829 ^ n12560 ;
  assign n12826 = x121 & n1058 ;
  assign n12819 = x118 & n1335 ;
  assign n12811 = n12543 ^ n12377 ;
  assign n12812 = ~n12549 & n12811 ;
  assign n12813 = n12812 ^ n12543 ;
  assign n12809 = x115 & n1666 ;
  assign n12802 = x112 & n2014 ;
  assign n12795 = x109 & n2429 ;
  assign n12788 = x106 & n2887 ;
  assign n12781 = x103 & n3383 ;
  assign n12770 = x99 & n3916 ;
  assign n12769 = x101 & n3919 ;
  assign n12771 = n12770 ^ n12769 ;
  assign n12772 = n12771 ^ x38 ;
  assign n12768 = n3920 & n4215 ;
  assign n12773 = n12772 ^ n12768 ;
  assign n12767 = x100 & n3924 ;
  assign n12774 = n12773 ^ n12767 ;
  assign n12764 = x97 & n4467 ;
  assign n12762 = n3660 & n4472 ;
  assign n12758 = x96 & n4474 ;
  assign n12757 = x98 & n4471 ;
  assign n12759 = n12758 ^ n12757 ;
  assign n12760 = n12759 ^ x41 ;
  assign n12754 = x94 & n5102 ;
  assign n12752 = n3159 & n5098 ;
  assign n12748 = x93 & n5094 ;
  assign n12747 = x95 & n5097 ;
  assign n12749 = n12748 ^ n12747 ;
  assign n12750 = n12749 ^ x44 ;
  assign n12740 = x90 & n5965 ;
  assign n12739 = x92 & n5729 ;
  assign n12741 = n12740 ^ n12739 ;
  assign n12742 = n12741 ^ x47 ;
  assign n12738 = n2684 & n5730 ;
  assign n12743 = n12742 ^ n12738 ;
  assign n12737 = x91 & n5736 ;
  assign n12744 = n12743 ^ n12737 ;
  assign n12730 = x87 & n6677 ;
  assign n12729 = x89 & n6428 ;
  assign n12731 = n12730 ^ n12729 ;
  assign n12732 = n12731 ^ x50 ;
  assign n12728 = n2249 & n6429 ;
  assign n12733 = n12732 ^ n12728 ;
  assign n12727 = x88 & n6433 ;
  assign n12734 = n12733 ^ n12727 ;
  assign n12719 = x81 & n7935 ;
  assign n12718 = x83 & n7938 ;
  assign n12720 = n12719 ^ n12718 ;
  assign n12721 = n12720 ^ x56 ;
  assign n12717 = n1512 & n7939 ;
  assign n12722 = n12721 ^ n12717 ;
  assign n12716 = x82 & n7931 ;
  assign n12723 = n12722 ^ n12716 ;
  assign n12709 = x78 & n8741 ;
  assign n12708 = x80 & n8744 ;
  assign n12710 = n12709 ^ n12708 ;
  assign n12711 = n12710 ^ x59 ;
  assign n12707 = n1206 & n8745 ;
  assign n12712 = n12711 ^ n12707 ;
  assign n12706 = x79 & n8737 ;
  assign n12713 = n12712 ^ n12706 ;
  assign n12700 = x75 & n9632 ;
  assign n12699 = x77 & n9635 ;
  assign n12701 = n12700 ^ n12699 ;
  assign n12702 = n12701 ^ x62 ;
  assign n12698 = ~n939 & n9636 ;
  assign n12703 = n12702 ^ n12698 ;
  assign n12697 = x76 & n9628 ;
  assign n12704 = n12703 ^ n12697 ;
  assign n12694 = x73 & n11875 ;
  assign n12693 = x74 & n9948 ;
  assign n12695 = n12694 ^ n12693 ;
  assign n12687 = x72 ^ x8 ;
  assign n12690 = n12420 & ~n12687 ;
  assign n12691 = n12690 ^ x72 ;
  assign n12692 = n12206 & n12691 ;
  assign n12696 = n12695 ^ n12692 ;
  assign n12705 = n12704 ^ n12696 ;
  assign n12714 = n12713 ^ n12705 ;
  assign n12684 = n12434 ^ n12429 ;
  assign n12685 = n12431 & ~n12684 ;
  assign n12686 = n12685 ^ n12434 ;
  assign n12715 = n12714 ^ n12686 ;
  assign n12724 = n12723 ^ n12715 ;
  assign n12681 = n12435 ^ n12412 ;
  assign n12682 = ~n12417 & n12681 ;
  assign n12683 = n12682 ^ n12412 ;
  assign n12725 = n12724 ^ n12683 ;
  assign n12678 = n12436 ^ n12404 ;
  assign n12679 = ~n12445 & ~n12678 ;
  assign n12671 = x84 & n7171 ;
  assign n12670 = x86 & n7174 ;
  assign n12672 = n12671 ^ n12670 ;
  assign n12673 = n12672 ^ x53 ;
  assign n12669 = n1857 & n7175 ;
  assign n12674 = n12673 ^ n12669 ;
  assign n12668 = x85 & n7179 ;
  assign n12675 = n12674 ^ n12668 ;
  assign n12676 = n12675 ^ n12436 ;
  assign n12680 = n12679 ^ n12676 ;
  assign n12726 = n12725 ^ n12680 ;
  assign n12735 = n12734 ^ n12726 ;
  assign n12665 = n12455 ^ n12446 ;
  assign n12666 = n12452 & ~n12665 ;
  assign n12667 = n12666 ^ n12455 ;
  assign n12736 = n12735 ^ n12667 ;
  assign n12745 = n12744 ^ n12736 ;
  assign n12662 = n12468 ^ n12464 ;
  assign n12663 = n12465 & n12662 ;
  assign n12664 = n12663 ^ n12468 ;
  assign n12746 = n12745 ^ n12664 ;
  assign n12751 = n12750 ^ n12746 ;
  assign n12753 = n12752 ^ n12751 ;
  assign n12755 = n12754 ^ n12753 ;
  assign n12659 = n12477 ^ n12398 ;
  assign n12660 = ~n12478 & ~n12659 ;
  assign n12661 = n12660 ^ n12477 ;
  assign n12756 = n12755 ^ n12661 ;
  assign n12761 = n12760 ^ n12756 ;
  assign n12763 = n12762 ^ n12761 ;
  assign n12765 = n12764 ^ n12763 ;
  assign n12656 = n12492 ^ n12479 ;
  assign n12657 = ~n12484 & n12656 ;
  assign n12658 = n12657 ^ n12479 ;
  assign n12766 = n12765 ^ n12658 ;
  assign n12775 = n12774 ^ n12766 ;
  assign n12653 = n12505 ^ n12501 ;
  assign n12654 = n12502 & n12653 ;
  assign n12655 = n12654 ^ n12505 ;
  assign n12776 = n12775 ^ n12655 ;
  assign n12777 = n12776 ^ x35 ;
  assign n12652 = x102 & n3375 ;
  assign n12778 = n12777 ^ n12652 ;
  assign n12651 = x104 & n3378 ;
  assign n12779 = n12778 ^ n12651 ;
  assign n12650 = n3379 & ~n4814 ;
  assign n12780 = n12779 ^ n12650 ;
  assign n12782 = n12781 ^ n12780 ;
  assign n12647 = n12515 ^ n12506 ;
  assign n12648 = n12512 & n12647 ;
  assign n12649 = n12648 ^ n12515 ;
  assign n12783 = n12782 ^ n12649 ;
  assign n12784 = n12783 ^ x32 ;
  assign n12646 = x105 & n2879 ;
  assign n12785 = n12784 ^ n12646 ;
  assign n12645 = x107 & n2882 ;
  assign n12786 = n12785 ^ n12645 ;
  assign n12644 = n2883 & ~n5448 ;
  assign n12787 = n12786 ^ n12644 ;
  assign n12789 = n12788 ^ n12787 ;
  assign n12641 = n12525 ^ n12516 ;
  assign n12642 = ~n12522 & ~n12641 ;
  assign n12643 = n12642 ^ n12525 ;
  assign n12790 = n12789 ^ n12643 ;
  assign n12791 = n12790 ^ x29 ;
  assign n12640 = x108 & n2581 ;
  assign n12792 = n12791 ^ n12640 ;
  assign n12639 = x110 & n2422 ;
  assign n12793 = n12792 ^ n12639 ;
  assign n12638 = n2423 & n6129 ;
  assign n12794 = n12793 ^ n12638 ;
  assign n12796 = n12795 ^ n12794 ;
  assign n12635 = n12535 ^ n12526 ;
  assign n12636 = n12532 & n12635 ;
  assign n12637 = n12636 ^ n12535 ;
  assign n12797 = n12796 ^ n12637 ;
  assign n12798 = n12797 ^ x26 ;
  assign n12634 = x111 & n2018 ;
  assign n12799 = n12798 ^ n12634 ;
  assign n12633 = x113 & n2021 ;
  assign n12800 = n12799 ^ n12633 ;
  assign n12632 = n2022 & ~n6839 ;
  assign n12801 = n12800 ^ n12632 ;
  assign n12803 = n12802 ^ n12801 ;
  assign n12629 = n12536 ^ n12383 ;
  assign n12630 = n12542 & ~n12629 ;
  assign n12631 = n12630 ^ n12536 ;
  assign n12804 = n12803 ^ n12631 ;
  assign n12805 = n12804 ^ x23 ;
  assign n12628 = x114 & n1658 ;
  assign n12806 = n12805 ^ n12628 ;
  assign n12627 = x116 & n1661 ;
  assign n12807 = n12806 ^ n12627 ;
  assign n12626 = n1662 & ~n7588 ;
  assign n12808 = n12807 ^ n12626 ;
  assign n12810 = n12809 ^ n12808 ;
  assign n12814 = n12813 ^ n12810 ;
  assign n12815 = n12814 ^ x20 ;
  assign n12625 = x117 & n1327 ;
  assign n12816 = n12815 ^ n12625 ;
  assign n12624 = x119 & n1330 ;
  assign n12817 = n12816 ^ n12624 ;
  assign n12623 = n1331 & n8394 ;
  assign n12818 = n12817 ^ n12623 ;
  assign n12820 = n12819 ^ n12818 ;
  assign n12620 = n12559 ^ n12550 ;
  assign n12621 = ~n12556 & n12620 ;
  assign n12622 = n12621 ^ n12559 ;
  assign n12821 = n12820 ^ n12622 ;
  assign n12822 = n12821 ^ x17 ;
  assign n12619 = x120 & n1050 ;
  assign n12823 = n12822 ^ n12619 ;
  assign n12618 = x122 & n1053 ;
  assign n12824 = n12823 ^ n12618 ;
  assign n12617 = n1054 & ~n9247 ;
  assign n12825 = n12824 ^ n12617 ;
  assign n12827 = n12826 ^ n12825 ;
  assign n12831 = n12830 ^ n12827 ;
  assign n12832 = n12831 ^ x14 ;
  assign n12616 = x123 & n877 ;
  assign n12833 = n12832 ^ n12616 ;
  assign n12615 = x125 & n782 ;
  assign n12834 = n12833 ^ n12615 ;
  assign n12614 = n783 & n10400 ;
  assign n12835 = n12834 ^ n12614 ;
  assign n12837 = n12836 ^ n12835 ;
  assign n12611 = n12576 ^ n12567 ;
  assign n12612 = n12573 & ~n12611 ;
  assign n12613 = n12612 ^ n12576 ;
  assign n12838 = n12837 ^ n12613 ;
  assign n12839 = n12838 ^ x11 ;
  assign n12610 = x126 & n647 ;
  assign n12840 = n12839 ^ n12610 ;
  assign n12609 = ~n573 & n10139 ;
  assign n12841 = n12840 ^ n12609 ;
  assign n12843 = n12842 ^ n12841 ;
  assign n12606 = n12586 ^ n12577 ;
  assign n12607 = n12583 & ~n12606 ;
  assign n12608 = n12607 ^ n12586 ;
  assign n12844 = n12843 ^ n12608 ;
  assign n12848 = n12847 ^ n12844 ;
  assign n12875 = n12874 ^ n12848 ;
  assign n13127 = n12874 ^ n12847 ;
  assign n13128 = n12848 & ~n13127 ;
  assign n13129 = n13128 ^ n12874 ;
  assign n13123 = n12838 ^ n12608 ;
  assign n13124 = ~n12843 & ~n13123 ;
  assign n13125 = n13124 ^ n12838 ;
  assign n13119 = n12831 ^ n12613 ;
  assign n13120 = ~n12837 & ~n13119 ;
  assign n13121 = n13120 ^ n12831 ;
  assign n13115 = x125 & n788 ;
  assign n13107 = n12814 ^ n12622 ;
  assign n13108 = ~n12820 & ~n13107 ;
  assign n13109 = n13108 ^ n12814 ;
  assign n13105 = x122 & n1058 ;
  assign n13098 = x119 & n1335 ;
  assign n13091 = x116 & n1666 ;
  assign n13083 = n12790 ^ n12637 ;
  assign n13084 = ~n12796 & n13083 ;
  assign n13085 = n13084 ^ n12790 ;
  assign n13081 = x113 & n2014 ;
  assign n13073 = n12783 ^ n12643 ;
  assign n13074 = n12789 & ~n13073 ;
  assign n13075 = n13074 ^ n12783 ;
  assign n13071 = x110 & n2429 ;
  assign n13063 = n12776 ^ n12649 ;
  assign n13064 = ~n12782 & n13063 ;
  assign n13065 = n13064 ^ n12776 ;
  assign n13061 = x107 & n2887 ;
  assign n13053 = n12774 ^ n12655 ;
  assign n13054 = ~n12775 & n13053 ;
  assign n13055 = n13054 ^ n12774 ;
  assign n13047 = x103 & n3375 ;
  assign n13046 = x105 & n3378 ;
  assign n13048 = n13047 ^ n13046 ;
  assign n13049 = n13048 ^ x35 ;
  assign n13045 = n3379 & ~n5023 ;
  assign n13050 = n13049 ^ n13045 ;
  assign n13044 = x104 & n3383 ;
  assign n13051 = n13050 ^ n13044 ;
  assign n13038 = x100 & n3916 ;
  assign n13037 = x102 & n3919 ;
  assign n13039 = n13038 ^ n13037 ;
  assign n13040 = n13039 ^ x38 ;
  assign n13036 = n3920 & n4410 ;
  assign n13041 = n13040 ^ n13036 ;
  assign n13035 = x101 & n3924 ;
  assign n13042 = n13041 ^ n13035 ;
  assign n13031 = n12756 ^ n12658 ;
  assign n13032 = ~n12765 & ~n13031 ;
  assign n13033 = n13032 ^ n12756 ;
  assign n13025 = x97 & n4474 ;
  assign n13024 = x99 & n4471 ;
  assign n13026 = n13025 ^ n13024 ;
  assign n13027 = n13026 ^ x41 ;
  assign n13023 = n3843 & n4472 ;
  assign n13028 = n13027 ^ n13023 ;
  assign n13022 = x98 & n4467 ;
  assign n13029 = n13028 ^ n13022 ;
  assign n13014 = x95 & n5102 ;
  assign n13012 = n3323 & n5098 ;
  assign n13008 = x94 & n5094 ;
  assign n13007 = x96 & n5097 ;
  assign n13009 = n13008 ^ n13007 ;
  assign n13010 = n13009 ^ x44 ;
  assign n13003 = n12734 ^ n12667 ;
  assign n13004 = ~n12735 & n13003 ;
  assign n13005 = n13004 ^ n12734 ;
  assign n12997 = x91 & n5965 ;
  assign n12996 = x93 & n5729 ;
  assign n12998 = n12997 ^ n12996 ;
  assign n12999 = n12998 ^ x47 ;
  assign n12995 = n2836 & n5730 ;
  assign n13000 = n12999 ^ n12995 ;
  assign n12994 = x92 & n5736 ;
  assign n13001 = n13000 ^ n12994 ;
  assign n12986 = x85 & n7171 ;
  assign n12985 = x87 & n7174 ;
  assign n12987 = n12986 ^ n12985 ;
  assign n12988 = n12987 ^ x53 ;
  assign n12984 = n1982 & n7175 ;
  assign n12989 = n12988 ^ n12984 ;
  assign n12983 = x86 & n7179 ;
  assign n12990 = n12989 ^ n12983 ;
  assign n12979 = n12713 ^ n12686 ;
  assign n12980 = ~n12714 & ~n12979 ;
  assign n12981 = n12980 ^ n12713 ;
  assign n12973 = x82 & n7935 ;
  assign n12972 = x84 & n7938 ;
  assign n12974 = n12973 ^ n12972 ;
  assign n12975 = n12974 ^ x56 ;
  assign n12971 = n1624 & n7939 ;
  assign n12976 = n12975 ^ n12971 ;
  assign n12970 = x83 & n7931 ;
  assign n12977 = n12976 ^ n12970 ;
  assign n12964 = x79 & n8741 ;
  assign n12963 = x81 & n8744 ;
  assign n12965 = n12964 ^ n12963 ;
  assign n12966 = n12965 ^ x59 ;
  assign n12962 = n1305 & n8745 ;
  assign n12967 = n12966 ^ n12962 ;
  assign n12961 = x80 & n8737 ;
  assign n12968 = n12967 ^ n12961 ;
  assign n12955 = x76 & n9632 ;
  assign n12954 = x78 & n9635 ;
  assign n12956 = n12955 ^ n12954 ;
  assign n12957 = n12956 ^ x62 ;
  assign n12953 = ~n1025 & n9636 ;
  assign n12958 = n12957 ^ n12953 ;
  assign n12952 = x77 & n9628 ;
  assign n12959 = n12958 ^ n12952 ;
  assign n537 = x74 ^ x73 ;
  assign n12947 = x63 & n537 ;
  assign n612 = x75 ^ x74 ;
  assign n12948 = n12947 ^ n612 ;
  assign n12949 = ~n9948 & n12948 ;
  assign n12950 = n12949 ^ n612 ;
  assign n12940 = n12704 ^ n12695 ;
  assign n12941 = n12696 & ~n12940 ;
  assign n12942 = n12941 ^ n12704 ;
  assign n12951 = n12950 ^ n12942 ;
  assign n12960 = n12959 ^ n12951 ;
  assign n12969 = n12968 ^ n12960 ;
  assign n12978 = n12977 ^ n12969 ;
  assign n12982 = n12981 ^ n12978 ;
  assign n12991 = n12990 ^ n12982 ;
  assign n12937 = n12723 ^ n12683 ;
  assign n12938 = n12724 & n12937 ;
  assign n12939 = n12938 ^ n12723 ;
  assign n12992 = n12991 ^ n12939 ;
  assign n12927 = x88 & n6677 ;
  assign n12926 = x90 & n6428 ;
  assign n12928 = n12927 ^ n12926 ;
  assign n12929 = n12928 ^ x50 ;
  assign n12925 = n2386 & n6429 ;
  assign n12930 = n12929 ^ n12925 ;
  assign n12924 = x89 & n6433 ;
  assign n12931 = n12930 ^ n12924 ;
  assign n12933 = n12931 ^ n12675 ;
  assign n12932 = n12931 ^ n12725 ;
  assign n12934 = n12933 ^ n12932 ;
  assign n12935 = ~n12680 & n12934 ;
  assign n12936 = n12935 ^ n12933 ;
  assign n12993 = n12992 ^ n12936 ;
  assign n13002 = n13001 ^ n12993 ;
  assign n13006 = n13005 ^ n13002 ;
  assign n13011 = n13010 ^ n13006 ;
  assign n13013 = n13012 ^ n13011 ;
  assign n13015 = n13014 ^ n13013 ;
  assign n12921 = n12744 ^ n12664 ;
  assign n12922 = ~n12745 & n12921 ;
  assign n12923 = n12922 ^ n12744 ;
  assign n13016 = n13015 ^ n12923 ;
  assign n13017 = n13016 ^ n12746 ;
  assign n13018 = n13017 ^ n12661 ;
  assign n13019 = n13018 ^ n13016 ;
  assign n13020 = ~n12755 & ~n13019 ;
  assign n13021 = n13020 ^ n13017 ;
  assign n13030 = n13029 ^ n13021 ;
  assign n13034 = n13033 ^ n13030 ;
  assign n13043 = n13042 ^ n13034 ;
  assign n13052 = n13051 ^ n13043 ;
  assign n13056 = n13055 ^ n13052 ;
  assign n13057 = n13056 ^ x32 ;
  assign n12920 = x106 & n2879 ;
  assign n13058 = n13057 ^ n12920 ;
  assign n12919 = x108 & n2882 ;
  assign n13059 = n13058 ^ n12919 ;
  assign n12918 = n2883 & n5670 ;
  assign n13060 = n13059 ^ n12918 ;
  assign n13062 = n13061 ^ n13060 ;
  assign n13066 = n13065 ^ n13062 ;
  assign n13067 = n13066 ^ x29 ;
  assign n12917 = x109 & n2581 ;
  assign n13068 = n13067 ^ n12917 ;
  assign n12916 = x111 & n2422 ;
  assign n13069 = n13068 ^ n12916 ;
  assign n12915 = n2423 & ~n6360 ;
  assign n13070 = n13069 ^ n12915 ;
  assign n13072 = n13071 ^ n13070 ;
  assign n13076 = n13075 ^ n13072 ;
  assign n13077 = n13076 ^ x26 ;
  assign n12914 = x112 & n2018 ;
  assign n13078 = n13077 ^ n12914 ;
  assign n12913 = x114 & n2021 ;
  assign n13079 = n13078 ^ n12913 ;
  assign n12912 = n2022 & ~n7092 ;
  assign n13080 = n13079 ^ n12912 ;
  assign n13082 = n13081 ^ n13080 ;
  assign n13086 = n13085 ^ n13082 ;
  assign n13087 = n13086 ^ x23 ;
  assign n12911 = x115 & n1658 ;
  assign n13088 = n13087 ^ n12911 ;
  assign n12910 = x117 & n1661 ;
  assign n13089 = n13088 ^ n12910 ;
  assign n12909 = n1662 & ~n7850 ;
  assign n13090 = n13089 ^ n12909 ;
  assign n13092 = n13091 ^ n13090 ;
  assign n12906 = n12797 ^ n12631 ;
  assign n12907 = n12803 & n12906 ;
  assign n12908 = n12907 ^ n12797 ;
  assign n13093 = n13092 ^ n12908 ;
  assign n13094 = n13093 ^ x20 ;
  assign n12905 = x118 & n1327 ;
  assign n13095 = n13094 ^ n12905 ;
  assign n12904 = x120 & n1330 ;
  assign n13096 = n13095 ^ n12904 ;
  assign n12903 = n1331 & n8891 ;
  assign n13097 = n13096 ^ n12903 ;
  assign n13099 = n13098 ^ n13097 ;
  assign n12900 = n12813 ^ n12804 ;
  assign n12901 = ~n12810 & ~n12900 ;
  assign n12902 = n12901 ^ n12813 ;
  assign n13100 = n13099 ^ n12902 ;
  assign n13101 = n13100 ^ x17 ;
  assign n12899 = x121 & n1050 ;
  assign n13102 = n13101 ^ n12899 ;
  assign n12898 = x123 & n1053 ;
  assign n13103 = n13102 ^ n12898 ;
  assign n12897 = n1054 & ~n9786 ;
  assign n13104 = n13103 ^ n12897 ;
  assign n13106 = n13105 ^ n13104 ;
  assign n13110 = n13109 ^ n13106 ;
  assign n13111 = n13110 ^ x14 ;
  assign n12896 = x124 & n877 ;
  assign n13112 = n13111 ^ n12896 ;
  assign n12895 = x126 & n782 ;
  assign n13113 = n13112 ^ n12895 ;
  assign n12894 = n783 & n10441 ;
  assign n13114 = n13113 ^ n12894 ;
  assign n13116 = n13115 ^ n13114 ;
  assign n12891 = n12830 ^ n12821 ;
  assign n12892 = n12827 & ~n12891 ;
  assign n12893 = n12892 ^ n12830 ;
  assign n13117 = n13116 ^ n12893 ;
  assign n12878 = ~x10 & x127 ;
  assign n12879 = n12878 ^ x11 ;
  assign n12880 = ~n10138 & ~n12879 ;
  assign n12881 = n12880 ^ x11 ;
  assign n12882 = n504 & ~n12881 ;
  assign n12883 = n503 ^ x11 ;
  assign n12886 = x127 & n569 ;
  assign n12887 = ~n12883 & n12886 ;
  assign n12888 = n12887 ^ n12883 ;
  assign n12889 = n12888 ^ n503 ;
  assign n12890 = ~n12882 & n12889 ;
  assign n13118 = n13117 ^ n12890 ;
  assign n13122 = n13121 ^ n13118 ;
  assign n13126 = n13125 ^ n13122 ;
  assign n13130 = n13129 ^ n13126 ;
  assign n13371 = n13110 ^ n12893 ;
  assign n13372 = ~n13116 & ~n13371 ;
  assign n13373 = n13372 ^ n13110 ;
  assign n13369 = x126 & n788 ;
  assign n13362 = x123 & n1058 ;
  assign n13354 = n13093 ^ n12902 ;
  assign n13355 = ~n13099 & n13354 ;
  assign n13356 = n13355 ^ n13093 ;
  assign n13352 = x120 & n1335 ;
  assign n13345 = x117 & n1666 ;
  assign n13338 = x114 & n2014 ;
  assign n13331 = x111 & n2429 ;
  assign n13324 = x108 & n2887 ;
  assign n13313 = x104 & n3375 ;
  assign n13312 = x106 & n3378 ;
  assign n13314 = n13313 ^ n13312 ;
  assign n13315 = n13314 ^ x35 ;
  assign n13311 = n3379 & ~n5240 ;
  assign n13316 = n13315 ^ n13311 ;
  assign n13310 = x105 & n3383 ;
  assign n13317 = n13316 ^ n13310 ;
  assign n13304 = x101 & n3916 ;
  assign n13303 = x103 & n3919 ;
  assign n13305 = n13304 ^ n13303 ;
  assign n13306 = n13305 ^ x38 ;
  assign n13302 = n3920 & ~n4615 ;
  assign n13307 = n13306 ^ n13302 ;
  assign n13301 = x102 & n3924 ;
  assign n13308 = n13307 ^ n13301 ;
  assign n13292 = n13029 ^ n13016 ;
  assign n13293 = n13021 & ~n13292 ;
  assign n13294 = n13293 ^ n13016 ;
  assign n13286 = x98 & n4474 ;
  assign n13285 = x100 & n4471 ;
  assign n13287 = n13286 ^ n13285 ;
  assign n13288 = n13287 ^ x41 ;
  assign n13284 = n4034 & n4472 ;
  assign n13289 = n13288 ^ n13284 ;
  assign n13283 = x99 & n4467 ;
  assign n13290 = n13289 ^ n13283 ;
  assign n13279 = n13006 ^ n12923 ;
  assign n13280 = ~n13015 & ~n13279 ;
  assign n13281 = n13280 ^ n13006 ;
  assign n13273 = x95 & n5094 ;
  assign n13272 = x97 & n5097 ;
  assign n13274 = n13273 ^ n13272 ;
  assign n13275 = n13274 ^ x44 ;
  assign n13271 = n3494 & n5098 ;
  assign n13276 = n13275 ^ n13271 ;
  assign n13270 = x96 & n5102 ;
  assign n13277 = n13276 ^ n13270 ;
  assign n13262 = x89 & n6677 ;
  assign n13261 = x91 & n6428 ;
  assign n13263 = n13262 ^ n13261 ;
  assign n13264 = n13263 ^ x50 ;
  assign n13260 = n2542 & n6429 ;
  assign n13265 = n13264 ^ n13260 ;
  assign n13259 = x90 & n6433 ;
  assign n13266 = n13265 ^ n13259 ;
  assign n13255 = n12990 ^ n12939 ;
  assign n13256 = ~n12991 & n13255 ;
  assign n13257 = n13256 ^ n12990 ;
  assign n13249 = x86 & n7171 ;
  assign n13248 = x88 & n7174 ;
  assign n13250 = n13249 ^ n13248 ;
  assign n13251 = n13250 ^ x53 ;
  assign n13247 = n2119 & n7175 ;
  assign n13252 = n13251 ^ n13247 ;
  assign n13246 = x87 & n7179 ;
  assign n13253 = n13252 ^ n13246 ;
  assign n13243 = x84 & n7931 ;
  assign n13236 = x81 & n8737 ;
  assign n13225 = x77 & n9632 ;
  assign n13224 = x79 & n9635 ;
  assign n13226 = n13225 ^ n13224 ;
  assign n13227 = n13226 ^ x62 ;
  assign n13223 = n1118 & n9636 ;
  assign n13228 = n13227 ^ n13223 ;
  assign n13222 = x78 & n9628 ;
  assign n13229 = n13228 ^ n13222 ;
  assign n13217 = x63 & x75 ;
  assign n13218 = n13217 ^ x76 ;
  assign n13219 = ~n9948 & n13218 ;
  assign n13211 = n12695 ^ x76 ;
  assign n13220 = n13219 ^ n13211 ;
  assign n13221 = n13220 ^ x11 ;
  assign n13230 = n13229 ^ n13221 ;
  assign n13205 = ~x75 & n12693 ;
  assign n13204 = ~x74 & n12694 ;
  assign n13206 = n13205 ^ n13204 ;
  assign n13207 = ~n12942 & ~n13206 ;
  assign n13208 = n13204 ^ n12950 ;
  assign n13209 = n13207 & ~n13208 ;
  assign n13210 = n13209 ^ n13206 ;
  assign n13231 = n13230 ^ n13210 ;
  assign n13232 = n13231 ^ x59 ;
  assign n13203 = x80 & n8741 ;
  assign n13233 = n13232 ^ n13203 ;
  assign n13202 = x82 & n8744 ;
  assign n13234 = n13233 ^ n13202 ;
  assign n13201 = n1411 & n8745 ;
  assign n13235 = n13234 ^ n13201 ;
  assign n13237 = n13236 ^ n13235 ;
  assign n13198 = n12968 ^ n12959 ;
  assign n13199 = n12960 & n13198 ;
  assign n13200 = n13199 ^ n12968 ;
  assign n13238 = n13237 ^ n13200 ;
  assign n13239 = n13238 ^ x56 ;
  assign n13197 = x83 & n7935 ;
  assign n13240 = n13239 ^ n13197 ;
  assign n13196 = x85 & n7938 ;
  assign n13241 = n13240 ^ n13196 ;
  assign n13195 = n1743 & n7939 ;
  assign n13242 = n13241 ^ n13195 ;
  assign n13244 = n13243 ^ n13242 ;
  assign n13192 = n12981 ^ n12977 ;
  assign n13193 = n12978 & n13192 ;
  assign n13194 = n13193 ^ n12981 ;
  assign n13245 = n13244 ^ n13194 ;
  assign n13254 = n13253 ^ n13245 ;
  assign n13258 = n13257 ^ n13254 ;
  assign n13267 = n13266 ^ n13258 ;
  assign n13189 = n12992 ^ n12931 ;
  assign n13190 = n12936 & ~n13189 ;
  assign n13191 = n13190 ^ n12931 ;
  assign n13268 = n13267 ^ n13191 ;
  assign n13179 = x92 & n5965 ;
  assign n13178 = x94 & n5729 ;
  assign n13180 = n13179 ^ n13178 ;
  assign n13181 = n13180 ^ x47 ;
  assign n13177 = n2997 & n5730 ;
  assign n13182 = n13181 ^ n13177 ;
  assign n13176 = x93 & n5736 ;
  assign n13183 = n13182 ^ n13176 ;
  assign n13184 = n13183 ^ n13005 ;
  assign n13185 = n13184 ^ n13001 ;
  assign n13186 = n13185 ^ n13183 ;
  assign n13187 = n13002 & n13186 ;
  assign n13188 = n13187 ^ n13184 ;
  assign n13269 = n13268 ^ n13188 ;
  assign n13278 = n13277 ^ n13269 ;
  assign n13282 = n13281 ^ n13278 ;
  assign n13291 = n13290 ^ n13282 ;
  assign n13295 = n13294 ^ n13291 ;
  assign n13296 = n13295 ^ n13042 ;
  assign n13297 = n13296 ^ n13033 ;
  assign n13298 = n13297 ^ n13295 ;
  assign n13299 = n13034 & ~n13298 ;
  assign n13300 = n13299 ^ n13296 ;
  assign n13309 = n13308 ^ n13300 ;
  assign n13318 = n13317 ^ n13309 ;
  assign n13173 = n13055 ^ n13051 ;
  assign n13174 = n13052 & n13173 ;
  assign n13175 = n13174 ^ n13055 ;
  assign n13319 = n13318 ^ n13175 ;
  assign n13320 = n13319 ^ x32 ;
  assign n13172 = x107 & n2879 ;
  assign n13321 = n13320 ^ n13172 ;
  assign n13171 = x109 & n2882 ;
  assign n13322 = n13321 ^ n13171 ;
  assign n13170 = n2883 & n5902 ;
  assign n13323 = n13322 ^ n13170 ;
  assign n13325 = n13324 ^ n13323 ;
  assign n13167 = n13065 ^ n13056 ;
  assign n13168 = n13062 & n13167 ;
  assign n13169 = n13168 ^ n13065 ;
  assign n13326 = n13325 ^ n13169 ;
  assign n13327 = n13326 ^ x29 ;
  assign n13166 = x110 & n2581 ;
  assign n13328 = n13327 ^ n13166 ;
  assign n13165 = x112 & n2422 ;
  assign n13329 = n13328 ^ n13165 ;
  assign n13164 = n2423 & ~n6600 ;
  assign n13330 = n13329 ^ n13164 ;
  assign n13332 = n13331 ^ n13330 ;
  assign n13161 = n13075 ^ n13066 ;
  assign n13162 = ~n13072 & n13161 ;
  assign n13163 = n13162 ^ n13075 ;
  assign n13333 = n13332 ^ n13163 ;
  assign n13334 = n13333 ^ x26 ;
  assign n13160 = x113 & n2018 ;
  assign n13335 = n13334 ^ n13160 ;
  assign n13159 = x115 & n2021 ;
  assign n13336 = n13335 ^ n13159 ;
  assign n13158 = n2022 & ~n7343 ;
  assign n13337 = n13336 ^ n13158 ;
  assign n13339 = n13338 ^ n13337 ;
  assign n13155 = n13085 ^ n13076 ;
  assign n13156 = ~n13082 & ~n13155 ;
  assign n13157 = n13156 ^ n13085 ;
  assign n13340 = n13339 ^ n13157 ;
  assign n13341 = n13340 ^ x23 ;
  assign n13154 = x116 & n1658 ;
  assign n13342 = n13341 ^ n13154 ;
  assign n13153 = x118 & n1661 ;
  assign n13343 = n13342 ^ n13153 ;
  assign n13152 = n1662 & ~n8123 ;
  assign n13344 = n13343 ^ n13152 ;
  assign n13346 = n13345 ^ n13344 ;
  assign n13149 = n13086 ^ n12908 ;
  assign n13150 = ~n13092 & ~n13149 ;
  assign n13151 = n13150 ^ n13086 ;
  assign n13347 = n13346 ^ n13151 ;
  assign n13348 = n13347 ^ x20 ;
  assign n13148 = x119 & n1327 ;
  assign n13349 = n13348 ^ n13148 ;
  assign n13147 = x121 & n1330 ;
  assign n13350 = n13349 ^ n13147 ;
  assign n13146 = n1331 & n8962 ;
  assign n13351 = n13350 ^ n13146 ;
  assign n13353 = n13352 ^ n13351 ;
  assign n13357 = n13356 ^ n13353 ;
  assign n13358 = n13357 ^ x17 ;
  assign n13145 = x122 & n1050 ;
  assign n13359 = n13358 ^ n13145 ;
  assign n13144 = x124 & n1053 ;
  assign n13360 = n13359 ^ n13144 ;
  assign n13143 = n1054 & n10095 ;
  assign n13361 = n13360 ^ n13143 ;
  assign n13363 = n13362 ^ n13361 ;
  assign n13140 = n13109 ^ n13100 ;
  assign n13141 = ~n13106 & ~n13140 ;
  assign n13142 = n13141 ^ n13109 ;
  assign n13364 = n13363 ^ n13142 ;
  assign n13365 = n13364 ^ x14 ;
  assign n13139 = x125 & n877 ;
  assign n13366 = n13365 ^ n13139 ;
  assign n13138 = x127 & n782 ;
  assign n13367 = n13366 ^ n13138 ;
  assign n13137 = n783 & n10972 ;
  assign n13368 = n13367 ^ n13137 ;
  assign n13370 = n13369 ^ n13368 ;
  assign n13374 = n13373 ^ n13370 ;
  assign n13134 = n13121 ^ n13117 ;
  assign n13135 = n13118 & n13134 ;
  assign n13136 = n13135 ^ n13121 ;
  assign n13375 = n13374 ^ n13136 ;
  assign n13131 = n13129 ^ n13125 ;
  assign n13132 = n13126 & n13131 ;
  assign n13133 = n13132 ^ n13129 ;
  assign n13376 = n13375 ^ n13133 ;
  assign n13604 = n13357 ^ n13142 ;
  assign n13605 = n13363 & ~n13604 ;
  assign n13606 = n13605 ^ n13357 ;
  assign n13602 = x127 & n788 ;
  assign n13596 = x124 & n1058 ;
  assign n13589 = x121 & n1335 ;
  assign n13581 = n13333 ^ n13157 ;
  assign n13582 = ~n13339 & n13581 ;
  assign n13583 = n13582 ^ n13333 ;
  assign n13579 = x118 & n1666 ;
  assign n13571 = n13326 ^ n13163 ;
  assign n13572 = ~n13332 & ~n13571 ;
  assign n13573 = n13572 ^ n13326 ;
  assign n13569 = x115 & n2014 ;
  assign n13559 = x111 & n2581 ;
  assign n13558 = x113 & n2422 ;
  assign n13560 = n13559 ^ n13558 ;
  assign n13561 = n13560 ^ x29 ;
  assign n13557 = n2423 & ~n6839 ;
  assign n13562 = n13561 ^ n13557 ;
  assign n13556 = x112 & n2429 ;
  assign n13563 = n13562 ^ n13556 ;
  assign n13544 = x108 & n2879 ;
  assign n13543 = x110 & n2882 ;
  assign n13545 = n13544 ^ n13543 ;
  assign n13546 = n13545 ^ x32 ;
  assign n13542 = n2883 & n6129 ;
  assign n13547 = n13546 ^ n13542 ;
  assign n13541 = x109 & n2887 ;
  assign n13548 = n13547 ^ n13541 ;
  assign n13535 = x105 & n3375 ;
  assign n13534 = x107 & n3378 ;
  assign n13536 = n13535 ^ n13534 ;
  assign n13537 = n13536 ^ x35 ;
  assign n13533 = n3379 & ~n5448 ;
  assign n13538 = n13537 ^ n13533 ;
  assign n13532 = x106 & n3383 ;
  assign n13539 = n13538 ^ n13532 ;
  assign n13528 = n13308 ^ n13295 ;
  assign n13529 = n13300 & n13528 ;
  assign n13530 = n13529 ^ n13295 ;
  assign n13522 = x102 & n3916 ;
  assign n13521 = x104 & n3919 ;
  assign n13523 = n13522 ^ n13521 ;
  assign n13524 = n13523 ^ x38 ;
  assign n13520 = n3920 & ~n4814 ;
  assign n13525 = n13524 ^ n13520 ;
  assign n13519 = x103 & n3924 ;
  assign n13526 = n13525 ^ n13519 ;
  assign n13512 = x99 & n4474 ;
  assign n13511 = x101 & n4471 ;
  assign n13513 = n13512 ^ n13511 ;
  assign n13514 = n13513 ^ x41 ;
  assign n13510 = n4215 & n4472 ;
  assign n13515 = n13514 ^ n13510 ;
  assign n13509 = x100 & n4467 ;
  assign n13516 = n13515 ^ n13509 ;
  assign n13505 = x97 & n5102 ;
  assign n13503 = n3660 & n5098 ;
  assign n13499 = x96 & n5094 ;
  assign n13498 = x98 & n5097 ;
  assign n13500 = n13499 ^ n13498 ;
  assign n13501 = n13500 ^ x44 ;
  assign n13491 = x93 & n5965 ;
  assign n13490 = x95 & n5729 ;
  assign n13492 = n13491 ^ n13490 ;
  assign n13493 = n13492 ^ x47 ;
  assign n13489 = n3159 & n5730 ;
  assign n13494 = n13493 ^ n13489 ;
  assign n13488 = x94 & n5736 ;
  assign n13495 = n13494 ^ n13488 ;
  assign n13481 = x90 & n6677 ;
  assign n13480 = x92 & n6428 ;
  assign n13482 = n13481 ^ n13480 ;
  assign n13483 = n13482 ^ x50 ;
  assign n13479 = n2684 & n6429 ;
  assign n13484 = n13483 ^ n13479 ;
  assign n13478 = x91 & n6433 ;
  assign n13485 = n13484 ^ n13478 ;
  assign n13474 = n13238 ^ n13194 ;
  assign n13475 = n13244 & n13474 ;
  assign n13476 = n13475 ^ n13238 ;
  assign n13468 = x87 & n7171 ;
  assign n13467 = x89 & n7174 ;
  assign n13469 = n13468 ^ n13467 ;
  assign n13470 = n13469 ^ x53 ;
  assign n13466 = n2249 & n7175 ;
  assign n13471 = n13470 ^ n13466 ;
  assign n13465 = x88 & n7179 ;
  assign n13472 = n13471 ^ n13465 ;
  assign n13457 = x81 & n8741 ;
  assign n13456 = x83 & n8744 ;
  assign n13458 = n13457 ^ n13456 ;
  assign n13459 = n13458 ^ x59 ;
  assign n13455 = n1512 & n8745 ;
  assign n13460 = n13459 ^ n13455 ;
  assign n13454 = x82 & n8737 ;
  assign n13461 = n13460 ^ n13454 ;
  assign n13448 = x78 & n9632 ;
  assign n13447 = x80 & n9635 ;
  assign n13449 = n13448 ^ n13447 ;
  assign n13450 = n13449 ^ x62 ;
  assign n13446 = n1206 & n9636 ;
  assign n13451 = n13450 ^ n13446 ;
  assign n13445 = x79 & n9628 ;
  assign n13452 = n13451 ^ n13445 ;
  assign n13441 = n12695 ^ x11 ;
  assign n13442 = ~n13220 & ~n13441 ;
  assign n13443 = n13442 ^ x11 ;
  assign n13437 = x63 & x76 ;
  assign n13438 = n13437 ^ x77 ;
  assign n13439 = ~n9948 & n13438 ;
  assign n13440 = n13439 ^ x77 ;
  assign n13444 = n13443 ^ n13440 ;
  assign n13453 = n13452 ^ n13444 ;
  assign n13462 = n13461 ^ n13453 ;
  assign n13434 = n13229 ^ n13210 ;
  assign n13435 = ~n13230 & ~n13434 ;
  assign n13436 = n13435 ^ n13229 ;
  assign n13463 = n13462 ^ n13436 ;
  assign n13431 = n13231 ^ n13200 ;
  assign n13432 = n13237 & n13431 ;
  assign n13424 = x84 & n7935 ;
  assign n13423 = x86 & n7938 ;
  assign n13425 = n13424 ^ n13423 ;
  assign n13426 = n13425 ^ x56 ;
  assign n13422 = n1857 & n7939 ;
  assign n13427 = n13426 ^ n13422 ;
  assign n13421 = x85 & n7931 ;
  assign n13428 = n13427 ^ n13421 ;
  assign n13429 = n13428 ^ n13231 ;
  assign n13433 = n13432 ^ n13429 ;
  assign n13464 = n13463 ^ n13433 ;
  assign n13473 = n13472 ^ n13464 ;
  assign n13477 = n13476 ^ n13473 ;
  assign n13486 = n13485 ^ n13477 ;
  assign n13418 = n13257 ^ n13253 ;
  assign n13419 = ~n13254 & n13418 ;
  assign n13420 = n13419 ^ n13257 ;
  assign n13487 = n13486 ^ n13420 ;
  assign n13496 = n13495 ^ n13487 ;
  assign n13415 = n13266 ^ n13191 ;
  assign n13416 = n13267 & n13415 ;
  assign n13417 = n13416 ^ n13266 ;
  assign n13497 = n13496 ^ n13417 ;
  assign n13502 = n13501 ^ n13497 ;
  assign n13504 = n13503 ^ n13502 ;
  assign n13506 = n13505 ^ n13504 ;
  assign n13412 = n13268 ^ n13183 ;
  assign n13413 = n13188 & n13412 ;
  assign n13414 = n13413 ^ n13183 ;
  assign n13507 = n13506 ^ n13414 ;
  assign n13409 = n13281 ^ n13277 ;
  assign n13410 = ~n13278 & ~n13409 ;
  assign n13411 = n13410 ^ n13281 ;
  assign n13508 = n13507 ^ n13411 ;
  assign n13517 = n13516 ^ n13508 ;
  assign n13406 = n13294 ^ n13290 ;
  assign n13407 = n13291 & ~n13406 ;
  assign n13408 = n13407 ^ n13294 ;
  assign n13518 = n13517 ^ n13408 ;
  assign n13527 = n13526 ^ n13518 ;
  assign n13531 = n13530 ^ n13527 ;
  assign n13540 = n13539 ^ n13531 ;
  assign n13549 = n13548 ^ n13540 ;
  assign n13403 = n13317 ^ n13175 ;
  assign n13404 = n13318 & n13403 ;
  assign n13405 = n13404 ^ n13317 ;
  assign n13550 = n13549 ^ n13405 ;
  assign n13551 = n13550 ^ n13319 ;
  assign n13552 = n13551 ^ n13550 ;
  assign n13553 = n13552 ^ n13169 ;
  assign n13554 = n13325 & ~n13553 ;
  assign n13555 = n13554 ^ n13551 ;
  assign n13564 = n13563 ^ n13555 ;
  assign n13565 = n13564 ^ x26 ;
  assign n13402 = x114 & n2018 ;
  assign n13566 = n13565 ^ n13402 ;
  assign n13401 = x116 & n2021 ;
  assign n13567 = n13566 ^ n13401 ;
  assign n13400 = n2022 & ~n7588 ;
  assign n13568 = n13567 ^ n13400 ;
  assign n13570 = n13569 ^ n13568 ;
  assign n13574 = n13573 ^ n13570 ;
  assign n13575 = n13574 ^ x23 ;
  assign n13399 = x117 & n1658 ;
  assign n13576 = n13575 ^ n13399 ;
  assign n13398 = x119 & n1661 ;
  assign n13577 = n13576 ^ n13398 ;
  assign n13397 = n1662 & n8394 ;
  assign n13578 = n13577 ^ n13397 ;
  assign n13580 = n13579 ^ n13578 ;
  assign n13584 = n13583 ^ n13580 ;
  assign n13585 = n13584 ^ x20 ;
  assign n13396 = x120 & n1327 ;
  assign n13586 = n13585 ^ n13396 ;
  assign n13395 = x122 & n1330 ;
  assign n13587 = n13586 ^ n13395 ;
  assign n13394 = n1331 & ~n9247 ;
  assign n13588 = n13587 ^ n13394 ;
  assign n13590 = n13589 ^ n13588 ;
  assign n13391 = n13340 ^ n13151 ;
  assign n13392 = n13346 & ~n13391 ;
  assign n13393 = n13392 ^ n13340 ;
  assign n13591 = n13590 ^ n13393 ;
  assign n13592 = n13591 ^ x17 ;
  assign n13390 = x123 & n1050 ;
  assign n13593 = n13592 ^ n13390 ;
  assign n13389 = x125 & n1053 ;
  assign n13594 = n13593 ^ n13389 ;
  assign n13388 = n1054 & n10400 ;
  assign n13595 = n13594 ^ n13388 ;
  assign n13597 = n13596 ^ n13595 ;
  assign n13385 = n13356 ^ n13347 ;
  assign n13386 = n13353 & n13385 ;
  assign n13387 = n13386 ^ n13356 ;
  assign n13598 = n13597 ^ n13387 ;
  assign n13599 = n13598 ^ x14 ;
  assign n13384 = x126 & n877 ;
  assign n13600 = n13599 ^ n13384 ;
  assign n13383 = n783 & n10139 ;
  assign n13601 = n13600 ^ n13383 ;
  assign n13603 = n13602 ^ n13601 ;
  assign n13607 = n13606 ^ n13603 ;
  assign n13380 = n13373 ^ n13364 ;
  assign n13381 = n13370 & n13380 ;
  assign n13382 = n13381 ^ n13373 ;
  assign n13608 = n13607 ^ n13382 ;
  assign n13377 = n13136 ^ n13133 ;
  assign n13378 = n13375 & n13377 ;
  assign n13379 = n13378 ^ n13133 ;
  assign n13609 = n13608 ^ n13379 ;
  assign n13844 = n13591 ^ n13387 ;
  assign n13845 = n13597 & ~n13844 ;
  assign n13846 = n13845 ^ n13591 ;
  assign n13837 = x124 & n1050 ;
  assign n13836 = x126 & n1053 ;
  assign n13838 = n13837 ^ n13836 ;
  assign n13839 = n13838 ^ x17 ;
  assign n13835 = n1054 & n10441 ;
  assign n13840 = n13839 ^ n13835 ;
  assign n13834 = x125 & n1058 ;
  assign n13841 = n13840 ^ n13834 ;
  assign n13827 = x121 & n1327 ;
  assign n13826 = x123 & n1330 ;
  assign n13828 = n13827 ^ n13826 ;
  assign n13829 = n13828 ^ x20 ;
  assign n13825 = n1331 & ~n9786 ;
  assign n13830 = n13829 ^ n13825 ;
  assign n13824 = x122 & n1335 ;
  assign n13831 = n13830 ^ n13824 ;
  assign n13820 = x119 & n1666 ;
  assign n13810 = x115 & n2018 ;
  assign n13809 = x117 & n2021 ;
  assign n13811 = n13810 ^ n13809 ;
  assign n13812 = n13811 ^ x26 ;
  assign n13808 = n2022 & ~n7850 ;
  assign n13813 = n13812 ^ n13808 ;
  assign n13807 = x116 & n2014 ;
  assign n13814 = n13813 ^ n13807 ;
  assign n13796 = x112 & n2581 ;
  assign n13795 = x114 & n2422 ;
  assign n13797 = n13796 ^ n13795 ;
  assign n13798 = n13797 ^ x29 ;
  assign n13794 = n2423 & ~n7092 ;
  assign n13799 = n13798 ^ n13794 ;
  assign n13793 = x113 & n2429 ;
  assign n13800 = n13799 ^ n13793 ;
  assign n13782 = x109 & n2879 ;
  assign n13781 = x111 & n2882 ;
  assign n13783 = n13782 ^ n13781 ;
  assign n13784 = n13783 ^ x32 ;
  assign n13780 = n2883 & ~n6360 ;
  assign n13785 = n13784 ^ n13780 ;
  assign n13779 = x110 & n2887 ;
  assign n13786 = n13785 ^ n13779 ;
  assign n13772 = x106 & n3375 ;
  assign n13771 = x108 & n3378 ;
  assign n13773 = n13772 ^ n13771 ;
  assign n13774 = n13773 ^ x35 ;
  assign n13770 = n3379 & n5670 ;
  assign n13775 = n13774 ^ n13770 ;
  assign n13769 = x107 & n3383 ;
  assign n13776 = n13775 ^ n13769 ;
  assign n13758 = x103 & n3916 ;
  assign n13757 = x105 & n3919 ;
  assign n13759 = n13758 ^ n13757 ;
  assign n13760 = n13759 ^ x38 ;
  assign n13756 = n3920 & ~n5023 ;
  assign n13761 = n13760 ^ n13756 ;
  assign n13755 = x104 & n3924 ;
  assign n13762 = n13761 ^ n13755 ;
  assign n13752 = n13516 ^ n13411 ;
  assign n13753 = n13508 & ~n13752 ;
  assign n13744 = x100 & n4474 ;
  assign n13743 = x102 & n4471 ;
  assign n13745 = n13744 ^ n13743 ;
  assign n13746 = n13745 ^ x41 ;
  assign n13742 = n4410 & n4472 ;
  assign n13747 = n13746 ^ n13742 ;
  assign n13741 = x101 & n4467 ;
  assign n13748 = n13747 ^ n13741 ;
  assign n13733 = x98 & n5102 ;
  assign n13731 = n3843 & n5098 ;
  assign n13727 = x97 & n5094 ;
  assign n13726 = x99 & n5097 ;
  assign n13728 = n13727 ^ n13726 ;
  assign n13729 = n13728 ^ x44 ;
  assign n13723 = x95 & n5736 ;
  assign n13721 = n3323 & n5730 ;
  assign n13717 = x94 & n5965 ;
  assign n13716 = x96 & n5729 ;
  assign n13718 = n13717 ^ n13716 ;
  assign n13719 = n13718 ^ x47 ;
  assign n13709 = x91 & n6677 ;
  assign n13708 = x93 & n6428 ;
  assign n13710 = n13709 ^ n13708 ;
  assign n13711 = n13710 ^ x50 ;
  assign n13707 = n2836 & n6429 ;
  assign n13712 = n13711 ^ n13707 ;
  assign n13706 = x92 & n6433 ;
  assign n13713 = n13712 ^ n13706 ;
  assign n13702 = x86 & n7931 ;
  assign n13700 = n1982 & n7939 ;
  assign n13696 = x85 & n7935 ;
  assign n13695 = x87 & n7938 ;
  assign n13697 = n13696 ^ n13695 ;
  assign n13698 = n13697 ^ x56 ;
  assign n13688 = n1305 & n9636 ;
  assign n13687 = x80 & n9628 ;
  assign n13689 = n13688 ^ n13687 ;
  assign n13685 = x79 & n9632 ;
  assign n13684 = x81 & n9635 ;
  assign n13686 = n13685 ^ n13684 ;
  assign n13690 = n13689 ^ n13686 ;
  assign n13683 = n837 ^ x62 ;
  assign n13691 = n13690 ^ n13683 ;
  assign n13680 = n13452 ^ n13443 ;
  assign n13681 = ~n13444 & ~n13680 ;
  assign n13682 = n13681 ^ n13452 ;
  assign n13692 = n13691 ^ n13682 ;
  assign n13677 = x63 & x78 ;
  assign n13675 = x63 & n837 ;
  assign n13674 = n13438 ^ x78 ;
  assign n13676 = n13675 ^ n13674 ;
  assign n13678 = n13677 ^ n13676 ;
  assign n13679 = ~n9948 & n13678 ;
  assign n13693 = n13692 ^ n13679 ;
  assign n13669 = x82 & n8741 ;
  assign n13668 = x84 & n8744 ;
  assign n13670 = n13669 ^ n13668 ;
  assign n13671 = n13670 ^ x59 ;
  assign n13667 = n1624 & n8745 ;
  assign n13672 = n13671 ^ n13667 ;
  assign n13666 = x83 & n8737 ;
  assign n13673 = n13672 ^ n13666 ;
  assign n13694 = n13693 ^ n13673 ;
  assign n13699 = n13698 ^ n13694 ;
  assign n13701 = n13700 ^ n13699 ;
  assign n13703 = n13702 ^ n13701 ;
  assign n13663 = n13461 ^ n13436 ;
  assign n13664 = n13462 & n13663 ;
  assign n13665 = n13664 ^ n13461 ;
  assign n13704 = n13703 ^ n13665 ;
  assign n13653 = x88 & n7171 ;
  assign n13652 = x90 & n7174 ;
  assign n13654 = n13653 ^ n13652 ;
  assign n13655 = n13654 ^ x53 ;
  assign n13651 = n2386 & n7175 ;
  assign n13656 = n13655 ^ n13651 ;
  assign n13650 = x89 & n7179 ;
  assign n13657 = n13656 ^ n13650 ;
  assign n13659 = n13657 ^ n13428 ;
  assign n13658 = n13657 ^ n13463 ;
  assign n13660 = n13659 ^ n13658 ;
  assign n13661 = n13433 & n13660 ;
  assign n13662 = n13661 ^ n13659 ;
  assign n13705 = n13704 ^ n13662 ;
  assign n13714 = n13713 ^ n13705 ;
  assign n13647 = n13476 ^ n13472 ;
  assign n13648 = ~n13473 & n13647 ;
  assign n13649 = n13648 ^ n13476 ;
  assign n13715 = n13714 ^ n13649 ;
  assign n13720 = n13719 ^ n13715 ;
  assign n13722 = n13721 ^ n13720 ;
  assign n13724 = n13723 ^ n13722 ;
  assign n13644 = n13485 ^ n13420 ;
  assign n13645 = n13486 & n13644 ;
  assign n13646 = n13645 ^ n13485 ;
  assign n13725 = n13724 ^ n13646 ;
  assign n13730 = n13729 ^ n13725 ;
  assign n13732 = n13731 ^ n13730 ;
  assign n13734 = n13733 ^ n13732 ;
  assign n13641 = n13495 ^ n13417 ;
  assign n13642 = n13496 & n13641 ;
  assign n13643 = n13642 ^ n13495 ;
  assign n13735 = n13734 ^ n13643 ;
  assign n13736 = n13735 ^ n13497 ;
  assign n13737 = n13736 ^ n13414 ;
  assign n13738 = n13737 ^ n13735 ;
  assign n13739 = n13506 & n13738 ;
  assign n13740 = n13739 ^ n13736 ;
  assign n13749 = n13748 ^ n13740 ;
  assign n13750 = n13749 ^ n13516 ;
  assign n13754 = n13753 ^ n13750 ;
  assign n13763 = n13762 ^ n13754 ;
  assign n13764 = n13763 ^ n13526 ;
  assign n13765 = n13764 ^ n13763 ;
  assign n13766 = n13765 ^ n13408 ;
  assign n13767 = ~n13518 & ~n13766 ;
  assign n13768 = n13767 ^ n13764 ;
  assign n13777 = n13776 ^ n13768 ;
  assign n13638 = n13539 ^ n13530 ;
  assign n13639 = ~n13531 & n13638 ;
  assign n13640 = n13639 ^ n13539 ;
  assign n13778 = n13777 ^ n13640 ;
  assign n13787 = n13786 ^ n13778 ;
  assign n13788 = n13787 ^ n13548 ;
  assign n13789 = n13788 ^ n13787 ;
  assign n13790 = n13789 ^ n13405 ;
  assign n13791 = n13549 & n13790 ;
  assign n13792 = n13791 ^ n13788 ;
  assign n13801 = n13800 ^ n13792 ;
  assign n13803 = n13801 ^ n13550 ;
  assign n13802 = n13801 ^ n13563 ;
  assign n13804 = n13803 ^ n13802 ;
  assign n13805 = n13555 & n13804 ;
  assign n13806 = n13805 ^ n13803 ;
  assign n13815 = n13814 ^ n13806 ;
  assign n13816 = n13815 ^ x23 ;
  assign n13637 = x118 & n1658 ;
  assign n13817 = n13816 ^ n13637 ;
  assign n13636 = x120 & n1661 ;
  assign n13818 = n13817 ^ n13636 ;
  assign n13635 = n1662 & n8891 ;
  assign n13819 = n13818 ^ n13635 ;
  assign n13821 = n13820 ^ n13819 ;
  assign n13632 = n13573 ^ n13564 ;
  assign n13633 = ~n13570 & ~n13632 ;
  assign n13634 = n13633 ^ n13573 ;
  assign n13822 = n13821 ^ n13634 ;
  assign n13629 = n13583 ^ n13574 ;
  assign n13630 = n13580 & n13629 ;
  assign n13631 = n13630 ^ n13583 ;
  assign n13823 = n13822 ^ n13631 ;
  assign n13832 = n13831 ^ n13823 ;
  assign n13626 = n13584 ^ n13393 ;
  assign n13627 = n13590 & n13626 ;
  assign n13628 = n13627 ^ n13584 ;
  assign n13833 = n13832 ^ n13628 ;
  assign n13842 = n13841 ^ n13833 ;
  assign n13616 = x127 & n876 ;
  assign n13617 = n13616 ^ n781 ;
  assign n13622 = n641 & n11265 ;
  assign n13623 = n13622 ^ n13616 ;
  assign n13624 = n13617 & ~n13623 ;
  assign n13625 = n13624 ^ x13 ;
  assign n13843 = n13842 ^ n13625 ;
  assign n13847 = n13846 ^ n13843 ;
  assign n13613 = n13606 ^ n13598 ;
  assign n13614 = n13603 & ~n13613 ;
  assign n13615 = n13614 ^ n13606 ;
  assign n13848 = n13847 ^ n13615 ;
  assign n13610 = n13382 ^ n13379 ;
  assign n13611 = n13608 & n13610 ;
  assign n13612 = n13611 ^ n13382 ;
  assign n13849 = n13848 ^ n13612 ;
  assign n14080 = n13846 ^ n13615 ;
  assign n14081 = n14080 ^ n13612 ;
  assign n14082 = ~n13848 & n14081 ;
  assign n14075 = x126 & n1058 ;
  assign n14068 = x123 & n1335 ;
  assign n14060 = n13815 ^ n13634 ;
  assign n14061 = ~n13821 & n14060 ;
  assign n14062 = n14061 ^ n13815 ;
  assign n14058 = x120 & n1666 ;
  assign n14050 = n13814 ^ n13801 ;
  assign n14051 = ~n13806 & ~n14050 ;
  assign n14052 = n14051 ^ n13801 ;
  assign n14044 = x116 & n2018 ;
  assign n14043 = x118 & n2021 ;
  assign n14045 = n14044 ^ n14043 ;
  assign n14046 = n14045 ^ x26 ;
  assign n14042 = n2022 & ~n8123 ;
  assign n14047 = n14046 ^ n14042 ;
  assign n14041 = x117 & n2014 ;
  assign n14048 = n14047 ^ n14041 ;
  assign n14037 = n13800 ^ n13787 ;
  assign n14038 = ~n13792 & ~n14037 ;
  assign n14039 = n14038 ^ n13787 ;
  assign n14031 = x113 & n2581 ;
  assign n14030 = x115 & n2422 ;
  assign n14032 = n14031 ^ n14030 ;
  assign n14033 = n14032 ^ x29 ;
  assign n14029 = n2423 & ~n7343 ;
  assign n14034 = n14033 ^ n14029 ;
  assign n14028 = x114 & n2429 ;
  assign n14035 = n14034 ^ n14028 ;
  assign n14021 = x110 & n2879 ;
  assign n14020 = x112 & n2882 ;
  assign n14022 = n14021 ^ n14020 ;
  assign n14023 = n14022 ^ x32 ;
  assign n14019 = n2883 & ~n6600 ;
  assign n14024 = n14023 ^ n14019 ;
  assign n14018 = x111 & n2887 ;
  assign n14025 = n14024 ^ n14018 ;
  assign n14014 = n13776 ^ n13763 ;
  assign n14015 = ~n13768 & ~n14014 ;
  assign n14016 = n14015 ^ n13763 ;
  assign n14008 = x107 & n3375 ;
  assign n14007 = x109 & n3378 ;
  assign n14009 = n14008 ^ n14007 ;
  assign n14010 = n14009 ^ x35 ;
  assign n14006 = n3379 & n5902 ;
  assign n14011 = n14010 ^ n14006 ;
  assign n14005 = x108 & n3383 ;
  assign n14012 = n14011 ^ n14005 ;
  assign n14001 = n13762 ^ n13749 ;
  assign n14002 = ~n13754 & ~n14001 ;
  assign n14003 = n14002 ^ n13749 ;
  assign n13995 = x104 & n3916 ;
  assign n13994 = x106 & n3919 ;
  assign n13996 = n13995 ^ n13994 ;
  assign n13997 = n13996 ^ x38 ;
  assign n13993 = n3920 & ~n5240 ;
  assign n13998 = n13997 ^ n13993 ;
  assign n13992 = x105 & n3924 ;
  assign n13999 = n13998 ^ n13992 ;
  assign n13989 = x102 & n4467 ;
  assign n13987 = n4472 & ~n4615 ;
  assign n13983 = x101 & n4474 ;
  assign n13982 = x103 & n4471 ;
  assign n13984 = n13983 ^ n13982 ;
  assign n13985 = n13984 ^ x41 ;
  assign n13978 = n13725 ^ n13643 ;
  assign n13979 = ~n13734 & ~n13978 ;
  assign n13980 = n13979 ^ n13725 ;
  assign n13972 = x98 & n5094 ;
  assign n13971 = x100 & n5097 ;
  assign n13973 = n13972 ^ n13971 ;
  assign n13974 = n13973 ^ x44 ;
  assign n13970 = n4034 & n5098 ;
  assign n13975 = n13974 ^ n13970 ;
  assign n13969 = x99 & n5102 ;
  assign n13976 = n13975 ^ n13969 ;
  assign n13965 = n13715 ^ n13646 ;
  assign n13966 = ~n13724 & ~n13965 ;
  assign n13967 = n13966 ^ n13715 ;
  assign n13959 = x95 & n5965 ;
  assign n13958 = x97 & n5729 ;
  assign n13960 = n13959 ^ n13958 ;
  assign n13961 = n13960 ^ x47 ;
  assign n13957 = n3494 & n5730 ;
  assign n13962 = n13961 ^ n13957 ;
  assign n13956 = x96 & n5736 ;
  assign n13963 = n13962 ^ n13956 ;
  assign n13949 = x92 & n6677 ;
  assign n13948 = x94 & n6428 ;
  assign n13950 = n13949 ^ n13948 ;
  assign n13951 = n13950 ^ x50 ;
  assign n13947 = n2997 & n6429 ;
  assign n13952 = n13951 ^ n13947 ;
  assign n13946 = x93 & n6433 ;
  assign n13953 = n13952 ^ n13946 ;
  assign n13939 = x89 & n7171 ;
  assign n13938 = x91 & n7174 ;
  assign n13940 = n13939 ^ n13938 ;
  assign n13941 = n13940 ^ x53 ;
  assign n13937 = n2542 & n7175 ;
  assign n13942 = n13941 ^ n13937 ;
  assign n13936 = x90 & n7179 ;
  assign n13943 = n13942 ^ n13936 ;
  assign n13932 = n13694 ^ n13665 ;
  assign n13933 = ~n13703 & ~n13932 ;
  assign n13934 = n13933 ^ n13694 ;
  assign n13926 = x86 & n7935 ;
  assign n13925 = x88 & n7938 ;
  assign n13927 = n13926 ^ n13925 ;
  assign n13928 = n13927 ^ x56 ;
  assign n13924 = n2119 & n7939 ;
  assign n13929 = n13928 ^ n13924 ;
  assign n13923 = x87 & n7931 ;
  assign n13930 = n13929 ^ n13923 ;
  assign n13916 = x83 & n8741 ;
  assign n13915 = x85 & n8744 ;
  assign n13917 = n13916 ^ n13915 ;
  assign n13918 = n13917 ^ x59 ;
  assign n13914 = n1743 & n8745 ;
  assign n13919 = n13918 ^ n13914 ;
  assign n13913 = x84 & n8737 ;
  assign n13920 = n13919 ^ n13913 ;
  assign n13906 = x80 & n9632 ;
  assign n13905 = x82 & n9635 ;
  assign n13907 = n13906 ^ n13905 ;
  assign n13908 = n13907 ^ x62 ;
  assign n13904 = n1411 & n9636 ;
  assign n13909 = n13908 ^ n13904 ;
  assign n13903 = x81 & n9628 ;
  assign n13910 = n13909 ^ n13903 ;
  assign n13898 = n13677 ^ x79 ;
  assign n13899 = ~n9948 & n13898 ;
  assign n13900 = n13899 ^ x79 ;
  assign n13901 = n13900 ^ x14 ;
  assign n13902 = n13901 ^ n13440 ;
  assign n13911 = n13910 ^ n13902 ;
  assign n13882 = n13690 ^ x78 ;
  assign n13892 = ~n13675 & n13882 ;
  assign n13893 = n13892 ^ x78 ;
  assign n753 = x77 ^ x76 ;
  assign n13888 = n13690 ^ x76 ;
  assign n13889 = ~n753 & n13888 ;
  assign n13890 = n13889 ^ x76 ;
  assign n13891 = x63 & n13890 ;
  assign n13894 = n13893 ^ n13891 ;
  assign n13895 = x62 & ~n13894 ;
  assign n13896 = n13895 ^ n13893 ;
  assign n13885 = ~n837 & ~n13882 ;
  assign n13886 = n13885 ^ x78 ;
  assign n13887 = n11874 & ~n13886 ;
  assign n13897 = n13896 ^ n13887 ;
  assign n13912 = n13911 ^ n13897 ;
  assign n13921 = n13920 ^ n13912 ;
  assign n13879 = n13682 ^ n13673 ;
  assign n13880 = n13693 & n13879 ;
  assign n13881 = n13880 ^ n13673 ;
  assign n13922 = n13921 ^ n13881 ;
  assign n13931 = n13930 ^ n13922 ;
  assign n13935 = n13934 ^ n13931 ;
  assign n13944 = n13943 ^ n13935 ;
  assign n13876 = n13704 ^ n13657 ;
  assign n13877 = n13662 & ~n13876 ;
  assign n13878 = n13877 ^ n13657 ;
  assign n13945 = n13944 ^ n13878 ;
  assign n13954 = n13953 ^ n13945 ;
  assign n13873 = n13705 ^ n13649 ;
  assign n13874 = ~n13714 & n13873 ;
  assign n13875 = n13874 ^ n13713 ;
  assign n13955 = n13954 ^ n13875 ;
  assign n13964 = n13963 ^ n13955 ;
  assign n13968 = n13967 ^ n13964 ;
  assign n13977 = n13976 ^ n13968 ;
  assign n13981 = n13980 ^ n13977 ;
  assign n13986 = n13985 ^ n13981 ;
  assign n13988 = n13987 ^ n13986 ;
  assign n13990 = n13989 ^ n13988 ;
  assign n13870 = n13748 ^ n13735 ;
  assign n13871 = ~n13740 & ~n13870 ;
  assign n13872 = n13871 ^ n13735 ;
  assign n13991 = n13990 ^ n13872 ;
  assign n14000 = n13999 ^ n13991 ;
  assign n14004 = n14003 ^ n14000 ;
  assign n14013 = n14012 ^ n14004 ;
  assign n14017 = n14016 ^ n14013 ;
  assign n14026 = n14025 ^ n14017 ;
  assign n13867 = n13786 ^ n13640 ;
  assign n13868 = n13778 & n13867 ;
  assign n13869 = n13868 ^ n13786 ;
  assign n14027 = n14026 ^ n13869 ;
  assign n14036 = n14035 ^ n14027 ;
  assign n14040 = n14039 ^ n14036 ;
  assign n14049 = n14048 ^ n14040 ;
  assign n14053 = n14052 ^ n14049 ;
  assign n14054 = n14053 ^ x23 ;
  assign n13866 = x119 & n1658 ;
  assign n14055 = n14054 ^ n13866 ;
  assign n13865 = x121 & n1661 ;
  assign n14056 = n14055 ^ n13865 ;
  assign n13864 = n1662 & n8962 ;
  assign n14057 = n14056 ^ n13864 ;
  assign n14059 = n14058 ^ n14057 ;
  assign n14063 = n14062 ^ n14059 ;
  assign n14064 = n14063 ^ x20 ;
  assign n13863 = x122 & n1327 ;
  assign n14065 = n14064 ^ n13863 ;
  assign n13862 = x124 & n1330 ;
  assign n14066 = n14065 ^ n13862 ;
  assign n13861 = n1331 & n10095 ;
  assign n14067 = n14066 ^ n13861 ;
  assign n14069 = n14068 ^ n14067 ;
  assign n13858 = n13831 ^ n13631 ;
  assign n13859 = n13823 & ~n13858 ;
  assign n13860 = n13859 ^ n13831 ;
  assign n14070 = n14069 ^ n13860 ;
  assign n14071 = n14070 ^ x17 ;
  assign n13857 = x125 & n1050 ;
  assign n14072 = n14071 ^ n13857 ;
  assign n13856 = x127 & n1053 ;
  assign n14073 = n14072 ^ n13856 ;
  assign n13855 = n1054 & n10972 ;
  assign n14074 = n14073 ^ n13855 ;
  assign n14076 = n14075 ^ n14074 ;
  assign n13852 = n13841 ^ n13628 ;
  assign n13853 = n13833 & n13852 ;
  assign n13854 = n13853 ^ n13841 ;
  assign n14077 = n14076 ^ n13854 ;
  assign n13851 = ~n13625 & n13842 ;
  assign n14078 = n14077 ^ n13851 ;
  assign n13850 = n13615 & n13846 ;
  assign n14079 = n14078 ^ n13850 ;
  assign n14083 = n14082 ^ n14079 ;
  assign n14319 = n1054 & n10139 ;
  assign n14318 = x126 & n1050 ;
  assign n14320 = n14319 ^ n14318 ;
  assign n14321 = n14320 ^ x17 ;
  assign n14317 = x127 & n1058 ;
  assign n14322 = n14321 ^ n14317 ;
  assign n14313 = n14063 ^ n13860 ;
  assign n14314 = n14069 & n14313 ;
  assign n14315 = n14314 ^ n14063 ;
  assign n14307 = x123 & n1327 ;
  assign n14306 = x125 & n1330 ;
  assign n14308 = n14307 ^ n14306 ;
  assign n14309 = n14308 ^ x20 ;
  assign n14305 = n1331 & n10400 ;
  assign n14310 = n14309 ^ n14305 ;
  assign n14304 = x124 & n1335 ;
  assign n14311 = n14310 ^ n14304 ;
  assign n14297 = x120 & n1658 ;
  assign n14296 = x122 & n1661 ;
  assign n14298 = n14297 ^ n14296 ;
  assign n14299 = n14298 ^ x23 ;
  assign n14295 = n1662 & ~n9247 ;
  assign n14300 = n14299 ^ n14295 ;
  assign n14294 = x121 & n1666 ;
  assign n14301 = n14300 ^ n14294 ;
  assign n14286 = x117 & n2018 ;
  assign n14285 = x119 & n2021 ;
  assign n14287 = n14286 ^ n14285 ;
  assign n14288 = n14287 ^ x26 ;
  assign n14284 = n2022 & n8394 ;
  assign n14289 = n14288 ^ n14284 ;
  assign n14283 = x118 & n2014 ;
  assign n14290 = n14289 ^ n14283 ;
  assign n14277 = x114 & n2581 ;
  assign n14276 = x116 & n2422 ;
  assign n14278 = n14277 ^ n14276 ;
  assign n14279 = n14278 ^ x29 ;
  assign n14275 = n2423 & ~n7588 ;
  assign n14280 = n14279 ^ n14275 ;
  assign n14274 = x115 & n2429 ;
  assign n14281 = n14280 ^ n14274 ;
  assign n14270 = n14025 ^ n13869 ;
  assign n14271 = ~n14026 & n14270 ;
  assign n14272 = n14271 ^ n14025 ;
  assign n14264 = x111 & n2879 ;
  assign n14263 = x113 & n2882 ;
  assign n14265 = n14264 ^ n14263 ;
  assign n14266 = n14265 ^ x32 ;
  assign n14262 = n2883 & ~n6839 ;
  assign n14267 = n14266 ^ n14262 ;
  assign n14261 = x112 & n2887 ;
  assign n14268 = n14267 ^ n14261 ;
  assign n14249 = x105 & n3916 ;
  assign n14248 = x107 & n3919 ;
  assign n14250 = n14249 ^ n14248 ;
  assign n14251 = n14250 ^ x38 ;
  assign n14247 = n3920 & ~n5448 ;
  assign n14252 = n14251 ^ n14247 ;
  assign n14246 = x106 & n3924 ;
  assign n14253 = n14252 ^ n14246 ;
  assign n14242 = n13981 ^ n13872 ;
  assign n14243 = n13990 & ~n14242 ;
  assign n14244 = n14243 ^ n13981 ;
  assign n14236 = x102 & n4474 ;
  assign n14235 = x104 & n4471 ;
  assign n14237 = n14236 ^ n14235 ;
  assign n14238 = n14237 ^ x41 ;
  assign n14234 = n4472 & ~n4814 ;
  assign n14239 = n14238 ^ n14234 ;
  assign n14233 = x103 & n4467 ;
  assign n14240 = n14239 ^ n14233 ;
  assign n14229 = x100 & n5102 ;
  assign n14227 = n4215 & n5098 ;
  assign n14223 = x99 & n5094 ;
  assign n14222 = x101 & n5097 ;
  assign n14224 = n14223 ^ n14222 ;
  assign n14225 = n14224 ^ x44 ;
  assign n14219 = n13967 ^ n13963 ;
  assign n14220 = ~n13964 & ~n14219 ;
  assign n14221 = n14220 ^ n13967 ;
  assign n14226 = n14225 ^ n14221 ;
  assign n14228 = n14227 ^ n14226 ;
  assign n14230 = n14229 ^ n14228 ;
  assign n14215 = n13953 ^ n13875 ;
  assign n14216 = n13954 & n14215 ;
  assign n14217 = n14216 ^ n13953 ;
  assign n14209 = x96 & n5965 ;
  assign n14208 = x98 & n5729 ;
  assign n14210 = n14209 ^ n14208 ;
  assign n14211 = n14210 ^ x47 ;
  assign n14207 = n3660 & n5730 ;
  assign n14212 = n14211 ^ n14207 ;
  assign n14206 = x97 & n5736 ;
  assign n14213 = n14212 ^ n14206 ;
  assign n14199 = x93 & n6677 ;
  assign n14198 = x95 & n6428 ;
  assign n14200 = n14199 ^ n14198 ;
  assign n14201 = n14200 ^ x50 ;
  assign n14197 = n3159 & n6429 ;
  assign n14202 = n14201 ^ n14197 ;
  assign n14196 = x94 & n6433 ;
  assign n14203 = n14202 ^ n14196 ;
  assign n14190 = n13910 ^ n13897 ;
  assign n14191 = ~n13911 & n14190 ;
  assign n14192 = n14191 ^ n13910 ;
  assign n14184 = ~x63 & n1009 ;
  assign n14185 = n14184 ^ x79 ;
  assign n14161 = x63 & x80 ;
  assign n14187 = n14185 ^ n14161 ;
  assign n14188 = x62 & ~n14187 ;
  assign n14180 = n1512 & n9636 ;
  assign n14179 = x82 & n9628 ;
  assign n14181 = n14180 ^ n14179 ;
  assign n14177 = x81 & n9632 ;
  assign n14176 = x83 & n9635 ;
  assign n14178 = n14177 ^ n14176 ;
  assign n14182 = n14181 ^ n14178 ;
  assign n14170 = x84 & n8741 ;
  assign n14169 = x86 & n8744 ;
  assign n14171 = n14170 ^ n14169 ;
  assign n14172 = n14171 ^ x59 ;
  assign n14168 = n1857 & n8745 ;
  assign n14173 = n14172 ^ n14168 ;
  assign n14167 = x85 & n8737 ;
  assign n14174 = n14173 ^ n14167 ;
  assign n14162 = n13440 ^ x14 ;
  assign n14163 = n13900 ^ n13440 ;
  assign n14164 = ~n14162 & ~n14163 ;
  assign n14165 = n14164 ^ x14 ;
  assign n14166 = n14165 ^ n14161 ;
  assign n14175 = n14174 ^ n14166 ;
  assign n14183 = n14182 ^ n14175 ;
  assign n14189 = n14188 ^ n14183 ;
  assign n14193 = n14192 ^ n14189 ;
  assign n14151 = x87 & n7935 ;
  assign n14150 = x89 & n7938 ;
  assign n14152 = n14151 ^ n14150 ;
  assign n14153 = n14152 ^ x56 ;
  assign n14149 = n2249 & n7939 ;
  assign n14154 = n14153 ^ n14149 ;
  assign n14148 = x88 & n7931 ;
  assign n14155 = n14154 ^ n14148 ;
  assign n14156 = n14155 ^ n13920 ;
  assign n14157 = n14156 ^ n13881 ;
  assign n14158 = n14157 ^ n14155 ;
  assign n14159 = ~n13921 & n14158 ;
  assign n14160 = n14159 ^ n14156 ;
  assign n14194 = n14193 ^ n14160 ;
  assign n14138 = x90 & n7171 ;
  assign n14137 = x92 & n7174 ;
  assign n14139 = n14138 ^ n14137 ;
  assign n14140 = n14139 ^ x53 ;
  assign n14136 = n2684 & n7175 ;
  assign n14141 = n14140 ^ n14136 ;
  assign n14135 = x91 & n7179 ;
  assign n14142 = n14141 ^ n14135 ;
  assign n14143 = n14142 ^ n13934 ;
  assign n14144 = n14143 ^ n13930 ;
  assign n14145 = n14144 ^ n14142 ;
  assign n14146 = n13931 & ~n14145 ;
  assign n14147 = n14146 ^ n14143 ;
  assign n14195 = n14194 ^ n14147 ;
  assign n14204 = n14203 ^ n14195 ;
  assign n14132 = n13943 ^ n13878 ;
  assign n14133 = n13944 & n14132 ;
  assign n14134 = n14133 ^ n13943 ;
  assign n14205 = n14204 ^ n14134 ;
  assign n14214 = n14213 ^ n14205 ;
  assign n14218 = n14217 ^ n14214 ;
  assign n14231 = n14230 ^ n14218 ;
  assign n14129 = n13980 ^ n13976 ;
  assign n14130 = n13977 & ~n14129 ;
  assign n14131 = n14130 ^ n13980 ;
  assign n14232 = n14231 ^ n14131 ;
  assign n14241 = n14240 ^ n14232 ;
  assign n14245 = n14244 ^ n14241 ;
  assign n14254 = n14253 ^ n14245 ;
  assign n14126 = n3379 & n6129 ;
  assign n14124 = x108 & n3375 ;
  assign n14120 = n14003 ^ n13999 ;
  assign n14121 = n14000 & ~n14120 ;
  assign n14122 = n14121 ^ n14003 ;
  assign n14118 = x110 & n3378 ;
  assign n14119 = n14118 ^ x35 ;
  assign n14123 = n14122 ^ n14119 ;
  assign n14125 = n14124 ^ n14123 ;
  assign n14127 = n14126 ^ n14125 ;
  assign n14117 = x109 & n3383 ;
  assign n14128 = n14127 ^ n14117 ;
  assign n14255 = n14254 ^ n14128 ;
  assign n14256 = n14255 ^ n14016 ;
  assign n14257 = n14256 ^ n14012 ;
  assign n14258 = n14257 ^ n14255 ;
  assign n14259 = ~n14013 & ~n14258 ;
  assign n14260 = n14259 ^ n14256 ;
  assign n14269 = n14268 ^ n14260 ;
  assign n14273 = n14272 ^ n14269 ;
  assign n14282 = n14281 ^ n14273 ;
  assign n14291 = n14290 ^ n14282 ;
  assign n14114 = n14039 ^ n14035 ;
  assign n14115 = n14036 & ~n14114 ;
  assign n14116 = n14115 ^ n14039 ;
  assign n14292 = n14291 ^ n14116 ;
  assign n14111 = n14052 ^ n14048 ;
  assign n14112 = ~n14049 & ~n14111 ;
  assign n14113 = n14112 ^ n14052 ;
  assign n14293 = n14292 ^ n14113 ;
  assign n14302 = n14301 ^ n14293 ;
  assign n14108 = n14062 ^ n14053 ;
  assign n14109 = n14059 & n14108 ;
  assign n14110 = n14109 ^ n14062 ;
  assign n14303 = n14302 ^ n14110 ;
  assign n14312 = n14311 ^ n14303 ;
  assign n14316 = n14315 ^ n14312 ;
  assign n14323 = n14322 ^ n14316 ;
  assign n14105 = n14070 ^ n13854 ;
  assign n14106 = n14076 & n14105 ;
  assign n14107 = n14106 ^ n14070 ;
  assign n14324 = n14323 ^ n14107 ;
  assign n14084 = n13851 ^ n13843 ;
  assign n14085 = n14077 ^ n13850 ;
  assign n14086 = n14085 ^ n14080 ;
  assign n14087 = ~n14084 & n14086 ;
  assign n14088 = ~n13612 & n14087 ;
  assign n14089 = n14085 ^ n14077 ;
  assign n14090 = n14085 ^ n13851 ;
  assign n14091 = n14090 ^ n14085 ;
  assign n14092 = n14089 & n14091 ;
  assign n14093 = n14092 ^ n14085 ;
  assign n14094 = n14088 & n14093 ;
  assign n14095 = n14094 ^ n14087 ;
  assign n14096 = n13846 ^ n13612 ;
  assign n14097 = n13615 ^ n13612 ;
  assign n14098 = ~n14096 & ~n14097 ;
  assign n14099 = n14098 ^ n13612 ;
  assign n14100 = ~n14095 & n14099 ;
  assign n14102 = ~n13851 & n14077 ;
  assign n14103 = n14100 & n14102 ;
  assign n14101 = n14100 ^ n14095 ;
  assign n14104 = n14103 ^ n14101 ;
  assign n14325 = n14324 ^ n14104 ;
  assign n14543 = x127 & n1049 ;
  assign n14544 = n14543 ^ n1047 ;
  assign n14549 = n869 & n11265 ;
  assign n14550 = n14549 ^ n14543 ;
  assign n14551 = n14544 & ~n14550 ;
  assign n14552 = n14551 ^ x16 ;
  assign n14537 = x124 & n1327 ;
  assign n14536 = x126 & n1330 ;
  assign n14538 = n14537 ^ n14536 ;
  assign n14539 = n14538 ^ x20 ;
  assign n14535 = n1331 & n10441 ;
  assign n14540 = n14539 ^ n14535 ;
  assign n14534 = x125 & n1335 ;
  assign n14541 = n14540 ^ n14534 ;
  assign n14527 = x121 & n1658 ;
  assign n14526 = x123 & n1661 ;
  assign n14528 = n14527 ^ n14526 ;
  assign n14529 = n14528 ^ x23 ;
  assign n14525 = n1662 & ~n9786 ;
  assign n14530 = n14529 ^ n14525 ;
  assign n14524 = x122 & n1666 ;
  assign n14531 = n14530 ^ n14524 ;
  assign n14517 = x118 & n2018 ;
  assign n14516 = x120 & n2021 ;
  assign n14518 = n14517 ^ n14516 ;
  assign n14519 = n14518 ^ x26 ;
  assign n14515 = n2022 & n8891 ;
  assign n14520 = n14519 ^ n14515 ;
  assign n14514 = x119 & n2014 ;
  assign n14521 = n14520 ^ n14514 ;
  assign n14503 = x115 & n2581 ;
  assign n14502 = x117 & n2422 ;
  assign n14504 = n14503 ^ n14502 ;
  assign n14505 = n14504 ^ x29 ;
  assign n14501 = n2423 & ~n7850 ;
  assign n14506 = n14505 ^ n14501 ;
  assign n14500 = x116 & n2429 ;
  assign n14507 = n14506 ^ n14500 ;
  assign n14489 = x112 & n2879 ;
  assign n14488 = x114 & n2882 ;
  assign n14490 = n14489 ^ n14488 ;
  assign n14491 = n14490 ^ x32 ;
  assign n14487 = n2883 & ~n7092 ;
  assign n14492 = n14491 ^ n14487 ;
  assign n14486 = x113 & n2887 ;
  assign n14493 = n14492 ^ n14486 ;
  assign n14475 = x109 & n3375 ;
  assign n14474 = x111 & n3378 ;
  assign n14476 = n14475 ^ n14474 ;
  assign n14477 = n14476 ^ x35 ;
  assign n14473 = n3379 & ~n6360 ;
  assign n14478 = n14477 ^ n14473 ;
  assign n14472 = x110 & n3383 ;
  assign n14479 = n14478 ^ n14472 ;
  assign n14465 = x106 & n3916 ;
  assign n14464 = x108 & n3919 ;
  assign n14466 = n14465 ^ n14464 ;
  assign n14467 = n14466 ^ x38 ;
  assign n14463 = n3920 & n5670 ;
  assign n14468 = n14467 ^ n14463 ;
  assign n14462 = x107 & n3924 ;
  assign n14469 = n14468 ^ n14462 ;
  assign n14459 = n14240 ^ n14131 ;
  assign n14460 = n14232 & ~n14459 ;
  assign n14451 = x103 & n4474 ;
  assign n14450 = x105 & n4471 ;
  assign n14452 = n14451 ^ n14450 ;
  assign n14453 = n14452 ^ x41 ;
  assign n14449 = n4472 & ~n5023 ;
  assign n14454 = n14453 ^ n14449 ;
  assign n14448 = x104 & n4467 ;
  assign n14455 = n14454 ^ n14448 ;
  assign n14444 = n14221 ^ n14218 ;
  assign n14445 = n14230 & n14444 ;
  assign n14446 = n14445 ^ n14218 ;
  assign n14441 = x101 & n5102 ;
  assign n14439 = n4410 & n5098 ;
  assign n14435 = x100 & n5094 ;
  assign n14434 = x102 & n5097 ;
  assign n14436 = n14435 ^ n14434 ;
  assign n14437 = n14436 ^ x44 ;
  assign n14429 = n14194 ^ n14142 ;
  assign n14430 = ~n14147 & n14429 ;
  assign n14431 = n14430 ^ n14142 ;
  assign n14427 = x95 & n6433 ;
  assign n14422 = x94 & n6677 ;
  assign n14421 = x96 & n6428 ;
  assign n14423 = n14422 ^ n14421 ;
  assign n14424 = n14423 ^ x50 ;
  assign n14420 = n3323 & n6429 ;
  assign n14425 = n14424 ^ n14420 ;
  assign n14416 = n14193 ^ n14155 ;
  assign n14417 = n14160 & n14416 ;
  assign n14418 = n14417 ^ n14155 ;
  assign n14414 = x92 & n7179 ;
  assign n14409 = x91 & n7171 ;
  assign n14408 = x93 & n7174 ;
  assign n14410 = n14409 ^ n14408 ;
  assign n14411 = n14410 ^ x53 ;
  assign n14407 = n2836 & n7175 ;
  assign n14412 = n14411 ^ n14407 ;
  assign n14401 = x88 & n7935 ;
  assign n14400 = x90 & n7938 ;
  assign n14402 = n14401 ^ n14400 ;
  assign n14403 = n14402 ^ x56 ;
  assign n14399 = n2386 & n7939 ;
  assign n14404 = n14403 ^ n14399 ;
  assign n14398 = x89 & n7931 ;
  assign n14405 = n14404 ^ n14398 ;
  assign n14394 = n14192 ^ n14174 ;
  assign n14395 = n14189 & n14394 ;
  assign n14396 = n14395 ^ n14174 ;
  assign n14381 = n14165 ^ x62 ;
  assign n14382 = n14381 ^ n14182 ;
  assign n14383 = n14185 ^ n14182 ;
  assign n14384 = n14383 ^ n14166 ;
  assign n14387 = n14187 & ~n14384 ;
  assign n14388 = n14387 ^ n14166 ;
  assign n14389 = ~n14382 & n14388 ;
  assign n14390 = n14389 ^ n14165 ;
  assign n14378 = x80 ^ x62 ;
  assign n14379 = n14378 ^ x81 ;
  assign n14375 = n1624 & n9636 ;
  assign n14374 = x83 & n9628 ;
  assign n14376 = n14375 ^ n14374 ;
  assign n14372 = x82 & n9632 ;
  assign n14371 = x84 & n9635 ;
  assign n14373 = n14372 ^ n14371 ;
  assign n14377 = n14376 ^ n14373 ;
  assign n14380 = n14379 ^ n14377 ;
  assign n14391 = n14390 ^ n14380 ;
  assign n14369 = n14185 ^ x81 ;
  assign n14370 = ~n9948 & n14369 ;
  assign n14392 = n14391 ^ n14370 ;
  assign n14364 = x85 & n8741 ;
  assign n14363 = x87 & n8744 ;
  assign n14365 = n14364 ^ n14363 ;
  assign n14366 = n14365 ^ x59 ;
  assign n14362 = n1982 & n8745 ;
  assign n14367 = n14366 ^ n14362 ;
  assign n14361 = x86 & n8737 ;
  assign n14368 = n14367 ^ n14361 ;
  assign n14393 = n14392 ^ n14368 ;
  assign n14397 = n14396 ^ n14393 ;
  assign n14406 = n14405 ^ n14397 ;
  assign n14413 = n14412 ^ n14406 ;
  assign n14415 = n14414 ^ n14413 ;
  assign n14419 = n14418 ^ n14415 ;
  assign n14426 = n14425 ^ n14419 ;
  assign n14428 = n14427 ^ n14426 ;
  assign n14432 = n14431 ^ n14428 ;
  assign n14358 = n3843 & n5730 ;
  assign n14356 = x97 & n5965 ;
  assign n14354 = x99 & n5729 ;
  assign n14350 = n14203 ^ n14134 ;
  assign n14351 = ~n14204 & n14350 ;
  assign n14352 = n14351 ^ n14203 ;
  assign n14353 = n14352 ^ x47 ;
  assign n14355 = n14354 ^ n14353 ;
  assign n14357 = n14356 ^ n14355 ;
  assign n14359 = n14358 ^ n14357 ;
  assign n14349 = x98 & n5736 ;
  assign n14360 = n14359 ^ n14349 ;
  assign n14433 = n14432 ^ n14360 ;
  assign n14438 = n14437 ^ n14433 ;
  assign n14440 = n14439 ^ n14438 ;
  assign n14442 = n14441 ^ n14440 ;
  assign n14346 = n14217 ^ n14213 ;
  assign n14347 = n14214 & n14346 ;
  assign n14348 = n14347 ^ n14217 ;
  assign n14443 = n14442 ^ n14348 ;
  assign n14447 = n14446 ^ n14443 ;
  assign n14456 = n14455 ^ n14447 ;
  assign n14457 = n14456 ^ n14240 ;
  assign n14461 = n14460 ^ n14457 ;
  assign n14470 = n14469 ^ n14461 ;
  assign n14343 = n14253 ^ n14244 ;
  assign n14344 = n14245 & n14343 ;
  assign n14345 = n14344 ^ n14253 ;
  assign n14471 = n14470 ^ n14345 ;
  assign n14480 = n14479 ^ n14471 ;
  assign n14481 = n14480 ^ n14254 ;
  assign n14482 = n14481 ^ n14480 ;
  assign n14483 = n14482 ^ n14122 ;
  assign n14484 = n14128 & n14483 ;
  assign n14485 = n14484 ^ n14481 ;
  assign n14494 = n14493 ^ n14485 ;
  assign n14496 = n14494 ^ n14255 ;
  assign n14495 = n14494 ^ n14268 ;
  assign n14497 = n14496 ^ n14495 ;
  assign n14498 = ~n14260 & n14497 ;
  assign n14499 = n14498 ^ n14496 ;
  assign n14508 = n14507 ^ n14499 ;
  assign n14509 = n14508 ^ n14281 ;
  assign n14510 = n14509 ^ n14272 ;
  assign n14511 = n14510 ^ n14508 ;
  assign n14512 = n14273 & n14511 ;
  assign n14513 = n14512 ^ n14509 ;
  assign n14522 = n14521 ^ n14513 ;
  assign n14340 = n14290 ^ n14116 ;
  assign n14341 = ~n14291 & ~n14340 ;
  assign n14342 = n14341 ^ n14290 ;
  assign n14523 = n14522 ^ n14342 ;
  assign n14532 = n14531 ^ n14523 ;
  assign n14337 = n14301 ^ n14113 ;
  assign n14338 = n14293 & ~n14337 ;
  assign n14339 = n14338 ^ n14301 ;
  assign n14533 = n14532 ^ n14339 ;
  assign n14542 = n14541 ^ n14533 ;
  assign n14553 = n14552 ^ n14542 ;
  assign n14334 = n14311 ^ n14110 ;
  assign n14335 = ~n14303 & ~n14334 ;
  assign n14336 = n14335 ^ n14311 ;
  assign n14554 = n14553 ^ n14336 ;
  assign n14329 = n14322 ^ n14312 ;
  assign n14331 = n14315 ^ n14107 ;
  assign n14330 = n14312 ^ n14104 ;
  assign n14332 = n14331 ^ n14330 ;
  assign n14333 = ~n14329 & ~n14332 ;
  assign n14555 = n14554 ^ n14333 ;
  assign n14326 = n14315 ^ n14104 ;
  assign n14327 = n14107 ^ n14104 ;
  assign n14328 = n14326 & n14327 ;
  assign n14556 = n14555 ^ n14328 ;
  assign n14808 = n14552 ^ n14336 ;
  assign n14809 = n14553 & n14808 ;
  assign n14810 = n14809 ^ n14552 ;
  assign n14801 = x125 & n1327 ;
  assign n14800 = x127 & n1330 ;
  assign n14802 = n14801 ^ n14800 ;
  assign n14803 = n14802 ^ x20 ;
  assign n14799 = n1331 & n10972 ;
  assign n14804 = n14803 ^ n14799 ;
  assign n14798 = x126 & n1335 ;
  assign n14805 = n14804 ^ n14798 ;
  assign n14791 = x122 & n1658 ;
  assign n14790 = x124 & n1661 ;
  assign n14792 = n14791 ^ n14790 ;
  assign n14793 = n14792 ^ x23 ;
  assign n14789 = n1662 & n10095 ;
  assign n14794 = n14793 ^ n14789 ;
  assign n14788 = x123 & n1666 ;
  assign n14795 = n14794 ^ n14788 ;
  assign n14782 = x119 & n2018 ;
  assign n14781 = x121 & n2021 ;
  assign n14783 = n14782 ^ n14781 ;
  assign n14784 = n14783 ^ x26 ;
  assign n14780 = n2022 & n8962 ;
  assign n14785 = n14784 ^ n14780 ;
  assign n14779 = x120 & n2014 ;
  assign n14786 = n14785 ^ n14779 ;
  assign n14770 = n14507 ^ n14494 ;
  assign n14771 = n14499 & n14770 ;
  assign n14772 = n14771 ^ n14494 ;
  assign n14764 = x116 & n2581 ;
  assign n14763 = x118 & n2422 ;
  assign n14765 = n14764 ^ n14763 ;
  assign n14766 = n14765 ^ x29 ;
  assign n14762 = n2423 & ~n8123 ;
  assign n14767 = n14766 ^ n14762 ;
  assign n14761 = x117 & n2429 ;
  assign n14768 = n14767 ^ n14761 ;
  assign n14757 = n14493 ^ n14480 ;
  assign n14758 = n14485 & ~n14757 ;
  assign n14759 = n14758 ^ n14480 ;
  assign n14751 = x113 & n2879 ;
  assign n14750 = x115 & n2882 ;
  assign n14752 = n14751 ^ n14750 ;
  assign n14753 = n14752 ^ x32 ;
  assign n14749 = n2883 & ~n7343 ;
  assign n14754 = n14753 ^ n14749 ;
  assign n14748 = x114 & n2887 ;
  assign n14755 = n14754 ^ n14748 ;
  assign n14744 = n14479 ^ n14345 ;
  assign n14745 = n14471 & n14744 ;
  assign n14746 = n14745 ^ n14479 ;
  assign n14742 = x111 & n3383 ;
  assign n14737 = x110 & n3375 ;
  assign n14736 = x112 & n3378 ;
  assign n14738 = n14737 ^ n14736 ;
  assign n14739 = n14738 ^ x35 ;
  assign n14735 = n3379 & ~n6600 ;
  assign n14740 = n14739 ^ n14735 ;
  assign n14731 = n14469 ^ n14456 ;
  assign n14732 = ~n14461 & ~n14731 ;
  assign n14733 = n14732 ^ n14456 ;
  assign n14725 = x107 & n3916 ;
  assign n14724 = x109 & n3919 ;
  assign n14726 = n14725 ^ n14724 ;
  assign n14727 = n14726 ^ x38 ;
  assign n14723 = n3920 & n5902 ;
  assign n14728 = n14727 ^ n14723 ;
  assign n14722 = x108 & n3924 ;
  assign n14729 = n14728 ^ n14722 ;
  assign n14715 = x104 & n4474 ;
  assign n14714 = x106 & n4471 ;
  assign n14716 = n14715 ^ n14714 ;
  assign n14717 = n14716 ^ x41 ;
  assign n14713 = n4472 & ~n5240 ;
  assign n14718 = n14717 ^ n14713 ;
  assign n14712 = x105 & n4467 ;
  assign n14719 = n14718 ^ n14712 ;
  assign n14708 = n14433 ^ n14348 ;
  assign n14709 = n14442 & n14708 ;
  assign n14710 = n14709 ^ n14433 ;
  assign n14702 = x101 & n5094 ;
  assign n14701 = x103 & n5097 ;
  assign n14703 = n14702 ^ n14701 ;
  assign n14704 = n14703 ^ x44 ;
  assign n14700 = ~n4615 & n5098 ;
  assign n14705 = n14704 ^ n14700 ;
  assign n14699 = x102 & n5102 ;
  assign n14706 = n14705 ^ n14699 ;
  assign n14695 = n14432 ^ n14352 ;
  assign n14696 = ~n14360 & n14695 ;
  assign n14697 = n14696 ^ n14432 ;
  assign n14689 = x98 & n5965 ;
  assign n14688 = x100 & n5729 ;
  assign n14690 = n14689 ^ n14688 ;
  assign n14691 = n14690 ^ x47 ;
  assign n14687 = n4034 & n5730 ;
  assign n14692 = n14691 ^ n14687 ;
  assign n14686 = x99 & n5736 ;
  assign n14693 = n14692 ^ n14686 ;
  assign n14679 = x95 & n6677 ;
  assign n14678 = x97 & n6428 ;
  assign n14680 = n14679 ^ n14678 ;
  assign n14681 = n14680 ^ x50 ;
  assign n14677 = n3494 & n6429 ;
  assign n14682 = n14681 ^ n14677 ;
  assign n14676 = x96 & n6433 ;
  assign n14683 = n14682 ^ n14676 ;
  assign n14669 = x92 & n7171 ;
  assign n14668 = x94 & n7174 ;
  assign n14670 = n14669 ^ n14668 ;
  assign n14671 = n14670 ^ x53 ;
  assign n14667 = n2997 & n7175 ;
  assign n14672 = n14671 ^ n14667 ;
  assign n14666 = x93 & n7179 ;
  assign n14673 = n14672 ^ n14666 ;
  assign n14662 = n14405 ^ n14396 ;
  assign n14663 = ~n14397 & n14662 ;
  assign n14664 = n14663 ^ n14405 ;
  assign n14656 = x89 & n7935 ;
  assign n14655 = x91 & n7938 ;
  assign n14657 = n14656 ^ n14655 ;
  assign n14658 = n14657 ^ x56 ;
  assign n14654 = n2542 & n7939 ;
  assign n14659 = n14658 ^ n14654 ;
  assign n14653 = x90 & n7931 ;
  assign n14660 = n14659 ^ n14653 ;
  assign n14625 = ~n1099 & ~n14377 ;
  assign n14640 = n14625 ^ n11874 ;
  assign n14631 = x81 ^ x79 ;
  assign n14629 = n14377 ^ x80 ;
  assign n14641 = n14631 ^ n14629 ;
  assign n14642 = n14641 ^ n14631 ;
  assign n14645 = n1009 & ~n14642 ;
  assign n14646 = n14645 ^ n14631 ;
  assign n14647 = n14640 & n14646 ;
  assign n14630 = n14377 ^ x62 ;
  assign n14648 = n14647 ^ n14630 ;
  assign n14632 = n14631 ^ n14630 ;
  assign n14633 = n14632 ^ n14630 ;
  assign n14634 = n14630 ^ x62 ;
  assign n14635 = ~x81 & ~n14634 ;
  assign n14636 = n14635 ^ n14630 ;
  assign n14637 = ~n14633 & ~n14636 ;
  assign n14638 = n14637 ^ n14630 ;
  assign n14639 = n14629 & ~n14638 ;
  assign n14649 = n14648 ^ n14639 ;
  assign n14623 = n14377 ^ x81 ;
  assign n14624 = n14377 ^ n1099 ;
  assign n14626 = n14625 ^ n14624 ;
  assign n14609 = ~x63 & n1099 ;
  assign n14627 = n14626 ^ n14609 ;
  assign n14628 = ~n14623 & ~n14627 ;
  assign n14650 = n14649 ^ n14628 ;
  assign n14616 = x83 & n9632 ;
  assign n14615 = x85 & n9635 ;
  assign n14617 = n14616 ^ n14615 ;
  assign n14618 = n14617 ^ x62 ;
  assign n14614 = n1743 & n9636 ;
  assign n14619 = n14618 ^ n14614 ;
  assign n14613 = x84 & n9628 ;
  assign n14620 = n14619 ^ n14613 ;
  assign n14612 = n1190 ^ x17 ;
  assign n14621 = n14620 ^ n14612 ;
  assign n14608 = n1190 ^ n1099 ;
  assign n14610 = n14609 ^ n14608 ;
  assign n14611 = ~n9948 & n14610 ;
  assign n14622 = n14621 ^ n14611 ;
  assign n14651 = n14650 ^ n14622 ;
  assign n14606 = x87 & n8737 ;
  assign n14604 = n2119 & n8745 ;
  assign n14602 = x86 & n8741 ;
  assign n14598 = n14390 ^ n14368 ;
  assign n14599 = n14392 & ~n14598 ;
  assign n14600 = n14599 ^ n14390 ;
  assign n14596 = x88 & n8744 ;
  assign n14597 = n14596 ^ x59 ;
  assign n14601 = n14600 ^ n14597 ;
  assign n14603 = n14602 ^ n14601 ;
  assign n14605 = n14604 ^ n14603 ;
  assign n14607 = n14606 ^ n14605 ;
  assign n14652 = n14651 ^ n14607 ;
  assign n14661 = n14660 ^ n14652 ;
  assign n14665 = n14664 ^ n14661 ;
  assign n14674 = n14673 ^ n14665 ;
  assign n14593 = n14418 ^ n14406 ;
  assign n14594 = n14415 & n14593 ;
  assign n14595 = n14594 ^ n14406 ;
  assign n14675 = n14674 ^ n14595 ;
  assign n14684 = n14683 ^ n14675 ;
  assign n14590 = n14431 ^ n14419 ;
  assign n14591 = n14428 & n14590 ;
  assign n14592 = n14591 ^ n14419 ;
  assign n14685 = n14684 ^ n14592 ;
  assign n14694 = n14693 ^ n14685 ;
  assign n14698 = n14697 ^ n14694 ;
  assign n14707 = n14706 ^ n14698 ;
  assign n14711 = n14710 ^ n14707 ;
  assign n14720 = n14719 ^ n14711 ;
  assign n14587 = n14455 ^ n14446 ;
  assign n14588 = n14447 & ~n14587 ;
  assign n14589 = n14588 ^ n14455 ;
  assign n14721 = n14720 ^ n14589 ;
  assign n14730 = n14729 ^ n14721 ;
  assign n14734 = n14733 ^ n14730 ;
  assign n14741 = n14740 ^ n14734 ;
  assign n14743 = n14742 ^ n14741 ;
  assign n14747 = n14746 ^ n14743 ;
  assign n14756 = n14755 ^ n14747 ;
  assign n14760 = n14759 ^ n14756 ;
  assign n14769 = n14768 ^ n14760 ;
  assign n14773 = n14772 ^ n14769 ;
  assign n14775 = n14773 ^ n14508 ;
  assign n14774 = n14773 ^ n14521 ;
  assign n14776 = n14775 ^ n14774 ;
  assign n14777 = n14513 & n14776 ;
  assign n14778 = n14777 ^ n14775 ;
  assign n14787 = n14786 ^ n14778 ;
  assign n14796 = n14795 ^ n14787 ;
  assign n14584 = n14531 ^ n14342 ;
  assign n14585 = ~n14523 & n14584 ;
  assign n14586 = n14585 ^ n14531 ;
  assign n14797 = n14796 ^ n14586 ;
  assign n14806 = n14805 ^ n14797 ;
  assign n14581 = n14541 ^ n14339 ;
  assign n14582 = ~n14533 & n14581 ;
  assign n14583 = n14582 ^ n14541 ;
  assign n14807 = n14806 ^ n14583 ;
  assign n14811 = n14810 ^ n14807 ;
  assign n14557 = n14312 & n14322 ;
  assign n14558 = n14557 ^ n14554 ;
  assign n14559 = n14107 & n14315 ;
  assign n14560 = n14559 ^ n14331 ;
  assign n14561 = n14558 ^ n14329 ;
  assign n14562 = n14561 ^ n14554 ;
  assign n14563 = n14559 ^ n14554 ;
  assign n14564 = n14563 ^ n14554 ;
  assign n14565 = ~n14562 & ~n14564 ;
  assign n14566 = n14565 ^ n14554 ;
  assign n14567 = n14104 & ~n14566 ;
  assign n14568 = n14560 & ~n14567 ;
  assign n14569 = n14558 & n14568 ;
  assign n14570 = n14330 ^ n14322 ;
  assign n14571 = n14570 ^ n14322 ;
  assign n14572 = n14329 ^ n14322 ;
  assign n14573 = n14572 ^ n14322 ;
  assign n14574 = n14571 & n14573 ;
  assign n14575 = n14574 ^ n14322 ;
  assign n14576 = ~n14569 & n14575 ;
  assign n14578 = ~n14554 & ~n14559 ;
  assign n14579 = n14576 & n14578 ;
  assign n14577 = n14576 ^ n14569 ;
  assign n14580 = n14579 ^ n14577 ;
  assign n14812 = n14811 ^ n14580 ;
  assign n15024 = n14583 & n14810 ;
  assign n15023 = ~n14797 & ~n14805 ;
  assign n15025 = n15024 ^ n15023 ;
  assign n15018 = n1331 & n10139 ;
  assign n15017 = x126 & n1327 ;
  assign n15019 = n15018 ^ n15017 ;
  assign n15020 = n15019 ^ x20 ;
  assign n15016 = x127 & n1335 ;
  assign n15021 = n15020 ^ n15016 ;
  assign n15009 = x123 & n1658 ;
  assign n15008 = x125 & n1661 ;
  assign n15010 = n15009 ^ n15008 ;
  assign n15011 = n15010 ^ x23 ;
  assign n15007 = n1662 & n10400 ;
  assign n15012 = n15011 ^ n15007 ;
  assign n15006 = x124 & n1666 ;
  assign n15013 = n15012 ^ n15006 ;
  assign n14995 = x120 & n2018 ;
  assign n14994 = x122 & n2021 ;
  assign n14996 = n14995 ^ n14994 ;
  assign n14997 = n14996 ^ x26 ;
  assign n14993 = n2022 & ~n9247 ;
  assign n14998 = n14997 ^ n14993 ;
  assign n14992 = x121 & n2014 ;
  assign n14999 = n14998 ^ n14992 ;
  assign n14984 = x117 & n2581 ;
  assign n14983 = x119 & n2422 ;
  assign n14985 = n14984 ^ n14983 ;
  assign n14986 = n14985 ^ x29 ;
  assign n14982 = n2423 & n8394 ;
  assign n14987 = n14986 ^ n14982 ;
  assign n14981 = x118 & n2429 ;
  assign n14988 = n14987 ^ n14981 ;
  assign n14975 = x114 & n2879 ;
  assign n14974 = x116 & n2882 ;
  assign n14976 = n14975 ^ n14974 ;
  assign n14977 = n14976 ^ x32 ;
  assign n14973 = n2883 & ~n7588 ;
  assign n14978 = n14977 ^ n14973 ;
  assign n14972 = x115 & n2887 ;
  assign n14979 = n14978 ^ n14972 ;
  assign n14965 = x111 & n3375 ;
  assign n14964 = x113 & n3378 ;
  assign n14966 = n14965 ^ n14964 ;
  assign n14967 = n14966 ^ x35 ;
  assign n14963 = n3379 & ~n6839 ;
  assign n14968 = n14967 ^ n14963 ;
  assign n14962 = x112 & n3383 ;
  assign n14969 = n14968 ^ n14962 ;
  assign n14951 = x108 & n3916 ;
  assign n14950 = x110 & n3919 ;
  assign n14952 = n14951 ^ n14950 ;
  assign n14953 = n14952 ^ x38 ;
  assign n14949 = n3920 & n6129 ;
  assign n14954 = n14953 ^ n14949 ;
  assign n14948 = x109 & n3924 ;
  assign n14955 = n14954 ^ n14948 ;
  assign n14937 = x105 & n4474 ;
  assign n14936 = x107 & n4471 ;
  assign n14938 = n14937 ^ n14936 ;
  assign n14939 = n14938 ^ x41 ;
  assign n14935 = n4472 & ~n5448 ;
  assign n14940 = n14939 ^ n14935 ;
  assign n14934 = x106 & n4467 ;
  assign n14941 = n14940 ^ n14934 ;
  assign n14927 = x102 & n5094 ;
  assign n14926 = x104 & n5097 ;
  assign n14928 = n14927 ^ n14926 ;
  assign n14929 = n14928 ^ x44 ;
  assign n14925 = ~n4814 & n5098 ;
  assign n14930 = n14929 ^ n14925 ;
  assign n14924 = x103 & n5102 ;
  assign n14931 = n14930 ^ n14924 ;
  assign n14913 = x99 & n5965 ;
  assign n14912 = x101 & n5729 ;
  assign n14914 = n14913 ^ n14912 ;
  assign n14915 = n14914 ^ x47 ;
  assign n14911 = n4215 & n5730 ;
  assign n14916 = n14915 ^ n14911 ;
  assign n14910 = x100 & n5736 ;
  assign n14917 = n14916 ^ n14910 ;
  assign n14906 = n14683 ^ n14592 ;
  assign n14907 = n14684 & n14906 ;
  assign n14908 = n14907 ^ n14683 ;
  assign n14900 = x96 & n6677 ;
  assign n14899 = x98 & n6428 ;
  assign n14901 = n14900 ^ n14899 ;
  assign n14902 = n14901 ^ x50 ;
  assign n14898 = n3660 & n6429 ;
  assign n14903 = n14902 ^ n14898 ;
  assign n14897 = x97 & n6433 ;
  assign n14904 = n14903 ^ n14897 ;
  assign n14893 = n14673 ^ n14595 ;
  assign n14894 = n14674 & n14893 ;
  assign n14895 = n14894 ^ n14673 ;
  assign n14887 = x93 & n7171 ;
  assign n14886 = x95 & n7174 ;
  assign n14888 = n14887 ^ n14886 ;
  assign n14889 = n14888 ^ x53 ;
  assign n14885 = n3159 & n7175 ;
  assign n14890 = n14889 ^ n14885 ;
  assign n14884 = x94 & n7179 ;
  assign n14891 = n14890 ^ n14884 ;
  assign n14875 = x87 & n8741 ;
  assign n14874 = x89 & n8744 ;
  assign n14876 = n14875 ^ n14874 ;
  assign n14877 = n14876 ^ x59 ;
  assign n14873 = n2249 & n8745 ;
  assign n14878 = n14877 ^ n14873 ;
  assign n14872 = x88 & n8737 ;
  assign n14879 = n14878 ^ n14872 ;
  assign n14866 = x84 & n9632 ;
  assign n14865 = x86 & n9635 ;
  assign n14867 = n14866 ^ n14865 ;
  assign n14868 = n14867 ^ x62 ;
  assign n14864 = n1857 & n9636 ;
  assign n14869 = n14868 ^ n14864 ;
  assign n14863 = x85 & n9628 ;
  assign n14870 = n14869 ^ n14863 ;
  assign n14854 = x81 ^ x17 ;
  assign n14857 = ~n11875 & n14608 ;
  assign n14858 = n14857 ^ n1099 ;
  assign n14859 = ~n14854 & ~n14858 ;
  assign n14860 = n14859 ^ x17 ;
  assign n14861 = n12206 & ~n14860 ;
  assign n14852 = x82 & n11875 ;
  assign n14851 = x83 & n9948 ;
  assign n14853 = n14852 ^ n14851 ;
  assign n14862 = n14861 ^ n14853 ;
  assign n14871 = n14870 ^ n14862 ;
  assign n14880 = n14879 ^ n14871 ;
  assign n14848 = n14650 ^ n14620 ;
  assign n14849 = n14622 & n14848 ;
  assign n14850 = n14849 ^ n14650 ;
  assign n14881 = n14880 ^ n14850 ;
  assign n14838 = x90 & n7935 ;
  assign n14837 = x92 & n7938 ;
  assign n14839 = n14838 ^ n14837 ;
  assign n14840 = n14839 ^ x56 ;
  assign n14836 = n2684 & n7939 ;
  assign n14841 = n14840 ^ n14836 ;
  assign n14835 = x91 & n7931 ;
  assign n14842 = n14841 ^ n14835 ;
  assign n14844 = n14842 ^ n14651 ;
  assign n14843 = n14842 ^ n14600 ;
  assign n14845 = n14844 ^ n14843 ;
  assign n14846 = n14607 & n14845 ;
  assign n14847 = n14846 ^ n14844 ;
  assign n14882 = n14881 ^ n14847 ;
  assign n14832 = n14664 ^ n14660 ;
  assign n14833 = ~n14661 & n14832 ;
  assign n14834 = n14833 ^ n14664 ;
  assign n14883 = n14882 ^ n14834 ;
  assign n14892 = n14891 ^ n14883 ;
  assign n14896 = n14895 ^ n14892 ;
  assign n14905 = n14904 ^ n14896 ;
  assign n14909 = n14908 ^ n14905 ;
  assign n14918 = n14917 ^ n14909 ;
  assign n14919 = n14918 ^ n14697 ;
  assign n14920 = n14919 ^ n14693 ;
  assign n14921 = n14920 ^ n14918 ;
  assign n14922 = ~n14694 & n14921 ;
  assign n14923 = n14922 ^ n14919 ;
  assign n14932 = n14931 ^ n14923 ;
  assign n14829 = n14710 ^ n14706 ;
  assign n14830 = ~n14707 & n14829 ;
  assign n14831 = n14830 ^ n14710 ;
  assign n14933 = n14932 ^ n14831 ;
  assign n14942 = n14941 ^ n14933 ;
  assign n14943 = n14942 ^ n14719 ;
  assign n14944 = n14943 ^ n14589 ;
  assign n14945 = n14944 ^ n14942 ;
  assign n14946 = n14720 & n14945 ;
  assign n14947 = n14946 ^ n14943 ;
  assign n14956 = n14955 ^ n14947 ;
  assign n14957 = n14956 ^ n14733 ;
  assign n14958 = n14957 ^ n14729 ;
  assign n14959 = n14958 ^ n14956 ;
  assign n14960 = ~n14730 & ~n14959 ;
  assign n14961 = n14960 ^ n14957 ;
  assign n14970 = n14969 ^ n14961 ;
  assign n14826 = n14746 ^ n14734 ;
  assign n14827 = ~n14743 & ~n14826 ;
  assign n14828 = n14827 ^ n14734 ;
  assign n14971 = n14970 ^ n14828 ;
  assign n14980 = n14979 ^ n14971 ;
  assign n14989 = n14988 ^ n14980 ;
  assign n14823 = n14759 ^ n14755 ;
  assign n14824 = n14756 & ~n14823 ;
  assign n14825 = n14824 ^ n14759 ;
  assign n14990 = n14989 ^ n14825 ;
  assign n14820 = n14772 ^ n14768 ;
  assign n14821 = ~n14769 & n14820 ;
  assign n14822 = n14821 ^ n14772 ;
  assign n14991 = n14990 ^ n14822 ;
  assign n15000 = n14999 ^ n14991 ;
  assign n15002 = n15000 ^ n14773 ;
  assign n15001 = n15000 ^ n14786 ;
  assign n15003 = n15002 ^ n15001 ;
  assign n15004 = n14778 & n15003 ;
  assign n15005 = n15004 ^ n15002 ;
  assign n15014 = n15013 ^ n15005 ;
  assign n14817 = n14795 ^ n14586 ;
  assign n14818 = n14796 & n14817 ;
  assign n14819 = n14818 ^ n14795 ;
  assign n15015 = n15014 ^ n14819 ;
  assign n15022 = n15021 ^ n15015 ;
  assign n15026 = n15025 ^ n15022 ;
  assign n14813 = n14806 ^ n14580 ;
  assign n14814 = n14810 ^ n14583 ;
  assign n14815 = n14814 ^ n14580 ;
  assign n14816 = n14813 & ~n14815 ;
  assign n15027 = n15026 ^ n14816 ;
  assign n15249 = x124 & n1658 ;
  assign n15248 = x126 & n1661 ;
  assign n15250 = n15249 ^ n15248 ;
  assign n15251 = n15250 ^ x23 ;
  assign n15247 = n1662 & n10441 ;
  assign n15252 = n15251 ^ n15247 ;
  assign n15246 = x125 & n1666 ;
  assign n15253 = n15252 ^ n15246 ;
  assign n15235 = x121 & n2018 ;
  assign n15234 = x123 & n2021 ;
  assign n15236 = n15235 ^ n15234 ;
  assign n15237 = n15236 ^ x26 ;
  assign n15233 = n2022 & ~n9786 ;
  assign n15238 = n15237 ^ n15233 ;
  assign n15232 = x122 & n2014 ;
  assign n15239 = n15238 ^ n15232 ;
  assign n15228 = n14988 ^ n14825 ;
  assign n15229 = n14989 & ~n15228 ;
  assign n15230 = n15229 ^ n14988 ;
  assign n15222 = x118 & n2581 ;
  assign n15221 = x120 & n2422 ;
  assign n15223 = n15222 ^ n15221 ;
  assign n15224 = n15223 ^ x29 ;
  assign n15220 = n2423 & n8891 ;
  assign n15225 = n15224 ^ n15220 ;
  assign n15219 = x119 & n2429 ;
  assign n15226 = n15225 ^ n15219 ;
  assign n15208 = x115 & n2879 ;
  assign n15207 = x117 & n2882 ;
  assign n15209 = n15208 ^ n15207 ;
  assign n15210 = n15209 ^ x32 ;
  assign n15206 = n2883 & ~n7850 ;
  assign n15211 = n15210 ^ n15206 ;
  assign n15205 = x116 & n2887 ;
  assign n15212 = n15211 ^ n15205 ;
  assign n15194 = x112 & n3375 ;
  assign n15193 = x114 & n3378 ;
  assign n15195 = n15194 ^ n15193 ;
  assign n15196 = n15195 ^ x35 ;
  assign n15192 = n3379 & ~n7092 ;
  assign n15197 = n15196 ^ n15192 ;
  assign n15191 = x113 & n3383 ;
  assign n15198 = n15197 ^ n15191 ;
  assign n15180 = x109 & n3916 ;
  assign n15179 = x111 & n3919 ;
  assign n15181 = n15180 ^ n15179 ;
  assign n15182 = n15181 ^ x38 ;
  assign n15178 = n3920 & ~n6360 ;
  assign n15183 = n15182 ^ n15178 ;
  assign n15177 = x110 & n3924 ;
  assign n15184 = n15183 ^ n15177 ;
  assign n15170 = x106 & n4474 ;
  assign n15169 = x108 & n4471 ;
  assign n15171 = n15170 ^ n15169 ;
  assign n15172 = n15171 ^ x41 ;
  assign n15168 = n4472 & n5670 ;
  assign n15173 = n15172 ^ n15168 ;
  assign n15167 = x107 & n4467 ;
  assign n15174 = n15173 ^ n15167 ;
  assign n15163 = n14931 ^ n14918 ;
  assign n15164 = n14923 & n15163 ;
  assign n15165 = n15164 ^ n14918 ;
  assign n15157 = x103 & n5094 ;
  assign n15156 = x105 & n5097 ;
  assign n15158 = n15157 ^ n15156 ;
  assign n15159 = n15158 ^ x44 ;
  assign n15155 = ~n5023 & n5098 ;
  assign n15160 = n15159 ^ n15155 ;
  assign n15154 = x104 & n5102 ;
  assign n15161 = n15160 ^ n15154 ;
  assign n15143 = x100 & n5965 ;
  assign n15142 = x102 & n5729 ;
  assign n15144 = n15143 ^ n15142 ;
  assign n15145 = n15144 ^ x47 ;
  assign n15141 = n4410 & n5730 ;
  assign n15146 = n15145 ^ n15141 ;
  assign n15140 = x101 & n5736 ;
  assign n15147 = n15146 ^ n15140 ;
  assign n15130 = n14881 ^ n14842 ;
  assign n15131 = ~n14847 & ~n15130 ;
  assign n15132 = n15131 ^ n14842 ;
  assign n15128 = x95 & n7179 ;
  assign n15123 = x94 & n7171 ;
  assign n15122 = x96 & n7174 ;
  assign n15124 = n15123 ^ n15122 ;
  assign n15125 = n15124 ^ x53 ;
  assign n15121 = n3323 & n7175 ;
  assign n15126 = n15125 ^ n15121 ;
  assign n15114 = x88 & n8741 ;
  assign n15113 = x90 & n8744 ;
  assign n15115 = n15114 ^ n15113 ;
  assign n15116 = n15115 ^ x59 ;
  assign n15112 = n2386 & n8745 ;
  assign n15117 = n15116 ^ n15112 ;
  assign n15111 = x89 & n8737 ;
  assign n15118 = n15117 ^ n15111 ;
  assign n15104 = x85 & n9632 ;
  assign n15103 = x87 & n9635 ;
  assign n15105 = n15104 ^ n15103 ;
  assign n15106 = n15105 ^ x62 ;
  assign n15102 = n1982 & n9636 ;
  assign n15107 = n15106 ^ n15102 ;
  assign n15101 = x86 & n9628 ;
  assign n15108 = n15107 ^ n15101 ;
  assign n15097 = ~x84 & n9948 ;
  assign n15098 = n15097 ^ n14852 ;
  assign n15099 = n15098 ^ n9948 ;
  assign n15096 = x83 & n12206 ;
  assign n15100 = n15099 ^ n15096 ;
  assign n15109 = n15108 ^ n15100 ;
  assign n15093 = n14870 ^ n14861 ;
  assign n15094 = n14862 & n15093 ;
  assign n15095 = n15094 ^ n14870 ;
  assign n15110 = n15109 ^ n15095 ;
  assign n15119 = n15118 ^ n15110 ;
  assign n15090 = n14879 ^ n14850 ;
  assign n15091 = ~n14880 & n15090 ;
  assign n15083 = x91 & n7935 ;
  assign n15082 = x93 & n7938 ;
  assign n15084 = n15083 ^ n15082 ;
  assign n15085 = n15084 ^ x56 ;
  assign n15081 = n2836 & n7939 ;
  assign n15086 = n15085 ^ n15081 ;
  assign n15080 = x92 & n7931 ;
  assign n15087 = n15086 ^ n15080 ;
  assign n15088 = n15087 ^ n14879 ;
  assign n15092 = n15091 ^ n15088 ;
  assign n15120 = n15119 ^ n15092 ;
  assign n15127 = n15126 ^ n15120 ;
  assign n15129 = n15128 ^ n15127 ;
  assign n15133 = n15132 ^ n15129 ;
  assign n15077 = n3843 & n6429 ;
  assign n15075 = x97 & n6677 ;
  assign n15071 = n14891 ^ n14834 ;
  assign n15072 = ~n14883 & n15071 ;
  assign n15073 = n15072 ^ n14891 ;
  assign n15069 = x99 & n6428 ;
  assign n15070 = n15069 ^ x50 ;
  assign n15074 = n15073 ^ n15070 ;
  assign n15076 = n15075 ^ n15074 ;
  assign n15078 = n15077 ^ n15076 ;
  assign n15068 = x98 & n6433 ;
  assign n15079 = n15078 ^ n15068 ;
  assign n15134 = n15133 ^ n15079 ;
  assign n15135 = n15134 ^ n14904 ;
  assign n15136 = n15135 ^ n14895 ;
  assign n15137 = n15136 ^ n15134 ;
  assign n15138 = ~n14896 & n15137 ;
  assign n15139 = n15138 ^ n15135 ;
  assign n15148 = n15147 ^ n15139 ;
  assign n15149 = n15148 ^ n14917 ;
  assign n15150 = n15149 ^ n14908 ;
  assign n15151 = n15150 ^ n15148 ;
  assign n15152 = ~n14909 & n15151 ;
  assign n15153 = n15152 ^ n15149 ;
  assign n15162 = n15161 ^ n15153 ;
  assign n15166 = n15165 ^ n15162 ;
  assign n15175 = n15174 ^ n15166 ;
  assign n15065 = n14941 ^ n14831 ;
  assign n15066 = ~n14933 & n15065 ;
  assign n15067 = n15066 ^ n14941 ;
  assign n15176 = n15175 ^ n15067 ;
  assign n15185 = n15184 ^ n15176 ;
  assign n15187 = n15185 ^ n14942 ;
  assign n15186 = n15185 ^ n14955 ;
  assign n15188 = n15187 ^ n15186 ;
  assign n15189 = n14947 & n15188 ;
  assign n15190 = n15189 ^ n15187 ;
  assign n15199 = n15198 ^ n15190 ;
  assign n15201 = n15199 ^ n14956 ;
  assign n15200 = n15199 ^ n14969 ;
  assign n15202 = n15201 ^ n15200 ;
  assign n15203 = ~n14961 & n15202 ;
  assign n15204 = n15203 ^ n15201 ;
  assign n15213 = n15212 ^ n15204 ;
  assign n15214 = n15213 ^ n14979 ;
  assign n15215 = n15214 ^ n15213 ;
  assign n15216 = n15215 ^ n14828 ;
  assign n15217 = ~n14971 & ~n15216 ;
  assign n15218 = n15217 ^ n15214 ;
  assign n15227 = n15226 ^ n15218 ;
  assign n15231 = n15230 ^ n15227 ;
  assign n15240 = n15239 ^ n15231 ;
  assign n15241 = n15240 ^ n14999 ;
  assign n15242 = n15241 ^ n15240 ;
  assign n15243 = n15242 ^ n14822 ;
  assign n15244 = n14991 & n15243 ;
  assign n15245 = n15244 ^ n15241 ;
  assign n15254 = n15253 ^ n15245 ;
  assign n15062 = n15021 ^ n14819 ;
  assign n15063 = n15015 & n15062 ;
  assign n15064 = n15063 ^ n15021 ;
  assign n15255 = n15254 ^ n15064 ;
  assign n15058 = n15013 ^ n15000 ;
  assign n15059 = ~n15005 & ~n15058 ;
  assign n15060 = n15059 ^ n15000 ;
  assign n15048 = x127 & n1326 ;
  assign n15049 = n15048 ^ n1324 ;
  assign n15054 = n1132 & n11265 ;
  assign n15055 = n15054 ^ n15048 ;
  assign n15056 = n15049 & ~n15055 ;
  assign n15057 = n15056 ^ x19 ;
  assign n15061 = n15060 ^ n15057 ;
  assign n15256 = n15255 ^ n15061 ;
  assign n15028 = n15023 ^ n15022 ;
  assign n15029 = n15022 ^ n14806 ;
  assign n15030 = n15029 ^ n15023 ;
  assign n15031 = n15030 ^ n15022 ;
  assign n15032 = n15024 ^ n14814 ;
  assign n15035 = ~n15031 & n15032 ;
  assign n15036 = n15035 ^ n15022 ;
  assign n15037 = n14580 & ~n15036 ;
  assign n15038 = ~n15024 & ~n15037 ;
  assign n15039 = n15028 & n15038 ;
  assign n15040 = n14797 ^ n14580 ;
  assign n15041 = n14806 & n15040 ;
  assign n15042 = n15041 ^ n14797 ;
  assign n15043 = ~n15039 & ~n15042 ;
  assign n15045 = ~n15022 & n15032 ;
  assign n15046 = n15043 & n15045 ;
  assign n15044 = n15043 ^ n15039 ;
  assign n15047 = n15046 ^ n15044 ;
  assign n15257 = n15256 ^ n15047 ;
  assign n15455 = n15057 ^ n15047 ;
  assign n15456 = n15061 & n15455 ;
  assign n15450 = n15253 ^ n15240 ;
  assign n15451 = ~n15245 & ~n15450 ;
  assign n15452 = n15451 ^ n15240 ;
  assign n15444 = x125 & n1658 ;
  assign n15443 = x127 & n1661 ;
  assign n15445 = n15444 ^ n15443 ;
  assign n15446 = n15445 ^ x23 ;
  assign n15442 = n1662 & n10972 ;
  assign n15447 = n15446 ^ n15442 ;
  assign n15441 = x126 & n1666 ;
  assign n15448 = n15447 ^ n15441 ;
  assign n15434 = x122 & n2018 ;
  assign n15433 = x124 & n2021 ;
  assign n15435 = n15434 ^ n15433 ;
  assign n15436 = n15435 ^ x26 ;
  assign n15432 = n2022 & n10095 ;
  assign n15437 = n15436 ^ n15432 ;
  assign n15431 = x123 & n2014 ;
  assign n15438 = n15437 ^ n15431 ;
  assign n15425 = x119 & n2581 ;
  assign n15424 = x121 & n2422 ;
  assign n15426 = n15425 ^ n15424 ;
  assign n15427 = n15426 ^ x29 ;
  assign n15423 = n2423 & n8962 ;
  assign n15428 = n15427 ^ n15423 ;
  assign n15422 = x120 & n2429 ;
  assign n15429 = n15428 ^ n15422 ;
  assign n15418 = n15226 ^ n15213 ;
  assign n15419 = ~n15218 & ~n15418 ;
  assign n15420 = n15419 ^ n15213 ;
  assign n15414 = n15212 ^ n15199 ;
  assign n15415 = ~n15204 & ~n15414 ;
  assign n15416 = n15415 ^ n15199 ;
  assign n15408 = x116 & n2879 ;
  assign n15407 = x118 & n2882 ;
  assign n15409 = n15408 ^ n15407 ;
  assign n15410 = n15409 ^ x32 ;
  assign n15406 = n2883 & ~n8123 ;
  assign n15411 = n15410 ^ n15406 ;
  assign n15405 = x117 & n2887 ;
  assign n15412 = n15411 ^ n15405 ;
  assign n15401 = n15198 ^ n15185 ;
  assign n15402 = ~n15190 & ~n15401 ;
  assign n15403 = n15402 ^ n15185 ;
  assign n15395 = x113 & n3375 ;
  assign n15394 = x115 & n3378 ;
  assign n15396 = n15395 ^ n15394 ;
  assign n15397 = n15396 ^ x35 ;
  assign n15393 = n3379 & ~n7343 ;
  assign n15398 = n15397 ^ n15393 ;
  assign n15392 = x114 & n3383 ;
  assign n15399 = n15398 ^ n15392 ;
  assign n15385 = x110 & n3916 ;
  assign n15384 = x112 & n3919 ;
  assign n15386 = n15385 ^ n15384 ;
  assign n15387 = n15386 ^ x38 ;
  assign n15383 = n3920 & ~n6600 ;
  assign n15388 = n15387 ^ n15383 ;
  assign n15382 = x111 & n3924 ;
  assign n15389 = n15388 ^ n15382 ;
  assign n15378 = n15174 ^ n15165 ;
  assign n15379 = n15166 & n15378 ;
  assign n15380 = n15379 ^ n15174 ;
  assign n15376 = x108 & n4467 ;
  assign n15371 = x107 & n4474 ;
  assign n15370 = x109 & n4471 ;
  assign n15372 = n15371 ^ n15370 ;
  assign n15373 = n15372 ^ x41 ;
  assign n15369 = n4472 & n5902 ;
  assign n15374 = n15373 ^ n15369 ;
  assign n15365 = n15161 ^ n15148 ;
  assign n15366 = ~n15153 & ~n15365 ;
  assign n15367 = n15366 ^ n15148 ;
  assign n15359 = x104 & n5094 ;
  assign n15358 = x106 & n5097 ;
  assign n15360 = n15359 ^ n15358 ;
  assign n15361 = n15360 ^ x44 ;
  assign n15357 = n5098 & ~n5240 ;
  assign n15362 = n15361 ^ n15357 ;
  assign n15356 = x105 & n5102 ;
  assign n15363 = n15362 ^ n15356 ;
  assign n15350 = x101 & n5965 ;
  assign n15349 = x103 & n5729 ;
  assign n15351 = n15350 ^ n15349 ;
  assign n15352 = n15351 ^ x47 ;
  assign n15348 = ~n4615 & n5730 ;
  assign n15353 = n15352 ^ n15348 ;
  assign n15347 = x102 & n5736 ;
  assign n15354 = n15353 ^ n15347 ;
  assign n15334 = x95 & n7171 ;
  assign n15333 = x97 & n7174 ;
  assign n15335 = n15334 ^ n15333 ;
  assign n15336 = n15335 ^ x53 ;
  assign n15332 = n3494 & n7175 ;
  assign n15337 = n15336 ^ n15332 ;
  assign n15331 = x96 & n7179 ;
  assign n15338 = n15337 ^ n15331 ;
  assign n15324 = x92 & n7935 ;
  assign n15323 = x94 & n7938 ;
  assign n15325 = n15324 ^ n15323 ;
  assign n15326 = n15325 ^ x56 ;
  assign n15322 = n2997 & n7939 ;
  assign n15327 = n15326 ^ n15322 ;
  assign n15321 = x93 & n7931 ;
  assign n15328 = n15327 ^ n15321 ;
  assign n15316 = ~n15100 & n15108 ;
  assign n15315 = x83 & n15098 ;
  assign n15317 = n15316 ^ n15315 ;
  assign n15318 = n15317 ^ n14852 ;
  assign n15308 = x86 & n9632 ;
  assign n15307 = x88 & n9635 ;
  assign n15309 = n15308 ^ n15307 ;
  assign n15310 = n15309 ^ x62 ;
  assign n15306 = n2119 & n9636 ;
  assign n15311 = n15310 ^ n15306 ;
  assign n15305 = x87 & n9628 ;
  assign n15312 = n15311 ^ n15305 ;
  assign n15313 = n15312 ^ x20 ;
  assign n15299 = x85 & n11875 ;
  assign n15300 = n15299 ^ n14851 ;
  assign n15301 = n15300 ^ n15096 ;
  assign n15302 = n15301 ^ x85 ;
  assign n15303 = n15302 ^ x84 ;
  assign n15304 = n12206 & n15303 ;
  assign n15314 = n15313 ^ n15304 ;
  assign n15319 = n15318 ^ n15314 ;
  assign n15296 = n15118 ^ n15095 ;
  assign n15297 = n15110 & n15296 ;
  assign n15289 = x89 & n8741 ;
  assign n15288 = x91 & n8744 ;
  assign n15290 = n15289 ^ n15288 ;
  assign n15291 = n15290 ^ x59 ;
  assign n15287 = n2542 & n8745 ;
  assign n15292 = n15291 ^ n15287 ;
  assign n15286 = x90 & n8737 ;
  assign n15293 = n15292 ^ n15286 ;
  assign n15294 = n15293 ^ n15118 ;
  assign n15298 = n15297 ^ n15294 ;
  assign n15320 = n15319 ^ n15298 ;
  assign n15329 = n15328 ^ n15320 ;
  assign n15283 = n15119 ^ n15087 ;
  assign n15284 = n15092 & ~n15283 ;
  assign n15285 = n15284 ^ n15087 ;
  assign n15330 = n15329 ^ n15285 ;
  assign n15339 = n15338 ^ n15330 ;
  assign n15280 = n15132 ^ n15120 ;
  assign n15281 = ~n15129 & ~n15280 ;
  assign n15282 = n15281 ^ n15120 ;
  assign n15340 = n15339 ^ n15282 ;
  assign n15270 = x98 & n6677 ;
  assign n15269 = x100 & n6428 ;
  assign n15271 = n15270 ^ n15269 ;
  assign n15272 = n15271 ^ x50 ;
  assign n15268 = n4034 & n6429 ;
  assign n15273 = n15272 ^ n15268 ;
  assign n15267 = x99 & n6433 ;
  assign n15274 = n15273 ^ n15267 ;
  assign n15275 = n15274 ^ n15133 ;
  assign n15276 = n15275 ^ n15073 ;
  assign n15277 = n15276 ^ n15274 ;
  assign n15278 = ~n15079 & ~n15277 ;
  assign n15279 = n15278 ^ n15275 ;
  assign n15341 = n15340 ^ n15279 ;
  assign n15343 = n15341 ^ n15134 ;
  assign n15342 = n15341 ^ n15147 ;
  assign n15344 = n15343 ^ n15342 ;
  assign n15345 = ~n15139 & ~n15344 ;
  assign n15346 = n15345 ^ n15343 ;
  assign n15355 = n15354 ^ n15346 ;
  assign n15364 = n15363 ^ n15355 ;
  assign n15368 = n15367 ^ n15364 ;
  assign n15375 = n15374 ^ n15368 ;
  assign n15377 = n15376 ^ n15375 ;
  assign n15381 = n15380 ^ n15377 ;
  assign n15390 = n15389 ^ n15381 ;
  assign n15264 = n15184 ^ n15067 ;
  assign n15265 = n15176 & n15264 ;
  assign n15266 = n15265 ^ n15184 ;
  assign n15391 = n15390 ^ n15266 ;
  assign n15400 = n15399 ^ n15391 ;
  assign n15404 = n15403 ^ n15400 ;
  assign n15413 = n15412 ^ n15404 ;
  assign n15417 = n15416 ^ n15413 ;
  assign n15421 = n15420 ^ n15417 ;
  assign n15430 = n15429 ^ n15421 ;
  assign n15439 = n15438 ^ n15430 ;
  assign n15261 = n15239 ^ n15230 ;
  assign n15262 = n15231 & n15261 ;
  assign n15263 = n15262 ^ n15239 ;
  assign n15440 = n15439 ^ n15263 ;
  assign n15449 = n15448 ^ n15440 ;
  assign n15453 = n15452 ^ n15449 ;
  assign n15258 = n15064 ^ n15061 ;
  assign n15259 = n15258 ^ n15047 ;
  assign n15260 = n15255 & n15259 ;
  assign n15454 = n15453 ^ n15260 ;
  assign n15457 = n15456 ^ n15454 ;
  assign n15649 = n15254 ^ n15060 ;
  assign n15650 = n15649 ^ n15057 ;
  assign n15651 = n15650 ^ n15064 ;
  assign n15652 = n15651 ^ n15061 ;
  assign n15653 = n15652 ^ n15453 ;
  assign n15654 = n15061 & ~n15653 ;
  assign n15655 = n15651 ^ n15057 ;
  assign n15656 = ~n15654 & ~n15655 ;
  assign n15657 = n15656 ^ n15057 ;
  assign n15658 = n15657 ^ n15654 ;
  assign n15661 = n15657 ^ n15652 ;
  assign n15662 = n15661 ^ n15657 ;
  assign n15663 = n15453 ^ n15064 ;
  assign n15666 = n15662 & n15663 ;
  assign n15667 = ~n15658 & n15666 ;
  assign n15668 = n15667 ^ n15658 ;
  assign n15669 = n15668 ^ n15654 ;
  assign n15670 = n15047 & ~n15669 ;
  assign n15671 = n15453 ^ n15060 ;
  assign n15672 = n15671 ^ n15453 ;
  assign n15673 = n15453 ^ n15057 ;
  assign n15674 = n15673 ^ n15453 ;
  assign n15675 = n15672 & ~n15674 ;
  assign n15676 = n15675 ^ n15453 ;
  assign n15683 = n15674 ^ n15672 ;
  assign n15684 = n15683 ^ n15453 ;
  assign n15677 = n15453 ^ n15254 ;
  assign n15678 = n15677 ^ n15663 ;
  assign n15679 = n15677 ^ n15673 ;
  assign n15680 = n15679 ^ n15671 ;
  assign n15681 = n15680 ^ n15453 ;
  assign n15682 = n15678 & ~n15681 ;
  assign n15685 = n15684 ^ n15682 ;
  assign n15686 = n15676 & ~n15685 ;
  assign n15687 = n15686 ^ n15453 ;
  assign n15690 = ~n15670 & ~n15687 ;
  assign n15643 = n1662 & n10139 ;
  assign n15642 = x126 & n1658 ;
  assign n15644 = n15643 ^ n15642 ;
  assign n15645 = n15644 ^ x23 ;
  assign n15641 = x127 & n1666 ;
  assign n15646 = n15645 ^ n15641 ;
  assign n15634 = x123 & n2018 ;
  assign n15633 = x125 & n2021 ;
  assign n15635 = n15634 ^ n15633 ;
  assign n15636 = n15635 ^ x26 ;
  assign n15632 = n2022 & n10400 ;
  assign n15637 = n15636 ^ n15632 ;
  assign n15631 = x124 & n2014 ;
  assign n15638 = n15637 ^ n15631 ;
  assign n15620 = x120 & n2581 ;
  assign n15619 = x122 & n2422 ;
  assign n15621 = n15620 ^ n15619 ;
  assign n15622 = n15621 ^ x29 ;
  assign n15618 = n2423 & ~n9247 ;
  assign n15623 = n15622 ^ n15618 ;
  assign n15617 = x121 & n2429 ;
  assign n15624 = n15623 ^ n15617 ;
  assign n15610 = x117 & n2879 ;
  assign n15609 = x119 & n2882 ;
  assign n15611 = n15610 ^ n15609 ;
  assign n15612 = n15611 ^ x32 ;
  assign n15608 = n2883 & n8394 ;
  assign n15613 = n15612 ^ n15608 ;
  assign n15607 = x118 & n2887 ;
  assign n15614 = n15613 ^ n15607 ;
  assign n15600 = x114 & n3375 ;
  assign n15599 = x116 & n3378 ;
  assign n15601 = n15600 ^ n15599 ;
  assign n15602 = n15601 ^ x35 ;
  assign n15598 = n3379 & ~n7588 ;
  assign n15603 = n15602 ^ n15598 ;
  assign n15597 = x115 & n3383 ;
  assign n15604 = n15603 ^ n15597 ;
  assign n15590 = x111 & n3916 ;
  assign n15589 = x113 & n3919 ;
  assign n15591 = n15590 ^ n15589 ;
  assign n15592 = n15591 ^ x38 ;
  assign n15588 = n3920 & ~n6839 ;
  assign n15593 = n15592 ^ n15588 ;
  assign n15587 = x112 & n3924 ;
  assign n15594 = n15593 ^ n15587 ;
  assign n15579 = x108 & n4474 ;
  assign n15578 = x110 & n4471 ;
  assign n15580 = n15579 ^ n15578 ;
  assign n15581 = n15580 ^ x41 ;
  assign n15577 = n4472 & n6129 ;
  assign n15582 = n15581 ^ n15577 ;
  assign n15576 = x109 & n4467 ;
  assign n15583 = n15582 ^ n15576 ;
  assign n15570 = x105 & n5094 ;
  assign n15569 = x107 & n5097 ;
  assign n15571 = n15570 ^ n15569 ;
  assign n15572 = n15571 ^ x44 ;
  assign n15568 = n5098 & ~n5448 ;
  assign n15573 = n15572 ^ n15568 ;
  assign n15567 = x106 & n5102 ;
  assign n15574 = n15573 ^ n15567 ;
  assign n15557 = n15338 ^ n15282 ;
  assign n15558 = ~n15339 & ~n15557 ;
  assign n15559 = n15558 ^ n15338 ;
  assign n15551 = x99 & n6677 ;
  assign n15550 = x101 & n6428 ;
  assign n15552 = n15551 ^ n15550 ;
  assign n15553 = n15552 ^ x50 ;
  assign n15549 = n4215 & n6429 ;
  assign n15554 = n15553 ^ n15549 ;
  assign n15548 = x100 & n6433 ;
  assign n15555 = n15554 ^ n15548 ;
  assign n15541 = x96 & n7171 ;
  assign n15540 = x98 & n7174 ;
  assign n15542 = n15541 ^ n15540 ;
  assign n15543 = n15542 ^ x53 ;
  assign n15539 = n3660 & n7175 ;
  assign n15544 = n15543 ^ n15539 ;
  assign n15538 = x97 & n7179 ;
  assign n15545 = n15544 ^ n15538 ;
  assign n15534 = n15319 ^ n15293 ;
  assign n15535 = n15298 & ~n15534 ;
  assign n15536 = n15535 ^ n15293 ;
  assign n15532 = x94 & n7931 ;
  assign n15527 = x93 & n7935 ;
  assign n15526 = x95 & n7938 ;
  assign n15528 = n15527 ^ n15526 ;
  assign n15529 = n15528 ^ x56 ;
  assign n15525 = n3159 & n7939 ;
  assign n15530 = n15529 ^ n15525 ;
  assign n15518 = x90 & n8741 ;
  assign n15517 = x92 & n8744 ;
  assign n15519 = n15518 ^ n15517 ;
  assign n15520 = n15519 ^ x59 ;
  assign n15516 = n2684 & n8745 ;
  assign n15521 = n15520 ^ n15516 ;
  assign n15515 = x91 & n8737 ;
  assign n15522 = n15521 ^ n15515 ;
  assign n15512 = x86 & n9948 ;
  assign n15513 = n15512 ^ n15299 ;
  assign n15509 = n2249 & n9636 ;
  assign n15507 = x87 & n9632 ;
  assign n15500 = x84 ^ x20 ;
  assign n15503 = n15303 & ~n15500 ;
  assign n15504 = n15503 ^ x84 ;
  assign n15505 = n12206 & n15504 ;
  assign n15498 = x89 & n9635 ;
  assign n15499 = n15498 ^ x62 ;
  assign n15506 = n15505 ^ n15499 ;
  assign n15508 = n15507 ^ n15506 ;
  assign n15510 = n15509 ^ n15508 ;
  assign n15497 = x88 & n9628 ;
  assign n15511 = n15510 ^ n15497 ;
  assign n15514 = n15513 ^ n15511 ;
  assign n15523 = n15522 ^ n15514 ;
  assign n15494 = n15318 ^ n15312 ;
  assign n15495 = n15314 & n15494 ;
  assign n15496 = n15495 ^ n15318 ;
  assign n15524 = n15523 ^ n15496 ;
  assign n15531 = n15530 ^ n15524 ;
  assign n15533 = n15532 ^ n15531 ;
  assign n15537 = n15536 ^ n15533 ;
  assign n15546 = n15545 ^ n15537 ;
  assign n15491 = n15328 ^ n15285 ;
  assign n15492 = ~n15329 & n15491 ;
  assign n15493 = n15492 ^ n15328 ;
  assign n15547 = n15546 ^ n15493 ;
  assign n15556 = n15555 ^ n15547 ;
  assign n15560 = n15559 ^ n15556 ;
  assign n15488 = ~n4814 & n5730 ;
  assign n15486 = x102 & n5965 ;
  assign n15482 = n15340 ^ n15274 ;
  assign n15483 = ~n15279 & n15482 ;
  assign n15484 = n15483 ^ n15274 ;
  assign n15480 = x104 & n5729 ;
  assign n15481 = n15480 ^ x47 ;
  assign n15485 = n15484 ^ n15481 ;
  assign n15487 = n15486 ^ n15485 ;
  assign n15489 = n15488 ^ n15487 ;
  assign n15479 = x103 & n5736 ;
  assign n15490 = n15489 ^ n15479 ;
  assign n15561 = n15560 ^ n15490 ;
  assign n15563 = n15561 ^ n15341 ;
  assign n15562 = n15561 ^ n15354 ;
  assign n15564 = n15563 ^ n15562 ;
  assign n15565 = n15346 & ~n15564 ;
  assign n15566 = n15565 ^ n15563 ;
  assign n15575 = n15574 ^ n15566 ;
  assign n15584 = n15583 ^ n15575 ;
  assign n15476 = n15367 ^ n15363 ;
  assign n15477 = ~n15364 & ~n15476 ;
  assign n15478 = n15477 ^ n15367 ;
  assign n15585 = n15584 ^ n15478 ;
  assign n15473 = n15380 ^ n15368 ;
  assign n15474 = ~n15377 & ~n15473 ;
  assign n15475 = n15474 ^ n15368 ;
  assign n15586 = n15585 ^ n15475 ;
  assign n15595 = n15594 ^ n15586 ;
  assign n15470 = n15381 ^ n15266 ;
  assign n15471 = ~n15390 & n15470 ;
  assign n15472 = n15471 ^ n15389 ;
  assign n15596 = n15595 ^ n15472 ;
  assign n15605 = n15604 ^ n15596 ;
  assign n15467 = n15403 ^ n15399 ;
  assign n15468 = n15400 & ~n15467 ;
  assign n15469 = n15468 ^ n15403 ;
  assign n15606 = n15605 ^ n15469 ;
  assign n15615 = n15614 ^ n15606 ;
  assign n15464 = n15416 ^ n15412 ;
  assign n15465 = ~n15413 & ~n15464 ;
  assign n15466 = n15465 ^ n15416 ;
  assign n15616 = n15615 ^ n15466 ;
  assign n15625 = n15624 ^ n15616 ;
  assign n15626 = n15625 ^ n15429 ;
  assign n15627 = n15626 ^ n15420 ;
  assign n15628 = n15627 ^ n15625 ;
  assign n15629 = ~n15421 & ~n15628 ;
  assign n15630 = n15629 ^ n15626 ;
  assign n15639 = n15638 ^ n15630 ;
  assign n15461 = n15438 ^ n15263 ;
  assign n15462 = n15439 & n15461 ;
  assign n15463 = n15462 ^ n15438 ;
  assign n15640 = n15639 ^ n15463 ;
  assign n15647 = n15646 ^ n15640 ;
  assign n15458 = n15452 ^ n15448 ;
  assign n15459 = ~n15449 & ~n15458 ;
  assign n15460 = n15459 ^ n15452 ;
  assign n15648 = n15647 ^ n15460 ;
  assign n15691 = n15690 ^ n15648 ;
  assign n15887 = n15690 ^ n15460 ;
  assign n15888 = n15648 & ~n15887 ;
  assign n15889 = n15888 ^ n15690 ;
  assign n15875 = x127 & n1657 ;
  assign n15876 = n15875 ^ n1655 ;
  assign n15881 = n1437 & n11265 ;
  assign n15882 = n15881 ^ n15875 ;
  assign n15883 = n15876 & ~n15882 ;
  assign n15884 = n15883 ^ x22 ;
  assign n15864 = x124 & n2018 ;
  assign n15863 = x126 & n2021 ;
  assign n15865 = n15864 ^ n15863 ;
  assign n15866 = n15865 ^ x26 ;
  assign n15862 = n2022 & n10441 ;
  assign n15867 = n15866 ^ n15862 ;
  assign n15861 = x125 & n2014 ;
  assign n15868 = n15867 ^ n15861 ;
  assign n15850 = x121 & n2581 ;
  assign n15849 = x123 & n2422 ;
  assign n15851 = n15850 ^ n15849 ;
  assign n15852 = n15851 ^ x29 ;
  assign n15848 = n2423 & ~n9786 ;
  assign n15853 = n15852 ^ n15848 ;
  assign n15847 = x122 & n2429 ;
  assign n15854 = n15853 ^ n15847 ;
  assign n15840 = x118 & n2879 ;
  assign n15839 = x120 & n2882 ;
  assign n15841 = n15840 ^ n15839 ;
  assign n15842 = n15841 ^ x32 ;
  assign n15838 = n2883 & n8891 ;
  assign n15843 = n15842 ^ n15838 ;
  assign n15837 = x119 & n2887 ;
  assign n15844 = n15843 ^ n15837 ;
  assign n15833 = n15604 ^ n15472 ;
  assign n15834 = ~n15596 & n15833 ;
  assign n15835 = n15834 ^ n15604 ;
  assign n15827 = x115 & n3375 ;
  assign n15826 = x117 & n3378 ;
  assign n15828 = n15827 ^ n15826 ;
  assign n15829 = n15828 ^ x35 ;
  assign n15825 = n3379 & ~n7850 ;
  assign n15830 = n15829 ^ n15825 ;
  assign n15824 = x116 & n3383 ;
  assign n15831 = n15830 ^ n15824 ;
  assign n15813 = x112 & n3916 ;
  assign n15812 = x114 & n3919 ;
  assign n15814 = n15813 ^ n15812 ;
  assign n15815 = n15814 ^ x38 ;
  assign n15811 = n3920 & ~n7092 ;
  assign n15816 = n15815 ^ n15811 ;
  assign n15810 = x113 & n3924 ;
  assign n15817 = n15816 ^ n15810 ;
  assign n15806 = n15583 ^ n15478 ;
  assign n15807 = n15584 & ~n15806 ;
  assign n15808 = n15807 ^ n15583 ;
  assign n15800 = x109 & n4474 ;
  assign n15799 = x111 & n4471 ;
  assign n15801 = n15800 ^ n15799 ;
  assign n15802 = n15801 ^ x41 ;
  assign n15798 = n4472 & ~n6360 ;
  assign n15803 = n15802 ^ n15798 ;
  assign n15797 = x110 & n4467 ;
  assign n15804 = n15803 ^ n15797 ;
  assign n15793 = n15574 ^ n15561 ;
  assign n15794 = n15566 & ~n15793 ;
  assign n15795 = n15794 ^ n15561 ;
  assign n15787 = x106 & n5094 ;
  assign n15786 = x108 & n5097 ;
  assign n15788 = n15787 ^ n15786 ;
  assign n15789 = n15788 ^ x44 ;
  assign n15785 = n5098 & n5670 ;
  assign n15790 = n15789 ^ n15785 ;
  assign n15784 = x107 & n5102 ;
  assign n15791 = n15790 ^ n15784 ;
  assign n15772 = x88 & n9632 ;
  assign n15771 = x90 & n9635 ;
  assign n15773 = n15772 ^ n15771 ;
  assign n15774 = n15773 ^ x62 ;
  assign n15770 = n2386 & n9636 ;
  assign n15775 = n15774 ^ n15770 ;
  assign n15769 = x89 & n9628 ;
  assign n15776 = n15775 ^ n15769 ;
  assign n15765 = x63 & n1608 ;
  assign n15766 = n15765 ^ n1724 ;
  assign n15767 = ~n9948 & n15766 ;
  assign n15768 = n15767 ^ n1724 ;
  assign n15777 = n15776 ^ n15768 ;
  assign n15758 = n2836 & n8745 ;
  assign n15756 = x91 & n8741 ;
  assign n15752 = n15513 ^ n15505 ;
  assign n15753 = ~n15511 & ~n15752 ;
  assign n15754 = n15753 ^ n15513 ;
  assign n15750 = x93 & n8744 ;
  assign n15751 = n15750 ^ x59 ;
  assign n15755 = n15754 ^ n15751 ;
  assign n15757 = n15756 ^ n15755 ;
  assign n15759 = n15758 ^ n15757 ;
  assign n15749 = x92 & n8737 ;
  assign n15760 = n15759 ^ n15749 ;
  assign n15778 = n15777 ^ n15760 ;
  assign n15747 = x95 & n7931 ;
  assign n15745 = n3323 & n7939 ;
  assign n15743 = x94 & n7935 ;
  assign n15739 = n15514 ^ n15496 ;
  assign n15740 = ~n15523 & n15739 ;
  assign n15741 = n15740 ^ n15522 ;
  assign n15737 = x96 & n7938 ;
  assign n15738 = n15737 ^ x56 ;
  assign n15742 = n15741 ^ n15738 ;
  assign n15744 = n15743 ^ n15742 ;
  assign n15746 = n15745 ^ n15744 ;
  assign n15748 = n15747 ^ n15746 ;
  assign n15779 = n15778 ^ n15748 ;
  assign n15735 = x98 & n7179 ;
  assign n15733 = n3843 & n7175 ;
  assign n15731 = x97 & n7171 ;
  assign n15727 = n15536 ^ n15524 ;
  assign n15728 = ~n15533 & ~n15727 ;
  assign n15729 = n15728 ^ n15524 ;
  assign n15725 = x99 & n7174 ;
  assign n15726 = n15725 ^ x53 ;
  assign n15730 = n15729 ^ n15726 ;
  assign n15732 = n15731 ^ n15730 ;
  assign n15734 = n15733 ^ n15732 ;
  assign n15736 = n15735 ^ n15734 ;
  assign n15780 = n15779 ^ n15736 ;
  assign n15722 = n4410 & n6429 ;
  assign n15720 = x100 & n6677 ;
  assign n15718 = x102 & n6428 ;
  assign n15714 = n15545 ^ n15493 ;
  assign n15715 = ~n15546 & n15714 ;
  assign n15716 = n15715 ^ n15545 ;
  assign n15717 = n15716 ^ x50 ;
  assign n15719 = n15718 ^ n15717 ;
  assign n15721 = n15720 ^ n15719 ;
  assign n15723 = n15722 ^ n15721 ;
  assign n15713 = x101 & n6433 ;
  assign n15724 = n15723 ^ n15713 ;
  assign n15781 = n15780 ^ n15724 ;
  assign n15710 = ~n5023 & n5730 ;
  assign n15708 = x103 & n5965 ;
  assign n15704 = n15559 ^ n15555 ;
  assign n15705 = n15556 & n15704 ;
  assign n15706 = n15705 ^ n15559 ;
  assign n15702 = x105 & n5729 ;
  assign n15703 = n15702 ^ x47 ;
  assign n15707 = n15706 ^ n15703 ;
  assign n15709 = n15708 ^ n15707 ;
  assign n15711 = n15710 ^ n15709 ;
  assign n15701 = x104 & n5736 ;
  assign n15712 = n15711 ^ n15701 ;
  assign n15782 = n15781 ^ n15712 ;
  assign n15698 = n15560 ^ n15484 ;
  assign n15699 = ~n15490 & ~n15698 ;
  assign n15700 = n15699 ^ n15560 ;
  assign n15783 = n15782 ^ n15700 ;
  assign n15792 = n15791 ^ n15783 ;
  assign n15796 = n15795 ^ n15792 ;
  assign n15805 = n15804 ^ n15796 ;
  assign n15809 = n15808 ^ n15805 ;
  assign n15818 = n15817 ^ n15809 ;
  assign n15819 = n15818 ^ n15594 ;
  assign n15820 = n15819 ^ n15818 ;
  assign n15821 = n15820 ^ n15475 ;
  assign n15822 = ~n15586 & ~n15821 ;
  assign n15823 = n15822 ^ n15819 ;
  assign n15832 = n15831 ^ n15823 ;
  assign n15836 = n15835 ^ n15832 ;
  assign n15845 = n15844 ^ n15836 ;
  assign n15695 = n15614 ^ n15469 ;
  assign n15696 = n15606 & ~n15695 ;
  assign n15697 = n15696 ^ n15614 ;
  assign n15846 = n15845 ^ n15697 ;
  assign n15855 = n15854 ^ n15846 ;
  assign n15856 = n15855 ^ n15624 ;
  assign n15857 = n15856 ^ n15855 ;
  assign n15858 = n15857 ^ n15466 ;
  assign n15859 = ~n15616 & ~n15858 ;
  assign n15860 = n15859 ^ n15856 ;
  assign n15869 = n15868 ^ n15860 ;
  assign n15871 = n15869 ^ n15625 ;
  assign n15870 = n15869 ^ n15638 ;
  assign n15872 = n15871 ^ n15870 ;
  assign n15873 = n15630 & n15872 ;
  assign n15874 = n15873 ^ n15871 ;
  assign n15885 = n15884 ^ n15874 ;
  assign n15692 = n15646 ^ n15463 ;
  assign n15693 = ~n15640 & n15692 ;
  assign n15694 = n15693 ^ n15646 ;
  assign n15886 = n15885 ^ n15694 ;
  assign n15890 = n15889 ^ n15886 ;
  assign n16072 = n15884 ^ n15869 ;
  assign n16073 = ~n15874 & ~n16072 ;
  assign n16074 = n16073 ^ n15869 ;
  assign n16068 = n15868 ^ n15855 ;
  assign n16069 = ~n15860 & ~n16068 ;
  assign n16070 = n16069 ^ n15855 ;
  assign n16062 = x125 & n2018 ;
  assign n16061 = x127 & n2021 ;
  assign n16063 = n16062 ^ n16061 ;
  assign n16064 = n16063 ^ x26 ;
  assign n16060 = n2022 & n10972 ;
  assign n16065 = n16064 ^ n16060 ;
  assign n16059 = x126 & n2014 ;
  assign n16066 = n16065 ^ n16059 ;
  assign n16052 = x122 & n2581 ;
  assign n16051 = x124 & n2422 ;
  assign n16053 = n16052 ^ n16051 ;
  assign n16054 = n16053 ^ x29 ;
  assign n16050 = n2423 & n10095 ;
  assign n16055 = n16054 ^ n16050 ;
  assign n16049 = x123 & n2429 ;
  assign n16056 = n16055 ^ n16049 ;
  assign n16043 = x119 & n2879 ;
  assign n16042 = x121 & n2882 ;
  assign n16044 = n16043 ^ n16042 ;
  assign n16045 = n16044 ^ x32 ;
  assign n16041 = n2883 & n8962 ;
  assign n16046 = n16045 ^ n16041 ;
  assign n16040 = x120 & n2887 ;
  assign n16047 = n16046 ^ n16040 ;
  assign n16031 = n15831 ^ n15818 ;
  assign n16032 = ~n15823 & ~n16031 ;
  assign n16033 = n16032 ^ n15818 ;
  assign n16025 = x116 & n3375 ;
  assign n16024 = x118 & n3378 ;
  assign n16026 = n16025 ^ n16024 ;
  assign n16027 = n16026 ^ x35 ;
  assign n16023 = n3379 & ~n8123 ;
  assign n16028 = n16027 ^ n16023 ;
  assign n16022 = x117 & n3383 ;
  assign n16029 = n16028 ^ n16022 ;
  assign n16015 = x113 & n3916 ;
  assign n16014 = x115 & n3919 ;
  assign n16016 = n16015 ^ n16014 ;
  assign n16017 = n16016 ^ x38 ;
  assign n16013 = n3920 & ~n7343 ;
  assign n16018 = n16017 ^ n16013 ;
  assign n16012 = x114 & n3924 ;
  assign n16019 = n16018 ^ n16012 ;
  assign n16008 = n15804 ^ n15795 ;
  assign n16009 = n15796 & ~n16008 ;
  assign n16010 = n16009 ^ n15804 ;
  assign n16006 = x111 & n4467 ;
  assign n16001 = x110 & n4474 ;
  assign n16000 = x112 & n4471 ;
  assign n16002 = n16001 ^ n16000 ;
  assign n16003 = n16002 ^ x41 ;
  assign n15999 = n4472 & ~n6600 ;
  assign n16004 = n16003 ^ n15999 ;
  assign n15995 = n15791 ^ n15700 ;
  assign n15996 = ~n15783 & ~n15995 ;
  assign n15997 = n15996 ^ n15791 ;
  assign n15993 = x108 & n5102 ;
  assign n15988 = x107 & n5094 ;
  assign n15987 = x109 & n5097 ;
  assign n15989 = n15988 ^ n15987 ;
  assign n15990 = n15989 ^ x44 ;
  assign n15986 = n5098 & n5902 ;
  assign n15991 = n15990 ^ n15986 ;
  assign n15980 = x104 & n5965 ;
  assign n15979 = x106 & n5729 ;
  assign n15981 = n15980 ^ n15979 ;
  assign n15982 = n15981 ^ x47 ;
  assign n15978 = ~n5240 & n5730 ;
  assign n15983 = n15982 ^ n15978 ;
  assign n15977 = x105 & n5736 ;
  assign n15984 = n15983 ^ n15977 ;
  assign n15973 = n15781 ^ n15706 ;
  assign n15974 = ~n15712 & ~n15973 ;
  assign n15975 = n15974 ^ n15781 ;
  assign n15968 = x96 & n7931 ;
  assign n15955 = x89 & n9632 ;
  assign n15954 = x91 & n9635 ;
  assign n15956 = n15955 ^ n15954 ;
  assign n15957 = n15956 ^ x62 ;
  assign n15953 = n2542 & n9636 ;
  assign n15958 = n15957 ^ n15953 ;
  assign n15952 = x90 & n9628 ;
  assign n15959 = n15958 ^ n15952 ;
  assign n15960 = n15959 ^ x23 ;
  assign n15948 = x88 ^ x86 ;
  assign n15949 = ~n11875 & n15948 ;
  assign n15950 = n15949 ^ n1724 ;
  assign n15951 = n12206 & n15950 ;
  assign n15961 = n15960 ^ n15951 ;
  assign n15944 = n15776 ^ n9948 ;
  assign n15945 = n15944 ^ x86 ;
  assign n15946 = n15768 & ~n15945 ;
  assign n15947 = n15946 ^ n15776 ;
  assign n15962 = n15961 ^ n15947 ;
  assign n15934 = x92 & n8741 ;
  assign n15933 = x94 & n8744 ;
  assign n15935 = n15934 ^ n15933 ;
  assign n15936 = n15935 ^ x59 ;
  assign n15932 = n2997 & n8745 ;
  assign n15937 = n15936 ^ n15932 ;
  assign n15931 = x93 & n8737 ;
  assign n15938 = n15937 ^ n15931 ;
  assign n15939 = n15938 ^ n15777 ;
  assign n15940 = n15939 ^ n15754 ;
  assign n15941 = n15940 ^ n15938 ;
  assign n15942 = n15760 & n15941 ;
  assign n15943 = n15942 ^ n15939 ;
  assign n15963 = n15962 ^ n15943 ;
  assign n15964 = n15963 ^ x56 ;
  assign n15930 = x95 & n7935 ;
  assign n15965 = n15964 ^ n15930 ;
  assign n15929 = x97 & n7938 ;
  assign n15966 = n15965 ^ n15929 ;
  assign n15928 = n3494 & n7939 ;
  assign n15967 = n15966 ^ n15928 ;
  assign n15969 = n15968 ^ n15967 ;
  assign n15925 = n15778 ^ n15741 ;
  assign n15926 = ~n15748 & n15925 ;
  assign n15927 = n15926 ^ n15778 ;
  assign n15970 = n15969 ^ n15927 ;
  assign n15915 = x98 & n7171 ;
  assign n15914 = x100 & n7174 ;
  assign n15916 = n15915 ^ n15914 ;
  assign n15917 = n15916 ^ x53 ;
  assign n15913 = n4034 & n7175 ;
  assign n15918 = n15917 ^ n15913 ;
  assign n15912 = x99 & n7179 ;
  assign n15919 = n15918 ^ n15912 ;
  assign n15921 = n15919 ^ n15779 ;
  assign n15920 = n15919 ^ n15729 ;
  assign n15922 = n15921 ^ n15920 ;
  assign n15923 = n15736 & ~n15922 ;
  assign n15924 = n15923 ^ n15921 ;
  assign n15971 = n15970 ^ n15924 ;
  assign n15909 = ~n4615 & n6429 ;
  assign n15907 = x101 & n6677 ;
  assign n15903 = n15780 ^ n15716 ;
  assign n15904 = ~n15724 & ~n15903 ;
  assign n15905 = n15904 ^ n15780 ;
  assign n15901 = x103 & n6428 ;
  assign n15902 = n15901 ^ x50 ;
  assign n15906 = n15905 ^ n15902 ;
  assign n15908 = n15907 ^ n15906 ;
  assign n15910 = n15909 ^ n15908 ;
  assign n15900 = x102 & n6433 ;
  assign n15911 = n15910 ^ n15900 ;
  assign n15972 = n15971 ^ n15911 ;
  assign n15976 = n15975 ^ n15972 ;
  assign n15985 = n15984 ^ n15976 ;
  assign n15992 = n15991 ^ n15985 ;
  assign n15994 = n15993 ^ n15992 ;
  assign n15998 = n15997 ^ n15994 ;
  assign n16005 = n16004 ^ n15998 ;
  assign n16007 = n16006 ^ n16005 ;
  assign n16011 = n16010 ^ n16007 ;
  assign n16020 = n16019 ^ n16011 ;
  assign n15897 = n15817 ^ n15808 ;
  assign n15898 = n15809 & n15897 ;
  assign n15899 = n15898 ^ n15817 ;
  assign n16021 = n16020 ^ n15899 ;
  assign n16030 = n16029 ^ n16021 ;
  assign n16034 = n16033 ^ n16030 ;
  assign n16035 = n16034 ^ n15844 ;
  assign n16036 = n16035 ^ n15835 ;
  assign n16037 = n16036 ^ n16034 ;
  assign n16038 = n15836 & n16037 ;
  assign n16039 = n16038 ^ n16035 ;
  assign n16048 = n16047 ^ n16039 ;
  assign n16057 = n16056 ^ n16048 ;
  assign n15894 = n15854 ^ n15697 ;
  assign n15895 = n15846 & n15894 ;
  assign n15896 = n15895 ^ n15854 ;
  assign n16058 = n16057 ^ n15896 ;
  assign n16067 = n16066 ^ n16058 ;
  assign n16071 = n16070 ^ n16067 ;
  assign n16075 = n16074 ^ n16071 ;
  assign n15891 = n15889 ^ n15694 ;
  assign n15892 = n15886 & n15891 ;
  assign n15893 = n15892 ^ n15889 ;
  assign n16076 = n16075 ^ n15893 ;
  assign n16260 = ~n16058 & n16071 ;
  assign n16256 = n16066 & ~n16070 ;
  assign n16255 = n16070 ^ n16066 ;
  assign n16257 = n16256 ^ n16255 ;
  assign n16250 = n2022 & n10139 ;
  assign n16249 = x126 & n2018 ;
  assign n16251 = n16250 ^ n16249 ;
  assign n16252 = n16251 ^ x26 ;
  assign n16248 = x127 & n2014 ;
  assign n16253 = n16252 ^ n16248 ;
  assign n16241 = x123 & n2581 ;
  assign n16240 = x125 & n2422 ;
  assign n16242 = n16241 ^ n16240 ;
  assign n16243 = n16242 ^ x29 ;
  assign n16239 = n2423 & n10400 ;
  assign n16244 = n16243 ^ n16239 ;
  assign n16238 = x124 & n2429 ;
  assign n16245 = n16244 ^ n16238 ;
  assign n16227 = x120 & n2879 ;
  assign n16226 = x122 & n2882 ;
  assign n16228 = n16227 ^ n16226 ;
  assign n16229 = n16228 ^ x32 ;
  assign n16225 = n2883 & ~n9247 ;
  assign n16230 = n16229 ^ n16225 ;
  assign n16224 = x121 & n2887 ;
  assign n16231 = n16230 ^ n16224 ;
  assign n16216 = x114 & n3916 ;
  assign n16215 = x116 & n3919 ;
  assign n16217 = n16216 ^ n16215 ;
  assign n16218 = n16217 ^ x38 ;
  assign n16214 = n3920 & ~n7588 ;
  assign n16219 = n16218 ^ n16214 ;
  assign n16213 = x115 & n3924 ;
  assign n16220 = n16219 ^ n16213 ;
  assign n16206 = x111 & n4474 ;
  assign n16205 = x113 & n4471 ;
  assign n16207 = n16206 ^ n16205 ;
  assign n16208 = n16207 ^ x41 ;
  assign n16204 = n4472 & ~n6839 ;
  assign n16209 = n16208 ^ n16204 ;
  assign n16203 = x112 & n4467 ;
  assign n16210 = n16209 ^ n16203 ;
  assign n16195 = x108 & n5094 ;
  assign n16194 = x110 & n5097 ;
  assign n16196 = n16195 ^ n16194 ;
  assign n16197 = n16196 ^ x44 ;
  assign n16193 = n5098 & n6129 ;
  assign n16198 = n16197 ^ n16193 ;
  assign n16192 = x109 & n5102 ;
  assign n16199 = n16198 ^ n16192 ;
  assign n16186 = x105 & n5965 ;
  assign n16185 = x107 & n5729 ;
  assign n16187 = n16186 ^ n16185 ;
  assign n16188 = n16187 ^ x47 ;
  assign n16184 = ~n5448 & n5730 ;
  assign n16189 = n16188 ^ n16184 ;
  assign n16183 = x106 & n5736 ;
  assign n16190 = n16189 ^ n16183 ;
  assign n16173 = x97 & n7931 ;
  assign n16171 = n3660 & n7939 ;
  assign n16167 = x96 & n7935 ;
  assign n16166 = x98 & n7938 ;
  assign n16168 = n16167 ^ n16166 ;
  assign n16169 = n16168 ^ x56 ;
  assign n16163 = x94 & n8737 ;
  assign n16161 = n3159 & n8745 ;
  assign n16157 = x93 & n8741 ;
  assign n16156 = x95 & n8744 ;
  assign n16158 = n16157 ^ n16156 ;
  assign n16159 = n16158 ^ x59 ;
  assign n16150 = x90 & n9632 ;
  assign n16149 = x92 & n9635 ;
  assign n16151 = n16150 ^ n16149 ;
  assign n16152 = n16151 ^ x62 ;
  assign n16148 = n2684 & n9636 ;
  assign n16153 = n16152 ^ n16148 ;
  assign n16147 = x91 & n9628 ;
  assign n16154 = n16153 ^ n16147 ;
  assign n16144 = x88 & n11875 ;
  assign n16138 = x87 ^ x23 ;
  assign n16141 = n15950 & ~n16138 ;
  assign n16142 = n16141 ^ x87 ;
  assign n16143 = n12206 & n16142 ;
  assign n16145 = n16144 ^ n16143 ;
  assign n16137 = x89 & n9948 ;
  assign n16146 = n16145 ^ n16137 ;
  assign n16155 = n16154 ^ n16146 ;
  assign n16160 = n16159 ^ n16155 ;
  assign n16162 = n16161 ^ n16160 ;
  assign n16164 = n16163 ^ n16162 ;
  assign n16134 = n15959 ^ n15947 ;
  assign n16135 = ~n15961 & n16134 ;
  assign n16136 = n16135 ^ n15959 ;
  assign n16165 = n16164 ^ n16136 ;
  assign n16170 = n16169 ^ n16165 ;
  assign n16172 = n16171 ^ n16170 ;
  assign n16174 = n16173 ^ n16172 ;
  assign n16131 = n15962 ^ n15938 ;
  assign n16132 = ~n15943 & ~n16131 ;
  assign n16133 = n16132 ^ n15938 ;
  assign n16175 = n16174 ^ n16133 ;
  assign n16128 = n4215 & n7175 ;
  assign n16126 = x99 & n7171 ;
  assign n16122 = n15963 ^ n15927 ;
  assign n16123 = n15969 & n16122 ;
  assign n16124 = n16123 ^ n15963 ;
  assign n16120 = x101 & n7174 ;
  assign n16121 = n16120 ^ x53 ;
  assign n16125 = n16124 ^ n16121 ;
  assign n16127 = n16126 ^ n16125 ;
  assign n16129 = n16128 ^ n16127 ;
  assign n16119 = x100 & n7179 ;
  assign n16130 = n16129 ^ n16119 ;
  assign n16176 = n16175 ^ n16130 ;
  assign n16116 = ~n4814 & n6429 ;
  assign n16114 = x102 & n6677 ;
  assign n16110 = n15970 ^ n15919 ;
  assign n16111 = n15924 & n16110 ;
  assign n16112 = n16111 ^ n15919 ;
  assign n16108 = x104 & n6428 ;
  assign n16109 = n16108 ^ x50 ;
  assign n16113 = n16112 ^ n16109 ;
  assign n16115 = n16114 ^ n16113 ;
  assign n16117 = n16116 ^ n16115 ;
  assign n16107 = x103 & n6433 ;
  assign n16118 = n16117 ^ n16107 ;
  assign n16177 = n16176 ^ n16118 ;
  assign n16178 = n16177 ^ n15971 ;
  assign n16179 = n16178 ^ n15905 ;
  assign n16180 = n16179 ^ n16177 ;
  assign n16181 = n15911 & ~n16180 ;
  assign n16182 = n16181 ^ n16178 ;
  assign n16191 = n16190 ^ n16182 ;
  assign n16200 = n16199 ^ n16191 ;
  assign n16104 = n15984 ^ n15975 ;
  assign n16105 = ~n15976 & ~n16104 ;
  assign n16106 = n16105 ^ n15984 ;
  assign n16201 = n16200 ^ n16106 ;
  assign n16101 = n15997 ^ n15985 ;
  assign n16102 = n15994 & n16101 ;
  assign n16103 = n16102 ^ n15985 ;
  assign n16202 = n16201 ^ n16103 ;
  assign n16211 = n16210 ^ n16202 ;
  assign n16098 = n16010 ^ n15998 ;
  assign n16099 = n16007 & n16098 ;
  assign n16100 = n16099 ^ n15998 ;
  assign n16212 = n16211 ^ n16100 ;
  assign n16221 = n16220 ^ n16212 ;
  assign n16088 = x117 & n3375 ;
  assign n16087 = x119 & n3378 ;
  assign n16089 = n16088 ^ n16087 ;
  assign n16090 = n16089 ^ x35 ;
  assign n16086 = n3379 & n8394 ;
  assign n16091 = n16090 ^ n16086 ;
  assign n16085 = x118 & n3383 ;
  assign n16092 = n16091 ^ n16085 ;
  assign n16093 = n16092 ^ n16019 ;
  assign n16094 = n16093 ^ n15899 ;
  assign n16095 = n16094 ^ n16092 ;
  assign n16096 = n16020 & n16095 ;
  assign n16097 = n16096 ^ n16093 ;
  assign n16222 = n16221 ^ n16097 ;
  assign n16082 = n16033 ^ n16029 ;
  assign n16083 = ~n16030 & ~n16082 ;
  assign n16084 = n16083 ^ n16033 ;
  assign n16223 = n16222 ^ n16084 ;
  assign n16232 = n16231 ^ n16223 ;
  assign n16234 = n16232 ^ n16034 ;
  assign n16233 = n16232 ^ n16047 ;
  assign n16235 = n16234 ^ n16233 ;
  assign n16236 = ~n16039 & ~n16235 ;
  assign n16237 = n16236 ^ n16234 ;
  assign n16246 = n16245 ^ n16237 ;
  assign n16079 = n16056 ^ n15896 ;
  assign n16080 = ~n16057 & n16079 ;
  assign n16081 = n16080 ^ n16056 ;
  assign n16247 = n16246 ^ n16081 ;
  assign n16254 = n16253 ^ n16247 ;
  assign n16258 = n16257 ^ n16254 ;
  assign n16077 = n16074 ^ n15893 ;
  assign n16078 = ~n16075 & n16077 ;
  assign n16259 = n16258 ^ n16078 ;
  assign n16261 = n16260 ^ n16259 ;
  assign n16436 = n16058 & n16074 ;
  assign n16435 = n16074 ^ n16058 ;
  assign n16437 = n16436 ^ n16435 ;
  assign n16438 = n16437 ^ n16254 ;
  assign n16439 = n15893 & ~n16257 ;
  assign n16440 = n16438 & n16439 ;
  assign n16441 = ~n16254 & ~n16440 ;
  assign n16442 = n16436 ^ n16070 ;
  assign n16443 = ~n16255 & n16442 ;
  assign n16444 = n16443 ^ n16070 ;
  assign n16445 = n16441 & ~n16444 ;
  assign n16446 = n16445 ^ n16440 ;
  assign n16447 = n16256 ^ n16254 ;
  assign n16448 = n16058 ^ n15893 ;
  assign n16449 = n16435 & ~n16448 ;
  assign n16450 = n16449 ^ n16058 ;
  assign n16451 = ~n16447 & ~n16450 ;
  assign n16452 = ~n16446 & ~n16451 ;
  assign n16430 = n16245 ^ n16232 ;
  assign n16431 = ~n16237 & n16430 ;
  assign n16432 = n16431 ^ n16232 ;
  assign n16423 = x124 & n2581 ;
  assign n16422 = x126 & n2422 ;
  assign n16424 = n16423 ^ n16422 ;
  assign n16425 = n16424 ^ x29 ;
  assign n16421 = n2423 & n10441 ;
  assign n16426 = n16425 ^ n16421 ;
  assign n16420 = x125 & n2429 ;
  assign n16427 = n16426 ^ n16420 ;
  assign n16413 = x121 & n2879 ;
  assign n16412 = x123 & n2882 ;
  assign n16414 = n16413 ^ n16412 ;
  assign n16415 = n16414 ^ x32 ;
  assign n16411 = n2883 & ~n9786 ;
  assign n16416 = n16415 ^ n16411 ;
  assign n16410 = x122 & n2887 ;
  assign n16417 = n16416 ^ n16410 ;
  assign n16403 = x118 & n3375 ;
  assign n16402 = x120 & n3378 ;
  assign n16404 = n16403 ^ n16402 ;
  assign n16405 = n16404 ^ x35 ;
  assign n16401 = n3379 & n8891 ;
  assign n16406 = n16405 ^ n16401 ;
  assign n16400 = x119 & n3383 ;
  assign n16407 = n16406 ^ n16400 ;
  assign n16396 = n16220 ^ n16100 ;
  assign n16397 = n16212 & n16396 ;
  assign n16398 = n16397 ^ n16220 ;
  assign n16390 = x115 & n3916 ;
  assign n16389 = x117 & n3919 ;
  assign n16391 = n16390 ^ n16389 ;
  assign n16392 = n16391 ^ x38 ;
  assign n16388 = n3920 & ~n7850 ;
  assign n16393 = n16392 ^ n16388 ;
  assign n16387 = x116 & n3924 ;
  assign n16394 = n16393 ^ n16387 ;
  assign n16376 = x112 & n4474 ;
  assign n16375 = x114 & n4471 ;
  assign n16377 = n16376 ^ n16375 ;
  assign n16378 = n16377 ^ x41 ;
  assign n16374 = n4472 & ~n7092 ;
  assign n16379 = n16378 ^ n16374 ;
  assign n16373 = x113 & n4467 ;
  assign n16380 = n16379 ^ n16373 ;
  assign n16370 = n16199 ^ n16106 ;
  assign n16371 = ~n16200 & n16370 ;
  assign n16362 = x109 & n5094 ;
  assign n16361 = x111 & n5097 ;
  assign n16363 = n16362 ^ n16361 ;
  assign n16364 = n16363 ^ x44 ;
  assign n16360 = n5098 & ~n6360 ;
  assign n16365 = n16364 ^ n16360 ;
  assign n16359 = x110 & n5102 ;
  assign n16366 = n16365 ^ n16359 ;
  assign n16355 = n16190 ^ n16177 ;
  assign n16356 = ~n16182 & ~n16355 ;
  assign n16357 = n16356 ^ n16177 ;
  assign n16348 = x106 & n5965 ;
  assign n16347 = x108 & n5729 ;
  assign n16349 = n16348 ^ n16347 ;
  assign n16350 = n16349 ^ x47 ;
  assign n16346 = n5670 & n5730 ;
  assign n16351 = n16350 ^ n16346 ;
  assign n16345 = x107 & n5736 ;
  assign n16352 = n16351 ^ n16345 ;
  assign n16339 = x103 & n6677 ;
  assign n16338 = x105 & n6428 ;
  assign n16340 = n16339 ^ n16338 ;
  assign n16341 = n16340 ^ x50 ;
  assign n16337 = ~n5023 & n6429 ;
  assign n16342 = n16341 ^ n16337 ;
  assign n16336 = x104 & n6433 ;
  assign n16343 = n16342 ^ n16336 ;
  assign n16333 = n16175 ^ n16124 ;
  assign n16334 = ~n16130 & ~n16333 ;
  assign n16324 = x100 & n7171 ;
  assign n16323 = x102 & n7174 ;
  assign n16325 = n16324 ^ n16323 ;
  assign n16326 = n16325 ^ x53 ;
  assign n16322 = n4410 & n7175 ;
  assign n16327 = n16326 ^ n16322 ;
  assign n16321 = x101 & n7179 ;
  assign n16328 = n16327 ^ n16321 ;
  assign n16317 = n16155 ^ n16136 ;
  assign n16318 = ~n16164 & ~n16317 ;
  assign n16319 = n16318 ^ n16155 ;
  assign n16311 = x97 & n7935 ;
  assign n16310 = x99 & n7938 ;
  assign n16312 = n16311 ^ n16310 ;
  assign n16313 = n16312 ^ x56 ;
  assign n16309 = n3843 & n7939 ;
  assign n16314 = n16313 ^ n16309 ;
  assign n16308 = x98 & n7931 ;
  assign n16315 = n16314 ^ n16308 ;
  assign n16302 = x94 & n8741 ;
  assign n16301 = x96 & n8744 ;
  assign n16303 = n16302 ^ n16301 ;
  assign n16304 = n16303 ^ x59 ;
  assign n16300 = n3323 & n8745 ;
  assign n16305 = n16304 ^ n16300 ;
  assign n16299 = x95 & n8737 ;
  assign n16306 = n16305 ^ n16299 ;
  assign n16292 = x91 & n9632 ;
  assign n16291 = x93 & n9635 ;
  assign n16293 = n16292 ^ n16291 ;
  assign n16294 = n16293 ^ x62 ;
  assign n16290 = n2836 & n9636 ;
  assign n16295 = n16294 ^ n16290 ;
  assign n16289 = x92 & n9628 ;
  assign n16296 = n16295 ^ n16289 ;
  assign n16285 = ~x90 & n9948 ;
  assign n16286 = n16285 ^ n16144 ;
  assign n16287 = n16286 ^ n9948 ;
  assign n16284 = x89 & n12206 ;
  assign n16288 = n16287 ^ n16284 ;
  assign n16297 = n16296 ^ n16288 ;
  assign n16281 = n16154 ^ n16143 ;
  assign n16282 = n16146 & n16281 ;
  assign n16283 = n16282 ^ n16154 ;
  assign n16298 = n16297 ^ n16283 ;
  assign n16307 = n16306 ^ n16298 ;
  assign n16316 = n16315 ^ n16307 ;
  assign n16320 = n16319 ^ n16316 ;
  assign n16329 = n16328 ^ n16320 ;
  assign n16278 = n16165 ^ n16133 ;
  assign n16279 = ~n16174 & ~n16278 ;
  assign n16280 = n16279 ^ n16165 ;
  assign n16330 = n16329 ^ n16280 ;
  assign n16331 = n16330 ^ n16175 ;
  assign n16335 = n16334 ^ n16331 ;
  assign n16344 = n16343 ^ n16335 ;
  assign n16353 = n16352 ^ n16344 ;
  assign n16275 = n16176 ^ n16112 ;
  assign n16276 = ~n16118 & ~n16275 ;
  assign n16277 = n16276 ^ n16176 ;
  assign n16354 = n16353 ^ n16277 ;
  assign n16358 = n16357 ^ n16354 ;
  assign n16367 = n16366 ^ n16358 ;
  assign n16368 = n16367 ^ n16199 ;
  assign n16372 = n16371 ^ n16368 ;
  assign n16381 = n16380 ^ n16372 ;
  assign n16382 = n16381 ^ n16210 ;
  assign n16383 = n16382 ^ n16381 ;
  assign n16384 = n16383 ^ n16103 ;
  assign n16385 = n16202 & n16384 ;
  assign n16386 = n16385 ^ n16382 ;
  assign n16395 = n16394 ^ n16386 ;
  assign n16399 = n16398 ^ n16395 ;
  assign n16408 = n16407 ^ n16399 ;
  assign n16272 = n16221 ^ n16092 ;
  assign n16273 = n16097 & ~n16272 ;
  assign n16274 = n16273 ^ n16092 ;
  assign n16409 = n16408 ^ n16274 ;
  assign n16418 = n16417 ^ n16409 ;
  assign n16269 = n16231 ^ n16084 ;
  assign n16270 = ~n16223 & ~n16269 ;
  assign n16271 = n16270 ^ n16231 ;
  assign n16419 = n16418 ^ n16271 ;
  assign n16428 = n16427 ^ n16419 ;
  assign n2023 = n2022 ^ n2018 ;
  assign n16266 = x127 & n2023 ;
  assign n16265 = n2022 & n10138 ;
  assign n16267 = n16266 ^ n16265 ;
  assign n16268 = n16267 ^ x26 ;
  assign n16429 = n16428 ^ n16268 ;
  assign n16433 = n16432 ^ n16429 ;
  assign n16262 = n16253 ^ n16081 ;
  assign n16263 = n16247 & n16262 ;
  assign n16264 = n16263 ^ n16253 ;
  assign n16434 = n16433 ^ n16264 ;
  assign n16453 = n16452 ^ n16434 ;
  assign n16617 = x125 & n2581 ;
  assign n16616 = x127 & n2422 ;
  assign n16618 = n16617 ^ n16616 ;
  assign n16619 = n16618 ^ x29 ;
  assign n16615 = n2423 & n10972 ;
  assign n16620 = n16619 ^ n16615 ;
  assign n16614 = x126 & n2429 ;
  assign n16621 = n16620 ^ n16614 ;
  assign n16607 = x122 & n2879 ;
  assign n16606 = x124 & n2882 ;
  assign n16608 = n16607 ^ n16606 ;
  assign n16609 = n16608 ^ x32 ;
  assign n16605 = n2883 & n10095 ;
  assign n16610 = n16609 ^ n16605 ;
  assign n16604 = x123 & n2887 ;
  assign n16611 = n16610 ^ n16604 ;
  assign n16598 = x119 & n3375 ;
  assign n16597 = x121 & n3378 ;
  assign n16599 = n16598 ^ n16597 ;
  assign n16600 = n16599 ^ x35 ;
  assign n16596 = n3379 & n8962 ;
  assign n16601 = n16600 ^ n16596 ;
  assign n16595 = x120 & n3383 ;
  assign n16602 = n16601 ^ n16595 ;
  assign n16590 = n16394 ^ n16381 ;
  assign n16591 = n16386 & n16590 ;
  assign n16592 = n16591 ^ n16381 ;
  assign n16584 = x116 & n3916 ;
  assign n16583 = x118 & n3919 ;
  assign n16585 = n16584 ^ n16583 ;
  assign n16586 = n16585 ^ x38 ;
  assign n16582 = n3920 & ~n8123 ;
  assign n16587 = n16586 ^ n16582 ;
  assign n16581 = x117 & n3924 ;
  assign n16588 = n16587 ^ n16581 ;
  assign n16577 = n16380 ^ n16367 ;
  assign n16578 = n16372 & n16577 ;
  assign n16579 = n16578 ^ n16367 ;
  assign n16571 = x113 & n4474 ;
  assign n16570 = x115 & n4471 ;
  assign n16572 = n16571 ^ n16570 ;
  assign n16573 = n16572 ^ x41 ;
  assign n16569 = n4472 & ~n7343 ;
  assign n16574 = n16573 ^ n16569 ;
  assign n16568 = x114 & n4467 ;
  assign n16575 = n16574 ^ n16568 ;
  assign n16564 = n16366 ^ n16357 ;
  assign n16565 = ~n16358 & ~n16564 ;
  assign n16566 = n16565 ^ n16366 ;
  assign n16562 = x111 & n5102 ;
  assign n16557 = x110 & n5094 ;
  assign n16556 = x112 & n5097 ;
  assign n16558 = n16557 ^ n16556 ;
  assign n16559 = n16558 ^ x44 ;
  assign n16555 = n5098 & ~n6600 ;
  assign n16560 = n16559 ^ n16555 ;
  assign n16551 = n16352 ^ n16277 ;
  assign n16552 = n16353 & ~n16551 ;
  assign n16553 = n16552 ^ n16352 ;
  assign n16545 = x107 & n5965 ;
  assign n16544 = x109 & n5729 ;
  assign n16546 = n16545 ^ n16544 ;
  assign n16547 = n16546 ^ x47 ;
  assign n16543 = n5730 & n5902 ;
  assign n16548 = n16547 ^ n16543 ;
  assign n16542 = x108 & n5736 ;
  assign n16549 = n16548 ^ n16542 ;
  assign n16537 = ~n4615 & n7175 ;
  assign n16535 = x101 & n7171 ;
  assign n16533 = x103 & n7174 ;
  assign n16529 = n16328 ^ n16280 ;
  assign n16530 = n16329 & ~n16529 ;
  assign n16531 = n16530 ^ n16328 ;
  assign n16532 = n16531 ^ x53 ;
  assign n16534 = n16533 ^ n16532 ;
  assign n16536 = n16535 ^ n16534 ;
  assign n16538 = n16537 ^ n16536 ;
  assign n16528 = x102 & n7179 ;
  assign n16539 = n16538 ^ n16528 ;
  assign n16521 = x98 & n7935 ;
  assign n16520 = x100 & n7938 ;
  assign n16522 = n16521 ^ n16520 ;
  assign n16523 = n16522 ^ x56 ;
  assign n16519 = n4034 & n7939 ;
  assign n16524 = n16523 ^ n16519 ;
  assign n16518 = x99 & n7931 ;
  assign n16525 = n16524 ^ n16518 ;
  assign n16515 = x96 & n8737 ;
  assign n16513 = n3494 & n8745 ;
  assign n16509 = x95 & n8741 ;
  assign n16508 = x97 & n8744 ;
  assign n16510 = n16509 ^ n16508 ;
  assign n16511 = n16510 ^ x59 ;
  assign n16502 = ~n16288 & n16296 ;
  assign n16501 = x89 & n16286 ;
  assign n16503 = n16502 ^ n16501 ;
  assign n16504 = n16503 ^ n16144 ;
  assign n16505 = n16504 ^ x26 ;
  assign n16497 = x91 ^ x89 ;
  assign n16498 = ~n11875 & n16497 ;
  assign n16499 = n16498 ^ n2103 ;
  assign n16500 = n12206 & n16499 ;
  assign n16506 = n16505 ^ n16500 ;
  assign n16492 = x92 & n9632 ;
  assign n16491 = x94 & n9635 ;
  assign n16493 = n16492 ^ n16491 ;
  assign n16494 = n16493 ^ x62 ;
  assign n16490 = n2997 & n9636 ;
  assign n16495 = n16494 ^ n16490 ;
  assign n16489 = x93 & n9628 ;
  assign n16496 = n16495 ^ n16489 ;
  assign n16507 = n16506 ^ n16496 ;
  assign n16512 = n16511 ^ n16507 ;
  assign n16514 = n16513 ^ n16512 ;
  assign n16516 = n16515 ^ n16514 ;
  assign n16486 = n16306 ^ n16283 ;
  assign n16487 = n16298 & n16486 ;
  assign n16488 = n16487 ^ n16306 ;
  assign n16517 = n16516 ^ n16488 ;
  assign n16526 = n16525 ^ n16517 ;
  assign n16483 = n16319 ^ n16315 ;
  assign n16484 = n16316 & ~n16483 ;
  assign n16485 = n16484 ^ n16319 ;
  assign n16527 = n16526 ^ n16485 ;
  assign n16540 = n16539 ^ n16527 ;
  assign n16473 = x104 & n6677 ;
  assign n16472 = x106 & n6428 ;
  assign n16474 = n16473 ^ n16472 ;
  assign n16475 = n16474 ^ x50 ;
  assign n16471 = ~n5240 & n6429 ;
  assign n16476 = n16475 ^ n16471 ;
  assign n16470 = x105 & n6433 ;
  assign n16477 = n16476 ^ n16470 ;
  assign n16479 = n16477 ^ n16330 ;
  assign n16478 = n16477 ^ n16343 ;
  assign n16480 = n16479 ^ n16478 ;
  assign n16481 = n16335 & ~n16480 ;
  assign n16482 = n16481 ^ n16479 ;
  assign n16541 = n16540 ^ n16482 ;
  assign n16550 = n16549 ^ n16541 ;
  assign n16554 = n16553 ^ n16550 ;
  assign n16561 = n16560 ^ n16554 ;
  assign n16563 = n16562 ^ n16561 ;
  assign n16567 = n16566 ^ n16563 ;
  assign n16576 = n16575 ^ n16567 ;
  assign n16580 = n16579 ^ n16576 ;
  assign n16589 = n16588 ^ n16580 ;
  assign n16593 = n16592 ^ n16589 ;
  assign n16467 = n16407 ^ n16398 ;
  assign n16468 = ~n16399 & n16467 ;
  assign n16469 = n16468 ^ n16407 ;
  assign n16594 = n16593 ^ n16469 ;
  assign n16603 = n16602 ^ n16594 ;
  assign n16612 = n16611 ^ n16603 ;
  assign n16464 = n16417 ^ n16274 ;
  assign n16465 = ~n16409 & n16464 ;
  assign n16466 = n16465 ^ n16417 ;
  assign n16613 = n16612 ^ n16466 ;
  assign n16622 = n16621 ^ n16613 ;
  assign n16461 = n16427 ^ n16271 ;
  assign n16462 = ~n16419 & n16461 ;
  assign n16463 = n16462 ^ n16427 ;
  assign n16623 = n16622 ^ n16463 ;
  assign n16460 = ~n16264 & ~n16432 ;
  assign n16624 = n16623 ^ n16460 ;
  assign n16455 = n16432 ^ n16264 ;
  assign n16454 = n16452 ^ n16428 ;
  assign n16458 = n16455 ^ n16454 ;
  assign n16459 = n16268 & ~n16458 ;
  assign n16625 = n16624 ^ n16459 ;
  assign n16456 = n16455 ^ n16428 ;
  assign n16457 = n16454 & n16456 ;
  assign n16626 = n16625 ^ n16457 ;
  assign n16813 = n2423 & n10139 ;
  assign n16812 = x126 & n2581 ;
  assign n16814 = n16813 ^ n16812 ;
  assign n16815 = n16814 ^ x29 ;
  assign n16811 = x127 & n2429 ;
  assign n16816 = n16815 ^ n16811 ;
  assign n16807 = n16611 ^ n16466 ;
  assign n16808 = ~n16612 & n16807 ;
  assign n16809 = n16808 ^ n16611 ;
  assign n16801 = x123 & n2879 ;
  assign n16800 = x125 & n2882 ;
  assign n16802 = n16801 ^ n16800 ;
  assign n16803 = n16802 ^ x32 ;
  assign n16799 = n2883 & n10400 ;
  assign n16804 = n16803 ^ n16799 ;
  assign n16798 = x124 & n2887 ;
  assign n16805 = n16804 ^ n16798 ;
  assign n16787 = x120 & n3375 ;
  assign n16786 = x122 & n3378 ;
  assign n16788 = n16787 ^ n16786 ;
  assign n16789 = n16788 ^ x35 ;
  assign n16785 = n3379 & ~n9247 ;
  assign n16790 = n16789 ^ n16785 ;
  assign n16784 = x121 & n3383 ;
  assign n16791 = n16790 ^ n16784 ;
  assign n16777 = x117 & n3916 ;
  assign n16776 = x119 & n3919 ;
  assign n16778 = n16777 ^ n16776 ;
  assign n16779 = n16778 ^ x38 ;
  assign n16775 = n3920 & n8394 ;
  assign n16780 = n16779 ^ n16775 ;
  assign n16774 = x118 & n3924 ;
  assign n16781 = n16780 ^ n16774 ;
  assign n16767 = x114 & n4474 ;
  assign n16766 = x116 & n4471 ;
  assign n16768 = n16767 ^ n16766 ;
  assign n16769 = n16768 ^ x41 ;
  assign n16765 = n4472 & ~n7588 ;
  assign n16770 = n16769 ^ n16765 ;
  assign n16764 = x115 & n4467 ;
  assign n16771 = n16770 ^ n16764 ;
  assign n16757 = x111 & n5094 ;
  assign n16756 = x113 & n5097 ;
  assign n16758 = n16757 ^ n16756 ;
  assign n16759 = n16758 ^ x44 ;
  assign n16755 = n5098 & ~n6839 ;
  assign n16760 = n16759 ^ n16755 ;
  assign n16754 = x112 & n5102 ;
  assign n16761 = n16760 ^ n16754 ;
  assign n16743 = x108 & n5965 ;
  assign n16742 = x110 & n5729 ;
  assign n16744 = n16743 ^ n16742 ;
  assign n16745 = n16744 ^ x47 ;
  assign n16741 = n5730 & n6129 ;
  assign n16746 = n16745 ^ n16741 ;
  assign n16740 = x109 & n5736 ;
  assign n16747 = n16746 ^ n16740 ;
  assign n16729 = x105 & n6677 ;
  assign n16728 = x107 & n6428 ;
  assign n16730 = n16729 ^ n16728 ;
  assign n16731 = n16730 ^ x50 ;
  assign n16727 = ~n5448 & n6429 ;
  assign n16732 = n16731 ^ n16727 ;
  assign n16726 = x106 & n6433 ;
  assign n16733 = n16732 ^ n16726 ;
  assign n16721 = n16525 ^ n16485 ;
  assign n16722 = ~n16526 & ~n16721 ;
  assign n16723 = n16722 ^ n16525 ;
  assign n16715 = x102 & n7171 ;
  assign n16714 = x104 & n7174 ;
  assign n16716 = n16715 ^ n16714 ;
  assign n16717 = n16716 ^ x53 ;
  assign n16713 = ~n4814 & n7175 ;
  assign n16718 = n16717 ^ n16713 ;
  assign n16712 = x103 & n7179 ;
  assign n16719 = n16718 ^ n16712 ;
  assign n16708 = x97 & n8737 ;
  assign n16706 = n3660 & n8745 ;
  assign n16702 = x96 & n8741 ;
  assign n16701 = x98 & n8744 ;
  assign n16703 = n16702 ^ n16701 ;
  assign n16704 = n16703 ^ x59 ;
  assign n16695 = x93 & n9632 ;
  assign n16694 = x95 & n9635 ;
  assign n16696 = n16695 ^ n16694 ;
  assign n16697 = n16696 ^ x62 ;
  assign n16693 = n3159 & n9636 ;
  assign n16698 = n16697 ^ n16693 ;
  assign n16692 = x94 & n9628 ;
  assign n16699 = n16698 ^ n16692 ;
  assign n16688 = ~x63 & x91 ;
  assign n16689 = n16688 ^ n2370 ;
  assign n16690 = ~n9948 & n16689 ;
  assign n16677 = x90 ^ x26 ;
  assign n16680 = n16499 & ~n16677 ;
  assign n16681 = n16680 ^ x90 ;
  assign n16682 = n12206 & n16681 ;
  assign n16683 = n16682 ^ x92 ;
  assign n16691 = n16690 ^ n16683 ;
  assign n16700 = n16699 ^ n16691 ;
  assign n16705 = n16704 ^ n16700 ;
  assign n16707 = n16706 ^ n16705 ;
  assign n16709 = n16708 ^ n16707 ;
  assign n16674 = n16504 ^ n16496 ;
  assign n16675 = ~n16506 & n16674 ;
  assign n16676 = n16675 ^ n16504 ;
  assign n16710 = n16709 ^ n16676 ;
  assign n16671 = n4215 & n7939 ;
  assign n16669 = x99 & n7935 ;
  assign n16665 = n16507 ^ n16488 ;
  assign n16666 = ~n16516 & ~n16665 ;
  assign n16667 = n16666 ^ n16507 ;
  assign n16663 = x101 & n7938 ;
  assign n16664 = n16663 ^ x56 ;
  assign n16668 = n16667 ^ n16664 ;
  assign n16670 = n16669 ^ n16668 ;
  assign n16672 = n16671 ^ n16670 ;
  assign n16662 = x100 & n7931 ;
  assign n16673 = n16672 ^ n16662 ;
  assign n16711 = n16710 ^ n16673 ;
  assign n16720 = n16719 ^ n16711 ;
  assign n16724 = n16723 ^ n16720 ;
  assign n16659 = n16531 ^ n16527 ;
  assign n16660 = n16539 & n16659 ;
  assign n16661 = n16660 ^ n16531 ;
  assign n16725 = n16724 ^ n16661 ;
  assign n16734 = n16733 ^ n16725 ;
  assign n16736 = n16734 ^ n16477 ;
  assign n16735 = n16734 ^ n16540 ;
  assign n16737 = n16736 ^ n16735 ;
  assign n16738 = ~n16482 & n16737 ;
  assign n16739 = n16738 ^ n16736 ;
  assign n16748 = n16747 ^ n16739 ;
  assign n16749 = n16748 ^ n16553 ;
  assign n16750 = n16749 ^ n16541 ;
  assign n16751 = n16750 ^ n16748 ;
  assign n16752 = n16550 & ~n16751 ;
  assign n16753 = n16752 ^ n16749 ;
  assign n16762 = n16761 ^ n16753 ;
  assign n16656 = n16566 ^ n16554 ;
  assign n16657 = ~n16563 & ~n16656 ;
  assign n16658 = n16657 ^ n16554 ;
  assign n16763 = n16762 ^ n16658 ;
  assign n16772 = n16771 ^ n16763 ;
  assign n16653 = n16579 ^ n16575 ;
  assign n16654 = n16576 & n16653 ;
  assign n16655 = n16654 ^ n16579 ;
  assign n16773 = n16772 ^ n16655 ;
  assign n16782 = n16781 ^ n16773 ;
  assign n16650 = n16592 ^ n16588 ;
  assign n16651 = n16589 & n16650 ;
  assign n16652 = n16651 ^ n16592 ;
  assign n16783 = n16782 ^ n16652 ;
  assign n16792 = n16791 ^ n16783 ;
  assign n16793 = n16792 ^ n16602 ;
  assign n16794 = n16793 ^ n16792 ;
  assign n16795 = n16794 ^ n16469 ;
  assign n16796 = n16594 & n16795 ;
  assign n16797 = n16796 ^ n16793 ;
  assign n16806 = n16805 ^ n16797 ;
  assign n16810 = n16809 ^ n16806 ;
  assign n16817 = n16816 ^ n16810 ;
  assign n16647 = n16621 ^ n16463 ;
  assign n16648 = ~n16622 & n16647 ;
  assign n16649 = n16648 ^ n16621 ;
  assign n16818 = n16817 ^ n16649 ;
  assign n16627 = ~n16268 & ~n16428 ;
  assign n16628 = n16627 ^ n16429 ;
  assign n16629 = n16628 ^ n16623 ;
  assign n16634 = ~n16452 & ~n16627 ;
  assign n16630 = n16460 ^ n16268 ;
  assign n16631 = n16429 & ~n16630 ;
  assign n16632 = n16631 ^ n16268 ;
  assign n16633 = ~n16623 & n16632 ;
  assign n16635 = n16624 ^ n16455 ;
  assign n16636 = ~n16633 & n16635 ;
  assign n16637 = n16634 & n16636 ;
  assign n16638 = n16637 ^ n16633 ;
  assign n16639 = n16452 ^ n16432 ;
  assign n16642 = n16455 & ~n16639 ;
  assign n16643 = n16642 ^ n16432 ;
  assign n16644 = ~n16638 & n16643 ;
  assign n16645 = n16629 & n16644 ;
  assign n16646 = n16645 ^ n16638 ;
  assign n16819 = n16818 ^ n16646 ;
  assign n16991 = n16649 ^ n16646 ;
  assign n16992 = n16818 & n16991 ;
  assign n16993 = n16992 ^ n16646 ;
  assign n16979 = x127 & n2580 ;
  assign n16980 = n16979 ^ n2421 ;
  assign n16985 = n2164 & n11265 ;
  assign n16986 = n16985 ^ n16979 ;
  assign n16987 = n16980 & ~n16986 ;
  assign n16988 = n16987 ^ x28 ;
  assign n16968 = x124 & n2879 ;
  assign n16967 = x126 & n2882 ;
  assign n16969 = n16968 ^ n16967 ;
  assign n16970 = n16969 ^ x32 ;
  assign n16966 = n2883 & n10441 ;
  assign n16971 = n16970 ^ n16966 ;
  assign n16965 = x125 & n2887 ;
  assign n16972 = n16971 ^ n16965 ;
  assign n16954 = x121 & n3375 ;
  assign n16953 = x123 & n3378 ;
  assign n16955 = n16954 ^ n16953 ;
  assign n16956 = n16955 ^ x35 ;
  assign n16952 = n3379 & ~n9786 ;
  assign n16957 = n16956 ^ n16952 ;
  assign n16951 = x122 & n3383 ;
  assign n16958 = n16957 ^ n16951 ;
  assign n16947 = n16781 ^ n16655 ;
  assign n16948 = n16773 & n16947 ;
  assign n16949 = n16948 ^ n16781 ;
  assign n16941 = x118 & n3916 ;
  assign n16940 = x120 & n3919 ;
  assign n16942 = n16941 ^ n16940 ;
  assign n16943 = n16942 ^ x38 ;
  assign n16939 = n3920 & n8891 ;
  assign n16944 = n16943 ^ n16939 ;
  assign n16938 = x119 & n3924 ;
  assign n16945 = n16944 ^ n16938 ;
  assign n16935 = n16771 ^ n16658 ;
  assign n16936 = n16763 & ~n16935 ;
  assign n16927 = x115 & n4474 ;
  assign n16926 = x117 & n4471 ;
  assign n16928 = n16927 ^ n16926 ;
  assign n16929 = n16928 ^ x41 ;
  assign n16925 = n4472 & ~n7850 ;
  assign n16930 = n16929 ^ n16925 ;
  assign n16924 = x116 & n4467 ;
  assign n16931 = n16930 ^ n16924 ;
  assign n16913 = x112 & n5094 ;
  assign n16912 = x114 & n5097 ;
  assign n16914 = n16913 ^ n16912 ;
  assign n16915 = n16914 ^ x44 ;
  assign n16911 = n5098 & ~n7092 ;
  assign n16916 = n16915 ^ n16911 ;
  assign n16910 = x113 & n5102 ;
  assign n16917 = n16916 ^ n16910 ;
  assign n16899 = x109 & n5965 ;
  assign n16898 = x111 & n5729 ;
  assign n16900 = n16899 ^ n16898 ;
  assign n16901 = n16900 ^ x47 ;
  assign n16897 = n5730 & ~n6360 ;
  assign n16902 = n16901 ^ n16897 ;
  assign n16896 = x110 & n5736 ;
  assign n16903 = n16902 ^ n16896 ;
  assign n16886 = x97 & n8741 ;
  assign n16885 = x99 & n8744 ;
  assign n16887 = n16886 ^ n16885 ;
  assign n16888 = n16887 ^ x59 ;
  assign n16884 = n3843 & n8745 ;
  assign n16889 = n16888 ^ n16884 ;
  assign n16883 = x98 & n8737 ;
  assign n16890 = n16889 ^ n16883 ;
  assign n16881 = x95 & n9628 ;
  assign n16872 = x63 & n2370 ;
  assign n16873 = n16872 ^ n2520 ;
  assign n16874 = ~n9948 & n16873 ;
  assign n16875 = n16874 ^ n2520 ;
  assign n16865 = n16699 ^ n16682 ;
  assign n16866 = n16691 & n16865 ;
  assign n16867 = n16866 ^ n16699 ;
  assign n16876 = n16875 ^ n16867 ;
  assign n16877 = n16876 ^ x62 ;
  assign n16864 = x94 & n9632 ;
  assign n16878 = n16877 ^ n16864 ;
  assign n16863 = x96 & n9635 ;
  assign n16879 = n16878 ^ n16863 ;
  assign n16862 = n3323 & n9636 ;
  assign n16880 = n16879 ^ n16862 ;
  assign n16882 = n16881 ^ n16880 ;
  assign n16891 = n16890 ^ n16882 ;
  assign n16859 = n4410 & n7939 ;
  assign n16857 = x100 & n7935 ;
  assign n16853 = n16700 ^ n16676 ;
  assign n16854 = ~n16709 & ~n16853 ;
  assign n16855 = n16854 ^ n16700 ;
  assign n16851 = x102 & n7938 ;
  assign n16852 = n16851 ^ x56 ;
  assign n16856 = n16855 ^ n16852 ;
  assign n16858 = n16857 ^ n16856 ;
  assign n16860 = n16859 ^ n16858 ;
  assign n16850 = x101 & n7931 ;
  assign n16861 = n16860 ^ n16850 ;
  assign n16892 = n16891 ^ n16861 ;
  assign n16847 = ~n5023 & n7175 ;
  assign n16845 = x103 & n7171 ;
  assign n16841 = n16710 ^ n16667 ;
  assign n16842 = n16673 & n16841 ;
  assign n16843 = n16842 ^ n16710 ;
  assign n16839 = x105 & n7174 ;
  assign n16840 = n16839 ^ x53 ;
  assign n16844 = n16843 ^ n16840 ;
  assign n16846 = n16845 ^ n16844 ;
  assign n16848 = n16847 ^ n16846 ;
  assign n16838 = x104 & n7179 ;
  assign n16849 = n16848 ^ n16838 ;
  assign n16893 = n16892 ^ n16849 ;
  assign n16835 = n5670 & n6429 ;
  assign n16833 = x106 & n6677 ;
  assign n16829 = n16723 ^ n16719 ;
  assign n16830 = ~n16720 & n16829 ;
  assign n16831 = n16830 ^ n16723 ;
  assign n16827 = x108 & n6428 ;
  assign n16828 = n16827 ^ x50 ;
  assign n16832 = n16831 ^ n16828 ;
  assign n16834 = n16833 ^ n16832 ;
  assign n16836 = n16835 ^ n16834 ;
  assign n16826 = x107 & n6433 ;
  assign n16837 = n16836 ^ n16826 ;
  assign n16894 = n16893 ^ n16837 ;
  assign n16823 = n16733 ^ n16661 ;
  assign n16824 = ~n16725 & n16823 ;
  assign n16825 = n16824 ^ n16733 ;
  assign n16895 = n16894 ^ n16825 ;
  assign n16904 = n16903 ^ n16895 ;
  assign n16906 = n16904 ^ n16734 ;
  assign n16905 = n16904 ^ n16747 ;
  assign n16907 = n16906 ^ n16905 ;
  assign n16908 = n16739 & n16907 ;
  assign n16909 = n16908 ^ n16906 ;
  assign n16918 = n16917 ^ n16909 ;
  assign n16920 = n16918 ^ n16748 ;
  assign n16919 = n16918 ^ n16761 ;
  assign n16921 = n16920 ^ n16919 ;
  assign n16922 = n16753 & n16921 ;
  assign n16923 = n16922 ^ n16920 ;
  assign n16932 = n16931 ^ n16923 ;
  assign n16933 = n16932 ^ n16771 ;
  assign n16937 = n16936 ^ n16933 ;
  assign n16946 = n16945 ^ n16937 ;
  assign n16950 = n16949 ^ n16946 ;
  assign n16959 = n16958 ^ n16950 ;
  assign n16960 = n16959 ^ n16791 ;
  assign n16961 = n16960 ^ n16959 ;
  assign n16962 = n16961 ^ n16652 ;
  assign n16963 = n16783 & n16962 ;
  assign n16964 = n16963 ^ n16960 ;
  assign n16973 = n16972 ^ n16964 ;
  assign n16975 = n16973 ^ n16792 ;
  assign n16974 = n16973 ^ n16805 ;
  assign n16976 = n16975 ^ n16974 ;
  assign n16977 = ~n16797 & ~n16976 ;
  assign n16978 = n16977 ^ n16975 ;
  assign n16989 = n16988 ^ n16978 ;
  assign n16820 = n16816 ^ n16809 ;
  assign n16821 = n16810 & n16820 ;
  assign n16822 = n16821 ^ n16816 ;
  assign n16990 = n16989 ^ n16822 ;
  assign n16994 = n16993 ^ n16990 ;
  assign n17153 = n16972 ^ n16959 ;
  assign n17154 = ~n16964 & ~n17153 ;
  assign n17155 = n17154 ^ n16959 ;
  assign n17150 = n16988 ^ n16973 ;
  assign n17151 = n16978 & ~n17150 ;
  assign n17152 = n17151 ^ n16973 ;
  assign n17156 = n17155 ^ n17152 ;
  assign n17144 = x125 & n2879 ;
  assign n17143 = x127 & n2882 ;
  assign n17145 = n17144 ^ n17143 ;
  assign n17146 = n17145 ^ x32 ;
  assign n17142 = n2883 & n10972 ;
  assign n17147 = n17146 ^ n17142 ;
  assign n17141 = x126 & n2887 ;
  assign n17148 = n17147 ^ n17141 ;
  assign n17134 = x122 & n3375 ;
  assign n17133 = x124 & n3378 ;
  assign n17135 = n17134 ^ n17133 ;
  assign n17136 = n17135 ^ x35 ;
  assign n17132 = n3379 & n10095 ;
  assign n17137 = n17136 ^ n17132 ;
  assign n17131 = x123 & n3383 ;
  assign n17138 = n17137 ^ n17131 ;
  assign n17125 = x119 & n3916 ;
  assign n17124 = x121 & n3919 ;
  assign n17126 = n17125 ^ n17124 ;
  assign n17127 = n17126 ^ x38 ;
  assign n17123 = n3920 & n8962 ;
  assign n17128 = n17127 ^ n17123 ;
  assign n17122 = x120 & n3924 ;
  assign n17129 = n17128 ^ n17122 ;
  assign n17113 = n16931 ^ n16918 ;
  assign n17114 = ~n16923 & ~n17113 ;
  assign n17115 = n17114 ^ n16918 ;
  assign n17107 = x116 & n4474 ;
  assign n17106 = x118 & n4471 ;
  assign n17108 = n17107 ^ n17106 ;
  assign n17109 = n17108 ^ x41 ;
  assign n17105 = n4472 & ~n8123 ;
  assign n17110 = n17109 ^ n17105 ;
  assign n17104 = x117 & n4467 ;
  assign n17111 = n17110 ^ n17104 ;
  assign n17100 = n16917 ^ n16904 ;
  assign n17101 = ~n16909 & ~n17100 ;
  assign n17102 = n17101 ^ n16904 ;
  assign n17094 = x113 & n5094 ;
  assign n17093 = x115 & n5097 ;
  assign n17095 = n17094 ^ n17093 ;
  assign n17096 = n17095 ^ x44 ;
  assign n17092 = n5098 & ~n7343 ;
  assign n17097 = n17096 ^ n17092 ;
  assign n17091 = x114 & n5102 ;
  assign n17098 = n17097 ^ n17091 ;
  assign n17084 = x110 & n5965 ;
  assign n17083 = x112 & n5729 ;
  assign n17085 = n17084 ^ n17083 ;
  assign n17086 = n17085 ^ x47 ;
  assign n17082 = n5730 & ~n6600 ;
  assign n17087 = n17086 ^ n17082 ;
  assign n17081 = x111 & n5736 ;
  assign n17088 = n17087 ^ n17081 ;
  assign n17069 = x95 & n9632 ;
  assign n17068 = x97 & n9635 ;
  assign n17070 = n17069 ^ n17068 ;
  assign n17071 = n17070 ^ x62 ;
  assign n17067 = n3494 & n9636 ;
  assign n17072 = n17071 ^ n17067 ;
  assign n17066 = x96 & n9628 ;
  assign n17073 = n17072 ^ n17066 ;
  assign n17074 = n17073 ^ x29 ;
  assign n17062 = x94 ^ x92 ;
  assign n17063 = ~n11875 & n17062 ;
  assign n17064 = n17063 ^ n2520 ;
  assign n17065 = n12206 & n17064 ;
  assign n17075 = n17074 ^ n17065 ;
  assign n17060 = ~n16867 & ~n16875 ;
  assign n17054 = n9948 ^ x92 ;
  assign n17055 = x63 & ~x91 ;
  assign n17056 = n17055 ^ x93 ;
  assign n17057 = x92 & n17056 ;
  assign n17058 = n17057 ^ x93 ;
  assign n17059 = n17054 & n17058 ;
  assign n17061 = n17060 ^ n17059 ;
  assign n17076 = n17075 ^ n17061 ;
  assign n17044 = x98 & n8741 ;
  assign n17043 = x100 & n8744 ;
  assign n17045 = n17044 ^ n17043 ;
  assign n17046 = n17045 ^ x59 ;
  assign n17042 = n4034 & n8745 ;
  assign n17047 = n17046 ^ n17042 ;
  assign n17041 = x99 & n8737 ;
  assign n17048 = n17047 ^ n17041 ;
  assign n17049 = n17048 ^ n16890 ;
  assign n17050 = n17049 ^ n16876 ;
  assign n17051 = n17050 ^ n17048 ;
  assign n17052 = n16882 & ~n17051 ;
  assign n17053 = n17052 ^ n17049 ;
  assign n17077 = n17076 ^ n17053 ;
  assign n17038 = ~n4615 & n7939 ;
  assign n17036 = x101 & n7935 ;
  assign n17032 = n16891 ^ n16855 ;
  assign n17033 = n16861 & n17032 ;
  assign n17034 = n17033 ^ n16891 ;
  assign n17030 = x103 & n7938 ;
  assign n17031 = n17030 ^ x56 ;
  assign n17035 = n17034 ^ n17031 ;
  assign n17037 = n17036 ^ n17035 ;
  assign n17039 = n17038 ^ n17037 ;
  assign n17029 = x102 & n7931 ;
  assign n17040 = n17039 ^ n17029 ;
  assign n17078 = n17077 ^ n17040 ;
  assign n17026 = n16892 ^ n16843 ;
  assign n17027 = n16849 & ~n17026 ;
  assign n17019 = x104 & n7171 ;
  assign n17018 = x106 & n7174 ;
  assign n17020 = n17019 ^ n17018 ;
  assign n17021 = n17020 ^ x53 ;
  assign n17017 = ~n5240 & n7175 ;
  assign n17022 = n17021 ^ n17017 ;
  assign n17016 = x105 & n7179 ;
  assign n17023 = n17022 ^ n17016 ;
  assign n17024 = n17023 ^ n16892 ;
  assign n17028 = n17027 ^ n17024 ;
  assign n17079 = n17078 ^ n17028 ;
  assign n17013 = n5902 & n6429 ;
  assign n17011 = x107 & n6677 ;
  assign n17009 = x109 & n6428 ;
  assign n17005 = n16893 ^ n16831 ;
  assign n17006 = ~n16837 & ~n17005 ;
  assign n17007 = n17006 ^ n16893 ;
  assign n17008 = n17007 ^ x50 ;
  assign n17010 = n17009 ^ n17008 ;
  assign n17012 = n17011 ^ n17010 ;
  assign n17014 = n17013 ^ n17012 ;
  assign n17004 = x108 & n6433 ;
  assign n17015 = n17014 ^ n17004 ;
  assign n17080 = n17079 ^ n17015 ;
  assign n17089 = n17088 ^ n17080 ;
  assign n17001 = n16903 ^ n16825 ;
  assign n17002 = n16895 & n17001 ;
  assign n17003 = n17002 ^ n16903 ;
  assign n17090 = n17089 ^ n17003 ;
  assign n17099 = n17098 ^ n17090 ;
  assign n17103 = n17102 ^ n17099 ;
  assign n17112 = n17111 ^ n17103 ;
  assign n17116 = n17115 ^ n17112 ;
  assign n17118 = n17116 ^ n16932 ;
  assign n17117 = n17116 ^ n16945 ;
  assign n17119 = n17118 ^ n17117 ;
  assign n17120 = ~n16937 & ~n17119 ;
  assign n17121 = n17120 ^ n17118 ;
  assign n17130 = n17129 ^ n17121 ;
  assign n17139 = n17138 ^ n17130 ;
  assign n16998 = n16958 ^ n16949 ;
  assign n16999 = n16950 & n16998 ;
  assign n17000 = n16999 ^ n16958 ;
  assign n17140 = n17139 ^ n17000 ;
  assign n17149 = n17148 ^ n17140 ;
  assign n17157 = n17156 ^ n17149 ;
  assign n16995 = n16993 ^ n16822 ;
  assign n16996 = ~n16990 & n16995 ;
  assign n16997 = n16996 ^ n16993 ;
  assign n17158 = n17157 ^ n16997 ;
  assign n17310 = n17140 & ~n17148 ;
  assign n17311 = n17310 ^ n17149 ;
  assign n17309 = n17152 & n17155 ;
  assign n17312 = n17311 ^ n17309 ;
  assign n17304 = n2883 & n10139 ;
  assign n17303 = x126 & n2879 ;
  assign n17305 = n17304 ^ n17303 ;
  assign n17306 = n17305 ^ x32 ;
  assign n17302 = x127 & n2887 ;
  assign n17307 = n17306 ^ n17302 ;
  assign n17298 = n17138 ^ n17000 ;
  assign n17299 = ~n17139 & n17298 ;
  assign n17300 = n17299 ^ n17138 ;
  assign n17292 = x123 & n3375 ;
  assign n17291 = x125 & n3378 ;
  assign n17293 = n17292 ^ n17291 ;
  assign n17294 = n17293 ^ x35 ;
  assign n17290 = n3379 & n10400 ;
  assign n17295 = n17294 ^ n17290 ;
  assign n17289 = x124 & n3383 ;
  assign n17296 = n17295 ^ n17289 ;
  assign n17285 = n17129 ^ n17116 ;
  assign n17286 = ~n17121 & n17285 ;
  assign n17287 = n17286 ^ n17116 ;
  assign n17279 = x120 & n3916 ;
  assign n17278 = x122 & n3919 ;
  assign n17280 = n17279 ^ n17278 ;
  assign n17281 = n17280 ^ x38 ;
  assign n17277 = n3920 & ~n9247 ;
  assign n17282 = n17281 ^ n17277 ;
  assign n17276 = x121 & n3924 ;
  assign n17283 = n17282 ^ n17276 ;
  assign n17269 = x117 & n4474 ;
  assign n17268 = x119 & n4471 ;
  assign n17270 = n17269 ^ n17268 ;
  assign n17271 = n17270 ^ x41 ;
  assign n17267 = n4472 & n8394 ;
  assign n17272 = n17271 ^ n17267 ;
  assign n17266 = x118 & n4467 ;
  assign n17273 = n17272 ^ n17266 ;
  assign n17259 = x114 & n5094 ;
  assign n17258 = x116 & n5097 ;
  assign n17260 = n17259 ^ n17258 ;
  assign n17261 = n17260 ^ x44 ;
  assign n17257 = n5098 & ~n7588 ;
  assign n17262 = n17261 ^ n17257 ;
  assign n17256 = x115 & n5102 ;
  assign n17263 = n17262 ^ n17256 ;
  assign n17249 = x111 & n5965 ;
  assign n17248 = x113 & n5729 ;
  assign n17250 = n17249 ^ n17248 ;
  assign n17251 = n17250 ^ x47 ;
  assign n17247 = n5730 & ~n6839 ;
  assign n17252 = n17251 ^ n17247 ;
  assign n17246 = x112 & n5736 ;
  assign n17253 = n17252 ^ n17246 ;
  assign n17236 = ~n5448 & n7175 ;
  assign n17234 = x105 & n7171 ;
  assign n17230 = n17077 ^ n17034 ;
  assign n17231 = n17040 & ~n17230 ;
  assign n17232 = n17231 ^ n17077 ;
  assign n17228 = x107 & n7174 ;
  assign n17229 = n17228 ^ x53 ;
  assign n17233 = n17232 ^ n17229 ;
  assign n17235 = n17234 ^ n17233 ;
  assign n17237 = n17236 ^ n17235 ;
  assign n17227 = x106 & n7179 ;
  assign n17238 = n17237 ^ n17227 ;
  assign n17224 = x103 & n7931 ;
  assign n17222 = ~n4814 & n7939 ;
  assign n17218 = x102 & n7935 ;
  assign n17217 = x104 & n7938 ;
  assign n17219 = n17218 ^ n17217 ;
  assign n17220 = n17219 ^ x56 ;
  assign n17213 = n4215 & n8745 ;
  assign n17211 = x99 & n8741 ;
  assign n17207 = x94 & n11875 ;
  assign n17206 = x95 & n9948 ;
  assign n17208 = n17207 ^ n17206 ;
  assign n17203 = n3660 & n9636 ;
  assign n17201 = x96 & n9632 ;
  assign n17194 = x93 ^ x29 ;
  assign n17197 = n17064 & ~n17194 ;
  assign n17198 = n17197 ^ x93 ;
  assign n17199 = n12206 & n17198 ;
  assign n17192 = x98 & n9635 ;
  assign n17193 = n17192 ^ x62 ;
  assign n17200 = n17199 ^ n17193 ;
  assign n17202 = n17201 ^ n17200 ;
  assign n17204 = n17203 ^ n17202 ;
  assign n17191 = x97 & n9628 ;
  assign n17205 = n17204 ^ n17191 ;
  assign n17209 = n17208 ^ n17205 ;
  assign n17189 = x101 & n8744 ;
  assign n17190 = n17189 ^ x59 ;
  assign n17210 = n17209 ^ n17190 ;
  assign n17212 = n17211 ^ n17210 ;
  assign n17214 = n17213 ^ n17212 ;
  assign n17188 = x100 & n8737 ;
  assign n17215 = n17214 ^ n17188 ;
  assign n17185 = n17073 ^ n17061 ;
  assign n17186 = ~n17075 & ~n17185 ;
  assign n17187 = n17186 ^ n17073 ;
  assign n17216 = n17215 ^ n17187 ;
  assign n17221 = n17220 ^ n17216 ;
  assign n17223 = n17222 ^ n17221 ;
  assign n17225 = n17224 ^ n17223 ;
  assign n17182 = n17076 ^ n17048 ;
  assign n17183 = n17053 & n17182 ;
  assign n17184 = n17183 ^ n17048 ;
  assign n17226 = n17225 ^ n17184 ;
  assign n17239 = n17238 ^ n17226 ;
  assign n17179 = n6129 & n6429 ;
  assign n17177 = x108 & n6677 ;
  assign n17173 = n17078 ^ n17023 ;
  assign n17174 = n17028 & ~n17173 ;
  assign n17175 = n17174 ^ n17023 ;
  assign n17171 = x110 & n6428 ;
  assign n17172 = n17171 ^ x50 ;
  assign n17176 = n17175 ^ n17172 ;
  assign n17178 = n17177 ^ n17176 ;
  assign n17180 = n17179 ^ n17178 ;
  assign n17170 = x109 & n6433 ;
  assign n17181 = n17180 ^ n17170 ;
  assign n17240 = n17239 ^ n17181 ;
  assign n17241 = n17240 ^ n17079 ;
  assign n17242 = n17241 ^ n17007 ;
  assign n17243 = n17242 ^ n17240 ;
  assign n17244 = n17015 & n17243 ;
  assign n17245 = n17244 ^ n17241 ;
  assign n17254 = n17253 ^ n17245 ;
  assign n17167 = n17088 ^ n17003 ;
  assign n17168 = n17089 & n17167 ;
  assign n17169 = n17168 ^ n17088 ;
  assign n17255 = n17254 ^ n17169 ;
  assign n17264 = n17263 ^ n17255 ;
  assign n17164 = n17102 ^ n17098 ;
  assign n17165 = ~n17099 & ~n17164 ;
  assign n17166 = n17165 ^ n17102 ;
  assign n17265 = n17264 ^ n17166 ;
  assign n17274 = n17273 ^ n17265 ;
  assign n17161 = n17115 ^ n17111 ;
  assign n17162 = n17112 & ~n17161 ;
  assign n17163 = n17162 ^ n17115 ;
  assign n17275 = n17274 ^ n17163 ;
  assign n17284 = n17283 ^ n17275 ;
  assign n17288 = n17287 ^ n17284 ;
  assign n17297 = n17296 ^ n17288 ;
  assign n17301 = n17300 ^ n17297 ;
  assign n17308 = n17307 ^ n17301 ;
  assign n17313 = n17312 ^ n17308 ;
  assign n17159 = n17149 ^ n16997 ;
  assign n17160 = ~n17157 & n17159 ;
  assign n17314 = n17313 ^ n17160 ;
  assign n17480 = n17308 ^ n17156 ;
  assign n17481 = ~n17310 & n17480 ;
  assign n17478 = n17308 ^ n17149 ;
  assign n17479 = ~n17309 & ~n17478 ;
  assign n17482 = n17481 ^ n17479 ;
  assign n17483 = n16997 & n17482 ;
  assign n17484 = n17308 ^ n17148 ;
  assign n17485 = n17484 ^ n17308 ;
  assign n17486 = n17308 ^ n17140 ;
  assign n17487 = n17486 ^ n17308 ;
  assign n17488 = n17485 & ~n17487 ;
  assign n17489 = n17488 ^ n17308 ;
  assign n17497 = n17487 ^ n17485 ;
  assign n17498 = n17497 ^ n17308 ;
  assign n17491 = n17308 ^ n17155 ;
  assign n17490 = n17308 ^ n17152 ;
  assign n17492 = n17491 ^ n17490 ;
  assign n17493 = n17491 ^ n17486 ;
  assign n17494 = n17493 ^ n17484 ;
  assign n17495 = n17494 ^ n17308 ;
  assign n17496 = ~n17492 & n17495 ;
  assign n17499 = n17498 ^ n17496 ;
  assign n17500 = n17489 & ~n17499 ;
  assign n17501 = n17500 ^ n17308 ;
  assign n17504 = ~n17483 & ~n17501 ;
  assign n17469 = x124 & n3375 ;
  assign n17468 = x126 & n3378 ;
  assign n17470 = n17469 ^ n17468 ;
  assign n17471 = n17470 ^ x35 ;
  assign n17467 = n3379 & n10441 ;
  assign n17472 = n17471 ^ n17467 ;
  assign n17466 = x125 & n3383 ;
  assign n17473 = n17472 ^ n17466 ;
  assign n17455 = x121 & n3916 ;
  assign n17454 = x123 & n3919 ;
  assign n17456 = n17455 ^ n17454 ;
  assign n17457 = n17456 ^ x38 ;
  assign n17453 = n3920 & ~n9786 ;
  assign n17458 = n17457 ^ n17453 ;
  assign n17452 = x122 & n3924 ;
  assign n17459 = n17458 ^ n17452 ;
  assign n17445 = x118 & n4474 ;
  assign n17444 = x120 & n4471 ;
  assign n17446 = n17445 ^ n17444 ;
  assign n17447 = n17446 ^ x41 ;
  assign n17443 = n4472 & n8891 ;
  assign n17448 = n17447 ^ n17443 ;
  assign n17442 = x119 & n4467 ;
  assign n17449 = n17448 ^ n17442 ;
  assign n17439 = n17263 ^ n17169 ;
  assign n17440 = ~n17255 & n17439 ;
  assign n17431 = x115 & n5094 ;
  assign n17430 = x117 & n5097 ;
  assign n17432 = n17431 ^ n17430 ;
  assign n17433 = n17432 ^ x44 ;
  assign n17429 = n5098 & ~n7850 ;
  assign n17434 = n17433 ^ n17429 ;
  assign n17428 = x116 & n5102 ;
  assign n17435 = n17434 ^ n17428 ;
  assign n17417 = x112 & n5965 ;
  assign n17416 = x114 & n5729 ;
  assign n17418 = n17417 ^ n17416 ;
  assign n17419 = n17418 ^ x47 ;
  assign n17415 = n5730 & ~n7092 ;
  assign n17420 = n17419 ^ n17415 ;
  assign n17414 = x113 & n5736 ;
  assign n17421 = n17420 ^ n17414 ;
  assign n17407 = x109 & n6677 ;
  assign n17406 = x111 & n6428 ;
  assign n17408 = n17407 ^ n17406 ;
  assign n17409 = n17408 ^ x50 ;
  assign n17405 = ~n6360 & n6429 ;
  assign n17410 = n17409 ^ n17405 ;
  assign n17404 = x110 & n6433 ;
  assign n17411 = n17410 ^ n17404 ;
  assign n17400 = n17232 ^ n17226 ;
  assign n17401 = ~n17238 & ~n17400 ;
  assign n17402 = n17401 ^ n17226 ;
  assign n17396 = n5670 & n7175 ;
  assign n17394 = x106 & n7171 ;
  assign n17390 = n17216 ^ n17184 ;
  assign n17391 = ~n17225 & ~n17390 ;
  assign n17392 = n17391 ^ n17216 ;
  assign n17388 = x108 & n7174 ;
  assign n17389 = n17388 ^ x53 ;
  assign n17393 = n17392 ^ n17389 ;
  assign n17395 = n17394 ^ n17393 ;
  assign n17397 = n17396 ^ n17395 ;
  assign n17387 = x107 & n7179 ;
  assign n17398 = n17397 ^ n17387 ;
  assign n17380 = x100 & n8741 ;
  assign n17379 = x102 & n8744 ;
  assign n17381 = n17380 ^ n17379 ;
  assign n17382 = n17381 ^ x59 ;
  assign n17378 = n4410 & n8745 ;
  assign n17383 = n17382 ^ n17378 ;
  assign n17377 = x101 & n8737 ;
  assign n17384 = n17383 ^ n17377 ;
  assign n17371 = x97 & n9632 ;
  assign n17370 = x99 & n9635 ;
  assign n17372 = n17371 ^ n17370 ;
  assign n17373 = n17372 ^ x62 ;
  assign n17369 = n3843 & n9636 ;
  assign n17374 = n17373 ^ n17369 ;
  assign n17368 = x98 & n9628 ;
  assign n17375 = n17374 ^ n17368 ;
  assign n17364 = n17208 ^ n17199 ;
  assign n17365 = ~n17205 & ~n17364 ;
  assign n17366 = n17365 ^ n17208 ;
  assign n17358 = n9948 ^ x95 ;
  assign n17354 = ~x96 & n9948 ;
  assign n17355 = n17354 ^ n17207 ;
  assign n17359 = n17355 ^ n12206 ;
  assign n17360 = n17358 & n17359 ;
  assign n17361 = n17360 ^ n2978 ;
  assign n17356 = x95 & n17355 ;
  assign n17357 = n17356 ^ n17207 ;
  assign n17362 = n17361 ^ n17357 ;
  assign n17363 = n17362 ^ n2978 ;
  assign n17367 = n17366 ^ n17363 ;
  assign n17376 = n17375 ^ n17367 ;
  assign n17385 = n17384 ^ n17376 ;
  assign n17351 = ~n5023 & n7939 ;
  assign n17349 = x103 & n7935 ;
  assign n17345 = n17209 ^ n17187 ;
  assign n17346 = ~n17215 & ~n17345 ;
  assign n17347 = n17346 ^ n17209 ;
  assign n17343 = x105 & n7938 ;
  assign n17344 = n17343 ^ x56 ;
  assign n17348 = n17347 ^ n17344 ;
  assign n17350 = n17349 ^ n17348 ;
  assign n17352 = n17351 ^ n17350 ;
  assign n17342 = x104 & n7931 ;
  assign n17353 = n17352 ^ n17342 ;
  assign n17386 = n17385 ^ n17353 ;
  assign n17399 = n17398 ^ n17386 ;
  assign n17403 = n17402 ^ n17399 ;
  assign n17412 = n17411 ^ n17403 ;
  assign n17339 = n17239 ^ n17175 ;
  assign n17340 = ~n17181 & ~n17339 ;
  assign n17341 = n17340 ^ n17239 ;
  assign n17413 = n17412 ^ n17341 ;
  assign n17422 = n17421 ^ n17413 ;
  assign n17424 = n17422 ^ n17240 ;
  assign n17423 = n17422 ^ n17253 ;
  assign n17425 = n17424 ^ n17423 ;
  assign n17426 = n17245 & ~n17425 ;
  assign n17427 = n17426 ^ n17424 ;
  assign n17436 = n17435 ^ n17427 ;
  assign n17437 = n17436 ^ n17263 ;
  assign n17441 = n17440 ^ n17437 ;
  assign n17450 = n17449 ^ n17441 ;
  assign n17336 = n17273 ^ n17166 ;
  assign n17337 = n17265 & ~n17336 ;
  assign n17338 = n17337 ^ n17273 ;
  assign n17451 = n17450 ^ n17338 ;
  assign n17460 = n17459 ^ n17451 ;
  assign n17461 = n17460 ^ n17283 ;
  assign n17462 = n17461 ^ n17460 ;
  assign n17463 = n17462 ^ n17163 ;
  assign n17464 = ~n17275 & ~n17463 ;
  assign n17465 = n17464 ^ n17461 ;
  assign n17474 = n17473 ^ n17465 ;
  assign n17323 = ~x31 & x127 ;
  assign n17324 = n17323 ^ x32 ;
  assign n17325 = ~n10138 & ~n17324 ;
  assign n17326 = n17325 ^ x32 ;
  assign n17327 = n2738 & ~n17326 ;
  assign n17328 = n2737 ^ x32 ;
  assign n17331 = x127 & n2877 ;
  assign n17332 = ~n17328 & n17331 ;
  assign n17333 = n17332 ^ n17328 ;
  assign n17334 = n17333 ^ n2737 ;
  assign n17335 = ~n17327 & n17334 ;
  assign n17475 = n17474 ^ n17335 ;
  assign n17318 = n17296 ^ n17287 ;
  assign n17319 = ~n17288 & n17318 ;
  assign n17320 = n17319 ^ n17296 ;
  assign n17476 = n17475 ^ n17320 ;
  assign n17315 = n17307 ^ n17300 ;
  assign n17316 = ~n17301 & n17315 ;
  assign n17317 = n17316 ^ n17307 ;
  assign n17477 = n17476 ^ n17317 ;
  assign n17505 = n17504 ^ n17477 ;
  assign n17649 = n17504 ^ n17317 ;
  assign n17650 = n17477 & ~n17649 ;
  assign n17651 = n17650 ^ n17504 ;
  assign n17644 = n17473 ^ n17460 ;
  assign n17645 = ~n17465 & ~n17644 ;
  assign n17646 = n17645 ^ n17460 ;
  assign n17638 = x125 & n3375 ;
  assign n17637 = x127 & n3378 ;
  assign n17639 = n17638 ^ n17637 ;
  assign n17640 = n17639 ^ x35 ;
  assign n17636 = n3379 & n10972 ;
  assign n17641 = n17640 ^ n17636 ;
  assign n17635 = x126 & n3383 ;
  assign n17642 = n17641 ^ n17635 ;
  assign n17628 = x122 & n3916 ;
  assign n17627 = x124 & n3919 ;
  assign n17629 = n17628 ^ n17627 ;
  assign n17630 = n17629 ^ x38 ;
  assign n17626 = n3920 & n10095 ;
  assign n17631 = n17630 ^ n17626 ;
  assign n17625 = x123 & n3924 ;
  assign n17632 = n17631 ^ n17625 ;
  assign n17619 = x119 & n4474 ;
  assign n17618 = x121 & n4471 ;
  assign n17620 = n17619 ^ n17618 ;
  assign n17621 = n17620 ^ x41 ;
  assign n17617 = n4472 & n8962 ;
  assign n17622 = n17621 ^ n17617 ;
  assign n17616 = x120 & n4467 ;
  assign n17623 = n17622 ^ n17616 ;
  assign n17612 = n17449 ^ n17436 ;
  assign n17613 = ~n17441 & ~n17612 ;
  assign n17614 = n17613 ^ n17436 ;
  assign n17606 = x116 & n5094 ;
  assign n17605 = x118 & n5097 ;
  assign n17607 = n17606 ^ n17605 ;
  assign n17608 = n17607 ^ x44 ;
  assign n17604 = n5098 & ~n8123 ;
  assign n17609 = n17608 ^ n17604 ;
  assign n17603 = x117 & n5102 ;
  assign n17610 = n17609 ^ n17603 ;
  assign n17594 = n17421 ^ n17341 ;
  assign n17595 = ~n17413 & ~n17594 ;
  assign n17596 = n17595 ^ n17421 ;
  assign n17592 = x114 & n5736 ;
  assign n17587 = x113 & n5965 ;
  assign n17586 = x115 & n5729 ;
  assign n17588 = n17587 ^ n17586 ;
  assign n17589 = n17588 ^ x47 ;
  assign n17585 = n5730 & ~n7343 ;
  assign n17590 = n17589 ^ n17585 ;
  assign n17577 = ~n17360 & n17366 ;
  assign n17578 = ~n17357 & n17577 ;
  assign n17579 = n17578 ^ n17360 ;
  assign n17570 = x98 & n9632 ;
  assign n17569 = x100 & n9635 ;
  assign n17571 = n17570 ^ n17569 ;
  assign n17572 = n17571 ^ x62 ;
  assign n17568 = n4034 & n9636 ;
  assign n17573 = n17572 ^ n17568 ;
  assign n17567 = x99 & n9628 ;
  assign n17574 = n17573 ^ n17567 ;
  assign n17575 = n17574 ^ x32 ;
  assign n17563 = x97 ^ x95 ;
  assign n17564 = ~n11875 & n17563 ;
  assign n17565 = n17564 ^ n2978 ;
  assign n17566 = n12206 & n17565 ;
  assign n17576 = n17575 ^ n17566 ;
  assign n17580 = n17579 ^ n17576 ;
  assign n17560 = ~n4615 & n8745 ;
  assign n17558 = x101 & n8741 ;
  assign n17554 = n17384 ^ n17375 ;
  assign n17555 = ~n17376 & n17554 ;
  assign n17556 = n17555 ^ n17384 ;
  assign n17552 = x103 & n8744 ;
  assign n17553 = n17552 ^ x59 ;
  assign n17557 = n17556 ^ n17553 ;
  assign n17559 = n17558 ^ n17557 ;
  assign n17561 = n17560 ^ n17559 ;
  assign n17551 = x102 & n8737 ;
  assign n17562 = n17561 ^ n17551 ;
  assign n17581 = n17580 ^ n17562 ;
  assign n17541 = x104 & n7935 ;
  assign n17540 = x106 & n7938 ;
  assign n17542 = n17541 ^ n17540 ;
  assign n17543 = n17542 ^ x56 ;
  assign n17539 = ~n5240 & n7939 ;
  assign n17544 = n17543 ^ n17539 ;
  assign n17538 = x105 & n7931 ;
  assign n17545 = n17544 ^ n17538 ;
  assign n17546 = n17545 ^ n17385 ;
  assign n17547 = n17546 ^ n17347 ;
  assign n17548 = n17547 ^ n17545 ;
  assign n17549 = n17353 & ~n17548 ;
  assign n17550 = n17549 ^ n17546 ;
  assign n17582 = n17581 ^ n17550 ;
  assign n17535 = n17392 ^ n17386 ;
  assign n17536 = n17398 & n17535 ;
  assign n17528 = x107 & n7171 ;
  assign n17527 = x109 & n7174 ;
  assign n17529 = n17528 ^ n17527 ;
  assign n17530 = n17529 ^ x53 ;
  assign n17526 = n5902 & n7175 ;
  assign n17531 = n17530 ^ n17526 ;
  assign n17525 = x108 & n7179 ;
  assign n17532 = n17531 ^ n17525 ;
  assign n17533 = n17532 ^ n17386 ;
  assign n17537 = n17536 ^ n17533 ;
  assign n17583 = n17582 ^ n17537 ;
  assign n17515 = x110 & n6677 ;
  assign n17514 = x112 & n6428 ;
  assign n17516 = n17515 ^ n17514 ;
  assign n17517 = n17516 ^ x50 ;
  assign n17513 = n6429 & ~n6600 ;
  assign n17518 = n17517 ^ n17513 ;
  assign n17512 = x111 & n6433 ;
  assign n17519 = n17518 ^ n17512 ;
  assign n17520 = n17519 ^ n17411 ;
  assign n17521 = n17520 ^ n17402 ;
  assign n17522 = n17521 ^ n17519 ;
  assign n17523 = n17403 & ~n17522 ;
  assign n17524 = n17523 ^ n17520 ;
  assign n17584 = n17583 ^ n17524 ;
  assign n17591 = n17590 ^ n17584 ;
  assign n17593 = n17592 ^ n17591 ;
  assign n17597 = n17596 ^ n17593 ;
  assign n17599 = n17597 ^ n17422 ;
  assign n17598 = n17597 ^ n17435 ;
  assign n17600 = n17599 ^ n17598 ;
  assign n17601 = ~n17427 & n17600 ;
  assign n17602 = n17601 ^ n17599 ;
  assign n17611 = n17610 ^ n17602 ;
  assign n17615 = n17614 ^ n17611 ;
  assign n17624 = n17623 ^ n17615 ;
  assign n17633 = n17632 ^ n17624 ;
  assign n17509 = n17459 ^ n17338 ;
  assign n17510 = n17451 & n17509 ;
  assign n17511 = n17510 ^ n17459 ;
  assign n17634 = n17633 ^ n17511 ;
  assign n17643 = n17642 ^ n17634 ;
  assign n17647 = n17646 ^ n17643 ;
  assign n17506 = n17474 ^ n17320 ;
  assign n17507 = ~n17475 & ~n17506 ;
  assign n17508 = n17507 ^ n17474 ;
  assign n17648 = n17647 ^ n17508 ;
  assign n17652 = n17651 ^ n17648 ;
  assign n17799 = n17651 ^ n17508 ;
  assign n17800 = ~n17648 & n17799 ;
  assign n17801 = n17800 ^ n17651 ;
  assign n17788 = n17632 ^ n17511 ;
  assign n17789 = n17633 & n17788 ;
  assign n17790 = n17789 ^ n17632 ;
  assign n17785 = n17646 ^ n17642 ;
  assign n17786 = ~n17643 & ~n17785 ;
  assign n17787 = n17786 ^ n17646 ;
  assign n17795 = n17790 ^ n17787 ;
  assign n17791 = n17787 & ~n17790 ;
  assign n17796 = n17795 ^ n17791 ;
  assign n17780 = n3379 & n10139 ;
  assign n17779 = x126 & n3375 ;
  assign n17781 = n17780 ^ n17779 ;
  assign n17782 = n17781 ^ x35 ;
  assign n17778 = x127 & n3383 ;
  assign n17783 = n17782 ^ n17778 ;
  assign n17772 = x123 & n3916 ;
  assign n17771 = x125 & n3919 ;
  assign n17773 = n17772 ^ n17771 ;
  assign n17774 = n17773 ^ x38 ;
  assign n17770 = n3920 & n10400 ;
  assign n17775 = n17774 ^ n17770 ;
  assign n17769 = x124 & n3924 ;
  assign n17776 = n17775 ^ n17769 ;
  assign n17758 = x120 & n4474 ;
  assign n17757 = x122 & n4471 ;
  assign n17759 = n17758 ^ n17757 ;
  assign n17760 = n17759 ^ x41 ;
  assign n17756 = n4472 & ~n9247 ;
  assign n17761 = n17760 ^ n17756 ;
  assign n17755 = x121 & n4467 ;
  assign n17762 = n17761 ^ n17755 ;
  assign n17751 = n17610 ^ n17597 ;
  assign n17752 = ~n17602 & ~n17751 ;
  assign n17753 = n17752 ^ n17597 ;
  assign n17745 = x117 & n5094 ;
  assign n17744 = x119 & n5097 ;
  assign n17746 = n17745 ^ n17744 ;
  assign n17747 = n17746 ^ x44 ;
  assign n17743 = n5098 & n8394 ;
  assign n17748 = n17747 ^ n17743 ;
  assign n17742 = x118 & n5102 ;
  assign n17749 = n17748 ^ n17742 ;
  assign n17730 = x114 & n5965 ;
  assign n17729 = x116 & n5729 ;
  assign n17731 = n17730 ^ n17729 ;
  assign n17732 = n17731 ^ x47 ;
  assign n17728 = n5730 & ~n7588 ;
  assign n17733 = n17732 ^ n17728 ;
  assign n17727 = x115 & n5736 ;
  assign n17734 = n17733 ^ n17727 ;
  assign n17721 = x103 & n8737 ;
  assign n17719 = ~n4814 & n8745 ;
  assign n17715 = x102 & n8741 ;
  assign n17714 = x104 & n8744 ;
  assign n17716 = n17715 ^ n17714 ;
  assign n17717 = n17716 ^ x59 ;
  assign n17711 = x97 & n11875 ;
  assign n17710 = x98 & n9948 ;
  assign n17712 = n17711 ^ n17710 ;
  assign n17707 = n4215 & n9636 ;
  assign n17705 = x99 & n9632 ;
  assign n17698 = x96 ^ x32 ;
  assign n17701 = n17565 & ~n17698 ;
  assign n17702 = n17701 ^ x96 ;
  assign n17703 = n12206 & n17702 ;
  assign n17696 = x101 & n9635 ;
  assign n17697 = n17696 ^ x62 ;
  assign n17704 = n17703 ^ n17697 ;
  assign n17706 = n17705 ^ n17704 ;
  assign n17708 = n17707 ^ n17706 ;
  assign n17695 = x100 & n9628 ;
  assign n17709 = n17708 ^ n17695 ;
  assign n17713 = n17712 ^ n17709 ;
  assign n17718 = n17717 ^ n17713 ;
  assign n17720 = n17719 ^ n17718 ;
  assign n17722 = n17721 ^ n17720 ;
  assign n17692 = n17579 ^ n17574 ;
  assign n17693 = n17576 & ~n17692 ;
  assign n17694 = n17693 ^ n17579 ;
  assign n17723 = n17722 ^ n17694 ;
  assign n17689 = ~n5448 & n7939 ;
  assign n17687 = x105 & n7935 ;
  assign n17683 = n17580 ^ n17556 ;
  assign n17684 = ~n17562 & n17683 ;
  assign n17685 = n17684 ^ n17580 ;
  assign n17681 = x107 & n7938 ;
  assign n17682 = n17681 ^ x56 ;
  assign n17686 = n17685 ^ n17682 ;
  assign n17688 = n17687 ^ n17686 ;
  assign n17690 = n17689 ^ n17688 ;
  assign n17680 = x106 & n7931 ;
  assign n17691 = n17690 ^ n17680 ;
  assign n17724 = n17723 ^ n17691 ;
  assign n17677 = n6129 & n7175 ;
  assign n17675 = x108 & n7171 ;
  assign n17671 = n17581 ^ n17545 ;
  assign n17672 = n17550 & n17671 ;
  assign n17673 = n17672 ^ n17545 ;
  assign n17669 = x110 & n7174 ;
  assign n17670 = n17669 ^ x53 ;
  assign n17674 = n17673 ^ n17670 ;
  assign n17676 = n17675 ^ n17674 ;
  assign n17678 = n17677 ^ n17676 ;
  assign n17668 = x109 & n7179 ;
  assign n17679 = n17678 ^ n17668 ;
  assign n17725 = n17724 ^ n17679 ;
  assign n17665 = n6429 & ~n6839 ;
  assign n17663 = x111 & n6677 ;
  assign n17659 = n17582 ^ n17532 ;
  assign n17660 = ~n17537 & n17659 ;
  assign n17661 = n17660 ^ n17532 ;
  assign n17657 = x113 & n6428 ;
  assign n17658 = n17657 ^ x50 ;
  assign n17662 = n17661 ^ n17658 ;
  assign n17664 = n17663 ^ n17662 ;
  assign n17666 = n17665 ^ n17664 ;
  assign n17656 = x112 & n6433 ;
  assign n17667 = n17666 ^ n17656 ;
  assign n17726 = n17725 ^ n17667 ;
  assign n17735 = n17734 ^ n17726 ;
  assign n17653 = n17583 ^ n17519 ;
  assign n17654 = n17524 & ~n17653 ;
  assign n17655 = n17654 ^ n17519 ;
  assign n17736 = n17735 ^ n17655 ;
  assign n17738 = n17736 ^ n17596 ;
  assign n17737 = n17736 ^ n17584 ;
  assign n17739 = n17738 ^ n17737 ;
  assign n17740 = ~n17593 & ~n17739 ;
  assign n17741 = n17740 ^ n17737 ;
  assign n17750 = n17749 ^ n17741 ;
  assign n17754 = n17753 ^ n17750 ;
  assign n17763 = n17762 ^ n17754 ;
  assign n17764 = n17763 ^ n17623 ;
  assign n17765 = n17764 ^ n17614 ;
  assign n17766 = n17765 ^ n17763 ;
  assign n17767 = ~n17615 & ~n17766 ;
  assign n17768 = n17767 ^ n17764 ;
  assign n17777 = n17776 ^ n17768 ;
  assign n17793 = n17783 ^ n17777 ;
  assign n17784 = n17777 & n17783 ;
  assign n17794 = n17793 ^ n17784 ;
  assign n17797 = n17796 ^ n17794 ;
  assign n17792 = n17791 ^ n17784 ;
  assign n17798 = n17797 ^ n17792 ;
  assign n17802 = n17801 ^ n17798 ;
  assign n17936 = x127 & n3374 ;
  assign n17937 = n17936 ^ n3372 ;
  assign n17942 = n3041 & n11265 ;
  assign n17943 = n17942 ^ n17936 ;
  assign n17944 = n17937 & ~n17943 ;
  assign n17945 = n17944 ^ x34 ;
  assign n17925 = x124 & n3916 ;
  assign n17924 = x126 & n3919 ;
  assign n17926 = n17925 ^ n17924 ;
  assign n17927 = n17926 ^ x38 ;
  assign n17923 = n3920 & n10441 ;
  assign n17928 = n17927 ^ n17923 ;
  assign n17922 = x125 & n3924 ;
  assign n17929 = n17928 ^ n17922 ;
  assign n17911 = x121 & n4474 ;
  assign n17910 = x123 & n4471 ;
  assign n17912 = n17911 ^ n17910 ;
  assign n17913 = n17912 ^ x41 ;
  assign n17909 = n4472 & ~n9786 ;
  assign n17914 = n17913 ^ n17909 ;
  assign n17908 = x122 & n4467 ;
  assign n17915 = n17914 ^ n17908 ;
  assign n17904 = n17749 ^ n17736 ;
  assign n17905 = ~n17741 & n17904 ;
  assign n17906 = n17905 ^ n17736 ;
  assign n17898 = x118 & n5094 ;
  assign n17897 = x120 & n5097 ;
  assign n17899 = n17898 ^ n17897 ;
  assign n17900 = n17899 ^ x44 ;
  assign n17896 = n5098 & n8891 ;
  assign n17901 = n17900 ^ n17896 ;
  assign n17895 = x119 & n5102 ;
  assign n17902 = n17901 ^ n17895 ;
  assign n17888 = x115 & n5965 ;
  assign n17887 = x117 & n5729 ;
  assign n17889 = n17888 ^ n17887 ;
  assign n17890 = n17889 ^ x47 ;
  assign n17886 = n5730 & ~n7850 ;
  assign n17891 = n17890 ^ n17886 ;
  assign n17885 = x116 & n5736 ;
  assign n17892 = n17891 ^ n17885 ;
  assign n17871 = x103 & n8741 ;
  assign n17870 = x105 & n8744 ;
  assign n17872 = n17871 ^ n17870 ;
  assign n17873 = n17872 ^ x59 ;
  assign n17869 = ~n5023 & n8745 ;
  assign n17874 = n17873 ^ n17869 ;
  assign n17868 = x104 & n8737 ;
  assign n17875 = n17874 ^ n17868 ;
  assign n17866 = x101 & n9628 ;
  assign n17858 = n17712 ^ n17703 ;
  assign n17859 = ~n17709 & ~n17858 ;
  assign n17860 = n17859 ^ n17712 ;
  assign n17852 = n9948 ^ x98 ;
  assign n17848 = ~x99 & n9948 ;
  assign n17849 = n17848 ^ n17711 ;
  assign n17853 = n17849 ^ n12206 ;
  assign n17854 = n17852 & n17853 ;
  assign n17855 = n17854 ^ n3475 ;
  assign n17850 = x98 & n17849 ;
  assign n17851 = n17850 ^ n17711 ;
  assign n17856 = n17855 ^ n17851 ;
  assign n17857 = n17856 ^ n3475 ;
  assign n17861 = n17860 ^ n17857 ;
  assign n17862 = n17861 ^ x62 ;
  assign n17847 = x100 & n9632 ;
  assign n17863 = n17862 ^ n17847 ;
  assign n17846 = x102 & n9635 ;
  assign n17864 = n17863 ^ n17846 ;
  assign n17845 = n4410 & n9636 ;
  assign n17865 = n17864 ^ n17845 ;
  assign n17867 = n17866 ^ n17865 ;
  assign n17876 = n17875 ^ n17867 ;
  assign n17842 = n5670 & n7939 ;
  assign n17840 = x106 & n7935 ;
  assign n17836 = n17713 ^ n17694 ;
  assign n17837 = ~n17722 & n17836 ;
  assign n17838 = n17837 ^ n17713 ;
  assign n17834 = x108 & n7938 ;
  assign n17835 = n17834 ^ x56 ;
  assign n17839 = n17838 ^ n17835 ;
  assign n17841 = n17840 ^ n17839 ;
  assign n17843 = n17842 ^ n17841 ;
  assign n17833 = x107 & n7931 ;
  assign n17844 = n17843 ^ n17833 ;
  assign n17877 = n17876 ^ n17844 ;
  assign n17831 = x110 & n7179 ;
  assign n17829 = ~n6360 & n7175 ;
  assign n17827 = x109 & n7171 ;
  assign n17823 = n17723 ^ n17685 ;
  assign n17824 = ~n17691 & n17823 ;
  assign n17825 = n17824 ^ n17723 ;
  assign n17821 = x111 & n7174 ;
  assign n17822 = n17821 ^ x53 ;
  assign n17826 = n17825 ^ n17822 ;
  assign n17828 = n17827 ^ n17826 ;
  assign n17830 = n17829 ^ n17828 ;
  assign n17832 = n17831 ^ n17830 ;
  assign n17878 = n17877 ^ n17832 ;
  assign n17819 = x113 & n6433 ;
  assign n17817 = n6429 & ~n7092 ;
  assign n17815 = x112 & n6677 ;
  assign n17811 = n17724 ^ n17673 ;
  assign n17812 = ~n17679 & n17811 ;
  assign n17813 = n17812 ^ n17724 ;
  assign n17809 = x114 & n6428 ;
  assign n17810 = n17809 ^ x50 ;
  assign n17814 = n17813 ^ n17810 ;
  assign n17816 = n17815 ^ n17814 ;
  assign n17818 = n17817 ^ n17816 ;
  assign n17820 = n17819 ^ n17818 ;
  assign n17879 = n17878 ^ n17820 ;
  assign n17880 = n17879 ^ n17725 ;
  assign n17881 = n17880 ^ n17661 ;
  assign n17882 = n17881 ^ n17879 ;
  assign n17883 = ~n17667 & n17882 ;
  assign n17884 = n17883 ^ n17880 ;
  assign n17893 = n17892 ^ n17884 ;
  assign n17806 = n17734 ^ n17655 ;
  assign n17807 = n17735 & n17806 ;
  assign n17808 = n17807 ^ n17734 ;
  assign n17894 = n17893 ^ n17808 ;
  assign n17903 = n17902 ^ n17894 ;
  assign n17907 = n17906 ^ n17903 ;
  assign n17916 = n17915 ^ n17907 ;
  assign n17917 = n17916 ^ n17762 ;
  assign n17918 = n17917 ^ n17753 ;
  assign n17919 = n17918 ^ n17916 ;
  assign n17920 = ~n17754 & ~n17919 ;
  assign n17921 = n17920 ^ n17917 ;
  assign n17930 = n17929 ^ n17921 ;
  assign n17932 = n17930 ^ n17763 ;
  assign n17931 = n17930 ^ n17776 ;
  assign n17933 = n17932 ^ n17931 ;
  assign n17934 = n17768 & n17933 ;
  assign n17935 = n17934 ^ n17932 ;
  assign n17946 = n17945 ^ n17935 ;
  assign n17947 = n17946 ^ n17792 ;
  assign n17803 = n17801 ^ n17787 ;
  assign n17804 = n17803 ^ n17790 ;
  assign n17805 = ~n17798 & n17804 ;
  assign n17948 = n17947 ^ n17805 ;
  assign n18078 = n17796 ^ n17791 ;
  assign n18079 = n18078 ^ n17946 ;
  assign n18080 = n18079 ^ n17796 ;
  assign n18081 = n18080 ^ n17946 ;
  assign n18082 = n18081 ^ n18080 ;
  assign n18085 = n17796 & ~n18082 ;
  assign n18091 = n18085 ^ n17796 ;
  assign n18083 = n18082 ^ n18080 ;
  assign n18087 = n18085 ^ n18083 ;
  assign n18088 = ~n17777 & ~n18087 ;
  assign n18089 = n18088 ^ n18080 ;
  assign n18090 = ~n17793 & n18089 ;
  assign n18092 = n18091 ^ n18090 ;
  assign n18093 = n18092 ^ n18081 ;
  assign n18094 = n17801 & n18093 ;
  assign n18095 = n17946 ^ n17777 ;
  assign n18096 = n18095 ^ n17946 ;
  assign n18097 = n17946 ^ n17783 ;
  assign n18098 = n18097 ^ n17946 ;
  assign n18099 = ~n18096 & ~n18098 ;
  assign n18100 = n18099 ^ n17946 ;
  assign n18108 = n18098 ^ n18096 ;
  assign n18109 = n18108 ^ n17946 ;
  assign n18102 = n17946 ^ n17787 ;
  assign n18101 = n17946 ^ n17790 ;
  assign n18103 = n18102 ^ n18101 ;
  assign n18104 = n18102 ^ n18095 ;
  assign n18105 = n18104 ^ n18097 ;
  assign n18106 = n18105 ^ n17946 ;
  assign n18107 = n18103 & n18106 ;
  assign n18110 = n18109 ^ n18107 ;
  assign n18111 = n18100 & n18110 ;
  assign n18112 = n18111 ^ n17946 ;
  assign n18115 = ~n18094 & ~n18112 ;
  assign n18074 = n17945 ^ n17930 ;
  assign n18075 = ~n17935 & ~n18074 ;
  assign n18076 = n18075 ^ n17930 ;
  assign n18070 = n17929 ^ n17916 ;
  assign n18071 = ~n17921 & ~n18070 ;
  assign n18072 = n18071 ^ n17916 ;
  assign n18064 = x125 & n3916 ;
  assign n18063 = x127 & n3919 ;
  assign n18065 = n18064 ^ n18063 ;
  assign n18066 = n18065 ^ x38 ;
  assign n18062 = n3920 & n10972 ;
  assign n18067 = n18066 ^ n18062 ;
  assign n18061 = x126 & n3924 ;
  assign n18068 = n18067 ^ n18061 ;
  assign n18054 = x122 & n4474 ;
  assign n18053 = x124 & n4471 ;
  assign n18055 = n18054 ^ n18053 ;
  assign n18056 = n18055 ^ x41 ;
  assign n18052 = n4472 & n10095 ;
  assign n18057 = n18056 ^ n18052 ;
  assign n18051 = x123 & n4467 ;
  assign n18058 = n18057 ^ n18051 ;
  assign n18044 = x119 & n5094 ;
  assign n18043 = x121 & n5097 ;
  assign n18045 = n18044 ^ n18043 ;
  assign n18046 = n18045 ^ x44 ;
  assign n18042 = n5098 & n8962 ;
  assign n18047 = n18046 ^ n18042 ;
  assign n18041 = x120 & n5102 ;
  assign n18048 = n18047 ^ n18041 ;
  assign n18037 = n17892 ^ n17879 ;
  assign n18038 = ~n17884 & ~n18037 ;
  assign n18039 = n18038 ^ n17879 ;
  assign n18031 = x116 & n5965 ;
  assign n18030 = x118 & n5729 ;
  assign n18032 = n18031 ^ n18030 ;
  assign n18033 = n18032 ^ x47 ;
  assign n18029 = n5730 & ~n8123 ;
  assign n18034 = n18033 ^ n18029 ;
  assign n18028 = x117 & n5736 ;
  assign n18035 = n18034 ^ n18028 ;
  assign n18022 = x113 & n6677 ;
  assign n18021 = x115 & n6428 ;
  assign n18023 = n18022 ^ n18021 ;
  assign n18024 = n18023 ^ x50 ;
  assign n18020 = n6429 & ~n7343 ;
  assign n18025 = n18024 ^ n18020 ;
  assign n18019 = x114 & n6433 ;
  assign n18026 = n18025 ^ n18019 ;
  assign n18007 = x110 & n7171 ;
  assign n18006 = x112 & n7174 ;
  assign n18008 = n18007 ^ n18006 ;
  assign n18009 = n18008 ^ x53 ;
  assign n18005 = ~n6600 & n7175 ;
  assign n18010 = n18009 ^ n18005 ;
  assign n18004 = x111 & n7179 ;
  assign n18011 = n18010 ^ n18004 ;
  assign n17994 = x101 & n9632 ;
  assign n17993 = x103 & n9635 ;
  assign n17995 = n17994 ^ n17993 ;
  assign n17996 = n17995 ^ x62 ;
  assign n17992 = ~n4615 & n9636 ;
  assign n17997 = n17996 ^ n17992 ;
  assign n17991 = x102 & n9628 ;
  assign n17998 = n17997 ^ n17991 ;
  assign n17999 = n17998 ^ x35 ;
  assign n17987 = x100 ^ x98 ;
  assign n17988 = ~n11875 & n17987 ;
  assign n17989 = n17988 ^ n3475 ;
  assign n17990 = n12206 & n17989 ;
  assign n18000 = n17999 ^ n17990 ;
  assign n17984 = ~n17854 & n17860 ;
  assign n17985 = ~n17851 & n17984 ;
  assign n17986 = n17985 ^ n17854 ;
  assign n18001 = n18000 ^ n17986 ;
  assign n17974 = x104 & n8741 ;
  assign n17973 = x106 & n8744 ;
  assign n17975 = n17974 ^ n17973 ;
  assign n17976 = n17975 ^ x59 ;
  assign n17972 = ~n5240 & n8745 ;
  assign n17977 = n17976 ^ n17972 ;
  assign n17971 = x105 & n8737 ;
  assign n17978 = n17977 ^ n17971 ;
  assign n17979 = n17978 ^ n17875 ;
  assign n17980 = n17979 ^ n17861 ;
  assign n17981 = n17980 ^ n17978 ;
  assign n17982 = ~n17867 & n17981 ;
  assign n17983 = n17982 ^ n17979 ;
  assign n18002 = n18001 ^ n17983 ;
  assign n17961 = x107 & n7935 ;
  assign n17960 = x109 & n7938 ;
  assign n17962 = n17961 ^ n17960 ;
  assign n17963 = n17962 ^ x56 ;
  assign n17959 = n5902 & n7939 ;
  assign n17964 = n17963 ^ n17959 ;
  assign n17958 = x108 & n7931 ;
  assign n17965 = n17964 ^ n17958 ;
  assign n17966 = n17965 ^ n17876 ;
  assign n17967 = n17966 ^ n17838 ;
  assign n17968 = n17967 ^ n17965 ;
  assign n17969 = n17844 & ~n17968 ;
  assign n17970 = n17969 ^ n17966 ;
  assign n18003 = n18002 ^ n17970 ;
  assign n18012 = n18011 ^ n18003 ;
  assign n17955 = n17877 ^ n17825 ;
  assign n17956 = ~n17832 & ~n17955 ;
  assign n17957 = n17956 ^ n17877 ;
  assign n18013 = n18012 ^ n17957 ;
  assign n18015 = n18013 ^ n17878 ;
  assign n18014 = n18013 ^ n17813 ;
  assign n18016 = n18015 ^ n18014 ;
  assign n18017 = ~n17820 & ~n18016 ;
  assign n18018 = n18017 ^ n18015 ;
  assign n18027 = n18026 ^ n18018 ;
  assign n18036 = n18035 ^ n18027 ;
  assign n18040 = n18039 ^ n18036 ;
  assign n18049 = n18048 ^ n18040 ;
  assign n17952 = n17902 ^ n17808 ;
  assign n17953 = n17894 & n17952 ;
  assign n17954 = n17953 ^ n17902 ;
  assign n18050 = n18049 ^ n17954 ;
  assign n18059 = n18058 ^ n18050 ;
  assign n17949 = n17915 ^ n17906 ;
  assign n17950 = n17907 & n17949 ;
  assign n17951 = n17950 ^ n17915 ;
  assign n18060 = n18059 ^ n17951 ;
  assign n18069 = n18068 ^ n18060 ;
  assign n18073 = n18072 ^ n18069 ;
  assign n18077 = n18076 ^ n18073 ;
  assign n18116 = n18115 ^ n18077 ;
  assign n18241 = n3920 & n10139 ;
  assign n18240 = x126 & n3916 ;
  assign n18242 = n18241 ^ n18240 ;
  assign n18243 = n18242 ^ x38 ;
  assign n18239 = x127 & n3924 ;
  assign n18244 = n18243 ^ n18239 ;
  assign n18232 = x123 & n4474 ;
  assign n18231 = x125 & n4471 ;
  assign n18233 = n18232 ^ n18231 ;
  assign n18234 = n18233 ^ x41 ;
  assign n18230 = n4472 & n10400 ;
  assign n18235 = n18234 ^ n18230 ;
  assign n18229 = x124 & n4467 ;
  assign n18236 = n18235 ^ n18229 ;
  assign n18222 = x120 & n5094 ;
  assign n18221 = x122 & n5097 ;
  assign n18223 = n18222 ^ n18221 ;
  assign n18224 = n18223 ^ x44 ;
  assign n18220 = n5098 & ~n9247 ;
  assign n18225 = n18224 ^ n18220 ;
  assign n18219 = x121 & n5102 ;
  assign n18226 = n18225 ^ n18219 ;
  assign n18212 = x117 & n5965 ;
  assign n18211 = x119 & n5729 ;
  assign n18213 = n18212 ^ n18211 ;
  assign n18214 = n18213 ^ x47 ;
  assign n18210 = n5730 & n8394 ;
  assign n18215 = n18214 ^ n18210 ;
  assign n18209 = x118 & n5736 ;
  assign n18216 = n18215 ^ n18209 ;
  assign n18194 = x102 & n9632 ;
  assign n18193 = x104 & n9635 ;
  assign n18195 = n18194 ^ n18193 ;
  assign n18196 = n18195 ^ x62 ;
  assign n18192 = ~n4814 & n9636 ;
  assign n18197 = n18196 ^ n18192 ;
  assign n18191 = x103 & n9628 ;
  assign n18198 = n18197 ^ n18191 ;
  assign n18188 = x100 & n11875 ;
  assign n18187 = x101 & n9948 ;
  assign n18189 = n18188 ^ n18187 ;
  assign n18181 = x99 ^ x35 ;
  assign n18184 = n17989 & ~n18181 ;
  assign n18185 = n18184 ^ x99 ;
  assign n18186 = n12206 & n18185 ;
  assign n18190 = n18189 ^ n18186 ;
  assign n18199 = n18198 ^ n18190 ;
  assign n18179 = x106 & n8737 ;
  assign n18177 = ~n5448 & n8745 ;
  assign n18175 = x105 & n8741 ;
  assign n18171 = n17998 ^ n17986 ;
  assign n18172 = ~n18000 & ~n18171 ;
  assign n18173 = n18172 ^ n17998 ;
  assign n18169 = x107 & n8744 ;
  assign n18170 = n18169 ^ x59 ;
  assign n18174 = n18173 ^ n18170 ;
  assign n18176 = n18175 ^ n18174 ;
  assign n18178 = n18177 ^ n18176 ;
  assign n18180 = n18179 ^ n18178 ;
  assign n18200 = n18199 ^ n18180 ;
  assign n18166 = n6129 & n7939 ;
  assign n18164 = x108 & n7935 ;
  assign n18160 = n18001 ^ n17978 ;
  assign n18161 = n17983 & n18160 ;
  assign n18162 = n18161 ^ n17978 ;
  assign n18158 = x110 & n7938 ;
  assign n18159 = n18158 ^ x56 ;
  assign n18163 = n18162 ^ n18159 ;
  assign n18165 = n18164 ^ n18163 ;
  assign n18167 = n18166 ^ n18165 ;
  assign n18157 = x109 & n7931 ;
  assign n18168 = n18167 ^ n18157 ;
  assign n18201 = n18200 ^ n18168 ;
  assign n18154 = ~n6839 & n7175 ;
  assign n18152 = x111 & n7171 ;
  assign n18148 = n18002 ^ n17965 ;
  assign n18149 = n17970 & n18148 ;
  assign n18150 = n18149 ^ n17965 ;
  assign n18146 = x113 & n7174 ;
  assign n18147 = n18146 ^ x53 ;
  assign n18151 = n18150 ^ n18147 ;
  assign n18153 = n18152 ^ n18151 ;
  assign n18155 = n18154 ^ n18153 ;
  assign n18145 = x112 & n7179 ;
  assign n18156 = n18155 ^ n18145 ;
  assign n18202 = n18201 ^ n18156 ;
  assign n18142 = n18011 ^ n17957 ;
  assign n18143 = n18012 & ~n18142 ;
  assign n18135 = x114 & n6677 ;
  assign n18134 = x116 & n6428 ;
  assign n18136 = n18135 ^ n18134 ;
  assign n18137 = n18136 ^ x50 ;
  assign n18133 = n6429 & ~n7588 ;
  assign n18138 = n18137 ^ n18133 ;
  assign n18132 = x115 & n6433 ;
  assign n18139 = n18138 ^ n18132 ;
  assign n18140 = n18139 ^ n18011 ;
  assign n18144 = n18143 ^ n18140 ;
  assign n18203 = n18202 ^ n18144 ;
  assign n18205 = n18203 ^ n18013 ;
  assign n18204 = n18203 ^ n18026 ;
  assign n18206 = n18205 ^ n18204 ;
  assign n18207 = n18018 & ~n18206 ;
  assign n18208 = n18207 ^ n18205 ;
  assign n18217 = n18216 ^ n18208 ;
  assign n18129 = n18039 ^ n18035 ;
  assign n18130 = ~n18036 & ~n18129 ;
  assign n18131 = n18130 ^ n18039 ;
  assign n18218 = n18217 ^ n18131 ;
  assign n18227 = n18226 ^ n18218 ;
  assign n18126 = n18048 ^ n17954 ;
  assign n18127 = ~n18049 & n18126 ;
  assign n18128 = n18127 ^ n18048 ;
  assign n18228 = n18227 ^ n18128 ;
  assign n18237 = n18236 ^ n18228 ;
  assign n18123 = n18058 ^ n17951 ;
  assign n18124 = ~n18059 & n18123 ;
  assign n18125 = n18124 ^ n18058 ;
  assign n18238 = n18237 ^ n18125 ;
  assign n18245 = n18244 ^ n18238 ;
  assign n18120 = n18072 ^ n18068 ;
  assign n18121 = n18069 & ~n18120 ;
  assign n18122 = n18121 ^ n18072 ;
  assign n18246 = n18245 ^ n18122 ;
  assign n18117 = n18115 ^ n18076 ;
  assign n18118 = n18077 & ~n18117 ;
  assign n18119 = n18118 ^ n18115 ;
  assign n18247 = n18246 ^ n18119 ;
  assign n18368 = x127 & n3915 ;
  assign n18369 = n18368 ^ n3913 ;
  assign n18374 = n3532 & n11265 ;
  assign n18375 = n18374 ^ n18368 ;
  assign n18376 = n18369 & ~n18375 ;
  assign n18377 = n18376 ^ x37 ;
  assign n18357 = x124 & n4474 ;
  assign n18356 = x126 & n4471 ;
  assign n18358 = n18357 ^ n18356 ;
  assign n18359 = n18358 ^ x41 ;
  assign n18355 = n4472 & n10441 ;
  assign n18360 = n18359 ^ n18355 ;
  assign n18354 = x125 & n4467 ;
  assign n18361 = n18360 ^ n18354 ;
  assign n18347 = x121 & n5094 ;
  assign n18346 = x123 & n5097 ;
  assign n18348 = n18347 ^ n18346 ;
  assign n18349 = n18348 ^ x44 ;
  assign n18345 = n5098 & ~n9786 ;
  assign n18350 = n18349 ^ n18345 ;
  assign n18344 = x122 & n5102 ;
  assign n18351 = n18350 ^ n18344 ;
  assign n18340 = n18216 ^ n18203 ;
  assign n18341 = n18208 & ~n18340 ;
  assign n18342 = n18341 ^ n18203 ;
  assign n18334 = x118 & n5965 ;
  assign n18333 = x120 & n5729 ;
  assign n18335 = n18334 ^ n18333 ;
  assign n18336 = n18335 ^ x47 ;
  assign n18332 = n5730 & n8891 ;
  assign n18337 = n18336 ^ n18332 ;
  assign n18331 = x119 & n5736 ;
  assign n18338 = n18337 ^ n18331 ;
  assign n18319 = x115 & n6677 ;
  assign n18318 = x117 & n6428 ;
  assign n18320 = n18319 ^ n18318 ;
  assign n18321 = n18320 ^ x50 ;
  assign n18317 = n6429 & ~n7850 ;
  assign n18322 = n18321 ^ n18317 ;
  assign n18316 = x116 & n6433 ;
  assign n18323 = n18322 ^ n18316 ;
  assign n18310 = x112 & n7171 ;
  assign n18309 = x114 & n7174 ;
  assign n18311 = n18310 ^ n18309 ;
  assign n18312 = n18311 ^ x53 ;
  assign n18308 = ~n7092 & n7175 ;
  assign n18313 = n18312 ^ n18308 ;
  assign n18307 = x113 & n7179 ;
  assign n18314 = n18313 ^ n18307 ;
  assign n18299 = x103 & n9632 ;
  assign n18298 = x105 & n9635 ;
  assign n18300 = n18299 ^ n18298 ;
  assign n18301 = n18300 ^ x62 ;
  assign n18297 = ~n5023 & n9636 ;
  assign n18302 = n18301 ^ n18297 ;
  assign n18296 = x104 & n9628 ;
  assign n18303 = n18302 ^ n18296 ;
  assign n18290 = x106 & n8741 ;
  assign n18289 = x108 & n8744 ;
  assign n18291 = n18290 ^ n18289 ;
  assign n18292 = n18291 ^ x59 ;
  assign n18288 = n5670 & n8745 ;
  assign n18293 = n18292 ^ n18288 ;
  assign n18287 = x107 & n8737 ;
  assign n18294 = n18293 ^ n18287 ;
  assign n18282 = x63 & n3818 ;
  assign n4014 = x102 ^ x101 ;
  assign n18283 = n18282 ^ n4014 ;
  assign n18284 = ~n9948 & n18283 ;
  assign n18285 = n18284 ^ n4014 ;
  assign n18275 = n18198 ^ n18189 ;
  assign n18276 = n18190 & ~n18275 ;
  assign n18277 = n18276 ^ n18198 ;
  assign n18286 = n18285 ^ n18277 ;
  assign n18295 = n18294 ^ n18286 ;
  assign n18304 = n18303 ^ n18295 ;
  assign n18272 = ~n6360 & n7939 ;
  assign n18270 = x109 & n7935 ;
  assign n18266 = n18199 ^ n18173 ;
  assign n18267 = ~n18180 & ~n18266 ;
  assign n18268 = n18267 ^ n18199 ;
  assign n18264 = x111 & n7938 ;
  assign n18265 = n18264 ^ x56 ;
  assign n18269 = n18268 ^ n18265 ;
  assign n18271 = n18270 ^ n18269 ;
  assign n18273 = n18272 ^ n18271 ;
  assign n18263 = x110 & n7931 ;
  assign n18274 = n18273 ^ n18263 ;
  assign n18305 = n18304 ^ n18274 ;
  assign n18260 = n18200 ^ n18162 ;
  assign n18261 = ~n18168 & ~n18260 ;
  assign n18262 = n18261 ^ n18200 ;
  assign n18306 = n18305 ^ n18262 ;
  assign n18315 = n18314 ^ n18306 ;
  assign n18324 = n18323 ^ n18315 ;
  assign n18257 = n18201 ^ n18150 ;
  assign n18258 = ~n18156 & ~n18257 ;
  assign n18259 = n18258 ^ n18201 ;
  assign n18325 = n18324 ^ n18259 ;
  assign n18327 = n18325 ^ n18139 ;
  assign n18326 = n18325 ^ n18202 ;
  assign n18328 = n18327 ^ n18326 ;
  assign n18329 = n18144 & ~n18328 ;
  assign n18330 = n18329 ^ n18327 ;
  assign n18339 = n18338 ^ n18330 ;
  assign n18343 = n18342 ^ n18339 ;
  assign n18352 = n18351 ^ n18343 ;
  assign n18254 = n18226 ^ n18131 ;
  assign n18255 = n18218 & ~n18254 ;
  assign n18256 = n18255 ^ n18226 ;
  assign n18353 = n18352 ^ n18256 ;
  assign n18362 = n18361 ^ n18353 ;
  assign n18363 = n18362 ^ n18236 ;
  assign n18364 = n18363 ^ n18362 ;
  assign n18365 = n18364 ^ n18128 ;
  assign n18366 = n18228 & n18365 ;
  assign n18367 = n18366 ^ n18363 ;
  assign n18378 = n18377 ^ n18367 ;
  assign n18251 = n18244 ^ n18125 ;
  assign n18252 = n18238 & n18251 ;
  assign n18253 = n18252 ^ n18244 ;
  assign n18379 = n18378 ^ n18253 ;
  assign n18248 = n18122 ^ n18119 ;
  assign n18249 = ~n18246 & ~n18248 ;
  assign n18250 = n18249 ^ n18119 ;
  assign n18380 = n18379 ^ n18250 ;
  assign n18512 = n18253 ^ n18250 ;
  assign n18513 = ~n18379 & n18512 ;
  assign n18514 = n18513 ^ n18253 ;
  assign n18507 = n18377 ^ n18362 ;
  assign n18508 = ~n18367 & ~n18507 ;
  assign n18509 = n18508 ^ n18362 ;
  assign n18501 = x122 & n5094 ;
  assign n18500 = x124 & n5097 ;
  assign n18502 = n18501 ^ n18500 ;
  assign n18503 = n18502 ^ x44 ;
  assign n18499 = n5098 & n10095 ;
  assign n18504 = n18503 ^ n18499 ;
  assign n18498 = x123 & n5102 ;
  assign n18505 = n18504 ^ n18498 ;
  assign n18489 = n18338 ^ n18325 ;
  assign n18490 = n18330 & n18489 ;
  assign n18491 = n18490 ^ n18325 ;
  assign n18483 = x119 & n5965 ;
  assign n18482 = x121 & n5729 ;
  assign n18484 = n18483 ^ n18482 ;
  assign n18485 = n18484 ^ x47 ;
  assign n18481 = n5730 & n8962 ;
  assign n18486 = n18485 ^ n18481 ;
  assign n18480 = x120 & n5736 ;
  assign n18487 = n18486 ^ n18480 ;
  assign n18473 = ~n18277 & ~n18285 ;
  assign n18469 = ~x102 & n9948 ;
  assign n18470 = n18469 ^ n18188 ;
  assign n18471 = x101 & n18470 ;
  assign n18472 = n18471 ^ n18188 ;
  assign n18474 = n18473 ^ n18472 ;
  assign n18459 = x104 & n9632 ;
  assign n18458 = x106 & n9635 ;
  assign n18460 = n18459 ^ n18458 ;
  assign n18461 = n18460 ^ x62 ;
  assign n18457 = ~n5240 & n9636 ;
  assign n18462 = n18461 ^ n18457 ;
  assign n18456 = x105 & n9628 ;
  assign n18463 = n18462 ^ n18456 ;
  assign n18451 = x63 & x102 ;
  assign n18452 = n18451 ^ x103 ;
  assign n18453 = ~n9948 & n18452 ;
  assign n18445 = n18189 ^ x103 ;
  assign n18454 = n18453 ^ n18445 ;
  assign n18455 = n18454 ^ x38 ;
  assign n18464 = n18463 ^ n18455 ;
  assign n18475 = n18474 ^ n18464 ;
  assign n18435 = x107 & n8741 ;
  assign n18434 = x109 & n8744 ;
  assign n18436 = n18435 ^ n18434 ;
  assign n18437 = n18436 ^ x59 ;
  assign n18433 = n5902 & n8745 ;
  assign n18438 = n18437 ^ n18433 ;
  assign n18432 = x108 & n8737 ;
  assign n18439 = n18438 ^ n18432 ;
  assign n18440 = n18439 ^ n18303 ;
  assign n18441 = n18440 ^ n18294 ;
  assign n18442 = n18441 ^ n18439 ;
  assign n18443 = n18295 & n18442 ;
  assign n18444 = n18443 ^ n18440 ;
  assign n18476 = n18475 ^ n18444 ;
  assign n18422 = x110 & n7935 ;
  assign n18421 = x112 & n7938 ;
  assign n18423 = n18422 ^ n18421 ;
  assign n18424 = n18423 ^ x56 ;
  assign n18420 = ~n6600 & n7939 ;
  assign n18425 = n18424 ^ n18420 ;
  assign n18419 = x111 & n7931 ;
  assign n18426 = n18425 ^ n18419 ;
  assign n18427 = n18426 ^ n18304 ;
  assign n18428 = n18427 ^ n18268 ;
  assign n18429 = n18428 ^ n18426 ;
  assign n18430 = n18274 & n18429 ;
  assign n18431 = n18430 ^ n18427 ;
  assign n18477 = n18476 ^ n18431 ;
  assign n18416 = n18314 ^ n18262 ;
  assign n18417 = n18306 & ~n18416 ;
  assign n18409 = x113 & n7171 ;
  assign n18408 = x115 & n7174 ;
  assign n18410 = n18409 ^ n18408 ;
  assign n18411 = n18410 ^ x53 ;
  assign n18407 = n7175 & ~n7343 ;
  assign n18412 = n18411 ^ n18407 ;
  assign n18406 = x114 & n7179 ;
  assign n18413 = n18412 ^ n18406 ;
  assign n18414 = n18413 ^ n18314 ;
  assign n18418 = n18417 ^ n18414 ;
  assign n18478 = n18477 ^ n18418 ;
  assign n18403 = n18323 ^ n18259 ;
  assign n18404 = ~n18324 & ~n18403 ;
  assign n18396 = x116 & n6677 ;
  assign n18395 = x118 & n6428 ;
  assign n18397 = n18396 ^ n18395 ;
  assign n18398 = n18397 ^ x50 ;
  assign n18394 = n6429 & ~n8123 ;
  assign n18399 = n18398 ^ n18394 ;
  assign n18393 = x117 & n6433 ;
  assign n18400 = n18399 ^ n18393 ;
  assign n18401 = n18400 ^ n18323 ;
  assign n18405 = n18404 ^ n18401 ;
  assign n18479 = n18478 ^ n18405 ;
  assign n18488 = n18487 ^ n18479 ;
  assign n18492 = n18491 ^ n18488 ;
  assign n18493 = n18492 ^ n18351 ;
  assign n18494 = n18493 ^ n18342 ;
  assign n18495 = n18494 ^ n18492 ;
  assign n18496 = n18343 & ~n18495 ;
  assign n18497 = n18496 ^ n18493 ;
  assign n18506 = n18505 ^ n18497 ;
  assign n18510 = n18509 ^ n18506 ;
  assign n18387 = x125 & n4474 ;
  assign n18386 = x127 & n4471 ;
  assign n18388 = n18387 ^ n18386 ;
  assign n18389 = n18388 ^ x41 ;
  assign n18385 = n4472 & n10972 ;
  assign n18390 = n18389 ^ n18385 ;
  assign n18384 = x126 & n4467 ;
  assign n18391 = n18390 ^ n18384 ;
  assign n18381 = n18361 ^ n18256 ;
  assign n18382 = n18353 & n18381 ;
  assign n18383 = n18382 ^ n18361 ;
  assign n18392 = n18391 ^ n18383 ;
  assign n18511 = n18510 ^ n18392 ;
  assign n18515 = n18514 ^ n18511 ;
  assign n18629 = n18383 & n18391 ;
  assign n18628 = n18506 & n18509 ;
  assign n18630 = n18629 ^ n18628 ;
  assign n18623 = n4472 & n10139 ;
  assign n18622 = x126 & n4474 ;
  assign n18624 = n18623 ^ n18622 ;
  assign n18625 = n18624 ^ x41 ;
  assign n18621 = x127 & n4467 ;
  assign n18626 = n18625 ^ n18621 ;
  assign n18612 = n5098 & n10400 ;
  assign n18610 = x123 & n5094 ;
  assign n18606 = x121 & n5736 ;
  assign n18604 = n5730 & ~n9247 ;
  assign n18600 = x120 & n5965 ;
  assign n18599 = x122 & n5729 ;
  assign n18601 = n18600 ^ n18599 ;
  assign n18602 = n18601 ^ x47 ;
  assign n18595 = n18477 ^ n18413 ;
  assign n18596 = n18418 & ~n18595 ;
  assign n18597 = n18596 ^ n18413 ;
  assign n18593 = x118 & n6433 ;
  assign n18588 = x117 & n6677 ;
  assign n18587 = x119 & n6428 ;
  assign n18589 = n18588 ^ n18587 ;
  assign n18590 = n18589 ^ x50 ;
  assign n18586 = n6429 & n8394 ;
  assign n18591 = n18590 ^ n18586 ;
  assign n18577 = x108 & n8741 ;
  assign n18576 = x110 & n8744 ;
  assign n18578 = n18577 ^ n18576 ;
  assign n18579 = n18578 ^ x59 ;
  assign n18575 = n6129 & n8745 ;
  assign n18580 = n18579 ^ n18575 ;
  assign n18574 = x109 & n8737 ;
  assign n18581 = n18580 ^ n18574 ;
  assign n18568 = x105 & n9632 ;
  assign n18567 = x107 & n9635 ;
  assign n18569 = n18568 ^ n18567 ;
  assign n18570 = n18569 ^ x62 ;
  assign n18566 = ~n5448 & n9636 ;
  assign n18571 = n18570 ^ n18566 ;
  assign n18565 = x106 & n9628 ;
  assign n18572 = n18571 ^ n18565 ;
  assign n18561 = n18189 ^ x38 ;
  assign n18562 = ~n18454 & ~n18561 ;
  assign n18563 = n18562 ^ x38 ;
  assign n18557 = x63 & x103 ;
  assign n18558 = n18557 ^ x104 ;
  assign n18559 = ~n9948 & n18558 ;
  assign n18560 = n18559 ^ x104 ;
  assign n18564 = n18563 ^ n18560 ;
  assign n18573 = n18572 ^ n18564 ;
  assign n18582 = n18581 ^ n18573 ;
  assign n18552 = n18474 ^ n18463 ;
  assign n18553 = n18464 & ~n18552 ;
  assign n18554 = n18553 ^ n18474 ;
  assign n18583 = n18582 ^ n18554 ;
  assign n18549 = ~n6839 & n7939 ;
  assign n18547 = x111 & n7935 ;
  assign n18543 = n18475 ^ n18439 ;
  assign n18544 = n18444 & n18543 ;
  assign n18545 = n18544 ^ n18439 ;
  assign n18541 = x113 & n7938 ;
  assign n18542 = n18541 ^ x56 ;
  assign n18546 = n18545 ^ n18542 ;
  assign n18548 = n18547 ^ n18546 ;
  assign n18550 = n18549 ^ n18548 ;
  assign n18540 = x112 & n7931 ;
  assign n18551 = n18550 ^ n18540 ;
  assign n18584 = n18583 ^ n18551 ;
  assign n18530 = x114 & n7171 ;
  assign n18529 = x116 & n7174 ;
  assign n18531 = n18530 ^ n18529 ;
  assign n18532 = n18531 ^ x53 ;
  assign n18528 = n7175 & ~n7588 ;
  assign n18533 = n18532 ^ n18528 ;
  assign n18527 = x115 & n7179 ;
  assign n18534 = n18533 ^ n18527 ;
  assign n18536 = n18534 ^ n18426 ;
  assign n18535 = n18534 ^ n18476 ;
  assign n18537 = n18536 ^ n18535 ;
  assign n18538 = ~n18431 & n18537 ;
  assign n18539 = n18538 ^ n18536 ;
  assign n18585 = n18584 ^ n18539 ;
  assign n18592 = n18591 ^ n18585 ;
  assign n18594 = n18593 ^ n18592 ;
  assign n18598 = n18597 ^ n18594 ;
  assign n18603 = n18602 ^ n18598 ;
  assign n18605 = n18604 ^ n18603 ;
  assign n18607 = n18606 ^ n18605 ;
  assign n18524 = n18478 ^ n18400 ;
  assign n18525 = n18405 & ~n18524 ;
  assign n18526 = n18525 ^ n18400 ;
  assign n18608 = n18607 ^ n18526 ;
  assign n18522 = x125 & n5097 ;
  assign n18523 = n18522 ^ x44 ;
  assign n18609 = n18608 ^ n18523 ;
  assign n18611 = n18610 ^ n18609 ;
  assign n18613 = n18612 ^ n18611 ;
  assign n18521 = x124 & n5102 ;
  assign n18614 = n18613 ^ n18521 ;
  assign n18518 = n18491 ^ n18487 ;
  assign n18519 = n18488 & n18518 ;
  assign n18520 = n18519 ^ n18491 ;
  assign n18615 = n18614 ^ n18520 ;
  assign n18617 = n18615 ^ n18492 ;
  assign n18616 = n18615 ^ n18505 ;
  assign n18618 = n18617 ^ n18616 ;
  assign n18619 = ~n18497 & ~n18618 ;
  assign n18620 = n18619 ^ n18617 ;
  assign n18627 = n18626 ^ n18620 ;
  assign n18631 = n18630 ^ n18627 ;
  assign n18516 = n18514 ^ n18510 ;
  assign n18517 = n18511 & n18516 ;
  assign n18632 = n18631 ^ n18517 ;
  assign n18744 = n18514 & ~n18628 ;
  assign n18739 = n18629 ^ n18392 ;
  assign n18740 = n18739 ^ n18506 ;
  assign n18741 = n18510 & ~n18740 ;
  assign n18742 = n18741 ^ n18506 ;
  assign n18743 = n18627 & ~n18742 ;
  assign n18745 = n18629 ^ n18627 ;
  assign n18746 = ~n18743 & n18745 ;
  assign n18747 = n18744 & n18746 ;
  assign n18748 = n18747 ^ n18743 ;
  assign n18749 = n18628 ^ n18510 ;
  assign n18750 = n18749 ^ n18627 ;
  assign n18751 = n18514 ^ n18391 ;
  assign n18754 = n18392 & n18751 ;
  assign n18755 = n18754 ^ n18391 ;
  assign n18756 = ~n18750 & n18755 ;
  assign n18757 = ~n18748 & ~n18756 ;
  assign n18735 = n18626 ^ n18615 ;
  assign n18736 = n18620 & ~n18735 ;
  assign n18737 = n18736 ^ n18615 ;
  assign n4475 = n4474 ^ n4472 ;
  assign n18730 = x127 & n4475 ;
  assign n18729 = n4472 & n10138 ;
  assign n18731 = n18730 ^ n18729 ;
  assign n18732 = n18731 ^ x41 ;
  assign n18726 = n18608 ^ n18520 ;
  assign n18727 = ~n18614 & ~n18726 ;
  assign n18728 = n18727 ^ n18608 ;
  assign n18733 = n18732 ^ n18728 ;
  assign n18720 = x124 & n5094 ;
  assign n18719 = x126 & n5097 ;
  assign n18721 = n18720 ^ n18719 ;
  assign n18722 = n18721 ^ x44 ;
  assign n18718 = n5098 & n10441 ;
  assign n18723 = n18722 ^ n18718 ;
  assign n18717 = x125 & n5102 ;
  assign n18724 = n18723 ^ n18717 ;
  assign n18710 = x121 & n5965 ;
  assign n18709 = x123 & n5729 ;
  assign n18711 = n18710 ^ n18709 ;
  assign n18712 = n18711 ^ x47 ;
  assign n18708 = n5730 & ~n9786 ;
  assign n18713 = n18712 ^ n18708 ;
  assign n18707 = x122 & n5736 ;
  assign n18714 = n18713 ^ n18707 ;
  assign n18697 = n7175 & ~n7850 ;
  assign n18695 = x115 & n7171 ;
  assign n18691 = n18583 ^ n18545 ;
  assign n18692 = ~n18551 & ~n18691 ;
  assign n18693 = n18692 ^ n18583 ;
  assign n18689 = x117 & n7174 ;
  assign n18690 = n18689 ^ x53 ;
  assign n18694 = n18693 ^ n18690 ;
  assign n18696 = n18695 ^ n18694 ;
  assign n18698 = n18697 ^ n18696 ;
  assign n18688 = x116 & n7179 ;
  assign n18699 = n18698 ^ n18688 ;
  assign n18681 = x109 & n8741 ;
  assign n18680 = x111 & n8744 ;
  assign n18682 = n18681 ^ n18680 ;
  assign n18683 = n18682 ^ x59 ;
  assign n18679 = ~n6360 & n8745 ;
  assign n18684 = n18683 ^ n18679 ;
  assign n18678 = x110 & n8737 ;
  assign n18685 = n18684 ^ n18678 ;
  assign n18676 = x107 & n9628 ;
  assign n18669 = n18572 ^ n18563 ;
  assign n18670 = n18564 & n18669 ;
  assign n18665 = x63 & x104 ;
  assign n18666 = n18665 ^ x105 ;
  assign n18667 = ~n9948 & n18666 ;
  assign n18668 = n18667 ^ x105 ;
  assign n18671 = n18670 ^ n18668 ;
  assign n18672 = n18671 ^ x62 ;
  assign n18662 = x106 & n9632 ;
  assign n18673 = n18672 ^ n18662 ;
  assign n18661 = x108 & n9635 ;
  assign n18674 = n18673 ^ n18661 ;
  assign n18660 = n5670 & n9636 ;
  assign n18675 = n18674 ^ n18660 ;
  assign n18677 = n18676 ^ n18675 ;
  assign n18686 = n18685 ^ n18677 ;
  assign n18658 = x113 & n7931 ;
  assign n18653 = x112 & n7935 ;
  assign n18652 = x114 & n7938 ;
  assign n18654 = n18653 ^ n18652 ;
  assign n18655 = n18654 ^ x56 ;
  assign n18651 = ~n7092 & n7939 ;
  assign n18656 = n18655 ^ n18651 ;
  assign n18648 = n18581 ^ n18554 ;
  assign n18649 = n18582 & ~n18648 ;
  assign n18650 = n18649 ^ n18581 ;
  assign n18657 = n18656 ^ n18650 ;
  assign n18659 = n18658 ^ n18657 ;
  assign n18687 = n18686 ^ n18659 ;
  assign n18700 = n18699 ^ n18687 ;
  assign n18645 = n6429 & n8891 ;
  assign n18643 = x118 & n6677 ;
  assign n18639 = n18584 ^ n18534 ;
  assign n18640 = n18539 & ~n18639 ;
  assign n18641 = n18640 ^ n18534 ;
  assign n18637 = x120 & n6428 ;
  assign n18638 = n18637 ^ x50 ;
  assign n18642 = n18641 ^ n18638 ;
  assign n18644 = n18643 ^ n18642 ;
  assign n18646 = n18645 ^ n18644 ;
  assign n18636 = x119 & n6433 ;
  assign n18647 = n18646 ^ n18636 ;
  assign n18701 = n18700 ^ n18647 ;
  assign n18703 = n18701 ^ n18597 ;
  assign n18702 = n18701 ^ n18585 ;
  assign n18704 = n18703 ^ n18702 ;
  assign n18705 = ~n18594 & ~n18704 ;
  assign n18706 = n18705 ^ n18702 ;
  assign n18715 = n18714 ^ n18706 ;
  assign n18633 = n18598 ^ n18526 ;
  assign n18634 = ~n18607 & ~n18633 ;
  assign n18635 = n18634 ^ n18598 ;
  assign n18716 = n18715 ^ n18635 ;
  assign n18725 = n18724 ^ n18716 ;
  assign n18734 = n18733 ^ n18725 ;
  assign n18738 = n18737 ^ n18734 ;
  assign n18758 = n18757 ^ n18738 ;
  assign n18876 = x125 & n5094 ;
  assign n18875 = x127 & n5097 ;
  assign n18877 = n18876 ^ n18875 ;
  assign n18878 = n18877 ^ x44 ;
  assign n18874 = n5098 & n10972 ;
  assign n18879 = n18878 ^ n18874 ;
  assign n18873 = x126 & n5102 ;
  assign n18880 = n18879 ^ n18873 ;
  assign n18869 = n18714 ^ n18701 ;
  assign n18870 = n18706 & ~n18869 ;
  assign n18871 = n18870 ^ n18701 ;
  assign n18863 = x122 & n5965 ;
  assign n18862 = x124 & n5729 ;
  assign n18864 = n18863 ^ n18862 ;
  assign n18865 = n18864 ^ x47 ;
  assign n18861 = n5730 & n10095 ;
  assign n18866 = n18865 ^ n18861 ;
  assign n18860 = x123 & n5736 ;
  assign n18867 = n18866 ^ n18860 ;
  assign n18851 = x113 & n7935 ;
  assign n18850 = x115 & n7938 ;
  assign n18852 = n18851 ^ n18850 ;
  assign n18853 = n18852 ^ x56 ;
  assign n18849 = ~n7343 & n7939 ;
  assign n18854 = n18853 ^ n18849 ;
  assign n18848 = x114 & n7931 ;
  assign n18855 = n18854 ^ n18848 ;
  assign n18841 = x110 & n8741 ;
  assign n18840 = x112 & n8744 ;
  assign n18842 = n18841 ^ n18840 ;
  assign n18843 = n18842 ^ x59 ;
  assign n18839 = ~n6600 & n8745 ;
  assign n18844 = n18843 ^ n18839 ;
  assign n18838 = x111 & n8737 ;
  assign n18845 = n18844 ^ n18838 ;
  assign n18832 = x63 & x105 ;
  assign n18833 = n18832 ^ x106 ;
  assign n18834 = ~n9948 & n18833 ;
  assign n18826 = n18560 ^ x106 ;
  assign n18835 = n18834 ^ n18826 ;
  assign n18836 = n18835 ^ x41 ;
  assign n18823 = n5902 & n9636 ;
  assign n18821 = x107 & n9632 ;
  assign n18817 = n18668 ^ n18560 ;
  assign n18818 = n18670 & ~n18817 ;
  assign n18819 = n18818 ^ n18560 ;
  assign n18815 = x109 & n9635 ;
  assign n18816 = n18815 ^ x62 ;
  assign n18820 = n18819 ^ n18816 ;
  assign n18822 = n18821 ^ n18820 ;
  assign n18824 = n18823 ^ n18822 ;
  assign n18814 = x108 & n9628 ;
  assign n18825 = n18824 ^ n18814 ;
  assign n18837 = n18836 ^ n18825 ;
  assign n18846 = n18845 ^ n18837 ;
  assign n18811 = n18685 ^ n18671 ;
  assign n18812 = ~n18677 & n18811 ;
  assign n18813 = n18812 ^ n18685 ;
  assign n18847 = n18846 ^ n18813 ;
  assign n18856 = n18855 ^ n18847 ;
  assign n18808 = n18686 ^ n18650 ;
  assign n18809 = n18659 & n18808 ;
  assign n18810 = n18809 ^ n18650 ;
  assign n18857 = n18856 ^ n18810 ;
  assign n18805 = n18693 ^ n18687 ;
  assign n18806 = n18699 & ~n18805 ;
  assign n18798 = x116 & n7171 ;
  assign n18797 = x118 & n7174 ;
  assign n18799 = n18798 ^ n18797 ;
  assign n18800 = n18799 ^ x53 ;
  assign n18796 = n7175 & ~n8123 ;
  assign n18801 = n18800 ^ n18796 ;
  assign n18795 = x117 & n7179 ;
  assign n18802 = n18801 ^ n18795 ;
  assign n18803 = n18802 ^ n18687 ;
  assign n18807 = n18806 ^ n18803 ;
  assign n18858 = n18857 ^ n18807 ;
  assign n18785 = x119 & n6677 ;
  assign n18784 = x121 & n6428 ;
  assign n18786 = n18785 ^ n18784 ;
  assign n18787 = n18786 ^ x50 ;
  assign n18783 = n6429 & n8962 ;
  assign n18788 = n18787 ^ n18783 ;
  assign n18782 = x120 & n6433 ;
  assign n18789 = n18788 ^ n18782 ;
  assign n18790 = n18789 ^ n18700 ;
  assign n18791 = n18790 ^ n18641 ;
  assign n18792 = n18791 ^ n18789 ;
  assign n18793 = ~n18647 & ~n18792 ;
  assign n18794 = n18793 ^ n18790 ;
  assign n18859 = n18858 ^ n18794 ;
  assign n18868 = n18867 ^ n18859 ;
  assign n18872 = n18871 ^ n18868 ;
  assign n18881 = n18880 ^ n18872 ;
  assign n18779 = n18724 ^ n18635 ;
  assign n18780 = n18716 & ~n18779 ;
  assign n18781 = n18780 ^ n18724 ;
  assign n18882 = n18881 ^ n18781 ;
  assign n18762 = n18732 ^ n18725 ;
  assign n18763 = ~n18733 & n18762 ;
  assign n18764 = n18763 ^ n18762 ;
  assign n18759 = ~n18728 & n18732 ;
  assign n18760 = ~n18725 & n18759 ;
  assign n18765 = n18764 ^ n18760 ;
  assign n18766 = n18737 & n18765 ;
  assign n18761 = ~n18737 & n18760 ;
  assign n18767 = n18766 ^ n18761 ;
  assign n18768 = n18763 ^ n18728 ;
  assign n18769 = n18760 ^ n18737 ;
  assign n18770 = n18769 ^ n18761 ;
  assign n18771 = ~n18768 & ~n18770 ;
  assign n18772 = n18771 ^ n18738 ;
  assign n18773 = n18772 ^ n18771 ;
  assign n18774 = n18771 ^ n18757 ;
  assign n18775 = n18774 ^ n18771 ;
  assign n18776 = ~n18773 & n18775 ;
  assign n18777 = n18776 ^ n18771 ;
  assign n18778 = ~n18767 & ~n18777 ;
  assign n18883 = n18882 ^ n18778 ;
  assign n18986 = n18772 ^ n18767 ;
  assign n18987 = ~n18757 & ~n18766 ;
  assign n18988 = n18882 ^ n18771 ;
  assign n18989 = ~n18761 & n18988 ;
  assign n18990 = n18987 & n18989 ;
  assign n18991 = n18990 ^ n18761 ;
  assign n18992 = n18882 & ~n18991 ;
  assign n18993 = n18986 & n18992 ;
  assign n18994 = n18993 ^ n18991 ;
  assign n18976 = n5098 & n10139 ;
  assign n18975 = x126 & n5094 ;
  assign n18977 = n18976 ^ n18975 ;
  assign n18978 = n18977 ^ x44 ;
  assign n18974 = x127 & n5102 ;
  assign n18979 = n18978 ^ n18974 ;
  assign n18966 = x120 & n6677 ;
  assign n18965 = x122 & n6428 ;
  assign n18967 = n18966 ^ n18965 ;
  assign n18968 = n18967 ^ x50 ;
  assign n18964 = n6429 & ~n9247 ;
  assign n18969 = n18968 ^ n18964 ;
  assign n18963 = x121 & n6433 ;
  assign n18970 = n18969 ^ n18963 ;
  assign n18954 = n18855 ^ n18810 ;
  assign n18955 = n18856 & n18954 ;
  assign n18956 = n18955 ^ n18855 ;
  assign n18948 = x117 & n7171 ;
  assign n18947 = x119 & n7174 ;
  assign n18949 = n18948 ^ n18947 ;
  assign n18950 = n18949 ^ x53 ;
  assign n18946 = n7175 & n8394 ;
  assign n18951 = n18950 ^ n18946 ;
  assign n18945 = x118 & n7179 ;
  assign n18952 = n18951 ^ n18945 ;
  assign n18937 = x108 & n9632 ;
  assign n18936 = x110 & n9635 ;
  assign n18938 = n18937 ^ n18936 ;
  assign n18939 = n18938 ^ x62 ;
  assign n18935 = n6129 & n9636 ;
  assign n18940 = n18939 ^ n18935 ;
  assign n18934 = x109 & n9628 ;
  assign n18941 = n18940 ^ n18934 ;
  assign n18930 = n18560 ^ x41 ;
  assign n18931 = ~n18835 & ~n18930 ;
  assign n18932 = n18931 ^ x41 ;
  assign n18926 = x63 & x106 ;
  assign n18927 = n18926 ^ x107 ;
  assign n18928 = ~n9948 & n18927 ;
  assign n18929 = n18928 ^ x107 ;
  assign n18933 = n18932 ^ n18929 ;
  assign n18942 = n18941 ^ n18933 ;
  assign n18921 = ~n6839 & n8745 ;
  assign n18919 = x111 & n8741 ;
  assign n18915 = n18836 ^ n18819 ;
  assign n18916 = n18825 & n18915 ;
  assign n18917 = n18916 ^ n18836 ;
  assign n18913 = x113 & n8744 ;
  assign n18914 = n18913 ^ x59 ;
  assign n18918 = n18917 ^ n18914 ;
  assign n18920 = n18919 ^ n18918 ;
  assign n18922 = n18921 ^ n18920 ;
  assign n18912 = x112 & n8737 ;
  assign n18923 = n18922 ^ n18912 ;
  assign n18943 = n18942 ^ n18923 ;
  assign n18909 = n18845 ^ n18813 ;
  assign n18910 = n18846 & n18909 ;
  assign n18902 = x114 & n7935 ;
  assign n18901 = x116 & n7938 ;
  assign n18903 = n18902 ^ n18901 ;
  assign n18904 = n18903 ^ x56 ;
  assign n18900 = ~n7588 & n7939 ;
  assign n18905 = n18904 ^ n18900 ;
  assign n18899 = x115 & n7931 ;
  assign n18906 = n18905 ^ n18899 ;
  assign n18907 = n18906 ^ n18845 ;
  assign n18911 = n18910 ^ n18907 ;
  assign n18944 = n18943 ^ n18911 ;
  assign n18953 = n18952 ^ n18944 ;
  assign n18957 = n18956 ^ n18953 ;
  assign n18959 = n18957 ^ n18802 ;
  assign n18958 = n18957 ^ n18857 ;
  assign n18960 = n18959 ^ n18958 ;
  assign n18961 = n18807 & n18960 ;
  assign n18962 = n18961 ^ n18959 ;
  assign n18971 = n18970 ^ n18962 ;
  assign n18896 = n5730 & n10400 ;
  assign n18894 = x123 & n5965 ;
  assign n18890 = n18858 ^ n18789 ;
  assign n18891 = ~n18794 & n18890 ;
  assign n18892 = n18891 ^ n18789 ;
  assign n18888 = x125 & n5729 ;
  assign n18889 = n18888 ^ x47 ;
  assign n18893 = n18892 ^ n18889 ;
  assign n18895 = n18894 ^ n18893 ;
  assign n18897 = n18896 ^ n18895 ;
  assign n18887 = x124 & n5736 ;
  assign n18898 = n18897 ^ n18887 ;
  assign n18972 = n18971 ^ n18898 ;
  assign n18884 = n18871 ^ n18867 ;
  assign n18885 = n18868 & ~n18884 ;
  assign n18886 = n18885 ^ n18871 ;
  assign n18973 = n18972 ^ n18886 ;
  assign n18980 = n18979 ^ n18973 ;
  assign n18981 = n18980 ^ n18880 ;
  assign n18982 = n18981 ^ n18781 ;
  assign n18983 = n18982 ^ n18980 ;
  assign n18984 = n18881 & n18983 ;
  assign n18985 = n18984 ^ n18981 ;
  assign n18995 = n18994 ^ n18985 ;
  assign n19087 = x127 & n5093 ;
  assign n19088 = n19087 ^ n5091 ;
  assign n19093 = n4670 & n11265 ;
  assign n19094 = n19093 ^ n19087 ;
  assign n19095 = n19088 & ~n19094 ;
  assign n19096 = n19095 ^ x43 ;
  assign n19084 = n18971 ^ n18892 ;
  assign n19085 = ~n18898 & ~n19084 ;
  assign n19086 = n19085 ^ n18971 ;
  assign n19097 = n19096 ^ n19086 ;
  assign n19081 = x125 & n5736 ;
  assign n19079 = n5730 & n10441 ;
  assign n19075 = x124 & n5965 ;
  assign n19074 = x126 & n5729 ;
  assign n19076 = n19075 ^ n19074 ;
  assign n19077 = n19076 ^ x47 ;
  assign n19071 = x122 & n6433 ;
  assign n19069 = n6429 & ~n9786 ;
  assign n19065 = x121 & n6677 ;
  assign n19064 = x123 & n6428 ;
  assign n19066 = n19065 ^ n19064 ;
  assign n19067 = n19066 ^ x50 ;
  assign n19061 = x119 & n7179 ;
  assign n19059 = n7175 & n8891 ;
  assign n19055 = x118 & n7171 ;
  assign n19054 = x120 & n7174 ;
  assign n19056 = n19055 ^ n19054 ;
  assign n19057 = n19056 ^ x53 ;
  assign n19047 = x115 & n7935 ;
  assign n19046 = x117 & n7938 ;
  assign n19048 = n19047 ^ n19046 ;
  assign n19049 = n19048 ^ x56 ;
  assign n19045 = ~n7850 & n7939 ;
  assign n19050 = n19049 ^ n19045 ;
  assign n19044 = x116 & n7931 ;
  assign n19051 = n19050 ^ n19044 ;
  assign n19038 = x112 & n8741 ;
  assign n19037 = x114 & n8744 ;
  assign n19039 = n19038 ^ n19037 ;
  assign n19040 = n19039 ^ x59 ;
  assign n19036 = ~n7092 & n8745 ;
  assign n19041 = n19040 ^ n19036 ;
  assign n19035 = x113 & n8737 ;
  assign n19042 = n19041 ^ n19035 ;
  assign n19029 = ~n6360 & n9636 ;
  assign n19028 = x110 & n9628 ;
  assign n19030 = n19029 ^ n19028 ;
  assign n19026 = x109 & n9632 ;
  assign n19025 = x111 & n9635 ;
  assign n19027 = n19026 ^ n19025 ;
  assign n19031 = n19030 ^ n19027 ;
  assign n19024 = n5218 ^ x62 ;
  assign n19032 = n19031 ^ n19024 ;
  assign n19021 = n18941 ^ n18932 ;
  assign n19022 = ~n18933 & ~n19021 ;
  assign n19023 = n19022 ^ n18941 ;
  assign n19033 = n19032 ^ n19023 ;
  assign n19018 = x63 & n4998 ;
  assign n19019 = n19018 ^ n5218 ;
  assign n19020 = ~n9948 & n19019 ;
  assign n19034 = n19033 ^ n19020 ;
  assign n19043 = n19042 ^ n19034 ;
  assign n19052 = n19051 ^ n19043 ;
  assign n19011 = n18942 ^ n18917 ;
  assign n19012 = n18923 & ~n19011 ;
  assign n19013 = n19012 ^ n18942 ;
  assign n19053 = n19052 ^ n19013 ;
  assign n19058 = n19057 ^ n19053 ;
  assign n19060 = n19059 ^ n19058 ;
  assign n19062 = n19061 ^ n19060 ;
  assign n19008 = n18943 ^ n18906 ;
  assign n19009 = n18911 & ~n19008 ;
  assign n19010 = n19009 ^ n18906 ;
  assign n19063 = n19062 ^ n19010 ;
  assign n19068 = n19067 ^ n19063 ;
  assign n19070 = n19069 ^ n19068 ;
  assign n19072 = n19071 ^ n19070 ;
  assign n19005 = n18956 ^ n18952 ;
  assign n19006 = n18953 & n19005 ;
  assign n19007 = n19006 ^ n18956 ;
  assign n19073 = n19072 ^ n19007 ;
  assign n19078 = n19077 ^ n19073 ;
  assign n19080 = n19079 ^ n19078 ;
  assign n19082 = n19081 ^ n19080 ;
  assign n19002 = n18970 ^ n18957 ;
  assign n19003 = ~n18962 & ~n19002 ;
  assign n19004 = n19003 ^ n18957 ;
  assign n19083 = n19082 ^ n19004 ;
  assign n19098 = n19097 ^ n19083 ;
  assign n18999 = n18979 ^ n18886 ;
  assign n19000 = ~n18973 & ~n18999 ;
  assign n19001 = n19000 ^ n18979 ;
  assign n19099 = n19098 ^ n19001 ;
  assign n18996 = n18994 ^ n18980 ;
  assign n18997 = n18985 & n18996 ;
  assign n18998 = n18997 ^ n18980 ;
  assign n19100 = n19099 ^ n18998 ;
  assign n19101 = n19096 ^ n19083 ;
  assign n19218 = n19083 ^ n18998 ;
  assign n19219 = ~n19101 & ~n19218 ;
  assign n19213 = n19073 ^ n19004 ;
  assign n19214 = ~n19082 & n19213 ;
  assign n19215 = n19214 ^ n19073 ;
  assign n19207 = x125 & n5965 ;
  assign n19206 = x127 & n5729 ;
  assign n19208 = n19207 ^ n19206 ;
  assign n19209 = n19208 ^ x47 ;
  assign n19205 = n5730 & n10972 ;
  assign n19210 = n19209 ^ n19205 ;
  assign n19204 = x126 & n5736 ;
  assign n19211 = n19210 ^ n19204 ;
  assign n19200 = n19063 ^ n19007 ;
  assign n19201 = ~n19072 & ~n19200 ;
  assign n19202 = n19201 ^ n19063 ;
  assign n19194 = x122 & n6677 ;
  assign n19193 = x124 & n6428 ;
  assign n19195 = n19194 ^ n19193 ;
  assign n19196 = n19195 ^ x50 ;
  assign n19192 = n6429 & n10095 ;
  assign n19197 = n19196 ^ n19192 ;
  assign n19191 = x123 & n6433 ;
  assign n19198 = n19197 ^ n19191 ;
  assign n19186 = n19051 ^ n19013 ;
  assign n19187 = ~n19052 & n19186 ;
  assign n19188 = n19187 ^ n19051 ;
  assign n19184 = x117 & n7931 ;
  assign n19165 = x108 ^ x63 ;
  assign n19166 = n19165 ^ n19031 ;
  assign n19169 = n5218 & ~n19166 ;
  assign n19170 = n19169 ^ n19031 ;
  assign n19171 = n9948 & n19170 ;
  assign n19154 = x107 & ~x108 ;
  assign n19156 = n19154 ^ x106 ;
  assign n19155 = n19154 ^ n19031 ;
  assign n19157 = n19156 ^ n19155 ;
  assign n19160 = ~n4998 & n19157 ;
  assign n19161 = n19160 ^ n19156 ;
  assign n19162 = x62 & n19161 ;
  assign n19163 = n19162 ^ n19154 ;
  assign n19164 = x63 & n19163 ;
  assign n19172 = n19171 ^ x62 ;
  assign n19173 = ~n19164 & ~n19172 ;
  assign n19174 = n19031 & n19173 ;
  assign n19175 = ~n19171 & n19174 ;
  assign n19176 = n19175 ^ n19173 ;
  assign n19177 = n19176 ^ n19164 ;
  assign n19148 = x110 & n9632 ;
  assign n19147 = x112 & n9635 ;
  assign n19149 = n19148 ^ n19147 ;
  assign n19150 = n19149 ^ x62 ;
  assign n19146 = ~n6600 & n9636 ;
  assign n19151 = n19150 ^ n19146 ;
  assign n19145 = x111 & n9628 ;
  assign n19152 = n19151 ^ n19145 ;
  assign n19140 = ~x63 & x108 ;
  assign n19141 = n19140 ^ n5427 ;
  assign n19142 = ~n9948 & n19141 ;
  assign n19135 = n18929 ^ x109 ;
  assign n19143 = n19142 ^ n19135 ;
  assign n19144 = n19143 ^ x44 ;
  assign n19153 = n19152 ^ n19144 ;
  assign n19178 = n19177 ^ n19153 ;
  assign n19132 = n19042 ^ n19023 ;
  assign n19133 = n19034 & n19132 ;
  assign n19125 = x113 & n8741 ;
  assign n19124 = x115 & n8744 ;
  assign n19126 = n19125 ^ n19124 ;
  assign n19127 = n19126 ^ x59 ;
  assign n19123 = ~n7343 & n8745 ;
  assign n19128 = n19127 ^ n19123 ;
  assign n19122 = x114 & n8737 ;
  assign n19129 = n19128 ^ n19122 ;
  assign n19130 = n19129 ^ n19042 ;
  assign n19134 = n19133 ^ n19130 ;
  assign n19179 = n19178 ^ n19134 ;
  assign n19180 = n19179 ^ x56 ;
  assign n19121 = x116 & n7935 ;
  assign n19181 = n19180 ^ n19121 ;
  assign n19120 = x118 & n7938 ;
  assign n19182 = n19181 ^ n19120 ;
  assign n19119 = n7939 & ~n8123 ;
  assign n19183 = n19182 ^ n19119 ;
  assign n19185 = n19184 ^ n19183 ;
  assign n19189 = n19188 ^ n19185 ;
  assign n19109 = x119 & n7171 ;
  assign n19108 = x121 & n7174 ;
  assign n19110 = n19109 ^ n19108 ;
  assign n19111 = n19110 ^ x53 ;
  assign n19107 = n7175 & n8962 ;
  assign n19112 = n19111 ^ n19107 ;
  assign n19106 = x120 & n7179 ;
  assign n19113 = n19112 ^ n19106 ;
  assign n19114 = n19113 ^ n19053 ;
  assign n19115 = n19114 ^ n19010 ;
  assign n19116 = n19115 ^ n19113 ;
  assign n19117 = ~n19062 & ~n19116 ;
  assign n19118 = n19117 ^ n19114 ;
  assign n19190 = n19189 ^ n19118 ;
  assign n19199 = n19198 ^ n19190 ;
  assign n19203 = n19202 ^ n19199 ;
  assign n19212 = n19211 ^ n19203 ;
  assign n19216 = n19215 ^ n19212 ;
  assign n19102 = n19101 ^ n18998 ;
  assign n19103 = n19102 ^ n19086 ;
  assign n19104 = n19086 ^ n19001 ;
  assign n19105 = ~n19103 & n19104 ;
  assign n19217 = n19216 ^ n19105 ;
  assign n19220 = n19219 ^ n19217 ;
  assign n19304 = n19001 & ~n19086 ;
  assign n19305 = n19304 ^ n19216 ;
  assign n19306 = n19305 ^ n19104 ;
  assign n19307 = ~n18998 & n19306 ;
  assign n19309 = n19307 ^ n19096 ;
  assign n19310 = n19309 ^ n19216 ;
  assign n19308 = n19307 ^ n19083 ;
  assign n19311 = n19310 ^ n19308 ;
  assign n19312 = n19307 & ~n19311 ;
  assign n19313 = n19312 ^ n19216 ;
  assign n19314 = n19308 ^ n19304 ;
  assign n19315 = n19312 ^ n19311 ;
  assign n19316 = n19314 & ~n19315 ;
  assign n19317 = n19316 ^ n19308 ;
  assign n19318 = n19313 & ~n19317 ;
  assign n19319 = n19318 ^ n19307 ;
  assign n19320 = ~n19083 & ~n19096 ;
  assign n19321 = n19320 ^ n19216 ;
  assign n19322 = n19001 ^ n18998 ;
  assign n19323 = n19104 ^ n18998 ;
  assign n19324 = n19323 ^ n18998 ;
  assign n19325 = n19322 & n19324 ;
  assign n19326 = n19325 ^ n18998 ;
  assign n19327 = n19321 & ~n19326 ;
  assign n19328 = ~n19319 & ~n19327 ;
  assign n19297 = n5730 & n10139 ;
  assign n19296 = x126 & n5965 ;
  assign n19298 = n19297 ^ n19296 ;
  assign n19299 = n19298 ^ x47 ;
  assign n19295 = x127 & n5736 ;
  assign n19300 = n19299 ^ n19295 ;
  assign n19292 = x124 & n6433 ;
  assign n19290 = n6429 & n10400 ;
  assign n19286 = x123 & n6677 ;
  assign n19285 = x125 & n6428 ;
  assign n19287 = n19286 ^ n19285 ;
  assign n19288 = n19287 ^ x50 ;
  assign n19278 = x120 & n7171 ;
  assign n19277 = x122 & n7174 ;
  assign n19279 = n19278 ^ n19277 ;
  assign n19280 = n19279 ^ x53 ;
  assign n19276 = n7175 & ~n9247 ;
  assign n19281 = n19280 ^ n19276 ;
  assign n19275 = x121 & n7179 ;
  assign n19282 = n19281 ^ n19275 ;
  assign n19271 = n19178 ^ n19129 ;
  assign n19272 = n19134 & n19271 ;
  assign n19273 = n19272 ^ n19129 ;
  assign n19265 = x117 & n7935 ;
  assign n19264 = x119 & n7938 ;
  assign n19266 = n19265 ^ n19264 ;
  assign n19267 = n19266 ^ x56 ;
  assign n19263 = n7939 & n8394 ;
  assign n19268 = n19267 ^ n19263 ;
  assign n19262 = x118 & n7931 ;
  assign n19269 = n19268 ^ n19262 ;
  assign n19255 = x114 & n8741 ;
  assign n19254 = x116 & n8744 ;
  assign n19256 = n19255 ^ n19254 ;
  assign n19257 = n19256 ^ x59 ;
  assign n19253 = ~n7588 & n8745 ;
  assign n19258 = n19257 ^ n19253 ;
  assign n19252 = x115 & n8737 ;
  assign n19259 = n19258 ^ n19252 ;
  assign n19249 = x109 & n11875 ;
  assign n19248 = x110 & n9948 ;
  assign n19250 = n19249 ^ n19248 ;
  assign n19245 = ~n6839 & n9636 ;
  assign n19243 = x111 & n9632 ;
  assign n19239 = n18929 ^ x44 ;
  assign n19240 = ~n19143 & ~n19239 ;
  assign n19241 = n19240 ^ x44 ;
  assign n19237 = x113 & n9635 ;
  assign n19238 = n19237 ^ x62 ;
  assign n19242 = n19241 ^ n19238 ;
  assign n19244 = n19243 ^ n19242 ;
  assign n19246 = n19245 ^ n19244 ;
  assign n19236 = x112 & n9628 ;
  assign n19247 = n19246 ^ n19236 ;
  assign n19251 = n19250 ^ n19247 ;
  assign n19260 = n19259 ^ n19251 ;
  assign n19233 = n19177 ^ n19152 ;
  assign n19234 = n19153 & ~n19233 ;
  assign n19235 = n19234 ^ n19177 ;
  assign n19261 = n19260 ^ n19235 ;
  assign n19270 = n19269 ^ n19261 ;
  assign n19274 = n19273 ^ n19270 ;
  assign n19283 = n19282 ^ n19274 ;
  assign n19230 = n19188 ^ n19179 ;
  assign n19231 = ~n19185 & n19230 ;
  assign n19232 = n19231 ^ n19188 ;
  assign n19284 = n19283 ^ n19232 ;
  assign n19289 = n19288 ^ n19284 ;
  assign n19291 = n19290 ^ n19289 ;
  assign n19293 = n19292 ^ n19291 ;
  assign n19227 = n19189 ^ n19113 ;
  assign n19228 = ~n19118 & n19227 ;
  assign n19229 = n19228 ^ n19113 ;
  assign n19294 = n19293 ^ n19229 ;
  assign n19301 = n19300 ^ n19294 ;
  assign n19224 = n19202 ^ n19198 ;
  assign n19225 = n19199 & ~n19224 ;
  assign n19226 = n19225 ^ n19202 ;
  assign n19302 = n19301 ^ n19226 ;
  assign n19221 = n19215 ^ n19211 ;
  assign n19222 = ~n19212 & ~n19221 ;
  assign n19223 = n19222 ^ n19215 ;
  assign n19303 = n19302 ^ n19223 ;
  assign n19329 = n19328 ^ n19303 ;
  assign n19422 = n19284 ^ n19229 ;
  assign n19423 = ~n19293 & ~n19422 ;
  assign n19424 = n19423 ^ n19284 ;
  assign n19342 = n5309 & n11265 ;
  assign n19337 = x127 & n5964 ;
  assign n19343 = n19342 ^ n19337 ;
  assign n19413 = x125 & n6433 ;
  assign n19411 = n6429 & n10441 ;
  assign n19407 = x124 & n6677 ;
  assign n19406 = x126 & n6428 ;
  assign n19408 = n19407 ^ n19406 ;
  assign n19409 = n19408 ^ x50 ;
  assign n19399 = x121 & n7171 ;
  assign n19398 = x123 & n7174 ;
  assign n19400 = n19399 ^ n19398 ;
  assign n19401 = n19400 ^ x53 ;
  assign n19397 = n7175 & ~n9786 ;
  assign n19402 = n19401 ^ n19397 ;
  assign n19396 = x122 & n7179 ;
  assign n19403 = n19402 ^ n19396 ;
  assign n19383 = ~x111 & n9948 ;
  assign n19384 = n19383 ^ n19249 ;
  assign n19385 = x110 & n19384 ;
  assign n19386 = n19385 ^ n19249 ;
  assign n19387 = n9948 ^ x110 ;
  assign n19388 = n19384 ^ n12206 ;
  assign n19389 = n19387 & n19388 ;
  assign n19478 = ~n19386 & ~n19389 ;
  assign n19380 = n19250 ^ n19241 ;
  assign n19381 = n19247 & n19380 ;
  assign n19382 = n19381 ^ n19250 ;
  assign n19393 = ~n19478 ^ n19382 ;
  assign n19377 = ~n7850 & n8745 ;
  assign n19375 = x115 & n8741 ;
  assign n19369 = x112 & n9632 ;
  assign n19368 = x114 & n9635 ;
  assign n19370 = n19369 ^ n19368 ;
  assign n19371 = n19370 ^ x62 ;
  assign n19367 = ~n7092 & n9636 ;
  assign n19372 = n19371 ^ n19367 ;
  assign n19366 = x113 & n9628 ;
  assign n19373 = n19372 ^ n19366 ;
  assign n19364 = x117 & n8744 ;
  assign n19365 = n19364 ^ x59 ;
  assign n19374 = n19373 ^ n19365 ;
  assign n19376 = n19375 ^ n19374 ;
  assign n19378 = n19377 ^ n19376 ;
  assign n19363 = x116 & n8737 ;
  assign n19379 = n19378 ^ n19363 ;
  assign n19394 = n19393 ^ n19379 ;
  assign n19360 = n19259 ^ n19235 ;
  assign n19361 = n19260 & ~n19360 ;
  assign n19353 = x118 & n7935 ;
  assign n19352 = x120 & n7938 ;
  assign n19354 = n19353 ^ n19352 ;
  assign n19355 = n19354 ^ x56 ;
  assign n19351 = n7939 & n8891 ;
  assign n19356 = n19355 ^ n19351 ;
  assign n19350 = x119 & n7931 ;
  assign n19357 = n19356 ^ n19350 ;
  assign n19358 = n19357 ^ n19259 ;
  assign n19362 = n19361 ^ n19358 ;
  assign n19395 = n19394 ^ n19362 ;
  assign n19404 = n19403 ^ n19395 ;
  assign n19347 = n19273 ^ n19269 ;
  assign n19348 = n19270 & n19347 ;
  assign n19349 = n19348 ^ n19273 ;
  assign n19405 = n19404 ^ n19349 ;
  assign n19410 = n19409 ^ n19405 ;
  assign n19412 = n19411 ^ n19410 ;
  assign n19414 = n19413 ^ n19412 ;
  assign n19344 = n19282 ^ n19232 ;
  assign n19345 = ~n19283 & n19344 ;
  assign n19346 = n19345 ^ n19282 ;
  assign n19415 = n19414 ^ n19346 ;
  assign n19418 = n19415 ^ x46 ;
  assign n19416 = n19415 ^ x47 ;
  assign n19417 = n19416 ^ n19337 ;
  assign n19419 = n19418 ^ n19417 ;
  assign n19420 = ~n19343 & n19419 ;
  assign n19421 = n19420 ^ n19418 ;
  assign n19425 = n19424 ^ n19421 ;
  assign n19333 = n19328 ^ n19294 ;
  assign n19330 = n19300 ^ n19226 ;
  assign n19334 = n19330 ^ n19294 ;
  assign n19335 = n19334 ^ n19223 ;
  assign n19336 = n19333 & ~n19335 ;
  assign n19426 = n19425 ^ n19336 ;
  assign n19331 = n19226 ^ n19223 ;
  assign n19332 = n19330 & ~n19331 ;
  assign n19427 = n19426 ^ n19332 ;
  assign n19518 = n19424 ^ n19415 ;
  assign n19519 = n19421 & ~n19518 ;
  assign n19520 = n19519 ^ n19415 ;
  assign n19515 = n19405 ^ n19346 ;
  assign n19516 = n19414 & n19515 ;
  assign n19517 = n19516 ^ n19405 ;
  assign n19521 = n19520 ^ n19517 ;
  assign n19509 = x125 & n6677 ;
  assign n19508 = x127 & n6428 ;
  assign n19510 = n19509 ^ n19508 ;
  assign n19511 = n19510 ^ x50 ;
  assign n19507 = n6429 & n10972 ;
  assign n19512 = n19511 ^ n19507 ;
  assign n19506 = x126 & n6433 ;
  assign n19513 = n19512 ^ n19506 ;
  assign n19499 = x122 & n7171 ;
  assign n19498 = x124 & n7174 ;
  assign n19500 = n19499 ^ n19498 ;
  assign n19501 = n19500 ^ x53 ;
  assign n19497 = n7175 & n10095 ;
  assign n19502 = n19501 ^ n19497 ;
  assign n19496 = x123 & n7179 ;
  assign n19503 = n19502 ^ n19496 ;
  assign n19492 = n19394 ^ n19357 ;
  assign n19493 = n19362 & n19492 ;
  assign n19494 = n19493 ^ n19357 ;
  assign n19490 = x120 & n7931 ;
  assign n19485 = x119 & n7935 ;
  assign n19484 = x121 & n7938 ;
  assign n19486 = n19485 ^ n19484 ;
  assign n19487 = n19486 ^ x56 ;
  assign n19483 = n7939 & n8962 ;
  assign n19488 = n19487 ^ n19483 ;
  assign n19479 = n19382 & n19478 ;
  assign n19480 = n19479 ^ n19389 ;
  assign n19471 = x113 & n9632 ;
  assign n19470 = x115 & n9635 ;
  assign n19472 = n19471 ^ n19470 ;
  assign n19473 = n19472 ^ x62 ;
  assign n19469 = ~n7343 & n9636 ;
  assign n19474 = n19473 ^ n19469 ;
  assign n19468 = x114 & n9628 ;
  assign n19475 = n19474 ^ n19468 ;
  assign n19476 = n19475 ^ x47 ;
  assign n19464 = x112 ^ x110 ;
  assign n19465 = ~n11875 & n19464 ;
  assign n5881 = x111 ^ x110 ;
  assign n19466 = n19465 ^ n5881 ;
  assign n19467 = n12206 & n19466 ;
  assign n19477 = n19476 ^ n19467 ;
  assign n19481 = n19480 ^ n19477 ;
  assign n19454 = x116 & n8741 ;
  assign n19453 = x118 & n8744 ;
  assign n19455 = n19454 ^ n19453 ;
  assign n19456 = n19455 ^ x59 ;
  assign n19452 = ~n8123 & n8745 ;
  assign n19457 = n19456 ^ n19452 ;
  assign n19451 = x117 & n8737 ;
  assign n19458 = n19457 ^ n19451 ;
  assign n19459 = n19458 ^ n19393 ;
  assign n19460 = n19459 ^ n19373 ;
  assign n19461 = n19460 ^ n19458 ;
  assign n19462 = ~n19379 & n19461 ;
  assign n19463 = n19462 ^ n19459 ;
  assign n19482 = n19481 ^ n19463 ;
  assign n19489 = n19488 ^ n19482 ;
  assign n19491 = n19490 ^ n19489 ;
  assign n19495 = n19494 ^ n19491 ;
  assign n19504 = n19503 ^ n19495 ;
  assign n19448 = n19395 ^ n19349 ;
  assign n19449 = n19404 & ~n19448 ;
  assign n19450 = n19449 ^ n19403 ;
  assign n19505 = n19504 ^ n19450 ;
  assign n19514 = n19513 ^ n19505 ;
  assign n19522 = n19521 ^ n19514 ;
  assign n19428 = n19223 & n19226 ;
  assign n19429 = n19428 ^ n19425 ;
  assign n19430 = n19294 & ~n19300 ;
  assign n19431 = n19430 ^ n19301 ;
  assign n19432 = n19431 ^ n19328 ;
  assign n19433 = n19428 ^ n19331 ;
  assign n19434 = ~n19430 & ~n19433 ;
  assign n19435 = n19434 ^ n19425 ;
  assign n19436 = n19432 & ~n19435 ;
  assign n19437 = ~n19431 & ~n19436 ;
  assign n19438 = n19429 & n19437 ;
  assign n19439 = n19328 ^ n19223 ;
  assign n19440 = n19328 ^ n19226 ;
  assign n19441 = ~n19439 & ~n19440 ;
  assign n19442 = n19441 ^ n19328 ;
  assign n19443 = ~n19438 & ~n19442 ;
  assign n19445 = ~n19425 & ~n19430 ;
  assign n19446 = n19443 & n19445 ;
  assign n19444 = n19443 ^ n19438 ;
  assign n19447 = n19446 ^ n19444 ;
  assign n19523 = n19522 ^ n19447 ;
  assign n19599 = ~n19517 & ~n19520 ;
  assign n19598 = n19505 & n19513 ;
  assign n19600 = n19599 ^ n19598 ;
  assign n19593 = n6429 & n10139 ;
  assign n19592 = x126 & n6677 ;
  assign n19594 = n19593 ^ n19592 ;
  assign n19595 = n19594 ^ x50 ;
  assign n19591 = x127 & n6433 ;
  assign n19596 = n19595 ^ n19591 ;
  assign n19587 = n19503 ^ n19450 ;
  assign n19588 = n19504 & n19587 ;
  assign n19589 = n19588 ^ n19503 ;
  assign n19578 = x117 & n8741 ;
  assign n19577 = x119 & n8744 ;
  assign n19579 = n19578 ^ n19577 ;
  assign n19580 = n19579 ^ x59 ;
  assign n19576 = n8394 & n8745 ;
  assign n19581 = n19580 ^ n19576 ;
  assign n19575 = x118 & n8737 ;
  assign n19582 = n19581 ^ n19575 ;
  assign n19569 = x114 & n9632 ;
  assign n19568 = x116 & n9635 ;
  assign n19570 = n19569 ^ n19568 ;
  assign n19571 = n19570 ^ x62 ;
  assign n19567 = ~n7588 & n9636 ;
  assign n19572 = n19571 ^ n19567 ;
  assign n19566 = x115 & n9628 ;
  assign n19573 = n19572 ^ n19566 ;
  assign n19559 = x111 ^ x47 ;
  assign n19562 = n19466 & ~n19559 ;
  assign n19563 = n19562 ^ x111 ;
  assign n19564 = n12206 & n19563 ;
  assign n19555 = x63 & x112 ;
  assign n19556 = n19555 ^ x113 ;
  assign n19557 = ~n9948 & n19556 ;
  assign n19558 = n19557 ^ x113 ;
  assign n19565 = n19564 ^ n19558 ;
  assign n19574 = n19573 ^ n19565 ;
  assign n19583 = n19582 ^ n19574 ;
  assign n19550 = n19480 ^ n19475 ;
  assign n19551 = n19477 & ~n19550 ;
  assign n19552 = n19551 ^ n19480 ;
  assign n19584 = n19583 ^ n19552 ;
  assign n19547 = n7939 & ~n9247 ;
  assign n19545 = x120 & n7935 ;
  assign n19541 = n19481 ^ n19458 ;
  assign n19542 = n19463 & n19541 ;
  assign n19543 = n19542 ^ n19458 ;
  assign n19539 = x122 & n7938 ;
  assign n19540 = n19539 ^ x56 ;
  assign n19544 = n19543 ^ n19540 ;
  assign n19546 = n19545 ^ n19544 ;
  assign n19548 = n19547 ^ n19546 ;
  assign n19538 = x121 & n7931 ;
  assign n19549 = n19548 ^ n19538 ;
  assign n19585 = n19584 ^ n19549 ;
  assign n19535 = n7175 & n10400 ;
  assign n19533 = x123 & n7171 ;
  assign n19529 = n19494 ^ n19482 ;
  assign n19530 = n19491 & n19529 ;
  assign n19531 = n19530 ^ n19482 ;
  assign n19527 = x125 & n7174 ;
  assign n19528 = n19527 ^ x53 ;
  assign n19532 = n19531 ^ n19528 ;
  assign n19534 = n19533 ^ n19532 ;
  assign n19536 = n19535 ^ n19534 ;
  assign n19526 = x124 & n7179 ;
  assign n19537 = n19536 ^ n19526 ;
  assign n19586 = n19585 ^ n19537 ;
  assign n19590 = n19589 ^ n19586 ;
  assign n19597 = n19596 ^ n19590 ;
  assign n19601 = n19600 ^ n19597 ;
  assign n19524 = n19514 ^ n19447 ;
  assign n19525 = n19522 & n19524 ;
  assign n19602 = n19601 ^ n19525 ;
  assign n19689 = n19582 ^ n19552 ;
  assign n19690 = ~n19583 & ~n19689 ;
  assign n19691 = n19690 ^ n19582 ;
  assign n19683 = x121 & n7935 ;
  assign n19682 = x123 & n7938 ;
  assign n19684 = n19683 ^ n19682 ;
  assign n19685 = n19684 ^ x56 ;
  assign n19681 = n7939 & ~n9786 ;
  assign n19686 = n19685 ^ n19681 ;
  assign n19680 = x122 & n7931 ;
  assign n19687 = n19686 ^ n19680 ;
  assign n19674 = x118 & n8741 ;
  assign n19673 = x120 & n8744 ;
  assign n19675 = n19674 ^ n19673 ;
  assign n19676 = n19675 ^ x59 ;
  assign n19672 = n8745 & n8891 ;
  assign n19677 = n19676 ^ n19672 ;
  assign n19671 = x119 & n8737 ;
  assign n19678 = n19677 ^ n19671 ;
  assign n19666 = n19573 ^ n19558 ;
  assign n19667 = n19565 & ~n19666 ;
  assign n19668 = n19667 ^ n19573 ;
  assign n19662 = ~n7850 & n9636 ;
  assign n19661 = x116 & n9628 ;
  assign n19663 = n19662 ^ n19661 ;
  assign n19659 = x115 & n9632 ;
  assign n19658 = x117 & n9635 ;
  assign n19660 = n19659 ^ n19658 ;
  assign n19664 = n19663 ^ n19660 ;
  assign n6582 = x114 ^ x113 ;
  assign n19657 = n6582 ^ x62 ;
  assign n19665 = n19664 ^ n19657 ;
  assign n19669 = n19668 ^ n19665 ;
  assign n6339 = x113 ^ x112 ;
  assign n19654 = x63 & n6339 ;
  assign n19655 = n19654 ^ n6582 ;
  assign n19656 = ~n9948 & n19655 ;
  assign n19670 = n19669 ^ n19656 ;
  assign n19679 = n19678 ^ n19670 ;
  assign n19688 = n19687 ^ n19679 ;
  assign n19692 = n19691 ^ n19688 ;
  assign n19648 = x125 & n7179 ;
  assign n19646 = n7175 & n10441 ;
  assign n19644 = x124 & n7171 ;
  assign n19640 = n19584 ^ n19543 ;
  assign n19641 = ~n19549 & n19640 ;
  assign n19642 = n19641 ^ n19584 ;
  assign n19638 = x126 & n7174 ;
  assign n19639 = n19638 ^ x53 ;
  assign n19643 = n19642 ^ n19639 ;
  assign n19645 = n19644 ^ n19643 ;
  assign n19647 = n19646 ^ n19645 ;
  assign n19649 = n19648 ^ n19647 ;
  assign n19693 = n19692 ^ n19649 ;
  assign n19635 = n19596 ^ n19589 ;
  assign n19636 = ~n19590 & n19635 ;
  assign n19637 = n19636 ^ n19596 ;
  assign n19694 = n19693 ^ n19637 ;
  assign n19631 = n19585 ^ n19531 ;
  assign n19632 = ~n19537 & n19631 ;
  assign n19633 = n19632 ^ n19585 ;
  assign n19621 = x127 & n6676 ;
  assign n19622 = n19621 ^ n6427 ;
  assign n19627 = n5972 & n11265 ;
  assign n19628 = n19627 ^ n19621 ;
  assign n19629 = n19622 & ~n19628 ;
  assign n19630 = n19629 ^ x49 ;
  assign n19634 = n19633 ^ n19630 ;
  assign n19695 = n19694 ^ n19634 ;
  assign n19603 = n19597 ^ n19521 ;
  assign n19604 = n19603 ^ n19599 ;
  assign n19610 = ~n19447 & ~n19599 ;
  assign n19605 = n19598 ^ n19514 ;
  assign n19606 = n19605 ^ n19517 ;
  assign n19607 = n19521 & n19606 ;
  assign n19608 = n19607 ^ n19517 ;
  assign n19609 = n19597 & n19608 ;
  assign n19611 = n19598 ^ n19597 ;
  assign n19612 = ~n19609 & n19611 ;
  assign n19613 = n19610 & n19612 ;
  assign n19614 = n19613 ^ n19609 ;
  assign n19615 = n19505 ^ n19447 ;
  assign n19616 = n19514 & ~n19615 ;
  assign n19617 = n19616 ^ n19505 ;
  assign n19618 = ~n19614 & n19617 ;
  assign n19619 = ~n19604 & n19618 ;
  assign n19620 = n19619 ^ n19614 ;
  assign n19696 = n19695 ^ n19620 ;
  assign n19782 = n19637 & ~n19693 ;
  assign n19781 = ~n19630 & ~n19633 ;
  assign n19783 = n19782 ^ n19781 ;
  assign n19777 = n19692 ^ n19642 ;
  assign n19778 = ~n19649 & ~n19777 ;
  assign n19779 = n19778 ^ n19692 ;
  assign n19771 = x125 & n7171 ;
  assign n19770 = x127 & n7174 ;
  assign n19772 = n19771 ^ n19770 ;
  assign n19773 = n19772 ^ x53 ;
  assign n19769 = n7175 & n10972 ;
  assign n19774 = n19773 ^ n19769 ;
  assign n19768 = x126 & n7179 ;
  assign n19775 = n19774 ^ n19768 ;
  assign n19761 = x122 & n7935 ;
  assign n19760 = x124 & n7938 ;
  assign n19762 = n19761 ^ n19760 ;
  assign n19763 = n19762 ^ x56 ;
  assign n19759 = n7939 & n10095 ;
  assign n19764 = n19763 ^ n19759 ;
  assign n19758 = x123 & n7931 ;
  assign n19765 = n19764 ^ n19758 ;
  assign n19743 = x114 ^ x63 ;
  assign n19744 = n19743 ^ n19664 ;
  assign n19747 = n6582 & ~n19744 ;
  assign n19748 = n19747 ^ n19664 ;
  assign n19749 = n9948 & n19748 ;
  assign n19732 = x113 & ~x114 ;
  assign n19734 = n19732 ^ x112 ;
  assign n19733 = n19732 ^ n19664 ;
  assign n19735 = n19734 ^ n19733 ;
  assign n19738 = ~n6339 & n19735 ;
  assign n19739 = n19738 ^ n19734 ;
  assign n19740 = x62 & n19739 ;
  assign n19741 = n19740 ^ n19732 ;
  assign n19742 = x63 & n19741 ;
  assign n19750 = n19749 ^ x62 ;
  assign n19751 = ~n19742 & ~n19750 ;
  assign n19752 = n19664 & n19751 ;
  assign n19753 = ~n19749 & n19752 ;
  assign n19754 = n19753 ^ n19751 ;
  assign n19755 = n19754 ^ n19742 ;
  assign n19726 = x116 & n9632 ;
  assign n19725 = x118 & n9635 ;
  assign n19727 = n19726 ^ n19725 ;
  assign n19728 = n19727 ^ x62 ;
  assign n19724 = ~n8123 & n9636 ;
  assign n19729 = n19728 ^ n19724 ;
  assign n19723 = x117 & n9628 ;
  assign n19730 = n19729 ^ n19723 ;
  assign n19717 = x63 & x114 ;
  assign n19718 = n19717 ^ x115 ;
  assign n19719 = ~n9948 & n19718 ;
  assign n19720 = n19719 ^ x115 ;
  assign n19721 = n19720 ^ x50 ;
  assign n19722 = n19721 ^ n19558 ;
  assign n19731 = n19730 ^ n19722 ;
  assign n19756 = n19755 ^ n19731 ;
  assign n19705 = x119 & n8741 ;
  assign n19704 = x121 & n8744 ;
  assign n19706 = n19705 ^ n19704 ;
  assign n19707 = n19706 ^ x59 ;
  assign n19703 = n8745 & n8962 ;
  assign n19708 = n19707 ^ n19703 ;
  assign n19702 = x120 & n8737 ;
  assign n19709 = n19708 ^ n19702 ;
  assign n19710 = n19709 ^ n19678 ;
  assign n19711 = n19710 ^ n19668 ;
  assign n19712 = n19711 ^ n19709 ;
  assign n19713 = n19670 & n19712 ;
  assign n19714 = n19713 ^ n19710 ;
  assign n19757 = n19756 ^ n19714 ;
  assign n19766 = n19765 ^ n19757 ;
  assign n19699 = n19691 ^ n19687 ;
  assign n19700 = n19688 & n19699 ;
  assign n19701 = n19700 ^ n19691 ;
  assign n19767 = n19766 ^ n19701 ;
  assign n19776 = n19775 ^ n19767 ;
  assign n19780 = n19779 ^ n19776 ;
  assign n19784 = n19783 ^ n19780 ;
  assign n19697 = n19634 ^ n19620 ;
  assign n19698 = ~n19695 & n19697 ;
  assign n19785 = n19784 ^ n19698 ;
  assign n19856 = n7175 & n10139 ;
  assign n19855 = x126 & n7171 ;
  assign n19857 = n19856 ^ n19855 ;
  assign n19858 = n19857 ^ x53 ;
  assign n19854 = x127 & n7179 ;
  assign n19859 = n19858 ^ n19854 ;
  assign n19850 = n19765 ^ n19701 ;
  assign n19851 = n19766 & n19850 ;
  assign n19852 = n19851 ^ n19765 ;
  assign n19842 = x120 & n8741 ;
  assign n19841 = x122 & n8744 ;
  assign n19843 = n19842 ^ n19841 ;
  assign n19844 = n19843 ^ x59 ;
  assign n19840 = n8745 & ~n9247 ;
  assign n19845 = n19844 ^ n19840 ;
  assign n19839 = x121 & n8737 ;
  assign n19846 = n19845 ^ n19839 ;
  assign n19836 = x115 & n11875 ;
  assign n19835 = x116 & n9948 ;
  assign n19837 = n19836 ^ n19835 ;
  assign n19832 = n8394 & n9636 ;
  assign n19830 = x117 & n9632 ;
  assign n19826 = n19720 ^ n19558 ;
  assign n19827 = ~n19721 & ~n19826 ;
  assign n19828 = n19827 ^ x50 ;
  assign n19824 = x119 & n9635 ;
  assign n19825 = n19824 ^ x62 ;
  assign n19829 = n19828 ^ n19825 ;
  assign n19831 = n19830 ^ n19829 ;
  assign n19833 = n19832 ^ n19831 ;
  assign n19823 = x118 & n9628 ;
  assign n19834 = n19833 ^ n19823 ;
  assign n19838 = n19837 ^ n19834 ;
  assign n19847 = n19846 ^ n19838 ;
  assign n19820 = n19755 ^ n19730 ;
  assign n19821 = n19731 & ~n19820 ;
  assign n19822 = n19821 ^ n19755 ;
  assign n19848 = n19847 ^ n19822 ;
  assign n19810 = x123 & n7935 ;
  assign n19809 = x125 & n7938 ;
  assign n19811 = n19810 ^ n19809 ;
  assign n19812 = n19811 ^ x56 ;
  assign n19808 = n7939 & n10400 ;
  assign n19813 = n19812 ^ n19808 ;
  assign n19807 = x124 & n7931 ;
  assign n19814 = n19813 ^ n19807 ;
  assign n19816 = n19814 ^ n19709 ;
  assign n19815 = n19814 ^ n19756 ;
  assign n19817 = n19816 ^ n19815 ;
  assign n19818 = n19714 & n19817 ;
  assign n19819 = n19818 ^ n19816 ;
  assign n19849 = n19848 ^ n19819 ;
  assign n19853 = n19852 ^ n19849 ;
  assign n19860 = n19859 ^ n19853 ;
  assign n19804 = n19779 ^ n19775 ;
  assign n19805 = ~n19776 & ~n19804 ;
  assign n19806 = n19805 ^ n19779 ;
  assign n19861 = n19860 ^ n19806 ;
  assign n19786 = n19780 ^ n19694 ;
  assign n19787 = n19786 ^ n19782 ;
  assign n19793 = ~n19620 & ~n19782 ;
  assign n19788 = n19781 ^ n19634 ;
  assign n19789 = n19788 ^ n19693 ;
  assign n19790 = ~n19694 & n19789 ;
  assign n19791 = n19790 ^ n19693 ;
  assign n19792 = n19780 & n19791 ;
  assign n19794 = n19781 ^ n19780 ;
  assign n19795 = ~n19792 & n19794 ;
  assign n19796 = n19793 & n19795 ;
  assign n19797 = n19796 ^ n19792 ;
  assign n19798 = n19630 ^ n19620 ;
  assign n19799 = n19634 & n19798 ;
  assign n19800 = n19799 ^ n19630 ;
  assign n19801 = ~n19797 & ~n19800 ;
  assign n19802 = n19787 & n19801 ;
  assign n19803 = n19802 ^ n19797 ;
  assign n19862 = n19861 ^ n19803 ;
  assign n19920 = x124 & n7935 ;
  assign n19919 = x126 & n7938 ;
  assign n19921 = n19920 ^ n19919 ;
  assign n19922 = n19921 ^ x56 ;
  assign n19918 = n7939 & n10441 ;
  assign n19923 = n19922 ^ n19918 ;
  assign n19917 = x125 & n7931 ;
  assign n19924 = n19923 ^ n19917 ;
  assign n19909 = n9948 ^ x116 ;
  assign n19906 = ~x117 & n9948 ;
  assign n19907 = n19906 ^ n19836 ;
  assign n19910 = n19907 ^ n12206 ;
  assign n19911 = n19909 & n19910 ;
  assign n19912 = n19911 ^ n19836 ;
  assign n19908 = x116 & n19907 ;
  assign n19913 = n19912 ^ n19908 ;
  assign n19903 = n19837 ^ n19828 ;
  assign n19904 = n19834 & n19903 ;
  assign n19905 = n19904 ^ n19837 ;
  assign n19914 = n19913 ^ n19905 ;
  assign n19900 = n8745 & ~n9786 ;
  assign n19898 = x121 & n8741 ;
  assign n19892 = x118 & n9632 ;
  assign n19891 = x120 & n9635 ;
  assign n19893 = n19892 ^ n19891 ;
  assign n19894 = n19893 ^ x62 ;
  assign n19890 = n8891 & n9636 ;
  assign n19895 = n19894 ^ n19890 ;
  assign n19889 = x119 & n9628 ;
  assign n19896 = n19895 ^ n19889 ;
  assign n19887 = x123 & n8744 ;
  assign n19888 = n19887 ^ x59 ;
  assign n19897 = n19896 ^ n19888 ;
  assign n19899 = n19898 ^ n19897 ;
  assign n19901 = n19900 ^ n19899 ;
  assign n19886 = x122 & n8737 ;
  assign n19902 = n19901 ^ n19886 ;
  assign n19915 = n19914 ^ n19902 ;
  assign n19883 = n19838 ^ n19822 ;
  assign n19884 = n19847 & n19883 ;
  assign n19885 = n19884 ^ n19846 ;
  assign n19916 = n19915 ^ n19885 ;
  assign n19925 = n19924 ^ n19916 ;
  assign n19873 = x127 & n7170 ;
  assign n19874 = n19873 ^ n7168 ;
  assign n19879 = n6670 & n11265 ;
  assign n19880 = n19879 ^ n19873 ;
  assign n19881 = n19874 & ~n19880 ;
  assign n19882 = n19881 ^ x52 ;
  assign n19926 = n19925 ^ n19882 ;
  assign n19870 = n19848 ^ n19814 ;
  assign n19871 = n19819 & ~n19870 ;
  assign n19872 = n19871 ^ n19814 ;
  assign n19927 = n19926 ^ n19872 ;
  assign n19867 = n19859 ^ n19852 ;
  assign n19868 = n19853 & n19867 ;
  assign n19869 = n19868 ^ n19859 ;
  assign n19928 = n19927 ^ n19869 ;
  assign n19863 = n19806 ^ n19803 ;
  assign n19864 = n19860 ^ n19803 ;
  assign n19865 = ~n19863 & n19864 ;
  assign n19866 = n19865 ^ n19860 ;
  assign n19929 = n19928 ^ n19866 ;
  assign n19977 = n19924 ^ n19885 ;
  assign n19978 = ~n19916 & n19977 ;
  assign n19979 = n19978 ^ n19924 ;
  assign n19974 = n19882 ^ n19872 ;
  assign n19975 = n19926 & n19974 ;
  assign n19976 = n19975 ^ n19882 ;
  assign n19980 = n19979 ^ n19976 ;
  assign n19968 = x125 & n7935 ;
  assign n19967 = x127 & n7938 ;
  assign n19969 = n19968 ^ n19967 ;
  assign n19970 = n19969 ^ x56 ;
  assign n19966 = n7939 & n10972 ;
  assign n19971 = n19970 ^ n19966 ;
  assign n19965 = x126 & n7931 ;
  assign n19972 = n19971 ^ n19965 ;
  assign n19956 = x119 & n9632 ;
  assign n19955 = x121 & n9635 ;
  assign n19957 = n19956 ^ n19955 ;
  assign n19958 = n19957 ^ x62 ;
  assign n19954 = n8962 & n9636 ;
  assign n19959 = n19958 ^ n19954 ;
  assign n19953 = x120 & n9628 ;
  assign n19960 = n19959 ^ n19953 ;
  assign n19961 = n19960 ^ x53 ;
  assign n19949 = x118 ^ x116 ;
  assign n19950 = ~n11875 & n19949 ;
  assign n7322 = x117 ^ x116 ;
  assign n19951 = n19950 ^ n7322 ;
  assign n19952 = n12206 & n19951 ;
  assign n19962 = n19961 ^ n19952 ;
  assign n19947 = n19905 & ~n19913 ;
  assign n19948 = n19947 ^ n19911 ;
  assign n19963 = n19962 ^ n19948 ;
  assign n19937 = x122 & n8741 ;
  assign n19936 = x124 & n8744 ;
  assign n19938 = n19937 ^ n19936 ;
  assign n19939 = n19938 ^ x59 ;
  assign n19935 = n8745 & n10095 ;
  assign n19940 = n19939 ^ n19935 ;
  assign n19934 = x123 & n8737 ;
  assign n19941 = n19940 ^ n19934 ;
  assign n19942 = n19941 ^ n19914 ;
  assign n19943 = n19942 ^ n19896 ;
  assign n19944 = n19943 ^ n19941 ;
  assign n19945 = ~n19902 & n19944 ;
  assign n19946 = n19945 ^ n19942 ;
  assign n19964 = n19963 ^ n19946 ;
  assign n19973 = n19972 ^ n19964 ;
  assign n19981 = n19980 ^ n19973 ;
  assign n19930 = n19927 ^ n19866 ;
  assign n19931 = n19869 ^ n19866 ;
  assign n19932 = ~n19930 & n19931 ;
  assign n19933 = n19932 ^ n19927 ;
  assign n19982 = n19981 ^ n19933 ;
  assign n19983 = n19979 ^ n19972 ;
  assign n19986 = ~n19973 & n19983 ;
  assign n19984 = n19976 ^ n19973 ;
  assign n19988 = n19986 ^ n19984 ;
  assign n19989 = ~n19933 & ~n19988 ;
  assign n19996 = n19989 ^ n19986 ;
  assign n19990 = n19989 ^ n19976 ;
  assign n19992 = n19976 ^ n19972 ;
  assign n19993 = n19992 ^ n19973 ;
  assign n19994 = n19993 ^ n19983 ;
  assign n19995 = n19990 & ~n19994 ;
  assign n19997 = n19996 ^ n19995 ;
  assign n19998 = n19997 ^ n19984 ;
  assign n20048 = ~n19964 & ~n19972 ;
  assign n20049 = n20048 ^ n19973 ;
  assign n20050 = ~n19933 & n20049 ;
  assign n20051 = n20048 ^ n19976 ;
  assign n20052 = n20048 ^ n19979 ;
  assign n20053 = n20051 & ~n20052 ;
  assign n20054 = n20053 ^ n19979 ;
  assign n20055 = n20050 & ~n20054 ;
  assign n20056 = n19998 & n20055 ;
  assign n20041 = n7939 & n10139 ;
  assign n20040 = x126 & n7935 ;
  assign n20042 = n20041 ^ n20040 ;
  assign n20043 = n20042 ^ x56 ;
  assign n20039 = x127 & n7931 ;
  assign n20044 = n20043 ^ n20039 ;
  assign n20027 = x120 & n9632 ;
  assign n20026 = x122 & n9635 ;
  assign n20028 = n20027 ^ n20026 ;
  assign n20029 = n20028 ^ x62 ;
  assign n20025 = ~n9247 & n9636 ;
  assign n20030 = n20029 ^ n20025 ;
  assign n20024 = x121 & n9628 ;
  assign n20031 = n20030 ^ n20024 ;
  assign n20019 = x63 & x118 ;
  assign n20020 = n20019 ^ x119 ;
  assign n20021 = ~n9948 & n20020 ;
  assign n20022 = n20021 ^ x119 ;
  assign n20011 = x117 ^ x53 ;
  assign n20014 = n19951 & ~n20011 ;
  assign n20015 = n20014 ^ x117 ;
  assign n20016 = n12206 & n20015 ;
  assign n20023 = n20022 ^ n20016 ;
  assign n20032 = n20031 ^ n20023 ;
  assign n20009 = x124 & n8737 ;
  assign n20007 = n8745 & n10400 ;
  assign n20005 = x123 & n8741 ;
  assign n20001 = n19960 ^ n19948 ;
  assign n20002 = ~n19962 & ~n20001 ;
  assign n20003 = n20002 ^ n19960 ;
  assign n19999 = x125 & n8744 ;
  assign n20000 = n19999 ^ x59 ;
  assign n20004 = n20003 ^ n20000 ;
  assign n20006 = n20005 ^ n20004 ;
  assign n20008 = n20007 ^ n20006 ;
  assign n20010 = n20009 ^ n20008 ;
  assign n20033 = n20032 ^ n20010 ;
  assign n20035 = n20033 ^ n19941 ;
  assign n20034 = n20033 ^ n19963 ;
  assign n20036 = n20035 ^ n20034 ;
  assign n20037 = n19946 & n20036 ;
  assign n20038 = n20037 ^ n20035 ;
  assign n20045 = n20044 ^ n20038 ;
  assign n20046 = n20045 ^ n19998 ;
  assign n20057 = n20056 ^ n20046 ;
  assign n20155 = n20044 ^ n20033 ;
  assign n20156 = ~n20038 & ~n20155 ;
  assign n20157 = n20156 ^ n20033 ;
  assign n20149 = x124 & n8741 ;
  assign n20148 = x126 & n8744 ;
  assign n20150 = n20149 ^ n20148 ;
  assign n20151 = n20150 ^ x59 ;
  assign n20147 = n8745 & n10441 ;
  assign n20152 = n20151 ^ n20147 ;
  assign n20146 = x125 & n8737 ;
  assign n20153 = n20152 ^ n20146 ;
  assign n20139 = x121 & n9632 ;
  assign n20138 = x123 & n9635 ;
  assign n20140 = n20139 ^ n20138 ;
  assign n20141 = n20140 ^ x62 ;
  assign n20137 = n9636 & ~n9786 ;
  assign n20142 = n20141 ^ n20137 ;
  assign n20136 = x122 & n9628 ;
  assign n20143 = n20142 ^ n20136 ;
  assign n20132 = x63 & n7825 ;
  assign n20133 = n20132 ^ n8100 ;
  assign n20134 = ~n9948 & n20133 ;
  assign n20135 = n20134 ^ n8100 ;
  assign n20144 = n20143 ^ n20135 ;
  assign n20125 = n20031 ^ n20022 ;
  assign n20126 = n20023 & ~n20125 ;
  assign n20127 = n20126 ^ n20031 ;
  assign n20145 = n20144 ^ n20127 ;
  assign n20154 = n20153 ^ n20145 ;
  assign n20158 = n20157 ^ n20154 ;
  assign n20121 = n20032 ^ n20003 ;
  assign n20122 = ~n20010 & ~n20121 ;
  assign n20123 = n20122 ^ n20032 ;
  assign n7940 = n7939 ^ n7935 ;
  assign n20118 = x127 & n7940 ;
  assign n20117 = n7939 & n10138 ;
  assign n20119 = n20118 ^ n20117 ;
  assign n20120 = n20119 ^ x56 ;
  assign n20124 = n20123 ^ n20120 ;
  assign n20159 = n20158 ^ n20124 ;
  assign n20061 = ~n19976 & ~n19979 ;
  assign n20113 = n20061 ^ n19980 ;
  assign n20058 = ~n20048 & ~n20050 ;
  assign n20067 = n20049 ^ n19933 ;
  assign n20065 = n20061 ^ n20049 ;
  assign n20059 = n20054 ^ n20045 ;
  assign n20066 = n20065 ^ n20059 ;
  assign n20103 = n20067 ^ n20066 ;
  assign n20060 = n20059 ^ n20049 ;
  assign n20104 = n20103 ^ n20060 ;
  assign n20105 = n20104 ^ n20054 ;
  assign n20107 = n20105 ^ n20103 ;
  assign n20076 = n20067 ^ n20045 ;
  assign n20089 = n20076 ^ n20049 ;
  assign n20080 = n20065 ^ n20054 ;
  assign n20092 = n20089 ^ n20080 ;
  assign n20088 = n20054 ^ n20049 ;
  assign n20093 = n20092 ^ n20088 ;
  assign n20094 = n20093 ^ n20059 ;
  assign n20096 = n20094 ^ n20092 ;
  assign n20077 = n20076 ^ n20061 ;
  assign n20078 = n20045 & n20059 ;
  assign n20081 = n20080 ^ n20078 ;
  assign n20082 = n20076 ^ n20059 ;
  assign n20083 = n20082 ^ n20078 ;
  assign n20084 = n20081 & ~n20083 ;
  assign n20085 = n19933 & n20084 ;
  assign n20086 = ~n20077 & ~n20085 ;
  assign n20087 = n20086 ^ n20078 ;
  assign n20097 = n20096 ^ n20087 ;
  assign n20098 = n20097 ^ n20076 ;
  assign n20099 = n20098 ^ n20094 ;
  assign n20068 = n20067 ^ n20059 ;
  assign n20075 = n20068 ^ n20045 ;
  assign n20100 = n20099 ^ n20075 ;
  assign n20069 = n20068 ^ n20066 ;
  assign n20101 = n20100 ^ n20069 ;
  assign n20108 = n20107 ^ n20101 ;
  assign n20109 = n20108 ^ n20045 ;
  assign n20110 = n20109 ^ n20105 ;
  assign n20111 = n20058 & n20110 ;
  assign n20114 = n20045 & n20111 ;
  assign n20115 = n20113 & n20114 ;
  assign n20112 = n20111 ^ n20110 ;
  assign n20116 = n20115 ^ n20112 ;
  assign n20160 = n20159 ^ n20116 ;
  assign n20209 = ~n20135 & n20143 ;
  assign n20203 = n9948 ^ x119 ;
  assign n20204 = x63 & ~x118 ;
  assign n20205 = n20204 ^ x120 ;
  assign n20206 = x119 & n20205 ;
  assign n20207 = n20206 ^ x120 ;
  assign n20208 = n20203 & n20207 ;
  assign n20210 = n20209 ^ n20208 ;
  assign n20197 = x122 & n9632 ;
  assign n20196 = x124 & n9635 ;
  assign n20198 = n20197 ^ n20196 ;
  assign n20199 = n20198 ^ x62 ;
  assign n20195 = n9636 & n10095 ;
  assign n20200 = n20199 ^ n20195 ;
  assign n20194 = x123 & n9628 ;
  assign n20201 = n20200 ^ n20194 ;
  assign n20188 = x63 & x120 ;
  assign n20189 = n20188 ^ x121 ;
  assign n20190 = ~n9948 & n20189 ;
  assign n20191 = n20190 ^ x121 ;
  assign n20192 = n20191 ^ x56 ;
  assign n20193 = n20192 ^ n20022 ;
  assign n20202 = n20201 ^ n20193 ;
  assign n20211 = n20210 ^ n20202 ;
  assign n20176 = x125 & n8741 ;
  assign n20175 = x127 & n8744 ;
  assign n20177 = n20176 ^ n20175 ;
  assign n20178 = n20177 ^ x59 ;
  assign n20174 = n8745 & n10972 ;
  assign n20179 = n20178 ^ n20174 ;
  assign n20173 = x126 & n8737 ;
  assign n20180 = n20179 ^ n20173 ;
  assign n20181 = n20180 ^ n20153 ;
  assign n20182 = n20181 ^ n20127 ;
  assign n20183 = n20182 ^ n20180 ;
  assign n20184 = n20145 & n20183 ;
  assign n20185 = n20184 ^ n20181 ;
  assign n20212 = n20211 ^ n20185 ;
  assign n20168 = ~n20120 & n20123 ;
  assign n20169 = n20168 ^ n20154 ;
  assign n20170 = n20158 & ~n20169 ;
  assign n20171 = n20170 ^ n20157 ;
  assign n20172 = n20171 ^ n20158 ;
  assign n20213 = n20212 ^ n20172 ;
  assign n20214 = n20213 ^ n20168 ;
  assign n20165 = ~n20123 & n20124 ;
  assign n20166 = n20165 ^ n20116 ;
  assign n20167 = ~n20159 & n20166 ;
  assign n20215 = n20214 ^ n20167 ;
  assign n20332 = n8745 & n10139 ;
  assign n20331 = x126 & n8741 ;
  assign n20333 = n20332 ^ n20331 ;
  assign n20334 = n20333 ^ x59 ;
  assign n20330 = x127 & n8737 ;
  assign n20335 = n20334 ^ n20330 ;
  assign n20326 = x121 & n11875 ;
  assign n20325 = x122 & n9948 ;
  assign n20327 = n20326 ^ n20325 ;
  assign n20322 = n9636 & n10400 ;
  assign n20320 = x123 & n9632 ;
  assign n20316 = n20191 ^ n20022 ;
  assign n20317 = ~n20192 & ~n20316 ;
  assign n20318 = n20317 ^ x56 ;
  assign n20314 = x125 & n9635 ;
  assign n20315 = n20314 ^ x62 ;
  assign n20319 = n20318 ^ n20315 ;
  assign n20321 = n20320 ^ n20319 ;
  assign n20323 = n20322 ^ n20321 ;
  assign n20313 = x124 & n9628 ;
  assign n20324 = n20323 ^ n20313 ;
  assign n20328 = n20327 ^ n20324 ;
  assign n20310 = n20210 ^ n20201 ;
  assign n20311 = n20202 & n20310 ;
  assign n20312 = n20311 ^ n20210 ;
  assign n20329 = n20328 ^ n20312 ;
  assign n20336 = n20335 ^ n20329 ;
  assign n20307 = n20211 ^ n20180 ;
  assign n20308 = n20185 & ~n20307 ;
  assign n20309 = n20308 ^ n20180 ;
  assign n20337 = n20336 ^ n20309 ;
  assign n20217 = n20154 & n20157 ;
  assign n20303 = n20217 ^ n20158 ;
  assign n20216 = n20168 ^ n20124 ;
  assign n20224 = n20216 ^ n20116 ;
  assign n20219 = n20212 ^ n20171 ;
  assign n20218 = n20217 ^ n20216 ;
  assign n20220 = n20219 ^ n20218 ;
  assign n20290 = n20224 ^ n20220 ;
  assign n20240 = n20219 ^ n20216 ;
  assign n20291 = n20290 ^ n20240 ;
  assign n20292 = n20291 ^ n20171 ;
  assign n20294 = n20292 ^ n20290 ;
  assign n20279 = n20240 ^ n20224 ;
  assign n20280 = n20279 ^ n20220 ;
  assign n20281 = n20280 ^ n20171 ;
  assign n20283 = n20281 ^ n20279 ;
  assign n20254 = n20171 & n20219 ;
  assign n20225 = n20224 ^ n20219 ;
  assign n20235 = n20225 ^ n20217 ;
  assign n20236 = n20235 ^ n20219 ;
  assign n20255 = n20254 ^ n20236 ;
  assign n20256 = n20255 ^ n20216 ;
  assign n20257 = n20256 ^ n20212 ;
  assign n20241 = n20240 ^ n20116 ;
  assign n20242 = n20241 ^ n20219 ;
  assign n20250 = n20242 ^ n20236 ;
  assign n20258 = n20250 ^ n20216 ;
  assign n20259 = n20258 ^ n20212 ;
  assign n20260 = n20257 & ~n20259 ;
  assign n20243 = n20242 ^ n20235 ;
  assign n20245 = n20243 ^ n20216 ;
  assign n20261 = n20245 ^ n20242 ;
  assign n20247 = n20245 ^ n20212 ;
  assign n20262 = n20261 ^ n20247 ;
  assign n20263 = n20245 ^ n20236 ;
  assign n20264 = n20263 ^ n20247 ;
  assign n20265 = ~n20262 & ~n20264 ;
  assign n20266 = n20260 & n20265 ;
  assign n20267 = n20266 ^ n20254 ;
  assign n20268 = n20267 ^ n20250 ;
  assign n20248 = n20247 ^ n20243 ;
  assign n20269 = n20268 ^ n20248 ;
  assign n20270 = n20269 ^ n20116 ;
  assign n20271 = n20270 ^ n20247 ;
  assign n20284 = n20283 ^ n20271 ;
  assign n20221 = n20220 ^ n20116 ;
  assign n20273 = n20225 ^ n20221 ;
  assign n20285 = n20284 ^ n20273 ;
  assign n20286 = n20285 ^ n20281 ;
  assign n20222 = n20221 ^ n20219 ;
  assign n20223 = n20222 ^ n20219 ;
  assign n20229 = n20224 ^ n20223 ;
  assign n20231 = n20229 ^ n20218 ;
  assign n20233 = n20231 ^ n20212 ;
  assign n20234 = n20233 ^ n20229 ;
  assign n20287 = n20286 ^ n20234 ;
  assign n20288 = n20287 ^ n20233 ;
  assign n20226 = n20225 ^ n20220 ;
  assign n20289 = n20288 ^ n20226 ;
  assign n20295 = n20294 ^ n20289 ;
  assign n20296 = n20295 ^ n20212 ;
  assign n20297 = n20296 ^ n20292 ;
  assign n20298 = n20120 ^ n20116 ;
  assign n20299 = ~n20124 & ~n20298 ;
  assign n20300 = n20299 ^ n20120 ;
  assign n20301 = n20297 & n20300 ;
  assign n20304 = n20212 & n20301 ;
  assign n20305 = n20303 & n20304 ;
  assign n20302 = n20301 ^ n20297 ;
  assign n20306 = n20305 ^ n20302 ;
  assign n20338 = n20337 ^ n20306 ;
  assign n8746 = n8745 ^ n8741 ;
  assign n20367 = x127 & n8746 ;
  assign n20366 = n8745 & n10138 ;
  assign n20368 = n20367 ^ n20366 ;
  assign n20369 = n20368 ^ x59 ;
  assign n20363 = n20335 ^ n20312 ;
  assign n20364 = ~n20329 & n20363 ;
  assign n20365 = n20364 ^ n20335 ;
  assign n20370 = n20369 ^ n20365 ;
  assign n20357 = x124 & n9632 ;
  assign n20356 = x126 & n9635 ;
  assign n20358 = n20357 ^ n20356 ;
  assign n20359 = n20358 ^ x62 ;
  assign n20355 = n9636 & n10441 ;
  assign n20360 = n20359 ^ n20355 ;
  assign n20354 = x125 & n9628 ;
  assign n20361 = n20360 ^ n20354 ;
  assign n20348 = n9948 ^ x122 ;
  assign n20345 = ~x123 & n9948 ;
  assign n20346 = n20345 ^ n20326 ;
  assign n20349 = n20346 ^ n12206 ;
  assign n20350 = n20348 & n20349 ;
  assign n20351 = n20350 ^ n20326 ;
  assign n20347 = x122 & n20346 ;
  assign n20352 = n20351 ^ n20347 ;
  assign n20342 = n20327 ^ n20318 ;
  assign n20343 = n20324 & n20342 ;
  assign n20344 = n20343 ^ n20327 ;
  assign n20353 = n20352 ^ n20344 ;
  assign n20362 = n20361 ^ n20353 ;
  assign n20371 = n20370 ^ n20362 ;
  assign n20339 = n20309 ^ n20306 ;
  assign n20340 = n20337 & ~n20339 ;
  assign n20341 = n20340 ^ n20309 ;
  assign n20372 = n20371 ^ n20341 ;
  assign n20387 = x125 & n9632 ;
  assign n20386 = x127 & n9635 ;
  assign n20388 = n20387 ^ n20386 ;
  assign n20389 = n20388 ^ x62 ;
  assign n20385 = n9636 & n10972 ;
  assign n20390 = n20389 ^ n20385 ;
  assign n20384 = x126 & n9628 ;
  assign n20391 = n20390 ^ n20384 ;
  assign n20392 = n20391 ^ x59 ;
  assign n20380 = x124 ^ x122 ;
  assign n20381 = ~n11875 & n20380 ;
  assign n20382 = n20381 ^ n8944 ;
  assign n20383 = n12206 & n20382 ;
  assign n20393 = n20392 ^ n20383 ;
  assign n20378 = n20344 & ~n20352 ;
  assign n20379 = n20378 ^ n20350 ;
  assign n20394 = n20393 ^ n20379 ;
  assign n20375 = n20370 ^ n20353 ;
  assign n20376 = n20375 ^ n20341 ;
  assign n20377 = ~n20362 & n20376 ;
  assign n20395 = n20394 ^ n20377 ;
  assign n20373 = n20365 ^ n20341 ;
  assign n20374 = ~n20370 & ~n20373 ;
  assign n20396 = n20395 ^ n20374 ;
  assign n20419 = n20394 ^ n20365 ;
  assign n20420 = n20419 ^ n20369 ;
  assign n20425 = ~n20353 & ~n20361 ;
  assign n20426 = n20420 & ~n20425 ;
  assign n20422 = n20394 ^ n20362 ;
  assign n20423 = ~n20369 & n20422 ;
  assign n20424 = ~n20370 & n20423 ;
  assign n20427 = n20426 ^ n20424 ;
  assign n20428 = n20427 ^ n20422 ;
  assign n20429 = n20341 & n20428 ;
  assign n20433 = n20353 & n20365 ;
  assign n20434 = n20433 ^ n20394 ;
  assign n20442 = n20365 ^ n20353 ;
  assign n20443 = n20442 ^ n20394 ;
  assign n20436 = n20394 ^ n20369 ;
  assign n20435 = n20394 ^ n20361 ;
  assign n20437 = n20436 ^ n20435 ;
  assign n20441 = n20375 & ~n20437 ;
  assign n20444 = n20443 ^ n20441 ;
  assign n20445 = n20434 & n20444 ;
  assign n20446 = n20445 ^ n20394 ;
  assign n20449 = ~n20429 & ~n20446 ;
  assign n20411 = n9520 & n11875 ;
  assign n20410 = x125 & n12206 ;
  assign n20412 = n20411 ^ n20410 ;
  assign n20407 = x126 & n9632 ;
  assign n20405 = n9636 & n10139 ;
  assign n20398 = x123 ^ x59 ;
  assign n20401 = n20382 & ~n20398 ;
  assign n20402 = n20401 ^ x123 ;
  assign n20403 = n12206 & n20402 ;
  assign n20404 = n20403 ^ x62 ;
  assign n20406 = n20405 ^ n20404 ;
  assign n20408 = n20407 ^ n20406 ;
  assign n20397 = x127 & n9628 ;
  assign n20409 = n20408 ^ n20397 ;
  assign n20413 = n20412 ^ n20409 ;
  assign n20414 = n20413 ^ n20391 ;
  assign n20415 = n20414 ^ n20379 ;
  assign n20416 = n20415 ^ n20413 ;
  assign n20417 = ~n20393 & ~n20416 ;
  assign n20418 = n20417 ^ n20414 ;
  assign n20450 = n20449 ^ n20418 ;
  assign n20462 = n20449 ^ n20413 ;
  assign n20463 = ~n20418 & n20462 ;
  assign n20464 = n20463 ^ n20413 ;
  assign n20460 = n9827 & n9948 ;
  assign n20456 = n20412 ^ n20403 ;
  assign n20457 = ~n20409 & ~n20456 ;
  assign n20458 = n20457 ^ n20412 ;
  assign n9637 = n9636 ^ n9632 ;
  assign n20453 = x127 & n9637 ;
  assign n20452 = n9636 & n10138 ;
  assign n20454 = n20453 ^ n20452 ;
  assign n20451 = n20411 ^ x62 ;
  assign n20455 = n20454 ^ n20451 ;
  assign n20459 = n20458 ^ n20455 ;
  assign n20461 = n20460 ^ n20459 ;
  assign n20465 = n20464 ^ n20461 ;
  assign n20469 = x126 ^ x124 ;
  assign n20475 = x63 & n20469 ;
  assign n20470 = x127 ^ x125 ;
  assign n20476 = n20475 ^ n20470 ;
  assign n20498 = ~n9948 & n20476 ;
  assign n20490 = n20454 ^ x126 ;
  assign n20491 = x63 & n9827 ;
  assign n20492 = n20490 & n20491 ;
  assign n20478 = x125 ^ x63 ;
  assign n20479 = n20478 ^ n20454 ;
  assign n20480 = n20469 ^ n20454 ;
  assign n20481 = n20480 ^ x125 ;
  assign n20482 = n20481 ^ n20469 ;
  assign n20485 = n9520 & n20482 ;
  assign n20486 = n20485 ^ n20469 ;
  assign n20487 = n20479 & n20486 ;
  assign n20488 = x62 & ~n20487 ;
  assign n20489 = n20488 ^ n20454 ;
  assign n20493 = n20492 ^ n20489 ;
  assign n20477 = n20470 ^ x62 ;
  assign n20494 = n20493 ^ n20477 ;
  assign n20499 = n20498 ^ n20494 ;
  assign n20466 = n20464 ^ n20458 ;
  assign n20467 = ~n20461 & n20466 ;
  assign n20468 = n20467 ^ n20464 ;
  assign n20500 = n20499 ^ n20468 ;
  assign n20521 = n20493 ^ n20468 ;
  assign n20522 = ~n20499 & ~n20521 ;
  assign n20512 = ~n20470 & n20478 ;
  assign n20504 = x124 & x126 ;
  assign n20505 = n20504 ^ x127 ;
  assign n20506 = x62 & ~n20505 ;
  assign n20513 = n20512 ^ n20506 ;
  assign n20515 = n20493 ^ x62 ;
  assign n20516 = n20515 ^ n20506 ;
  assign n20514 = n20493 ^ x63 ;
  assign n20517 = n20516 ^ n20514 ;
  assign n20518 = n20517 ^ n20512 ;
  assign n20519 = ~n20513 & n20518 ;
  assign n20520 = n20519 ^ n20516 ;
  assign n20523 = n20522 ^ n20520 ;
  assign y0 = n129 ;
  assign y1 = n132 ;
  assign y2 = ~n147 ;
  assign y3 = n180 ;
  assign y4 = n214 ;
  assign y5 = n268 ;
  assign y6 = n306 ;
  assign y7 = n355 ;
  assign y8 = ~n412 ;
  assign y9 = ~n468 ;
  assign y10 = n533 ;
  assign y11 = ~n611 ;
  assign y12 = n677 ;
  assign y13 = n752 ;
  assign y14 = n833 ;
  assign y15 = n913 ;
  assign y16 = n1005 ;
  assign y17 = n1098 ;
  assign y18 = n1186 ;
  assign y19 = n1285 ;
  assign y20 = n1391 ;
  assign y21 = n1492 ;
  assign y22 = n1604 ;
  assign y23 = n1723 ;
  assign y24 = n1837 ;
  assign y25 = n1962 ;
  assign y26 = n2099 ;
  assign y27 = n2229 ;
  assign y28 = n2366 ;
  assign y29 = ~n2519 ;
  assign y30 = ~n2664 ;
  assign y31 = n2816 ;
  assign y32 = ~n2974 ;
  assign y33 = n3130 ;
  assign y34 = n3303 ;
  assign y35 = ~n3474 ;
  assign y36 = ~n3640 ;
  assign y37 = n3817 ;
  assign y38 = n4010 ;
  assign y39 = n4193 ;
  assign y40 = n4388 ;
  assign y41 = n4593 ;
  assign y42 = n4792 ;
  assign y43 = n4997 ;
  assign y44 = n5214 ;
  assign y45 = n5426 ;
  assign y46 = n5646 ;
  assign y47 = ~n5880 ;
  assign y48 = ~n6107 ;
  assign y49 = ~n6338 ;
  assign y50 = ~n6578 ;
  assign y51 = n6817 ;
  assign y52 = ~n7070 ;
  assign y53 = n7321 ;
  assign y54 = ~n7568 ;
  assign y55 = n7824 ;
  assign y56 = n8096 ;
  assign y57 = n8368 ;
  assign y58 = ~n8638 ;
  assign y59 = ~n8922 ;
  assign y60 = ~n9215 ;
  assign y61 = ~n9513 ;
  assign y62 = n9823 ;
  assign y63 = n10121 ;
  assign y64 = ~n10424 ;
  assign y65 = n10711 ;
  assign y66 = ~n10986 ;
  assign y67 = n11256 ;
  assign y68 = n11530 ;
  assign y69 = ~n11807 ;
  assign y70 = n12084 ;
  assign y71 = n12353 ;
  assign y72 = ~n12605 ;
  assign y73 = n12875 ;
  assign y74 = n13130 ;
  assign y75 = n13376 ;
  assign y76 = ~n13609 ;
  assign y77 = n13849 ;
  assign y78 = ~n14083 ;
  assign y79 = ~n14325 ;
  assign y80 = ~n14556 ;
  assign y81 = n14812 ;
  assign y82 = n15027 ;
  assign y83 = ~n15257 ;
  assign y84 = n15457 ;
  assign y85 = ~n15691 ;
  assign y86 = ~n15890 ;
  assign y87 = ~n16076 ;
  assign y88 = n16261 ;
  assign y89 = ~n16453 ;
  assign y90 = n16626 ;
  assign y91 = ~n16819 ;
  assign y92 = n16994 ;
  assign y93 = ~n17158 ;
  assign y94 = ~n17314 ;
  assign y95 = n17505 ;
  assign y96 = ~n17652 ;
  assign y97 = n17802 ;
  assign y98 = n17948 ;
  assign y99 = ~n18116 ;
  assign y100 = n18247 ;
  assign y101 = ~n18380 ;
  assign y102 = n18515 ;
  assign y103 = ~n18632 ;
  assign y104 = n18758 ;
  assign y105 = n18883 ;
  assign y106 = n18995 ;
  assign y107 = ~n19100 ;
  assign y108 = n19220 ;
  assign y109 = ~n19329 ;
  assign y110 = n19427 ;
  assign y111 = ~n19523 ;
  assign y112 = ~n19602 ;
  assign y113 = ~n19696 ;
  assign y114 = n19785 ;
  assign y115 = ~n19862 ;
  assign y116 = ~n19929 ;
  assign y117 = n19982 ;
  assign y118 = ~n20057 ;
  assign y119 = n20160 ;
  assign y120 = ~n20215 ;
  assign y121 = ~n20338 ;
  assign y122 = n20372 ;
  assign y123 = ~n20396 ;
  assign y124 = n20450 ;
  assign y125 = ~n20465 ;
  assign y126 = n20500 ;
  assign y127 = ~n20523 ;
endmodule
