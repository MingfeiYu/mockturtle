module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n663 , n664 , n665 , n668 , n669 , n671 , n673 , n674 , n676 , n678 , n679 , n681 , n683 , n684 , n686 , n688 , n689 , n691 , n693 , n694 , n696 , n698 , n699 , n701 , n703 , n704 , n706 , n708 , n709 , n711 , n713 , n714 , n716 , n718 , n719 , n721 , n723 , n724 , n726 , n728 , n729 , n731 , n733 , n734 , n736 , n738 , n739 , n741 , n743 , n744 , n746 , n748 , n749 , n751 , n753 , n754 , n756 , n758 , n759 , n761 , n763 , n764 , n766 , n768 , n769 , n771 , n773 , n774 , n776 , n778 , n779 , n781 , n783 , n784 , n786 , n788 , n789 , n791 , n793 , n794 , n796 , n798 , n799 , n801 , n803 , n804 , n806 , n808 , n809 , n811 , n813 , n814 , n816 , n818 , n819 , n821 , n823 , n824 , n826 , n828 , n829 , n831 , n833 , n834 , n836 , n838 , n839 , n841 , n843 , n844 , n846 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n863 , n864 , n865 , n868 , n869 , n871 , n873 , n874 , n876 , n878 , n879 , n881 , n883 , n884 , n886 , n888 , n889 , n891 , n893 , n894 , n896 , n898 , n899 , n901 , n903 , n904 , n906 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n917 , n918 , n919 , n922 , n923 , n925 , n927 , n928 , n930 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n954 , n955 , n956 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n967 , n969 , n970 , n972 , n974 , n975 , n977 , n979 , n980 , n982 , n984 , n985 , n987 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1007 , n1009 , n1010 , n1012 , n1014 , n1015 , n1017 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1032 , n1034 , n1035 , n1037 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1052 , n1054 , n1055 , n1057 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1067 , n1069 , n1070 , n1072 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1082 , n1084 , n1085 , n1087 , n1089 , n1090 , n1092 , n1094 , n1095 , n1097 , n1099 , n1100 , n1102 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1117 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1132 , n1134 , n1135 , n1137 , n1139 , n1140 , n1142 , n1144 , n1145 , n1147 , n1149 , n1150 , n1152 , n1154 , n1155 , n1157 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1167 , n1168 , n1169 , n1170 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1318 , n1319 , n1320 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1336 , n1338 , n1339 , n1341 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1351 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1366 , n1368 , n1369 , n1371 , n1373 , n1374 , n1376 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1391 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1401 , n1403 , n1404 , n1406 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1416 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1436 , n1438 , n1439 , n1441 , n1443 , n1444 , n1446 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1456 , n1458 , n1459 , n1461 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1471 , n1473 , n1474 , n1476 , n1478 , n1479 , n1481 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1491 , n1493 , n1494 , n1496 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1523 , n1524 , n1525 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1536 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1546 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1563 , n1564 , n1565 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1577 , n1578 , n1579 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1595 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1620 , n1622 , n1623 , n1625 , n1627 , n1628 , n1630 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1660 , n1662 , n1663 , n1665 , n1667 , n1668 , n1670 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1690 , n1692 , n1693 , n1695 , n1697 , n1698 , n1700 , n1702 , n1703 , n1705 , n1707 , n1708 , n1710 , n1712 , n1713 , n1715 , n1717 , n1718 , n1720 , n1722 , n1723 , n1725 , n1727 , n1728 , n1730 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1740 , n1742 , n1743 , n1745 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1760 , n1762 , n1763 , n1765 , n1767 , n1768 , n1770 , n1772 , n1773 , n1775 , n1777 , n1778 , n1780 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1790 , n1792 , n1793 , n1795 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1820 , n1822 , n1823 , n1825 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1835 , n1836 , n1837 , n1838 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 ;
  assign n1183 = x384 ^ x256 ;
  assign n1184 = x511 ^ x383 ;
  assign n1185 = x509 ^ x381 ;
  assign n1186 = x510 ^ x382 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1188 = ~x380 & x508 ;
  assign n1190 = x507 ^ x379 ;
  assign n1189 = x379 & ~x507 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1192 = ~n1188 & ~n1191 ;
  assign n1193 = n1187 & n1192 ;
  assign n1194 = x506 ^ x378 ;
  assign n1198 = x455 ^ x327 ;
  assign n1197 = x327 & ~x455 ;
  assign n1199 = n1198 ^ n1197 ;
  assign n1200 = x454 ^ x326 ;
  assign n1202 = x324 & ~x452 ;
  assign n1201 = x454 ^ x453 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1204 = n1203 ^ x325 ;
  assign n1205 = n1204 ^ n1201 ;
  assign n1206 = n1202 ^ x454 ;
  assign n1207 = n1206 ^ n1201 ;
  assign n1208 = ~n1205 & ~n1207 ;
  assign n1209 = n1208 ^ n1201 ;
  assign n1210 = ~n1200 & ~n1209 ;
  assign n1211 = n1210 ^ x326 ;
  assign n1212 = ~n1197 & ~n1211 ;
  assign n1213 = x453 ^ x325 ;
  assign n1214 = ~n1200 & ~n1213 ;
  assign n1216 = x451 ^ x323 ;
  assign n1215 = x323 & ~x451 ;
  assign n1217 = n1216 ^ n1215 ;
  assign n1218 = x452 ^ x324 ;
  assign n1219 = n1218 ^ n1202 ;
  assign n1220 = ~n1217 & ~n1219 ;
  assign n1221 = n1214 & n1220 ;
  assign n1222 = x450 ^ x322 ;
  assign n1226 = x448 ^ x320 ;
  assign n1225 = x320 & ~x448 ;
  assign n1227 = n1226 ^ n1225 ;
  assign n1228 = x316 & ~x444 ;
  assign n1229 = x317 & ~x445 ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = ~x319 & x447 ;
  assign n1232 = x445 ^ x317 ;
  assign n1233 = n1232 ^ n1229 ;
  assign n1235 = x318 & ~x446 ;
  assign n1234 = x446 ^ x318 ;
  assign n1236 = n1235 ^ n1234 ;
  assign n1237 = ~n1233 & ~n1236 ;
  assign n1238 = ~n1231 & n1237 ;
  assign n1239 = n1230 & n1238 ;
  assign n1240 = n1239 ^ n1238 ;
  assign n1241 = x447 ^ x319 ;
  assign n1242 = n1235 ^ x447 ;
  assign n1243 = ~n1241 & ~n1242 ;
  assign n1244 = n1243 ^ x447 ;
  assign n1245 = ~n1225 & n1244 ;
  assign n1246 = ~n1240 & n1245 ;
  assign n1247 = x444 ^ x316 ;
  assign n1248 = n1247 ^ n1228 ;
  assign n1249 = n1238 & ~n1248 ;
  assign n1250 = x443 ^ x315 ;
  assign n1252 = x442 ^ x314 ;
  assign n1256 = x435 ^ x307 ;
  assign n1255 = x307 & ~x435 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1258 = x306 & ~x434 ;
  assign n1259 = ~n1255 & ~n1258 ;
  assign n1260 = ~x305 & x433 ;
  assign n1261 = x434 ^ x306 ;
  assign n1262 = n1261 ^ n1258 ;
  assign n1263 = ~n1260 & ~n1262 ;
  assign n1264 = x304 & ~x432 ;
  assign n1265 = x433 ^ x305 ;
  assign n1266 = n1265 ^ n1260 ;
  assign n1267 = ~n1264 & ~n1266 ;
  assign n1268 = x431 ^ x303 ;
  assign n1269 = x430 ^ x302 ;
  assign n1271 = x300 & ~x428 ;
  assign n1270 = x430 ^ x429 ;
  assign n1272 = n1271 ^ n1270 ;
  assign n1273 = n1272 ^ x301 ;
  assign n1274 = n1273 ^ n1270 ;
  assign n1275 = n1271 ^ x430 ;
  assign n1276 = n1275 ^ n1270 ;
  assign n1277 = ~n1274 & ~n1276 ;
  assign n1278 = n1277 ^ n1270 ;
  assign n1279 = ~n1269 & ~n1278 ;
  assign n1280 = n1279 ^ x302 ;
  assign n1281 = ~n1268 & ~n1280 ;
  assign n1282 = x429 ^ x301 ;
  assign n1283 = ~n1269 & ~n1282 ;
  assign n1284 = ~x299 & x427 ;
  assign n1285 = x428 ^ x300 ;
  assign n1286 = n1285 ^ n1271 ;
  assign n1287 = n1284 & ~n1286 ;
  assign n1288 = n1287 ^ n1286 ;
  assign n1289 = n1283 & ~n1288 ;
  assign n1290 = x427 ^ x299 ;
  assign n1291 = x426 ^ x298 ;
  assign n1293 = x296 & ~x424 ;
  assign n1292 = x426 ^ x425 ;
  assign n1294 = n1293 ^ n1292 ;
  assign n1295 = n1294 ^ x297 ;
  assign n1296 = n1295 ^ n1292 ;
  assign n1297 = n1293 ^ x426 ;
  assign n1298 = n1297 ^ n1292 ;
  assign n1299 = ~n1296 & ~n1298 ;
  assign n1300 = n1299 ^ n1292 ;
  assign n1301 = ~n1291 & ~n1300 ;
  assign n1302 = n1301 ^ x298 ;
  assign n1303 = ~n1290 & ~n1302 ;
  assign n1304 = x425 ^ x297 ;
  assign n1305 = ~n1291 & ~n1304 ;
  assign n1307 = x423 ^ x295 ;
  assign n1306 = x295 & ~x423 ;
  assign n1308 = n1307 ^ n1306 ;
  assign n1309 = x424 ^ x296 ;
  assign n1310 = n1309 ^ n1293 ;
  assign n1311 = ~n1308 & ~n1310 ;
  assign n1312 = n1305 & n1311 ;
  assign n1313 = x422 ^ x294 ;
  assign n1318 = x256 & ~x384 ;
  assign n1319 = n1318 ^ x385 ;
  assign n2208 = x385 ^ x257 ;
  assign n1323 = n1319 & ~n2208 ;
  assign n1320 = x386 ^ x257 ;
  assign n1324 = n1323 ^ n1320 ;
  assign n1326 = x387 ^ x258 ;
  assign n1325 = x387 ^ x386 ;
  assign n1327 = n1326 ^ n1325 ;
  assign n1328 = n1324 & ~n1327 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1331 = x388 ^ x259 ;
  assign n1330 = x388 ^ x387 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1333 = n1329 & ~n1332 ;
  assign n1334 = n1333 ^ n1331 ;
  assign n2201 = x388 ^ x260 ;
  assign n1338 = n1334 & ~n2201 ;
  assign n1336 = x389 ^ x260 ;
  assign n1339 = n1338 ^ n1336 ;
  assign n2194 = x389 ^ x261 ;
  assign n1343 = n1339 & ~n2194 ;
  assign n1341 = x390 ^ x261 ;
  assign n1344 = n1343 ^ n1341 ;
  assign n1346 = x391 ^ x262 ;
  assign n1345 = x391 ^ x390 ;
  assign n1347 = n1346 ^ n1345 ;
  assign n1348 = n1344 & ~n1347 ;
  assign n1349 = n1348 ^ n1346 ;
  assign n2187 = x391 ^ x263 ;
  assign n1353 = n1349 & ~n2187 ;
  assign n1351 = x392 ^ x263 ;
  assign n1354 = n1353 ^ n1351 ;
  assign n1356 = x393 ^ x264 ;
  assign n1355 = x393 ^ x392 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1358 = n1354 & ~n1357 ;
  assign n1359 = n1358 ^ n1356 ;
  assign n1361 = x394 ^ x265 ;
  assign n1360 = x394 ^ x393 ;
  assign n1362 = n1361 ^ n1360 ;
  assign n1363 = n1359 & ~n1362 ;
  assign n1364 = n1363 ^ n1361 ;
  assign n2180 = x394 ^ x266 ;
  assign n1368 = n1364 & ~n2180 ;
  assign n1366 = x395 ^ x266 ;
  assign n1369 = n1368 ^ n1366 ;
  assign n2173 = x395 ^ x267 ;
  assign n1373 = n1369 & ~n2173 ;
  assign n1371 = x396 ^ x267 ;
  assign n1374 = n1373 ^ n1371 ;
  assign n2166 = x396 ^ x268 ;
  assign n1378 = n1374 & ~n2166 ;
  assign n1376 = x397 ^ x268 ;
  assign n1379 = n1378 ^ n1376 ;
  assign n1381 = x398 ^ x269 ;
  assign n1380 = x398 ^ x397 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1383 = n1379 & ~n1382 ;
  assign n1384 = n1383 ^ n1381 ;
  assign n1386 = x399 ^ x270 ;
  assign n1385 = x399 ^ x398 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1388 = n1384 & ~n1387 ;
  assign n1389 = n1388 ^ n1386 ;
  assign n2159 = x399 ^ x271 ;
  assign n1393 = n1389 & ~n2159 ;
  assign n1391 = x400 ^ x271 ;
  assign n1394 = n1393 ^ n1391 ;
  assign n1396 = x401 ^ x272 ;
  assign n1395 = x401 ^ x400 ;
  assign n1397 = n1396 ^ n1395 ;
  assign n1398 = n1394 & ~n1397 ;
  assign n1399 = n1398 ^ n1396 ;
  assign n2152 = x401 ^ x273 ;
  assign n1403 = n1399 & ~n2152 ;
  assign n1401 = x402 ^ x273 ;
  assign n1404 = n1403 ^ n1401 ;
  assign n2145 = x402 ^ x274 ;
  assign n1408 = n1404 & ~n2145 ;
  assign n1406 = x403 ^ x274 ;
  assign n1409 = n1408 ^ n1406 ;
  assign n1411 = x404 ^ x275 ;
  assign n1410 = x404 ^ x403 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1413 = n1409 & ~n1412 ;
  assign n1414 = n1413 ^ n1411 ;
  assign n2138 = x404 ^ x276 ;
  assign n1418 = n1414 & ~n2138 ;
  assign n1416 = x405 ^ x276 ;
  assign n1419 = n1418 ^ n1416 ;
  assign n1421 = x406 ^ x277 ;
  assign n1420 = x406 ^ x405 ;
  assign n1422 = n1421 ^ n1420 ;
  assign n1423 = n1419 & ~n1422 ;
  assign n1424 = n1423 ^ n1421 ;
  assign n1426 = x407 ^ x278 ;
  assign n1425 = x407 ^ x406 ;
  assign n1427 = n1426 ^ n1425 ;
  assign n1428 = n1424 & ~n1427 ;
  assign n1429 = n1428 ^ n1426 ;
  assign n1431 = x408 ^ x279 ;
  assign n1430 = x408 ^ x407 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1433 = n1429 & ~n1432 ;
  assign n1434 = n1433 ^ n1431 ;
  assign n2131 = x408 ^ x280 ;
  assign n1438 = n1434 & ~n2131 ;
  assign n1436 = x409 ^ x280 ;
  assign n1439 = n1438 ^ n1436 ;
  assign n2124 = x409 ^ x281 ;
  assign n1443 = n1439 & ~n2124 ;
  assign n1441 = x410 ^ x281 ;
  assign n1444 = n1443 ^ n1441 ;
  assign n2117 = x410 ^ x282 ;
  assign n1448 = n1444 & ~n2117 ;
  assign n1446 = x411 ^ x282 ;
  assign n1449 = n1448 ^ n1446 ;
  assign n1451 = x412 ^ x283 ;
  assign n1450 = x412 ^ x411 ;
  assign n1452 = n1451 ^ n1450 ;
  assign n1453 = n1449 & ~n1452 ;
  assign n1454 = n1453 ^ n1451 ;
  assign n2110 = x412 ^ x284 ;
  assign n1458 = n1454 & ~n2110 ;
  assign n1456 = x413 ^ x284 ;
  assign n1459 = n1458 ^ n1456 ;
  assign n2103 = x413 ^ x285 ;
  assign n1463 = n1459 & ~n2103 ;
  assign n1461 = x414 ^ x285 ;
  assign n1464 = n1463 ^ n1461 ;
  assign n1466 = x415 ^ x286 ;
  assign n1465 = x415 ^ x414 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1468 = n1464 & ~n1467 ;
  assign n1469 = n1468 ^ n1466 ;
  assign n2096 = x415 ^ x287 ;
  assign n1473 = n1469 & ~n2096 ;
  assign n1471 = x416 ^ x287 ;
  assign n1474 = n1473 ^ n1471 ;
  assign n2089 = x416 ^ x288 ;
  assign n1478 = n1474 & ~n2089 ;
  assign n1476 = x417 ^ x288 ;
  assign n1479 = n1478 ^ n1476 ;
  assign n2082 = x417 ^ x289 ;
  assign n1483 = n1479 & ~n2082 ;
  assign n1481 = x418 ^ x289 ;
  assign n1484 = n1483 ^ n1481 ;
  assign n1486 = x419 ^ x290 ;
  assign n1485 = x419 ^ x418 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1488 = n1484 & ~n1487 ;
  assign n1489 = n1488 ^ n1486 ;
  assign n2075 = x419 ^ x291 ;
  assign n1493 = n1489 & ~n2075 ;
  assign n1491 = x420 ^ x291 ;
  assign n1494 = n1493 ^ n1491 ;
  assign n2068 = x420 ^ x292 ;
  assign n1498 = n1494 & ~n2068 ;
  assign n1496 = x421 ^ x292 ;
  assign n1499 = n1498 ^ n1496 ;
  assign n1501 = x422 ^ x293 ;
  assign n1500 = x422 ^ x421 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1503 = n1499 & ~n1502 ;
  assign n1504 = n1503 ^ n1501 ;
  assign n1505 = ~n1313 & n1504 ;
  assign n1506 = n1505 ^ x294 ;
  assign n1507 = ~n1306 & ~n1506 ;
  assign n1508 = n1312 & ~n1507 ;
  assign n1509 = n1303 & ~n1508 ;
  assign n1510 = n1289 & ~n1509 ;
  assign n1511 = n1281 & ~n1510 ;
  assign n1512 = ~x303 & x431 ;
  assign n1513 = x432 ^ x304 ;
  assign n1514 = n1513 ^ n1264 ;
  assign n1515 = n1512 & ~n1514 ;
  assign n1516 = n1515 ^ n1514 ;
  assign n1517 = ~n1511 & ~n1516 ;
  assign n1518 = n1267 & ~n1517 ;
  assign n1519 = n1263 & ~n1518 ;
  assign n1520 = n1259 & ~n1519 ;
  assign n1523 = ~n1257 & ~n1520 ;
  assign n1253 = x437 ^ x436 ;
  assign n1254 = n1253 ^ x308 ;
  assign n1524 = n1523 ^ n1254 ;
  assign n1525 = n1524 ^ n1253 ;
  assign n2015 = x436 ^ x308 ;
  assign n1528 = ~n1525 & ~n2015 ;
  assign n1529 = n1528 ^ n1253 ;
  assign n1531 = x438 ^ x309 ;
  assign n1530 = x438 ^ x437 ;
  assign n1532 = n1531 ^ n1530 ;
  assign n1533 = ~n1529 & ~n1532 ;
  assign n1534 = n1533 ^ n1531 ;
  assign n2008 = x438 ^ x310 ;
  assign n1538 = n1534 & ~n2008 ;
  assign n1536 = x439 ^ x310 ;
  assign n1539 = n1538 ^ n1536 ;
  assign n1541 = x440 ^ x311 ;
  assign n1540 = x440 ^ x439 ;
  assign n1542 = n1541 ^ n1540 ;
  assign n1543 = n1539 & ~n1542 ;
  assign n1544 = n1543 ^ n1541 ;
  assign n2001 = x440 ^ x312 ;
  assign n1548 = n1544 & ~n2001 ;
  assign n1546 = x441 ^ x312 ;
  assign n1549 = n1548 ^ n1546 ;
  assign n1551 = x442 ^ x313 ;
  assign n1550 = x442 ^ x441 ;
  assign n1552 = n1551 ^ n1550 ;
  assign n1553 = n1549 & ~n1552 ;
  assign n1554 = n1553 ^ n1551 ;
  assign n1555 = ~n1252 & n1554 ;
  assign n1251 = x443 ^ x314 ;
  assign n1556 = n1555 ^ n1251 ;
  assign n1557 = ~n1250 & n1556 ;
  assign n1558 = n1557 ^ x315 ;
  assign n1559 = n1249 & n1558 ;
  assign n1560 = n1246 & ~n1559 ;
  assign n1563 = ~n1227 & ~n1560 ;
  assign n1223 = x450 ^ x449 ;
  assign n1224 = n1223 ^ x321 ;
  assign n1564 = n1563 ^ n1224 ;
  assign n1565 = n1564 ^ n1223 ;
  assign n1973 = x449 ^ x321 ;
  assign n1568 = ~n1565 & ~n1973 ;
  assign n1569 = n1568 ^ n1223 ;
  assign n1570 = ~n1222 & ~n1569 ;
  assign n1571 = n1570 ^ x322 ;
  assign n1572 = ~n1215 & ~n1571 ;
  assign n1573 = n1221 & ~n1572 ;
  assign n1574 = n1212 & ~n1573 ;
  assign n1577 = ~n1199 & ~n1574 ;
  assign n1195 = x457 ^ x456 ;
  assign n1196 = n1195 ^ x328 ;
  assign n1578 = n1577 ^ n1196 ;
  assign n1579 = n1578 ^ n1195 ;
  assign n1941 = x456 ^ x328 ;
  assign n1582 = ~n1579 & ~n1941 ;
  assign n1583 = n1582 ^ n1195 ;
  assign n1585 = x458 ^ x329 ;
  assign n1584 = x458 ^ x457 ;
  assign n1586 = n1585 ^ n1584 ;
  assign n1587 = ~n1583 & ~n1586 ;
  assign n1588 = n1587 ^ n1585 ;
  assign n1590 = x459 ^ x330 ;
  assign n1589 = x459 ^ x458 ;
  assign n1591 = n1590 ^ n1589 ;
  assign n1592 = n1588 & ~n1591 ;
  assign n1593 = n1592 ^ n1590 ;
  assign n2654 = x459 ^ x331 ;
  assign n1597 = n1593 & ~n2654 ;
  assign n1595 = x460 ^ x331 ;
  assign n1598 = n1597 ^ n1595 ;
  assign n1600 = x461 ^ x332 ;
  assign n1599 = x461 ^ x460 ;
  assign n1601 = n1600 ^ n1599 ;
  assign n1602 = n1598 & ~n1601 ;
  assign n1603 = n1602 ^ n1600 ;
  assign n1605 = x462 ^ x333 ;
  assign n1604 = x462 ^ x461 ;
  assign n1606 = n1605 ^ n1604 ;
  assign n1607 = n1603 & ~n1606 ;
  assign n1608 = n1607 ^ n1605 ;
  assign n1610 = x463 ^ x334 ;
  assign n1609 = x463 ^ x462 ;
  assign n1611 = n1610 ^ n1609 ;
  assign n1612 = n1608 & ~n1611 ;
  assign n1613 = n1612 ^ n1610 ;
  assign n1615 = x464 ^ x335 ;
  assign n1614 = x464 ^ x463 ;
  assign n1616 = n1615 ^ n1614 ;
  assign n1617 = n1613 & ~n1616 ;
  assign n1618 = n1617 ^ n1615 ;
  assign n1935 = x464 ^ x336 ;
  assign n1622 = n1618 & ~n1935 ;
  assign n1620 = x465 ^ x336 ;
  assign n1623 = n1622 ^ n1620 ;
  assign n1928 = x465 ^ x337 ;
  assign n1627 = n1623 & ~n1928 ;
  assign n1625 = x466 ^ x337 ;
  assign n1628 = n1627 ^ n1625 ;
  assign n2711 = x466 ^ x338 ;
  assign n1632 = n1628 & ~n2711 ;
  assign n1630 = x467 ^ x338 ;
  assign n1633 = n1632 ^ n1630 ;
  assign n1635 = x468 ^ x339 ;
  assign n1634 = x468 ^ x467 ;
  assign n1636 = n1635 ^ n1634 ;
  assign n1637 = n1633 & ~n1636 ;
  assign n1638 = n1637 ^ n1635 ;
  assign n1640 = x469 ^ x340 ;
  assign n1639 = x469 ^ x468 ;
  assign n1641 = n1640 ^ n1639 ;
  assign n1642 = n1638 & ~n1641 ;
  assign n1643 = n1642 ^ n1640 ;
  assign n1645 = x470 ^ x341 ;
  assign n1644 = x470 ^ x469 ;
  assign n1646 = n1645 ^ n1644 ;
  assign n1647 = n1643 & ~n1646 ;
  assign n1648 = n1647 ^ n1645 ;
  assign n1650 = x471 ^ x342 ;
  assign n1649 = x471 ^ x470 ;
  assign n1651 = n1650 ^ n1649 ;
  assign n1652 = n1648 & ~n1651 ;
  assign n1653 = n1652 ^ n1650 ;
  assign n1655 = x472 ^ x343 ;
  assign n1654 = x472 ^ x471 ;
  assign n1656 = n1655 ^ n1654 ;
  assign n1657 = n1653 & ~n1656 ;
  assign n1658 = n1657 ^ n1655 ;
  assign n2777 = x472 ^ x344 ;
  assign n1662 = n1658 & ~n2777 ;
  assign n1660 = x473 ^ x344 ;
  assign n1663 = n1662 ^ n1660 ;
  assign n2788 = x473 ^ x345 ;
  assign n1667 = n1663 & ~n2788 ;
  assign n1665 = x474 ^ x345 ;
  assign n1668 = n1667 ^ n1665 ;
  assign n2799 = x474 ^ x346 ;
  assign n1672 = n1668 & ~n2799 ;
  assign n1670 = x475 ^ x346 ;
  assign n1673 = n1672 ^ n1670 ;
  assign n1675 = x476 ^ x347 ;
  assign n1674 = x476 ^ x475 ;
  assign n1676 = n1675 ^ n1674 ;
  assign n1677 = n1673 & ~n1676 ;
  assign n1678 = n1677 ^ n1675 ;
  assign n1680 = x477 ^ x348 ;
  assign n1679 = x477 ^ x476 ;
  assign n1681 = n1680 ^ n1679 ;
  assign n1682 = n1678 & ~n1681 ;
  assign n1683 = n1682 ^ n1680 ;
  assign n1685 = x478 ^ x349 ;
  assign n1684 = x478 ^ x477 ;
  assign n1686 = n1685 ^ n1684 ;
  assign n1687 = n1683 & ~n1686 ;
  assign n1688 = n1687 ^ n1685 ;
  assign n2843 = x478 ^ x350 ;
  assign n1692 = n1688 & ~n2843 ;
  assign n1690 = x479 ^ x350 ;
  assign n1693 = n1692 ^ n1690 ;
  assign n2854 = x479 ^ x351 ;
  assign n1697 = n1693 & ~n2854 ;
  assign n1695 = x480 ^ x351 ;
  assign n1698 = n1697 ^ n1695 ;
  assign n1921 = x480 ^ x352 ;
  assign n1702 = n1698 & ~n1921 ;
  assign n1700 = x481 ^ x352 ;
  assign n1703 = n1702 ^ n1700 ;
  assign n1914 = x481 ^ x353 ;
  assign n1707 = n1703 & ~n1914 ;
  assign n1705 = x482 ^ x353 ;
  assign n1708 = n1707 ^ n1705 ;
  assign n2871 = x482 ^ x354 ;
  assign n1712 = n1708 & ~n2871 ;
  assign n1710 = x483 ^ x354 ;
  assign n1713 = n1712 ^ n1710 ;
  assign n2882 = x483 ^ x355 ;
  assign n1717 = n1713 & ~n2882 ;
  assign n1715 = x484 ^ x355 ;
  assign n1718 = n1717 ^ n1715 ;
  assign n1907 = x484 ^ x356 ;
  assign n1722 = n1718 & ~n1907 ;
  assign n1720 = x485 ^ x356 ;
  assign n1723 = n1722 ^ n1720 ;
  assign n1900 = x485 ^ x357 ;
  assign n1727 = n1723 & ~n1900 ;
  assign n1725 = x486 ^ x357 ;
  assign n1728 = n1727 ^ n1725 ;
  assign n2899 = x486 ^ x358 ;
  assign n1732 = n1728 & ~n2899 ;
  assign n1730 = x487 ^ x358 ;
  assign n1733 = n1732 ^ n1730 ;
  assign n1735 = x488 ^ x359 ;
  assign n1734 = x488 ^ x487 ;
  assign n1736 = n1735 ^ n1734 ;
  assign n1737 = n1733 & ~n1736 ;
  assign n1738 = n1737 ^ n1735 ;
  assign n1893 = x488 ^ x360 ;
  assign n1742 = n1738 & ~n1893 ;
  assign n1740 = x489 ^ x360 ;
  assign n1743 = n1742 ^ n1740 ;
  assign n2924 = x489 ^ x361 ;
  assign n1747 = n1743 & ~n2924 ;
  assign n1745 = x490 ^ x361 ;
  assign n1748 = n1747 ^ n1745 ;
  assign n1750 = x491 ^ x362 ;
  assign n1749 = x491 ^ x490 ;
  assign n1751 = n1750 ^ n1749 ;
  assign n1752 = n1748 & ~n1751 ;
  assign n1753 = n1752 ^ n1750 ;
  assign n1755 = x492 ^ x363 ;
  assign n1754 = x492 ^ x491 ;
  assign n1756 = n1755 ^ n1754 ;
  assign n1757 = n1753 & ~n1756 ;
  assign n1758 = n1757 ^ n1755 ;
  assign n1886 = x492 ^ x364 ;
  assign n1762 = n1758 & ~n1886 ;
  assign n1760 = x493 ^ x364 ;
  assign n1763 = n1762 ^ n1760 ;
  assign n1879 = x493 ^ x365 ;
  assign n1767 = n1763 & ~n1879 ;
  assign n1765 = x494 ^ x365 ;
  assign n1768 = n1767 ^ n1765 ;
  assign n1872 = x494 ^ x366 ;
  assign n1772 = n1768 & ~n1872 ;
  assign n1770 = x495 ^ x366 ;
  assign n1773 = n1772 ^ n1770 ;
  assign n2966 = x495 ^ x367 ;
  assign n1777 = n1773 & ~n2966 ;
  assign n1775 = x496 ^ x367 ;
  assign n1778 = n1777 ^ n1775 ;
  assign n2977 = x496 ^ x368 ;
  assign n1782 = n1778 & ~n2977 ;
  assign n1780 = x497 ^ x368 ;
  assign n1783 = n1782 ^ n1780 ;
  assign n1785 = x498 ^ x369 ;
  assign n1784 = x498 ^ x497 ;
  assign n1786 = n1785 ^ n1784 ;
  assign n1787 = n1783 & ~n1786 ;
  assign n1788 = n1787 ^ n1785 ;
  assign n2999 = x498 ^ x370 ;
  assign n1792 = n1788 & ~n2999 ;
  assign n1790 = x499 ^ x370 ;
  assign n1793 = n1792 ^ n1790 ;
  assign n3010 = x499 ^ x371 ;
  assign n1797 = n1793 & ~n3010 ;
  assign n1795 = x500 ^ x371 ;
  assign n1798 = n1797 ^ n1795 ;
  assign n1800 = x501 ^ x372 ;
  assign n1799 = x501 ^ x500 ;
  assign n1801 = n1800 ^ n1799 ;
  assign n1802 = n1798 & ~n1801 ;
  assign n1803 = n1802 ^ n1800 ;
  assign n1805 = x502 ^ x373 ;
  assign n1804 = x502 ^ x501 ;
  assign n1806 = n1805 ^ n1804 ;
  assign n1807 = n1803 & ~n1806 ;
  assign n1808 = n1807 ^ n1805 ;
  assign n1810 = x503 ^ x374 ;
  assign n1809 = x503 ^ x502 ;
  assign n1811 = n1810 ^ n1809 ;
  assign n1812 = n1808 & ~n1811 ;
  assign n1813 = n1812 ^ n1810 ;
  assign n1815 = x504 ^ x375 ;
  assign n1814 = x504 ^ x503 ;
  assign n1816 = n1815 ^ n1814 ;
  assign n1817 = n1813 & ~n1816 ;
  assign n1818 = n1817 ^ n1815 ;
  assign n1865 = x504 ^ x376 ;
  assign n1822 = n1818 & ~n1865 ;
  assign n1820 = x505 ^ x376 ;
  assign n1823 = n1822 ^ n1820 ;
  assign n1858 = x505 ^ x377 ;
  assign n1827 = n1823 & ~n1858 ;
  assign n1825 = x506 ^ x377 ;
  assign n1828 = n1827 ^ n1825 ;
  assign n1829 = ~n1194 & n1828 ;
  assign n1830 = n1829 ^ x378 ;
  assign n1831 = ~n1189 & ~n1830 ;
  assign n1832 = n1193 & ~n1831 ;
  assign n1836 = n1188 ^ x509 ;
  assign n1835 = x508 ^ x380 ;
  assign n1837 = n1836 ^ n1835 ;
  assign n1841 = ~n1185 & n1837 ;
  assign n1838 = x510 ^ x381 ;
  assign n1842 = n1841 ^ n1838 ;
  assign n1843 = ~n1186 & n1842 ;
  assign n1844 = n1843 ^ x382 ;
  assign n1845 = ~n1832 & ~n1844 ;
  assign n1846 = n1845 ^ x511 ;
  assign n1847 = ~n1184 & n1846 ;
  assign n1848 = n1847 ^ x383 ;
  assign n1849 = n1183 & n1848 ;
  assign n1850 = n1849 ^ x256 ;
  assign n513 = x128 ^ x0 ;
  assign n514 = x255 ^ x127 ;
  assign n515 = x253 ^ x125 ;
  assign n516 = x254 ^ x126 ;
  assign n517 = ~n515 & ~n516 ;
  assign n518 = ~x124 & x252 ;
  assign n520 = x251 ^ x123 ;
  assign n519 = x123 & ~x251 ;
  assign n521 = n520 ^ n519 ;
  assign n522 = ~n518 & ~n521 ;
  assign n523 = n517 & n522 ;
  assign n524 = x250 ^ x122 ;
  assign n528 = x208 ^ x80 ;
  assign n527 = ~x80 & x208 ;
  assign n529 = n528 ^ n527 ;
  assign n530 = ~x79 & x207 ;
  assign n531 = ~n527 & ~n530 ;
  assign n532 = x78 & ~x206 ;
  assign n533 = x207 ^ x79 ;
  assign n534 = n533 ^ n530 ;
  assign n535 = ~n532 & ~n534 ;
  assign n536 = ~x77 & x205 ;
  assign n537 = x206 ^ x78 ;
  assign n538 = n537 ^ n532 ;
  assign n539 = ~n536 & ~n538 ;
  assign n540 = x76 & ~x204 ;
  assign n541 = x205 ^ x77 ;
  assign n542 = n541 ^ n536 ;
  assign n543 = ~n540 & ~n542 ;
  assign n544 = ~x75 & x203 ;
  assign n545 = x204 ^ x76 ;
  assign n546 = n545 ^ n540 ;
  assign n547 = ~n544 & ~n546 ;
  assign n548 = x74 & ~x202 ;
  assign n549 = x203 ^ x75 ;
  assign n550 = n549 ^ n544 ;
  assign n551 = ~n548 & ~n550 ;
  assign n552 = ~x73 & x201 ;
  assign n553 = x202 ^ x74 ;
  assign n554 = n553 ^ n548 ;
  assign n555 = ~n552 & ~n554 ;
  assign n556 = x72 & ~x200 ;
  assign n557 = x201 ^ x73 ;
  assign n558 = n557 ^ n552 ;
  assign n559 = ~n556 & ~n558 ;
  assign n560 = x199 ^ x71 ;
  assign n561 = x198 ^ x70 ;
  assign n563 = x68 & ~x196 ;
  assign n562 = x198 ^ x197 ;
  assign n564 = n563 ^ n562 ;
  assign n565 = n564 ^ x69 ;
  assign n566 = n565 ^ n562 ;
  assign n567 = n563 ^ x198 ;
  assign n568 = n567 ^ n562 ;
  assign n569 = ~n566 & ~n568 ;
  assign n570 = n569 ^ n562 ;
  assign n571 = ~n561 & ~n570 ;
  assign n572 = n571 ^ x70 ;
  assign n573 = ~n560 & ~n572 ;
  assign n574 = x196 ^ x68 ;
  assign n575 = n574 ^ n563 ;
  assign n576 = x197 ^ x69 ;
  assign n577 = ~n561 & ~n576 ;
  assign n578 = ~n575 & n577 ;
  assign n579 = x195 ^ x67 ;
  assign n583 = x191 ^ x63 ;
  assign n582 = x63 & ~x191 ;
  assign n584 = n583 ^ n582 ;
  assign n585 = x190 ^ x62 ;
  assign n587 = x60 & ~x188 ;
  assign n586 = x190 ^ x189 ;
  assign n588 = n587 ^ n586 ;
  assign n589 = n588 ^ x61 ;
  assign n590 = n589 ^ n586 ;
  assign n591 = n587 ^ x190 ;
  assign n592 = n591 ^ n586 ;
  assign n593 = ~n590 & ~n592 ;
  assign n594 = n593 ^ n586 ;
  assign n595 = ~n585 & ~n594 ;
  assign n596 = n595 ^ x62 ;
  assign n597 = ~n582 & ~n596 ;
  assign n598 = x189 ^ x61 ;
  assign n599 = ~n585 & ~n598 ;
  assign n601 = x187 ^ x59 ;
  assign n600 = x59 & ~x187 ;
  assign n602 = n601 ^ n600 ;
  assign n603 = x188 ^ x60 ;
  assign n604 = n603 ^ n587 ;
  assign n605 = ~n602 & ~n604 ;
  assign n606 = n599 & n605 ;
  assign n607 = x186 ^ x58 ;
  assign n611 = x176 ^ x48 ;
  assign n610 = ~x48 & x176 ;
  assign n612 = n611 ^ n610 ;
  assign n613 = x175 ^ x47 ;
  assign n614 = x174 ^ x46 ;
  assign n616 = x44 & ~x172 ;
  assign n615 = x174 ^ x173 ;
  assign n617 = n616 ^ n615 ;
  assign n618 = n617 ^ x45 ;
  assign n619 = n618 ^ n615 ;
  assign n620 = n616 ^ x174 ;
  assign n621 = n620 ^ n615 ;
  assign n622 = ~n619 & ~n621 ;
  assign n623 = n622 ^ n615 ;
  assign n624 = ~n614 & ~n623 ;
  assign n625 = n624 ^ x46 ;
  assign n626 = ~n613 & ~n625 ;
  assign n627 = x173 ^ x45 ;
  assign n628 = ~n614 & ~n627 ;
  assign n629 = ~x43 & x171 ;
  assign n630 = x172 ^ x44 ;
  assign n631 = n630 ^ n616 ;
  assign n632 = n629 & ~n631 ;
  assign n633 = n632 ^ n631 ;
  assign n634 = n628 & ~n633 ;
  assign n635 = x171 ^ x43 ;
  assign n636 = x170 ^ x42 ;
  assign n638 = x40 & ~x168 ;
  assign n637 = x170 ^ x169 ;
  assign n639 = n638 ^ n637 ;
  assign n640 = n639 ^ x41 ;
  assign n641 = n640 ^ n637 ;
  assign n642 = n638 ^ x170 ;
  assign n643 = n642 ^ n637 ;
  assign n644 = ~n641 & ~n643 ;
  assign n645 = n644 ^ n637 ;
  assign n646 = ~n636 & ~n645 ;
  assign n647 = n646 ^ x42 ;
  assign n648 = ~n635 & ~n647 ;
  assign n649 = x169 ^ x41 ;
  assign n650 = ~n636 & ~n649 ;
  assign n651 = ~x39 & x167 ;
  assign n652 = x168 ^ x40 ;
  assign n653 = n652 ^ n638 ;
  assign n654 = n651 & ~n653 ;
  assign n655 = n654 ^ n653 ;
  assign n656 = n650 & ~n655 ;
  assign n657 = x167 ^ x39 ;
  assign n658 = x166 ^ x38 ;
  assign n663 = x0 & ~x128 ;
  assign n664 = n663 ^ x129 ;
  assign n2211 = x129 ^ x1 ;
  assign n668 = n664 & ~n2211 ;
  assign n665 = x130 ^ x1 ;
  assign n669 = n668 ^ n665 ;
  assign n2222 = x130 ^ x2 ;
  assign n673 = n669 & ~n2222 ;
  assign n671 = x131 ^ x2 ;
  assign n674 = n673 ^ n671 ;
  assign n2233 = x131 ^ x3 ;
  assign n678 = n674 & ~n2233 ;
  assign n676 = x132 ^ x3 ;
  assign n679 = n678 ^ n676 ;
  assign n2204 = x132 ^ x4 ;
  assign n683 = n679 & ~n2204 ;
  assign n681 = x133 ^ x4 ;
  assign n684 = n683 ^ n681 ;
  assign n2197 = x133 ^ x5 ;
  assign n688 = n684 & ~n2197 ;
  assign n686 = x134 ^ x5 ;
  assign n689 = n688 ^ n686 ;
  assign n2250 = x134 ^ x6 ;
  assign n693 = n689 & ~n2250 ;
  assign n691 = x135 ^ x6 ;
  assign n694 = n693 ^ n691 ;
  assign n2190 = x135 ^ x7 ;
  assign n698 = n694 & ~n2190 ;
  assign n696 = x136 ^ x7 ;
  assign n699 = n698 ^ n696 ;
  assign n2264 = x136 ^ x8 ;
  assign n703 = n699 & ~n2264 ;
  assign n701 = x137 ^ x8 ;
  assign n704 = n703 ^ n701 ;
  assign n2275 = x137 ^ x9 ;
  assign n708 = n704 & ~n2275 ;
  assign n706 = x138 ^ x9 ;
  assign n709 = n708 ^ n706 ;
  assign n2183 = x138 ^ x10 ;
  assign n713 = n709 & ~n2183 ;
  assign n711 = x139 ^ x10 ;
  assign n714 = n713 ^ n711 ;
  assign n2176 = x139 ^ x11 ;
  assign n718 = n714 & ~n2176 ;
  assign n716 = x140 ^ x11 ;
  assign n719 = n718 ^ n716 ;
  assign n2169 = x140 ^ x12 ;
  assign n723 = n719 & ~n2169 ;
  assign n721 = x141 ^ x12 ;
  assign n724 = n723 ^ n721 ;
  assign n2295 = x141 ^ x13 ;
  assign n728 = n724 & ~n2295 ;
  assign n726 = x142 ^ x13 ;
  assign n729 = n728 ^ n726 ;
  assign n2306 = x142 ^ x14 ;
  assign n733 = n729 & ~n2306 ;
  assign n731 = x143 ^ x14 ;
  assign n734 = n733 ^ n731 ;
  assign n2162 = x143 ^ x15 ;
  assign n738 = n734 & ~n2162 ;
  assign n736 = x144 ^ x15 ;
  assign n739 = n738 ^ n736 ;
  assign n2320 = x144 ^ x16 ;
  assign n743 = n739 & ~n2320 ;
  assign n741 = x145 ^ x16 ;
  assign n744 = n743 ^ n741 ;
  assign n2155 = x145 ^ x17 ;
  assign n748 = n744 & ~n2155 ;
  assign n746 = x146 ^ x17 ;
  assign n749 = n748 ^ n746 ;
  assign n2148 = x146 ^ x18 ;
  assign n753 = n749 & ~n2148 ;
  assign n751 = x147 ^ x18 ;
  assign n754 = n753 ^ n751 ;
  assign n2337 = x147 ^ x19 ;
  assign n758 = n754 & ~n2337 ;
  assign n756 = x148 ^ x19 ;
  assign n759 = n758 ^ n756 ;
  assign n2141 = x148 ^ x20 ;
  assign n763 = n759 & ~n2141 ;
  assign n761 = x149 ^ x20 ;
  assign n764 = n763 ^ n761 ;
  assign n2351 = x149 ^ x21 ;
  assign n768 = n764 & ~n2351 ;
  assign n766 = x150 ^ x21 ;
  assign n769 = n768 ^ n766 ;
  assign n2362 = x150 ^ x22 ;
  assign n773 = n769 & ~n2362 ;
  assign n771 = x151 ^ x22 ;
  assign n774 = n773 ^ n771 ;
  assign n2373 = x151 ^ x23 ;
  assign n778 = n774 & ~n2373 ;
  assign n776 = x152 ^ x23 ;
  assign n779 = n778 ^ n776 ;
  assign n2134 = x152 ^ x24 ;
  assign n783 = n779 & ~n2134 ;
  assign n781 = x153 ^ x24 ;
  assign n784 = n783 ^ n781 ;
  assign n2127 = x153 ^ x25 ;
  assign n788 = n784 & ~n2127 ;
  assign n786 = x154 ^ x25 ;
  assign n789 = n788 ^ n786 ;
  assign n2120 = x154 ^ x26 ;
  assign n793 = n789 & ~n2120 ;
  assign n791 = x155 ^ x26 ;
  assign n794 = n793 ^ n791 ;
  assign n2393 = x155 ^ x27 ;
  assign n798 = n794 & ~n2393 ;
  assign n796 = x156 ^ x27 ;
  assign n799 = n798 ^ n796 ;
  assign n2113 = x156 ^ x28 ;
  assign n803 = n799 & ~n2113 ;
  assign n801 = x157 ^ x28 ;
  assign n804 = n803 ^ n801 ;
  assign n2106 = x157 ^ x29 ;
  assign n808 = n804 & ~n2106 ;
  assign n806 = x158 ^ x29 ;
  assign n809 = n808 ^ n806 ;
  assign n2410 = x158 ^ x30 ;
  assign n813 = n809 & ~n2410 ;
  assign n811 = x159 ^ x30 ;
  assign n814 = n813 ^ n811 ;
  assign n2099 = x159 ^ x31 ;
  assign n818 = n814 & ~n2099 ;
  assign n816 = x160 ^ x31 ;
  assign n819 = n818 ^ n816 ;
  assign n2092 = x160 ^ x32 ;
  assign n823 = n819 & ~n2092 ;
  assign n821 = x161 ^ x32 ;
  assign n824 = n823 ^ n821 ;
  assign n2085 = x161 ^ x33 ;
  assign n828 = n824 & ~n2085 ;
  assign n826 = x162 ^ x33 ;
  assign n829 = n828 ^ n826 ;
  assign n2430 = x162 ^ x34 ;
  assign n833 = n829 & ~n2430 ;
  assign n831 = x163 ^ x34 ;
  assign n834 = n833 ^ n831 ;
  assign n2078 = x163 ^ x35 ;
  assign n838 = n834 & ~n2078 ;
  assign n836 = x164 ^ x35 ;
  assign n839 = n838 ^ n836 ;
  assign n2071 = x164 ^ x36 ;
  assign n843 = n839 & ~n2071 ;
  assign n841 = x165 ^ x36 ;
  assign n844 = n843 ^ n841 ;
  assign n2447 = x165 ^ x37 ;
  assign n848 = n844 & ~n2447 ;
  assign n846 = x166 ^ x37 ;
  assign n849 = n848 ^ n846 ;
  assign n850 = ~n658 & n849 ;
  assign n851 = n850 ^ x38 ;
  assign n852 = ~n657 & ~n851 ;
  assign n853 = n656 & ~n852 ;
  assign n854 = n648 & ~n853 ;
  assign n855 = n634 & ~n854 ;
  assign n856 = n626 & ~n855 ;
  assign n857 = ~x47 & x175 ;
  assign n858 = ~n610 & n857 ;
  assign n859 = n858 ^ n610 ;
  assign n860 = ~n856 & ~n859 ;
  assign n863 = ~n612 & ~n860 ;
  assign n608 = x178 ^ x177 ;
  assign n609 = n608 ^ x49 ;
  assign n864 = n863 ^ n609 ;
  assign n865 = n864 ^ n608 ;
  assign n2024 = x177 ^ x49 ;
  assign n868 = n865 & ~n2024 ;
  assign n869 = n868 ^ n608 ;
  assign n2509 = x178 ^ x50 ;
  assign n873 = ~n869 & ~n2509 ;
  assign n871 = x179 ^ x50 ;
  assign n874 = n873 ^ n871 ;
  assign n2518 = x179 ^ x51 ;
  assign n878 = n874 & ~n2518 ;
  assign n876 = x180 ^ x51 ;
  assign n879 = n878 ^ n876 ;
  assign n2018 = x180 ^ x52 ;
  assign n883 = n879 & ~n2018 ;
  assign n881 = x181 ^ x52 ;
  assign n884 = n883 ^ n881 ;
  assign n2530 = x181 ^ x53 ;
  assign n888 = n884 & ~n2530 ;
  assign n886 = x182 ^ x53 ;
  assign n889 = n888 ^ n886 ;
  assign n2011 = x182 ^ x54 ;
  assign n893 = n889 & ~n2011 ;
  assign n891 = x183 ^ x54 ;
  assign n894 = n893 ^ n891 ;
  assign n2544 = x183 ^ x55 ;
  assign n898 = n894 & ~n2544 ;
  assign n896 = x184 ^ x55 ;
  assign n899 = n898 ^ n896 ;
  assign n2004 = x184 ^ x56 ;
  assign n903 = n899 & ~n2004 ;
  assign n901 = x185 ^ x56 ;
  assign n904 = n903 ^ n901 ;
  assign n2558 = x185 ^ x57 ;
  assign n908 = n904 & ~n2558 ;
  assign n906 = x186 ^ x57 ;
  assign n909 = n908 ^ n906 ;
  assign n910 = ~n607 & n909 ;
  assign n911 = n910 ^ x58 ;
  assign n912 = ~n600 & ~n911 ;
  assign n913 = n606 & ~n912 ;
  assign n914 = n597 & ~n913 ;
  assign n917 = ~n584 & ~n914 ;
  assign n580 = x193 ^ x192 ;
  assign n581 = n580 ^ x64 ;
  assign n918 = n917 ^ n581 ;
  assign n919 = n918 ^ n580 ;
  assign n1982 = x192 ^ x64 ;
  assign n922 = ~n919 & ~n1982 ;
  assign n923 = n922 ^ n580 ;
  assign n1976 = x193 ^ x65 ;
  assign n927 = ~n923 & ~n1976 ;
  assign n925 = x194 ^ x65 ;
  assign n928 = n927 ^ n925 ;
  assign n1969 = x194 ^ x66 ;
  assign n932 = n928 & ~n1969 ;
  assign n930 = x195 ^ x66 ;
  assign n933 = n932 ^ n930 ;
  assign n934 = ~n579 & n933 ;
  assign n935 = n934 ^ x67 ;
  assign n936 = n578 & n935 ;
  assign n937 = n573 & ~n936 ;
  assign n938 = ~x71 & x199 ;
  assign n939 = x200 ^ x72 ;
  assign n940 = n939 ^ n556 ;
  assign n941 = n938 & ~n940 ;
  assign n942 = n941 ^ n940 ;
  assign n943 = ~n937 & ~n942 ;
  assign n944 = n559 & ~n943 ;
  assign n945 = n555 & ~n944 ;
  assign n946 = n551 & ~n945 ;
  assign n947 = n547 & ~n946 ;
  assign n948 = n543 & ~n947 ;
  assign n949 = n539 & ~n948 ;
  assign n950 = n535 & ~n949 ;
  assign n951 = n531 & ~n950 ;
  assign n954 = ~n529 & ~n951 ;
  assign n525 = x210 ^ x209 ;
  assign n526 = n525 ^ x81 ;
  assign n955 = n954 ^ n526 ;
  assign n956 = n955 ^ n525 ;
  assign n1931 = x209 ^ x81 ;
  assign n959 = n956 & ~n1931 ;
  assign n960 = n959 ^ n525 ;
  assign n962 = x211 ^ x82 ;
  assign n961 = x211 ^ x210 ;
  assign n963 = n962 ^ n961 ;
  assign n964 = ~n960 & ~n963 ;
  assign n965 = n964 ^ n962 ;
  assign n2722 = x211 ^ x83 ;
  assign n969 = n965 & ~n2722 ;
  assign n967 = x212 ^ x83 ;
  assign n970 = n969 ^ n967 ;
  assign n2733 = x212 ^ x84 ;
  assign n974 = n970 & ~n2733 ;
  assign n972 = x213 ^ x84 ;
  assign n975 = n974 ^ n972 ;
  assign n2744 = x213 ^ x85 ;
  assign n979 = n975 & ~n2744 ;
  assign n977 = x214 ^ x85 ;
  assign n980 = n979 ^ n977 ;
  assign n2755 = x214 ^ x86 ;
  assign n984 = n980 & ~n2755 ;
  assign n982 = x215 ^ x86 ;
  assign n985 = n984 ^ n982 ;
  assign n2766 = x215 ^ x87 ;
  assign n989 = n985 & ~n2766 ;
  assign n987 = x216 ^ x87 ;
  assign n990 = n989 ^ n987 ;
  assign n992 = x217 ^ x88 ;
  assign n991 = x217 ^ x216 ;
  assign n993 = n992 ^ n991 ;
  assign n994 = n990 & ~n993 ;
  assign n995 = n994 ^ n992 ;
  assign n997 = x218 ^ x89 ;
  assign n996 = x218 ^ x217 ;
  assign n998 = n997 ^ n996 ;
  assign n999 = n995 & ~n998 ;
  assign n1000 = n999 ^ n997 ;
  assign n1002 = x219 ^ x90 ;
  assign n1001 = x219 ^ x218 ;
  assign n1003 = n1002 ^ n1001 ;
  assign n1004 = n1000 & ~n1003 ;
  assign n1005 = n1004 ^ n1002 ;
  assign n2810 = x219 ^ x91 ;
  assign n1009 = n1005 & ~n2810 ;
  assign n1007 = x220 ^ x91 ;
  assign n1010 = n1009 ^ n1007 ;
  assign n2821 = x220 ^ x92 ;
  assign n1014 = n1010 & ~n2821 ;
  assign n1012 = x221 ^ x92 ;
  assign n1015 = n1014 ^ n1012 ;
  assign n2832 = x221 ^ x93 ;
  assign n1019 = n1015 & ~n2832 ;
  assign n1017 = x222 ^ x93 ;
  assign n1020 = n1019 ^ n1017 ;
  assign n1022 = x223 ^ x94 ;
  assign n1021 = x223 ^ x222 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = n1024 ^ n1022 ;
  assign n1027 = x224 ^ x95 ;
  assign n1026 = x224 ^ x223 ;
  assign n1028 = n1027 ^ n1026 ;
  assign n1029 = n1025 & ~n1028 ;
  assign n1030 = n1029 ^ n1027 ;
  assign n1924 = x224 ^ x96 ;
  assign n1034 = n1030 & ~n1924 ;
  assign n1032 = x225 ^ x96 ;
  assign n1035 = n1034 ^ n1032 ;
  assign n1917 = x225 ^ x97 ;
  assign n1039 = n1035 & ~n1917 ;
  assign n1037 = x226 ^ x97 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n1042 = x227 ^ x98 ;
  assign n1041 = x227 ^ x226 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1044 = n1040 & ~n1043 ;
  assign n1045 = n1044 ^ n1042 ;
  assign n1047 = x228 ^ x99 ;
  assign n1046 = x228 ^ x227 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1049 = n1045 & ~n1048 ;
  assign n1050 = n1049 ^ n1047 ;
  assign n1910 = x228 ^ x100 ;
  assign n1054 = n1050 & ~n1910 ;
  assign n1052 = x229 ^ x100 ;
  assign n1055 = n1054 ^ n1052 ;
  assign n1903 = x229 ^ x101 ;
  assign n1059 = n1055 & ~n1903 ;
  assign n1057 = x230 ^ x101 ;
  assign n1060 = n1059 ^ n1057 ;
  assign n1062 = x231 ^ x102 ;
  assign n1061 = x231 ^ x230 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1064 = n1060 & ~n1063 ;
  assign n1065 = n1064 ^ n1062 ;
  assign n2910 = x231 ^ x103 ;
  assign n1069 = n1065 & ~n2910 ;
  assign n1067 = x232 ^ x103 ;
  assign n1070 = n1069 ^ n1067 ;
  assign n1896 = x232 ^ x104 ;
  assign n1074 = n1070 & ~n1896 ;
  assign n1072 = x233 ^ x104 ;
  assign n1075 = n1074 ^ n1072 ;
  assign n1077 = x234 ^ x105 ;
  assign n1076 = x234 ^ x233 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1079 = n1075 & ~n1078 ;
  assign n1080 = n1079 ^ n1077 ;
  assign n2935 = x234 ^ x106 ;
  assign n1084 = n1080 & ~n2935 ;
  assign n1082 = x235 ^ x106 ;
  assign n1085 = n1084 ^ n1082 ;
  assign n2946 = x235 ^ x107 ;
  assign n1089 = n1085 & ~n2946 ;
  assign n1087 = x236 ^ x107 ;
  assign n1090 = n1089 ^ n1087 ;
  assign n1889 = x236 ^ x108 ;
  assign n1094 = n1090 & ~n1889 ;
  assign n1092 = x237 ^ x108 ;
  assign n1095 = n1094 ^ n1092 ;
  assign n1882 = x237 ^ x109 ;
  assign n1099 = n1095 & ~n1882 ;
  assign n1097 = x238 ^ x109 ;
  assign n1100 = n1099 ^ n1097 ;
  assign n1875 = x238 ^ x110 ;
  assign n1104 = n1100 & ~n1875 ;
  assign n1102 = x239 ^ x110 ;
  assign n1105 = n1104 ^ n1102 ;
  assign n1107 = x240 ^ x111 ;
  assign n1106 = x240 ^ x239 ;
  assign n1108 = n1107 ^ n1106 ;
  assign n1109 = n1105 & ~n1108 ;
  assign n1110 = n1109 ^ n1107 ;
  assign n1112 = x241 ^ x112 ;
  assign n1111 = x241 ^ x240 ;
  assign n1113 = n1112 ^ n1111 ;
  assign n1114 = n1110 & ~n1113 ;
  assign n1115 = n1114 ^ n1112 ;
  assign n2988 = x241 ^ x113 ;
  assign n1119 = n1115 & ~n2988 ;
  assign n1117 = x242 ^ x113 ;
  assign n1120 = n1119 ^ n1117 ;
  assign n1122 = x243 ^ x114 ;
  assign n1121 = x243 ^ x242 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1124 = n1120 & ~n1123 ;
  assign n1125 = n1124 ^ n1122 ;
  assign n1127 = x244 ^ x115 ;
  assign n1126 = x244 ^ x243 ;
  assign n1128 = n1127 ^ n1126 ;
  assign n1129 = n1125 & ~n1128 ;
  assign n1130 = n1129 ^ n1127 ;
  assign n3021 = x244 ^ x116 ;
  assign n1134 = n1130 & ~n3021 ;
  assign n1132 = x245 ^ x116 ;
  assign n1135 = n1134 ^ n1132 ;
  assign n3032 = x245 ^ x117 ;
  assign n1139 = n1135 & ~n3032 ;
  assign n1137 = x246 ^ x117 ;
  assign n1140 = n1139 ^ n1137 ;
  assign n3043 = x246 ^ x118 ;
  assign n1144 = n1140 & ~n3043 ;
  assign n1142 = x247 ^ x118 ;
  assign n1145 = n1144 ^ n1142 ;
  assign n3054 = x247 ^ x119 ;
  assign n1149 = n1145 & ~n3054 ;
  assign n1147 = x248 ^ x119 ;
  assign n1150 = n1149 ^ n1147 ;
  assign n1868 = x248 ^ x120 ;
  assign n1154 = n1150 & ~n1868 ;
  assign n1152 = x249 ^ x120 ;
  assign n1155 = n1154 ^ n1152 ;
  assign n1861 = x249 ^ x121 ;
  assign n1159 = n1155 & ~n1861 ;
  assign n1157 = x250 ^ x121 ;
  assign n1160 = n1159 ^ n1157 ;
  assign n1161 = ~n524 & n1160 ;
  assign n1162 = n1161 ^ x122 ;
  assign n1163 = ~n519 & ~n1162 ;
  assign n1164 = n523 & ~n1163 ;
  assign n1168 = n518 ^ x253 ;
  assign n1167 = x252 ^ x124 ;
  assign n1169 = n1168 ^ n1167 ;
  assign n1173 = ~n515 & n1169 ;
  assign n1170 = x254 ^ x125 ;
  assign n1174 = n1173 ^ n1170 ;
  assign n1175 = ~n516 & n1174 ;
  assign n1176 = n1175 ^ x126 ;
  assign n1177 = ~n1164 & ~n1176 ;
  assign n1178 = n1177 ^ x255 ;
  assign n1179 = ~n514 & n1178 ;
  assign n1180 = n1179 ^ x127 ;
  assign n1181 = n513 & n1180 ;
  assign n1182 = n1181 ^ x0 ;
  assign n1851 = n1850 ^ n1182 ;
  assign n1853 = x383 & x511 ;
  assign n1852 = x127 & x255 ;
  assign n1854 = n1853 ^ n1852 ;
  assign n3099 = n515 & n1180 ;
  assign n3100 = n3099 ^ x125 ;
  assign n1855 = n516 & n1180 ;
  assign n1856 = n1855 ^ x126 ;
  assign n3109 = n3100 ^ n1856 ;
  assign n3089 = n1835 & n1848 ;
  assign n3090 = n3089 ^ x380 ;
  assign n3101 = n3100 ^ n3090 ;
  assign n3079 = n1190 & n1848 ;
  assign n3080 = n3079 ^ x379 ;
  assign n3091 = n3090 ^ n3080 ;
  assign n3071 = n524 & n1180 ;
  assign n3072 = n3071 ^ x122 ;
  assign n3081 = n3080 ^ n3072 ;
  assign n1862 = n1180 & n1861 ;
  assign n1863 = n1862 ^ x121 ;
  assign n3073 = n3072 ^ n1863 ;
  assign n1859 = n1848 & n1858 ;
  assign n1860 = n1859 ^ x377 ;
  assign n1864 = n1863 ^ n1860 ;
  assign n1869 = n1180 & n1868 ;
  assign n1870 = n1869 ^ x120 ;
  assign n3068 = n1870 ^ n1860 ;
  assign n1866 = n1848 & n1865 ;
  assign n1867 = n1866 ^ x376 ;
  assign n1871 = n1870 ^ n1867 ;
  assign n3055 = n1180 & n3054 ;
  assign n3056 = n3055 ^ x119 ;
  assign n3065 = n3056 ^ n1867 ;
  assign n3044 = n1180 & n3043 ;
  assign n3045 = n3044 ^ x118 ;
  assign n3057 = n3056 ^ n3045 ;
  assign n3033 = n1180 & n3032 ;
  assign n3034 = n3033 ^ x117 ;
  assign n3046 = n3045 ^ n3034 ;
  assign n3022 = n1180 & n3021 ;
  assign n3023 = n3022 ^ x116 ;
  assign n3035 = n3034 ^ n3023 ;
  assign n3011 = n1848 & n3010 ;
  assign n3012 = n3011 ^ x371 ;
  assign n3024 = n3023 ^ n3012 ;
  assign n3000 = n1848 & n2999 ;
  assign n3001 = n3000 ^ x370 ;
  assign n3013 = n3012 ^ n3001 ;
  assign n2989 = n1180 & n2988 ;
  assign n2990 = n2989 ^ x113 ;
  assign n3002 = n3001 ^ n2990 ;
  assign n2978 = n1848 & n2977 ;
  assign n2979 = n2978 ^ x368 ;
  assign n2991 = n2990 ^ n2979 ;
  assign n2967 = n1848 & n2966 ;
  assign n2968 = n2967 ^ x367 ;
  assign n2980 = n2979 ^ n2968 ;
  assign n1876 = n1180 & n1875 ;
  assign n1877 = n1876 ^ x110 ;
  assign n2969 = n2968 ^ n1877 ;
  assign n1873 = n1848 & n1872 ;
  assign n1874 = n1873 ^ x366 ;
  assign n1878 = n1877 ^ n1874 ;
  assign n1883 = n1180 & n1882 ;
  assign n1884 = n1883 ^ x109 ;
  assign n2963 = n1884 ^ n1874 ;
  assign n1880 = n1848 & n1879 ;
  assign n1881 = n1880 ^ x365 ;
  assign n1885 = n1884 ^ n1881 ;
  assign n1890 = n1180 & n1889 ;
  assign n1891 = n1890 ^ x108 ;
  assign n2960 = n1891 ^ n1881 ;
  assign n1887 = n1848 & n1886 ;
  assign n1888 = n1887 ^ x364 ;
  assign n1892 = n1891 ^ n1888 ;
  assign n2947 = n1180 & n2946 ;
  assign n2948 = n2947 ^ x107 ;
  assign n2957 = n2948 ^ n1888 ;
  assign n2936 = n1180 & n2935 ;
  assign n2937 = n2936 ^ x106 ;
  assign n2949 = n2948 ^ n2937 ;
  assign n2925 = n1848 & n2924 ;
  assign n2926 = n2925 ^ x361 ;
  assign n2938 = n2937 ^ n2926 ;
  assign n1897 = n1180 & n1896 ;
  assign n1898 = n1897 ^ x104 ;
  assign n2927 = n2926 ^ n1898 ;
  assign n1894 = n1848 & n1893 ;
  assign n1895 = n1894 ^ x360 ;
  assign n1899 = n1898 ^ n1895 ;
  assign n2911 = n1180 & n2910 ;
  assign n2912 = n2911 ^ x103 ;
  assign n2921 = n2912 ^ n1895 ;
  assign n2900 = n1848 & n2899 ;
  assign n2901 = n2900 ^ x358 ;
  assign n2913 = n2912 ^ n2901 ;
  assign n1904 = n1180 & n1903 ;
  assign n1905 = n1904 ^ x101 ;
  assign n2902 = n2901 ^ n1905 ;
  assign n1901 = n1848 & n1900 ;
  assign n1902 = n1901 ^ x357 ;
  assign n1906 = n1905 ^ n1902 ;
  assign n1911 = n1180 & n1910 ;
  assign n1912 = n1911 ^ x100 ;
  assign n2896 = n1912 ^ n1902 ;
  assign n1908 = n1848 & n1907 ;
  assign n1909 = n1908 ^ x356 ;
  assign n1913 = n1912 ^ n1909 ;
  assign n2883 = n1848 & n2882 ;
  assign n2884 = n2883 ^ x355 ;
  assign n2893 = n2884 ^ n1909 ;
  assign n2872 = n1848 & n2871 ;
  assign n2873 = n2872 ^ x354 ;
  assign n2885 = n2884 ^ n2873 ;
  assign n1918 = n1180 & n1917 ;
  assign n1919 = n1918 ^ x97 ;
  assign n2874 = n2873 ^ n1919 ;
  assign n1915 = n1848 & n1914 ;
  assign n1916 = n1915 ^ x353 ;
  assign n1920 = n1919 ^ n1916 ;
  assign n1925 = n1180 & n1924 ;
  assign n1926 = n1925 ^ x96 ;
  assign n2868 = n1926 ^ n1916 ;
  assign n1922 = n1848 & n1921 ;
  assign n1923 = n1922 ^ x352 ;
  assign n1927 = n1926 ^ n1923 ;
  assign n2855 = n1848 & n2854 ;
  assign n2856 = n2855 ^ x351 ;
  assign n2865 = n2856 ^ n1923 ;
  assign n2844 = n1848 & n2843 ;
  assign n2845 = n2844 ^ x350 ;
  assign n2857 = n2856 ^ n2845 ;
  assign n2833 = n1180 & n2832 ;
  assign n2834 = n2833 ^ x93 ;
  assign n2846 = n2845 ^ n2834 ;
  assign n2822 = n1180 & n2821 ;
  assign n2823 = n2822 ^ x92 ;
  assign n2835 = n2834 ^ n2823 ;
  assign n2811 = n1180 & n2810 ;
  assign n2812 = n2811 ^ x91 ;
  assign n2824 = n2823 ^ n2812 ;
  assign n2800 = n1848 & n2799 ;
  assign n2801 = n2800 ^ x346 ;
  assign n2813 = n2812 ^ n2801 ;
  assign n2789 = n1848 & n2788 ;
  assign n2790 = n2789 ^ x345 ;
  assign n2802 = n2801 ^ n2790 ;
  assign n2778 = n1848 & n2777 ;
  assign n2779 = n2778 ^ x344 ;
  assign n2791 = n2790 ^ n2779 ;
  assign n2767 = n1180 & n2766 ;
  assign n2768 = n2767 ^ x87 ;
  assign n2780 = n2779 ^ n2768 ;
  assign n2756 = n1180 & n2755 ;
  assign n2757 = n2756 ^ x86 ;
  assign n2769 = n2768 ^ n2757 ;
  assign n2745 = n1180 & n2744 ;
  assign n2746 = n2745 ^ x85 ;
  assign n2758 = n2757 ^ n2746 ;
  assign n2734 = n1180 & n2733 ;
  assign n2735 = n2734 ^ x84 ;
  assign n2747 = n2746 ^ n2735 ;
  assign n2723 = n1180 & n2722 ;
  assign n2724 = n2723 ^ x83 ;
  assign n2736 = n2735 ^ n2724 ;
  assign n2712 = n1848 & n2711 ;
  assign n2713 = n2712 ^ x338 ;
  assign n2725 = n2724 ^ n2713 ;
  assign n1932 = n1180 & n1931 ;
  assign n1933 = n1932 ^ x81 ;
  assign n2714 = n2713 ^ n1933 ;
  assign n1929 = n1848 & n1928 ;
  assign n1930 = n1929 ^ x337 ;
  assign n1934 = n1933 ^ n1930 ;
  assign n1938 = n528 & n1180 ;
  assign n1939 = n1938 ^ x80 ;
  assign n2708 = n1939 ^ n1930 ;
  assign n1936 = n1848 & n1935 ;
  assign n1937 = n1936 ^ x336 ;
  assign n1940 = n1939 ^ n1937 ;
  assign n2695 = n533 & n1180 ;
  assign n2696 = n2695 ^ x79 ;
  assign n2705 = n2696 ^ n1937 ;
  assign n2685 = n537 & n1180 ;
  assign n2686 = n2685 ^ x78 ;
  assign n2697 = n2696 ^ n2686 ;
  assign n2675 = n541 & n1180 ;
  assign n2676 = n2675 ^ x77 ;
  assign n2687 = n2686 ^ n2676 ;
  assign n2665 = n545 & n1180 ;
  assign n2666 = n2665 ^ x76 ;
  assign n2677 = n2676 ^ n2666 ;
  assign n2655 = n1848 & n2654 ;
  assign n2656 = n2655 ^ x331 ;
  assign n2667 = n2666 ^ n2656 ;
  assign n2644 = n553 & n1180 ;
  assign n2645 = n2644 ^ x74 ;
  assign n2657 = n2656 ^ n2645 ;
  assign n2634 = n557 & n1180 ;
  assign n2635 = n2634 ^ x73 ;
  assign n2646 = n2645 ^ n2635 ;
  assign n1944 = n939 & n1180 ;
  assign n1945 = n1944 ^ x72 ;
  assign n2636 = n2635 ^ n1945 ;
  assign n1942 = n1848 & n1941 ;
  assign n1943 = n1942 ^ x328 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1949 = n560 & n1180 ;
  assign n1950 = n1949 ^ x71 ;
  assign n2631 = n1950 ^ n1943 ;
  assign n1947 = n1198 & n1848 ;
  assign n1948 = n1947 ^ x327 ;
  assign n1951 = n1950 ^ n1948 ;
  assign n1954 = n561 & n1180 ;
  assign n1955 = n1954 ^ x70 ;
  assign n2628 = n1955 ^ n1948 ;
  assign n1952 = n1200 & n1848 ;
  assign n1953 = n1952 ^ x326 ;
  assign n1956 = n1955 ^ n1953 ;
  assign n1959 = n576 & n1180 ;
  assign n1960 = n1959 ^ x69 ;
  assign n2625 = n1960 ^ n1953 ;
  assign n1957 = n1213 & n1848 ;
  assign n1958 = n1957 ^ x325 ;
  assign n1961 = n1960 ^ n1958 ;
  assign n2614 = n574 & n1180 ;
  assign n2615 = n2614 ^ x68 ;
  assign n2622 = n2615 ^ n1958 ;
  assign n1964 = n579 & n1180 ;
  assign n1965 = n1964 ^ x67 ;
  assign n2616 = n2615 ^ n1965 ;
  assign n1962 = n1216 & n1848 ;
  assign n1963 = n1962 ^ x323 ;
  assign n1966 = n1965 ^ n1963 ;
  assign n1970 = n1180 & n1969 ;
  assign n1971 = n1970 ^ x66 ;
  assign n2611 = n1971 ^ n1963 ;
  assign n1967 = n1222 & n1848 ;
  assign n1968 = n1967 ^ x322 ;
  assign n1972 = n1971 ^ n1968 ;
  assign n1977 = n1180 & n1976 ;
  assign n1978 = n1977 ^ x65 ;
  assign n2608 = n1978 ^ n1968 ;
  assign n1974 = n1848 & n1973 ;
  assign n1975 = n1974 ^ x321 ;
  assign n1979 = n1978 ^ n1975 ;
  assign n1983 = n1180 & n1982 ;
  assign n1984 = n1983 ^ x64 ;
  assign n2605 = n1984 ^ n1975 ;
  assign n1980 = n1226 & n1848 ;
  assign n1981 = n1980 ^ x320 ;
  assign n1985 = n1984 ^ n1981 ;
  assign n1988 = n583 & n1180 ;
  assign n1989 = n1988 ^ x63 ;
  assign n2602 = n1989 ^ n1981 ;
  assign n1986 = n1241 & n1848 ;
  assign n1987 = n1986 ^ x319 ;
  assign n1990 = n1989 ^ n1987 ;
  assign n1993 = n585 & n1180 ;
  assign n1994 = n1993 ^ x62 ;
  assign n2599 = n1994 ^ n1987 ;
  assign n1991 = n1234 & n1848 ;
  assign n1992 = n1991 ^ x318 ;
  assign n1995 = n1994 ^ n1992 ;
  assign n2588 = n598 & n1180 ;
  assign n2589 = n2588 ^ x61 ;
  assign n2596 = n2589 ^ n1992 ;
  assign n1998 = n603 & n1180 ;
  assign n1999 = n1998 ^ x60 ;
  assign n2590 = n2589 ^ n1999 ;
  assign n1996 = n1247 & n1848 ;
  assign n1997 = n1996 ^ x316 ;
  assign n2000 = n1999 ^ n1997 ;
  assign n2577 = n601 & n1180 ;
  assign n2578 = n2577 ^ x59 ;
  assign n2585 = n2578 ^ n1997 ;
  assign n2569 = n607 & n1180 ;
  assign n2570 = n2569 ^ x58 ;
  assign n2579 = n2578 ^ n2570 ;
  assign n2559 = n1180 & n2558 ;
  assign n2560 = n2559 ^ x57 ;
  assign n2571 = n2570 ^ n2560 ;
  assign n2005 = n1180 & n2004 ;
  assign n2006 = n2005 ^ x56 ;
  assign n2561 = n2560 ^ n2006 ;
  assign n2002 = n1848 & n2001 ;
  assign n2003 = n2002 ^ x312 ;
  assign n2007 = n2006 ^ n2003 ;
  assign n2545 = n1180 & n2544 ;
  assign n2546 = n2545 ^ x55 ;
  assign n2555 = n2546 ^ n2003 ;
  assign n2012 = n1180 & n2011 ;
  assign n2013 = n2012 ^ x54 ;
  assign n2547 = n2546 ^ n2013 ;
  assign n2009 = n1848 & n2008 ;
  assign n2010 = n2009 ^ x310 ;
  assign n2014 = n2013 ^ n2010 ;
  assign n2531 = n1180 & n2530 ;
  assign n2532 = n2531 ^ x53 ;
  assign n2541 = n2532 ^ n2010 ;
  assign n2019 = n1180 & n2018 ;
  assign n2020 = n2019 ^ x52 ;
  assign n2533 = n2532 ^ n2020 ;
  assign n2016 = n1848 & n2015 ;
  assign n2017 = n2016 ^ x308 ;
  assign n2021 = n2020 ^ n2017 ;
  assign n2519 = n1180 & n2518 ;
  assign n2520 = n2519 ^ x51 ;
  assign n2527 = n2520 ^ n2017 ;
  assign n2510 = n1180 & n2509 ;
  assign n2511 = n2510 ^ x50 ;
  assign n2521 = n2520 ^ n2511 ;
  assign n2025 = n1180 & n2024 ;
  assign n2026 = n2025 ^ x49 ;
  assign n2512 = n2511 ^ n2026 ;
  assign n2022 = n1265 & n1848 ;
  assign n2023 = n2022 ^ x305 ;
  assign n2027 = n2026 ^ n2023 ;
  assign n2498 = n611 & n1180 ;
  assign n2499 = n2498 ^ x48 ;
  assign n2506 = n2499 ^ n2023 ;
  assign n2030 = n613 & n1180 ;
  assign n2031 = n2030 ^ x47 ;
  assign n2500 = n2499 ^ n2031 ;
  assign n2028 = n1268 & n1848 ;
  assign n2029 = n2028 ^ x303 ;
  assign n2032 = n2031 ^ n2029 ;
  assign n2035 = n614 & n1180 ;
  assign n2036 = n2035 ^ x46 ;
  assign n2495 = n2036 ^ n2029 ;
  assign n2033 = n1269 & n1848 ;
  assign n2034 = n2033 ^ x302 ;
  assign n2037 = n2036 ^ n2034 ;
  assign n2040 = n627 & n1180 ;
  assign n2041 = n2040 ^ x45 ;
  assign n2492 = n2041 ^ n2034 ;
  assign n2038 = n1282 & n1848 ;
  assign n2039 = n2038 ^ x301 ;
  assign n2042 = n2041 ^ n2039 ;
  assign n2481 = n630 & n1180 ;
  assign n2482 = n2481 ^ x44 ;
  assign n2489 = n2482 ^ n2039 ;
  assign n2473 = n635 & n1180 ;
  assign n2474 = n2473 ^ x43 ;
  assign n2483 = n2482 ^ n2474 ;
  assign n2045 = n636 & n1180 ;
  assign n2046 = n2045 ^ x42 ;
  assign n2475 = n2474 ^ n2046 ;
  assign n2043 = n1291 & n1848 ;
  assign n2044 = n2043 ^ x298 ;
  assign n2047 = n2046 ^ n2044 ;
  assign n2050 = n649 & n1180 ;
  assign n2051 = n2050 ^ x41 ;
  assign n2470 = n2051 ^ n2044 ;
  assign n2048 = n1304 & n1848 ;
  assign n2049 = n2048 ^ x297 ;
  assign n2052 = n2051 ^ n2049 ;
  assign n2055 = n652 & n1180 ;
  assign n2056 = n2055 ^ x40 ;
  assign n2467 = n2056 ^ n2049 ;
  assign n2053 = n1309 & n1848 ;
  assign n2054 = n2053 ^ x296 ;
  assign n2057 = n2056 ^ n2054 ;
  assign n2060 = n657 & n1180 ;
  assign n2061 = n2060 ^ x39 ;
  assign n2464 = n2061 ^ n2054 ;
  assign n2058 = n1307 & n1848 ;
  assign n2059 = n2058 ^ x295 ;
  assign n2062 = n2061 ^ n2059 ;
  assign n2065 = n658 & n1180 ;
  assign n2066 = n2065 ^ x38 ;
  assign n2461 = n2066 ^ n2059 ;
  assign n2063 = n1313 & n1848 ;
  assign n2064 = n2063 ^ x294 ;
  assign n2067 = n2066 ^ n2064 ;
  assign n2448 = n1180 & n2447 ;
  assign n2449 = n2448 ^ x37 ;
  assign n2458 = n2449 ^ n2064 ;
  assign n2072 = n1180 & n2071 ;
  assign n2073 = n2072 ^ x36 ;
  assign n2450 = n2449 ^ n2073 ;
  assign n2069 = n1848 & n2068 ;
  assign n2070 = n2069 ^ x292 ;
  assign n2074 = n2073 ^ n2070 ;
  assign n2079 = n1180 & n2078 ;
  assign n2080 = n2079 ^ x35 ;
  assign n2444 = n2080 ^ n2070 ;
  assign n2076 = n1848 & n2075 ;
  assign n2077 = n2076 ^ x291 ;
  assign n2081 = n2080 ^ n2077 ;
  assign n2431 = n1180 & n2430 ;
  assign n2432 = n2431 ^ x34 ;
  assign n2441 = n2432 ^ n2077 ;
  assign n2086 = n1180 & n2085 ;
  assign n2087 = n2086 ^ x33 ;
  assign n2433 = n2432 ^ n2087 ;
  assign n2083 = n1848 & n2082 ;
  assign n2084 = n2083 ^ x289 ;
  assign n2088 = n2087 ^ n2084 ;
  assign n2093 = n1180 & n2092 ;
  assign n2094 = n2093 ^ x32 ;
  assign n2427 = n2094 ^ n2084 ;
  assign n2090 = n1848 & n2089 ;
  assign n2091 = n2090 ^ x288 ;
  assign n2095 = n2094 ^ n2091 ;
  assign n2100 = n1180 & n2099 ;
  assign n2101 = n2100 ^ x31 ;
  assign n2424 = n2101 ^ n2091 ;
  assign n2097 = n1848 & n2096 ;
  assign n2098 = n2097 ^ x287 ;
  assign n2102 = n2101 ^ n2098 ;
  assign n2411 = n1180 & n2410 ;
  assign n2412 = n2411 ^ x30 ;
  assign n2421 = n2412 ^ n2098 ;
  assign n2107 = n1180 & n2106 ;
  assign n2108 = n2107 ^ x29 ;
  assign n2413 = n2412 ^ n2108 ;
  assign n2104 = n1848 & n2103 ;
  assign n2105 = n2104 ^ x285 ;
  assign n2109 = n2108 ^ n2105 ;
  assign n2114 = n1180 & n2113 ;
  assign n2115 = n2114 ^ x28 ;
  assign n2407 = n2115 ^ n2105 ;
  assign n2111 = n1848 & n2110 ;
  assign n2112 = n2111 ^ x284 ;
  assign n2116 = n2115 ^ n2112 ;
  assign n2394 = n1180 & n2393 ;
  assign n2395 = n2394 ^ x27 ;
  assign n2404 = n2395 ^ n2112 ;
  assign n2121 = n1180 & n2120 ;
  assign n2122 = n2121 ^ x26 ;
  assign n2396 = n2395 ^ n2122 ;
  assign n2118 = n1848 & n2117 ;
  assign n2119 = n2118 ^ x282 ;
  assign n2123 = n2122 ^ n2119 ;
  assign n2128 = n1180 & n2127 ;
  assign n2129 = n2128 ^ x25 ;
  assign n2390 = n2129 ^ n2119 ;
  assign n2125 = n1848 & n2124 ;
  assign n2126 = n2125 ^ x281 ;
  assign n2130 = n2129 ^ n2126 ;
  assign n2135 = n1180 & n2134 ;
  assign n2136 = n2135 ^ x24 ;
  assign n2387 = n2136 ^ n2126 ;
  assign n2132 = n1848 & n2131 ;
  assign n2133 = n2132 ^ x280 ;
  assign n2137 = n2136 ^ n2133 ;
  assign n2374 = n1180 & n2373 ;
  assign n2375 = n2374 ^ x23 ;
  assign n2384 = n2375 ^ n2133 ;
  assign n2363 = n1180 & n2362 ;
  assign n2364 = n2363 ^ x22 ;
  assign n2376 = n2375 ^ n2364 ;
  assign n2352 = n1180 & n2351 ;
  assign n2353 = n2352 ^ x21 ;
  assign n2365 = n2364 ^ n2353 ;
  assign n2142 = n1180 & n2141 ;
  assign n2143 = n2142 ^ x20 ;
  assign n2354 = n2353 ^ n2143 ;
  assign n2139 = n1848 & n2138 ;
  assign n2140 = n2139 ^ x276 ;
  assign n2144 = n2143 ^ n2140 ;
  assign n2338 = n1180 & n2337 ;
  assign n2339 = n2338 ^ x19 ;
  assign n2348 = n2339 ^ n2140 ;
  assign n2149 = n1180 & n2148 ;
  assign n2150 = n2149 ^ x18 ;
  assign n2340 = n2339 ^ n2150 ;
  assign n2146 = n1848 & n2145 ;
  assign n2147 = n2146 ^ x274 ;
  assign n2151 = n2150 ^ n2147 ;
  assign n2156 = n1180 & n2155 ;
  assign n2157 = n2156 ^ x17 ;
  assign n2334 = n2157 ^ n2147 ;
  assign n2153 = n1848 & n2152 ;
  assign n2154 = n2153 ^ x273 ;
  assign n2158 = n2157 ^ n2154 ;
  assign n2321 = n1180 & n2320 ;
  assign n2322 = n2321 ^ x16 ;
  assign n2331 = n2322 ^ n2154 ;
  assign n2163 = n1180 & n2162 ;
  assign n2164 = n2163 ^ x15 ;
  assign n2323 = n2322 ^ n2164 ;
  assign n2160 = n1848 & n2159 ;
  assign n2161 = n2160 ^ x271 ;
  assign n2165 = n2164 ^ n2161 ;
  assign n2307 = n1180 & n2306 ;
  assign n2308 = n2307 ^ x14 ;
  assign n2317 = n2308 ^ n2161 ;
  assign n2296 = n1180 & n2295 ;
  assign n2297 = n2296 ^ x13 ;
  assign n2309 = n2308 ^ n2297 ;
  assign n2170 = n1180 & n2169 ;
  assign n2171 = n2170 ^ x12 ;
  assign n2298 = n2297 ^ n2171 ;
  assign n2167 = n1848 & n2166 ;
  assign n2168 = n2167 ^ x268 ;
  assign n2172 = n2171 ^ n2168 ;
  assign n2177 = n1180 & n2176 ;
  assign n2178 = n2177 ^ x11 ;
  assign n2292 = n2178 ^ n2168 ;
  assign n2174 = n1848 & n2173 ;
  assign n2175 = n2174 ^ x267 ;
  assign n2179 = n2178 ^ n2175 ;
  assign n2184 = n1180 & n2183 ;
  assign n2185 = n2184 ^ x10 ;
  assign n2289 = n2185 ^ n2175 ;
  assign n2181 = n1848 & n2180 ;
  assign n2182 = n2181 ^ x266 ;
  assign n2186 = n2185 ^ n2182 ;
  assign n2276 = n1180 & n2275 ;
  assign n2277 = n2276 ^ x9 ;
  assign n2286 = n2277 ^ n2182 ;
  assign n2265 = n1180 & n2264 ;
  assign n2266 = n2265 ^ x8 ;
  assign n2278 = n2277 ^ n2266 ;
  assign n2191 = n1180 & n2190 ;
  assign n2192 = n2191 ^ x7 ;
  assign n2267 = n2266 ^ n2192 ;
  assign n2188 = n1848 & n2187 ;
  assign n2189 = n2188 ^ x263 ;
  assign n2193 = n2192 ^ n2189 ;
  assign n2251 = n1180 & n2250 ;
  assign n2252 = n2251 ^ x6 ;
  assign n2261 = n2252 ^ n2189 ;
  assign n2198 = n1180 & n2197 ;
  assign n2199 = n2198 ^ x5 ;
  assign n2253 = n2252 ^ n2199 ;
  assign n2195 = n1848 & n2194 ;
  assign n2196 = n2195 ^ x261 ;
  assign n2200 = n2199 ^ n2196 ;
  assign n2205 = n1180 & n2204 ;
  assign n2206 = n2205 ^ x4 ;
  assign n2247 = n2206 ^ n2196 ;
  assign n2202 = n1848 & n2201 ;
  assign n2203 = n2202 ^ x260 ;
  assign n2207 = n2206 ^ n2203 ;
  assign n2234 = n1180 & n2233 ;
  assign n2235 = n2234 ^ x3 ;
  assign n2244 = n2235 ^ n2203 ;
  assign n2223 = n1180 & n2222 ;
  assign n2224 = n2223 ^ x2 ;
  assign n2236 = n2235 ^ n2224 ;
  assign n2212 = n1180 & n2211 ;
  assign n2213 = n2212 ^ x1 ;
  assign n2225 = n2224 ^ n2213 ;
  assign n2209 = n1848 & n2208 ;
  assign n2210 = n2209 ^ x257 ;
  assign n2214 = n2213 ^ n2210 ;
  assign n2219 = n1182 & ~n1850 ;
  assign n2220 = n2219 ^ n2210 ;
  assign n2221 = ~n2214 & n2220 ;
  assign n2226 = n2225 ^ n2221 ;
  assign n2227 = n2224 ^ x258 ;
  assign n2228 = n2227 ^ x386 ;
  assign n2229 = n2228 ^ n2224 ;
  assign n2230 = n1848 & n2229 ;
  assign n2231 = n2230 ^ n2227 ;
  assign n2232 = n2226 & ~n2231 ;
  assign n2237 = n2236 ^ n2232 ;
  assign n2238 = n2235 ^ x259 ;
  assign n2239 = n2238 ^ x387 ;
  assign n2240 = n2239 ^ n2235 ;
  assign n2241 = n1848 & n2240 ;
  assign n2242 = n2241 ^ n2238 ;
  assign n2243 = n2237 & ~n2242 ;
  assign n2245 = n2244 ^ n2243 ;
  assign n2246 = ~n2207 & n2245 ;
  assign n2248 = n2247 ^ n2246 ;
  assign n2249 = ~n2200 & n2248 ;
  assign n2254 = n2253 ^ n2249 ;
  assign n2255 = n2252 ^ x262 ;
  assign n2256 = n2255 ^ x390 ;
  assign n2257 = n2256 ^ n2252 ;
  assign n2258 = n1848 & n2257 ;
  assign n2259 = n2258 ^ n2255 ;
  assign n2260 = n2254 & ~n2259 ;
  assign n2262 = n2261 ^ n2260 ;
  assign n2263 = ~n2193 & n2262 ;
  assign n2268 = n2267 ^ n2263 ;
  assign n2269 = n2266 ^ x264 ;
  assign n2270 = n2269 ^ x392 ;
  assign n2271 = n2270 ^ n2266 ;
  assign n2272 = n1848 & n2271 ;
  assign n2273 = n2272 ^ n2269 ;
  assign n2274 = n2268 & ~n2273 ;
  assign n2279 = n2278 ^ n2274 ;
  assign n2280 = n2277 ^ x265 ;
  assign n2281 = n2280 ^ x393 ;
  assign n2282 = n2281 ^ n2277 ;
  assign n2283 = n1848 & n2282 ;
  assign n2284 = n2283 ^ n2280 ;
  assign n2285 = n2279 & ~n2284 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2288 = ~n2186 & n2287 ;
  assign n2290 = n2289 ^ n2288 ;
  assign n2291 = ~n2179 & n2290 ;
  assign n2293 = n2292 ^ n2291 ;
  assign n2294 = ~n2172 & n2293 ;
  assign n2299 = n2298 ^ n2294 ;
  assign n2300 = n2297 ^ x269 ;
  assign n2301 = n2300 ^ x397 ;
  assign n2302 = n2301 ^ n2297 ;
  assign n2303 = n1848 & n2302 ;
  assign n2304 = n2303 ^ n2300 ;
  assign n2305 = n2299 & ~n2304 ;
  assign n2310 = n2309 ^ n2305 ;
  assign n2311 = n2308 ^ x270 ;
  assign n2312 = n2311 ^ x398 ;
  assign n2313 = n2312 ^ n2308 ;
  assign n2314 = n1848 & n2313 ;
  assign n2315 = n2314 ^ n2311 ;
  assign n2316 = n2310 & ~n2315 ;
  assign n2318 = n2317 ^ n2316 ;
  assign n2319 = ~n2165 & n2318 ;
  assign n2324 = n2323 ^ n2319 ;
  assign n2325 = n2322 ^ x272 ;
  assign n2326 = n2325 ^ x400 ;
  assign n2327 = n2326 ^ n2322 ;
  assign n2328 = n1848 & n2327 ;
  assign n2329 = n2328 ^ n2325 ;
  assign n2330 = n2324 & ~n2329 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2333 = ~n2158 & n2332 ;
  assign n2335 = n2334 ^ n2333 ;
  assign n2336 = ~n2151 & n2335 ;
  assign n2341 = n2340 ^ n2336 ;
  assign n2342 = n2339 ^ x275 ;
  assign n2343 = n2342 ^ x403 ;
  assign n2344 = n2343 ^ n2339 ;
  assign n2345 = n1848 & n2344 ;
  assign n2346 = n2345 ^ n2342 ;
  assign n2347 = n2341 & ~n2346 ;
  assign n2349 = n2348 ^ n2347 ;
  assign n2350 = ~n2144 & n2349 ;
  assign n2355 = n2354 ^ n2350 ;
  assign n2356 = n2353 ^ x277 ;
  assign n2357 = n2356 ^ x405 ;
  assign n2358 = n2357 ^ n2353 ;
  assign n2359 = n1848 & n2358 ;
  assign n2360 = n2359 ^ n2356 ;
  assign n2361 = n2355 & ~n2360 ;
  assign n2366 = n2365 ^ n2361 ;
  assign n2367 = n2364 ^ x278 ;
  assign n2368 = n2367 ^ x406 ;
  assign n2369 = n2368 ^ n2364 ;
  assign n2370 = n1848 & n2369 ;
  assign n2371 = n2370 ^ n2367 ;
  assign n2372 = n2366 & ~n2371 ;
  assign n2377 = n2376 ^ n2372 ;
  assign n2378 = n2375 ^ x279 ;
  assign n2379 = n2378 ^ x407 ;
  assign n2380 = n2379 ^ n2375 ;
  assign n2381 = n1848 & n2380 ;
  assign n2382 = n2381 ^ n2378 ;
  assign n2383 = n2377 & ~n2382 ;
  assign n2385 = n2384 ^ n2383 ;
  assign n2386 = ~n2137 & n2385 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2389 = ~n2130 & n2388 ;
  assign n2391 = n2390 ^ n2389 ;
  assign n2392 = ~n2123 & n2391 ;
  assign n2397 = n2396 ^ n2392 ;
  assign n2398 = n2395 ^ x283 ;
  assign n2399 = n2398 ^ x411 ;
  assign n2400 = n2399 ^ n2395 ;
  assign n2401 = n1848 & n2400 ;
  assign n2402 = n2401 ^ n2398 ;
  assign n2403 = n2397 & ~n2402 ;
  assign n2405 = n2404 ^ n2403 ;
  assign n2406 = ~n2116 & n2405 ;
  assign n2408 = n2407 ^ n2406 ;
  assign n2409 = ~n2109 & n2408 ;
  assign n2414 = n2413 ^ n2409 ;
  assign n2415 = n2412 ^ x286 ;
  assign n2416 = n2415 ^ x414 ;
  assign n2417 = n2416 ^ n2412 ;
  assign n2418 = n1848 & n2417 ;
  assign n2419 = n2418 ^ n2415 ;
  assign n2420 = n2414 & ~n2419 ;
  assign n2422 = n2421 ^ n2420 ;
  assign n2423 = ~n2102 & n2422 ;
  assign n2425 = n2424 ^ n2423 ;
  assign n2426 = ~n2095 & n2425 ;
  assign n2428 = n2427 ^ n2426 ;
  assign n2429 = ~n2088 & n2428 ;
  assign n2434 = n2433 ^ n2429 ;
  assign n2435 = n2432 ^ x290 ;
  assign n2436 = n2435 ^ x418 ;
  assign n2437 = n2436 ^ n2432 ;
  assign n2438 = n1848 & n2437 ;
  assign n2439 = n2438 ^ n2435 ;
  assign n2440 = n2434 & ~n2439 ;
  assign n2442 = n2441 ^ n2440 ;
  assign n2443 = ~n2081 & n2442 ;
  assign n2445 = n2444 ^ n2443 ;
  assign n2446 = ~n2074 & n2445 ;
  assign n2451 = n2450 ^ n2446 ;
  assign n2452 = n2449 ^ x293 ;
  assign n2453 = n2452 ^ x421 ;
  assign n2454 = n2453 ^ n2449 ;
  assign n2455 = n1848 & n2454 ;
  assign n2456 = n2455 ^ n2452 ;
  assign n2457 = n2451 & ~n2456 ;
  assign n2459 = n2458 ^ n2457 ;
  assign n2460 = ~n2067 & n2459 ;
  assign n2462 = n2461 ^ n2460 ;
  assign n2463 = ~n2062 & n2462 ;
  assign n2465 = n2464 ^ n2463 ;
  assign n2466 = ~n2057 & n2465 ;
  assign n2468 = n2467 ^ n2466 ;
  assign n2469 = ~n2052 & n2468 ;
  assign n2471 = n2470 ^ n2469 ;
  assign n2472 = ~n2047 & n2471 ;
  assign n2476 = n2475 ^ n2472 ;
  assign n2478 = n1290 & n1848 ;
  assign n2477 = n2474 ^ x299 ;
  assign n2479 = n2478 ^ n2477 ;
  assign n2480 = n2476 & ~n2479 ;
  assign n2484 = n2483 ^ n2480 ;
  assign n2486 = n1285 & n1848 ;
  assign n2485 = n2482 ^ x300 ;
  assign n2487 = n2486 ^ n2485 ;
  assign n2488 = n2484 & ~n2487 ;
  assign n2490 = n2489 ^ n2488 ;
  assign n2491 = ~n2042 & n2490 ;
  assign n2493 = n2492 ^ n2491 ;
  assign n2494 = ~n2037 & n2493 ;
  assign n2496 = n2495 ^ n2494 ;
  assign n2497 = ~n2032 & n2496 ;
  assign n2501 = n2500 ^ n2497 ;
  assign n2503 = n1513 & n1848 ;
  assign n2502 = n2499 ^ x304 ;
  assign n2504 = n2503 ^ n2502 ;
  assign n2505 = n2501 & ~n2504 ;
  assign n2507 = n2506 ^ n2505 ;
  assign n2508 = ~n2027 & n2507 ;
  assign n2513 = n2512 ^ n2508 ;
  assign n2515 = n1261 & n1848 ;
  assign n2514 = n2511 ^ x306 ;
  assign n2516 = n2515 ^ n2514 ;
  assign n2517 = n2513 & ~n2516 ;
  assign n2522 = n2521 ^ n2517 ;
  assign n2524 = n1256 & n1848 ;
  assign n2523 = n2520 ^ x307 ;
  assign n2525 = n2524 ^ n2523 ;
  assign n2526 = n2522 & ~n2525 ;
  assign n2528 = n2527 ^ n2526 ;
  assign n2529 = ~n2021 & n2528 ;
  assign n2534 = n2533 ^ n2529 ;
  assign n2535 = n2532 ^ x309 ;
  assign n2536 = n2535 ^ x437 ;
  assign n2537 = n2536 ^ n2532 ;
  assign n2538 = n1848 & n2537 ;
  assign n2539 = n2538 ^ n2535 ;
  assign n2540 = n2534 & ~n2539 ;
  assign n2542 = n2541 ^ n2540 ;
  assign n2543 = ~n2014 & n2542 ;
  assign n2548 = n2547 ^ n2543 ;
  assign n2549 = n2546 ^ x311 ;
  assign n2550 = n2549 ^ x439 ;
  assign n2551 = n2550 ^ n2546 ;
  assign n2552 = n1848 & n2551 ;
  assign n2553 = n2552 ^ n2549 ;
  assign n2554 = n2548 & ~n2553 ;
  assign n2556 = n2555 ^ n2554 ;
  assign n2557 = ~n2007 & n2556 ;
  assign n2562 = n2561 ^ n2557 ;
  assign n2563 = n2560 ^ x313 ;
  assign n2564 = n2563 ^ x441 ;
  assign n2565 = n2564 ^ n2560 ;
  assign n2566 = n1848 & n2565 ;
  assign n2567 = n2566 ^ n2563 ;
  assign n2568 = n2562 & ~n2567 ;
  assign n2572 = n2571 ^ n2568 ;
  assign n2574 = n1252 & n1848 ;
  assign n2573 = n2570 ^ x314 ;
  assign n2575 = n2574 ^ n2573 ;
  assign n2576 = n2572 & ~n2575 ;
  assign n2580 = n2579 ^ n2576 ;
  assign n2582 = n1250 & n1848 ;
  assign n2581 = n2578 ^ x315 ;
  assign n2583 = n2582 ^ n2581 ;
  assign n2584 = n2580 & ~n2583 ;
  assign n2586 = n2585 ^ n2584 ;
  assign n2587 = ~n2000 & n2586 ;
  assign n2591 = n2590 ^ n2587 ;
  assign n2593 = n1232 & n1848 ;
  assign n2592 = n2589 ^ x317 ;
  assign n2594 = n2593 ^ n2592 ;
  assign n2595 = n2591 & ~n2594 ;
  assign n2597 = n2596 ^ n2595 ;
  assign n2598 = ~n1995 & n2597 ;
  assign n2600 = n2599 ^ n2598 ;
  assign n2601 = ~n1990 & n2600 ;
  assign n2603 = n2602 ^ n2601 ;
  assign n2604 = ~n1985 & n2603 ;
  assign n2606 = n2605 ^ n2604 ;
  assign n2607 = ~n1979 & n2606 ;
  assign n2609 = n2608 ^ n2607 ;
  assign n2610 = ~n1972 & n2609 ;
  assign n2612 = n2611 ^ n2610 ;
  assign n2613 = ~n1966 & n2612 ;
  assign n2617 = n2616 ^ n2613 ;
  assign n2619 = n1218 & n1848 ;
  assign n2618 = n2615 ^ x324 ;
  assign n2620 = n2619 ^ n2618 ;
  assign n2621 = n2617 & ~n2620 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2624 = ~n1961 & n2623 ;
  assign n2626 = n2625 ^ n2624 ;
  assign n2627 = ~n1956 & n2626 ;
  assign n2629 = n2628 ^ n2627 ;
  assign n2630 = ~n1951 & n2629 ;
  assign n2632 = n2631 ^ n2630 ;
  assign n2633 = ~n1946 & n2632 ;
  assign n2637 = n2636 ^ n2633 ;
  assign n2638 = n2635 ^ x329 ;
  assign n2639 = n2638 ^ x457 ;
  assign n2640 = n2639 ^ n2635 ;
  assign n2641 = n1848 & n2640 ;
  assign n2642 = n2641 ^ n2638 ;
  assign n2643 = n2637 & ~n2642 ;
  assign n2647 = n2646 ^ n2643 ;
  assign n2648 = n2645 ^ x330 ;
  assign n2649 = n2648 ^ x458 ;
  assign n2650 = n2649 ^ n2645 ;
  assign n2651 = n1848 & n2650 ;
  assign n2652 = n2651 ^ n2648 ;
  assign n2653 = n2647 & ~n2652 ;
  assign n2658 = n2657 ^ n2653 ;
  assign n2659 = n2656 ^ x75 ;
  assign n2660 = n2659 ^ x203 ;
  assign n2661 = n2660 ^ n2656 ;
  assign n2662 = n1180 & n2661 ;
  assign n2663 = n2662 ^ n2659 ;
  assign n2664 = ~n2658 & ~n2663 ;
  assign n2668 = n2667 ^ n2664 ;
  assign n2669 = n2666 ^ x332 ;
  assign n2670 = n2669 ^ x460 ;
  assign n2671 = n2670 ^ n2666 ;
  assign n2672 = n1848 & n2671 ;
  assign n2673 = n2672 ^ n2669 ;
  assign n2674 = ~n2668 & ~n2673 ;
  assign n2678 = n2677 ^ n2674 ;
  assign n2679 = n2676 ^ x333 ;
  assign n2680 = n2679 ^ x461 ;
  assign n2681 = n2680 ^ n2676 ;
  assign n2682 = n1848 & n2681 ;
  assign n2683 = n2682 ^ n2679 ;
  assign n2684 = n2678 & ~n2683 ;
  assign n2688 = n2687 ^ n2684 ;
  assign n2689 = n2686 ^ x334 ;
  assign n2690 = n2689 ^ x462 ;
  assign n2691 = n2690 ^ n2686 ;
  assign n2692 = n1848 & n2691 ;
  assign n2693 = n2692 ^ n2689 ;
  assign n2694 = n2688 & ~n2693 ;
  assign n2698 = n2697 ^ n2694 ;
  assign n2699 = n2696 ^ x335 ;
  assign n2700 = n2699 ^ x463 ;
  assign n2701 = n2700 ^ n2696 ;
  assign n2702 = n1848 & n2701 ;
  assign n2703 = n2702 ^ n2699 ;
  assign n2704 = n2698 & ~n2703 ;
  assign n2706 = n2705 ^ n2704 ;
  assign n2707 = ~n1940 & n2706 ;
  assign n2709 = n2708 ^ n2707 ;
  assign n2710 = ~n1934 & n2709 ;
  assign n2715 = n2714 ^ n2710 ;
  assign n2716 = n2713 ^ x82 ;
  assign n2717 = n2716 ^ x210 ;
  assign n2718 = n2717 ^ n2713 ;
  assign n2719 = n1180 & n2718 ;
  assign n2720 = n2719 ^ n2716 ;
  assign n2721 = ~n2715 & ~n2720 ;
  assign n2726 = n2725 ^ n2721 ;
  assign n2727 = n2724 ^ x339 ;
  assign n2728 = n2727 ^ x467 ;
  assign n2729 = n2728 ^ n2724 ;
  assign n2730 = n1848 & n2729 ;
  assign n2731 = n2730 ^ n2727 ;
  assign n2732 = ~n2726 & ~n2731 ;
  assign n2737 = n2736 ^ n2732 ;
  assign n2738 = n2735 ^ x340 ;
  assign n2739 = n2738 ^ x468 ;
  assign n2740 = n2739 ^ n2735 ;
  assign n2741 = n1848 & n2740 ;
  assign n2742 = n2741 ^ n2738 ;
  assign n2743 = n2737 & ~n2742 ;
  assign n2748 = n2747 ^ n2743 ;
  assign n2749 = n2746 ^ x341 ;
  assign n2750 = n2749 ^ x469 ;
  assign n2751 = n2750 ^ n2746 ;
  assign n2752 = n1848 & n2751 ;
  assign n2753 = n2752 ^ n2749 ;
  assign n2754 = n2748 & ~n2753 ;
  assign n2759 = n2758 ^ n2754 ;
  assign n2760 = n2757 ^ x342 ;
  assign n2761 = n2760 ^ x470 ;
  assign n2762 = n2761 ^ n2757 ;
  assign n2763 = n1848 & n2762 ;
  assign n2764 = n2763 ^ n2760 ;
  assign n2765 = n2759 & ~n2764 ;
  assign n2770 = n2769 ^ n2765 ;
  assign n2771 = n2768 ^ x343 ;
  assign n2772 = n2771 ^ x471 ;
  assign n2773 = n2772 ^ n2768 ;
  assign n2774 = n1848 & n2773 ;
  assign n2775 = n2774 ^ n2771 ;
  assign n2776 = n2770 & ~n2775 ;
  assign n2781 = n2780 ^ n2776 ;
  assign n2782 = n2779 ^ x88 ;
  assign n2783 = n2782 ^ x216 ;
  assign n2784 = n2783 ^ n2779 ;
  assign n2785 = n1180 & n2784 ;
  assign n2786 = n2785 ^ n2782 ;
  assign n2787 = ~n2781 & ~n2786 ;
  assign n2792 = n2791 ^ n2787 ;
  assign n2793 = n2790 ^ x89 ;
  assign n2794 = n2793 ^ x217 ;
  assign n2795 = n2794 ^ n2790 ;
  assign n2796 = n1180 & n2795 ;
  assign n2797 = n2796 ^ n2793 ;
  assign n2798 = n2792 & ~n2797 ;
  assign n2803 = n2802 ^ n2798 ;
  assign n2804 = n2801 ^ x90 ;
  assign n2805 = n2804 ^ x218 ;
  assign n2806 = n2805 ^ n2801 ;
  assign n2807 = n1180 & n2806 ;
  assign n2808 = n2807 ^ n2804 ;
  assign n2809 = n2803 & ~n2808 ;
  assign n2814 = n2813 ^ n2809 ;
  assign n2815 = n2812 ^ x347 ;
  assign n2816 = n2815 ^ x475 ;
  assign n2817 = n2816 ^ n2812 ;
  assign n2818 = n1848 & n2817 ;
  assign n2819 = n2818 ^ n2815 ;
  assign n2820 = ~n2814 & ~n2819 ;
  assign n2825 = n2824 ^ n2820 ;
  assign n2826 = n2823 ^ x348 ;
  assign n2827 = n2826 ^ x476 ;
  assign n2828 = n2827 ^ n2823 ;
  assign n2829 = n1848 & n2828 ;
  assign n2830 = n2829 ^ n2826 ;
  assign n2831 = n2825 & ~n2830 ;
  assign n2836 = n2835 ^ n2831 ;
  assign n2837 = n2834 ^ x349 ;
  assign n2838 = n2837 ^ x477 ;
  assign n2839 = n2838 ^ n2834 ;
  assign n2840 = n1848 & n2839 ;
  assign n2841 = n2840 ^ n2837 ;
  assign n2842 = n2836 & ~n2841 ;
  assign n2847 = n2846 ^ n2842 ;
  assign n2848 = n2845 ^ x94 ;
  assign n2849 = n2848 ^ x222 ;
  assign n2850 = n2849 ^ n2845 ;
  assign n2851 = n1180 & n2850 ;
  assign n2852 = n2851 ^ n2848 ;
  assign n2853 = ~n2847 & ~n2852 ;
  assign n2858 = n2857 ^ n2853 ;
  assign n2859 = n2856 ^ x95 ;
  assign n2860 = n2859 ^ x223 ;
  assign n2861 = n2860 ^ n2856 ;
  assign n2862 = n1180 & n2861 ;
  assign n2863 = n2862 ^ n2859 ;
  assign n2864 = n2858 & ~n2863 ;
  assign n2866 = n2865 ^ n2864 ;
  assign n2867 = ~n1927 & ~n2866 ;
  assign n2869 = n2868 ^ n2867 ;
  assign n2870 = ~n1920 & n2869 ;
  assign n2875 = n2874 ^ n2870 ;
  assign n2876 = n2873 ^ x98 ;
  assign n2877 = n2876 ^ x226 ;
  assign n2878 = n2877 ^ n2873 ;
  assign n2879 = n1180 & n2878 ;
  assign n2880 = n2879 ^ n2876 ;
  assign n2881 = ~n2875 & ~n2880 ;
  assign n2886 = n2885 ^ n2881 ;
  assign n2887 = n2884 ^ x99 ;
  assign n2888 = n2887 ^ x227 ;
  assign n2889 = n2888 ^ n2884 ;
  assign n2890 = n1180 & n2889 ;
  assign n2891 = n2890 ^ n2887 ;
  assign n2892 = n2886 & ~n2891 ;
  assign n2894 = n2893 ^ n2892 ;
  assign n2895 = ~n1913 & ~n2894 ;
  assign n2897 = n2896 ^ n2895 ;
  assign n2898 = ~n1906 & n2897 ;
  assign n2903 = n2902 ^ n2898 ;
  assign n2904 = n2901 ^ x102 ;
  assign n2905 = n2904 ^ x230 ;
  assign n2906 = n2905 ^ n2901 ;
  assign n2907 = n1180 & n2906 ;
  assign n2908 = n2907 ^ n2904 ;
  assign n2909 = ~n2903 & ~n2908 ;
  assign n2914 = n2913 ^ n2909 ;
  assign n2915 = n2912 ^ x359 ;
  assign n2916 = n2915 ^ x487 ;
  assign n2917 = n2916 ^ n2912 ;
  assign n2918 = n1848 & n2917 ;
  assign n2919 = n2918 ^ n2915 ;
  assign n2920 = ~n2914 & ~n2919 ;
  assign n2922 = n2921 ^ n2920 ;
  assign n2923 = ~n1899 & n2922 ;
  assign n2928 = n2927 ^ n2923 ;
  assign n2929 = n2926 ^ x105 ;
  assign n2930 = n2929 ^ x233 ;
  assign n2931 = n2930 ^ n2926 ;
  assign n2932 = n1180 & n2931 ;
  assign n2933 = n2932 ^ n2929 ;
  assign n2934 = ~n2928 & ~n2933 ;
  assign n2939 = n2938 ^ n2934 ;
  assign n2940 = n2937 ^ x362 ;
  assign n2941 = n2940 ^ x490 ;
  assign n2942 = n2941 ^ n2937 ;
  assign n2943 = n1848 & n2942 ;
  assign n2944 = n2943 ^ n2940 ;
  assign n2945 = ~n2939 & ~n2944 ;
  assign n2950 = n2949 ^ n2945 ;
  assign n2951 = n2948 ^ x363 ;
  assign n2952 = n2951 ^ x491 ;
  assign n2953 = n2952 ^ n2948 ;
  assign n2954 = n1848 & n2953 ;
  assign n2955 = n2954 ^ n2951 ;
  assign n2956 = n2950 & ~n2955 ;
  assign n2958 = n2957 ^ n2956 ;
  assign n2959 = ~n1892 & n2958 ;
  assign n2961 = n2960 ^ n2959 ;
  assign n2962 = ~n1885 & n2961 ;
  assign n2964 = n2963 ^ n2962 ;
  assign n2965 = ~n1878 & n2964 ;
  assign n2970 = n2969 ^ n2965 ;
  assign n2971 = n2968 ^ x111 ;
  assign n2972 = n2971 ^ x239 ;
  assign n2973 = n2972 ^ n2968 ;
  assign n2974 = n1180 & n2973 ;
  assign n2975 = n2974 ^ n2971 ;
  assign n2976 = ~n2970 & ~n2975 ;
  assign n2981 = n2980 ^ n2976 ;
  assign n2982 = n2979 ^ x112 ;
  assign n2983 = n2982 ^ x240 ;
  assign n2984 = n2983 ^ n2979 ;
  assign n2985 = n1180 & n2984 ;
  assign n2986 = n2985 ^ n2982 ;
  assign n2987 = n2981 & ~n2986 ;
  assign n2992 = n2991 ^ n2987 ;
  assign n2993 = n2990 ^ x369 ;
  assign n2994 = n2993 ^ x497 ;
  assign n2995 = n2994 ^ n2990 ;
  assign n2996 = n1848 & n2995 ;
  assign n2997 = n2996 ^ n2993 ;
  assign n2998 = ~n2992 & ~n2997 ;
  assign n3003 = n3002 ^ n2998 ;
  assign n3004 = n3001 ^ x114 ;
  assign n3005 = n3004 ^ x242 ;
  assign n3006 = n3005 ^ n3001 ;
  assign n3007 = n1180 & n3006 ;
  assign n3008 = n3007 ^ n3004 ;
  assign n3009 = ~n3003 & ~n3008 ;
  assign n3014 = n3013 ^ n3009 ;
  assign n3015 = n3012 ^ x115 ;
  assign n3016 = n3015 ^ x243 ;
  assign n3017 = n3016 ^ n3012 ;
  assign n3018 = n1180 & n3017 ;
  assign n3019 = n3018 ^ n3015 ;
  assign n3020 = n3014 & ~n3019 ;
  assign n3025 = n3024 ^ n3020 ;
  assign n3026 = n3023 ^ x372 ;
  assign n3027 = n3026 ^ x500 ;
  assign n3028 = n3027 ^ n3023 ;
  assign n3029 = n1848 & n3028 ;
  assign n3030 = n3029 ^ n3026 ;
  assign n3031 = ~n3025 & ~n3030 ;
  assign n3036 = n3035 ^ n3031 ;
  assign n3037 = n3034 ^ x373 ;
  assign n3038 = n3037 ^ x501 ;
  assign n3039 = n3038 ^ n3034 ;
  assign n3040 = n1848 & n3039 ;
  assign n3041 = n3040 ^ n3037 ;
  assign n3042 = n3036 & ~n3041 ;
  assign n3047 = n3046 ^ n3042 ;
  assign n3048 = n3045 ^ x374 ;
  assign n3049 = n3048 ^ x502 ;
  assign n3050 = n3049 ^ n3045 ;
  assign n3051 = n1848 & n3050 ;
  assign n3052 = n3051 ^ n3048 ;
  assign n3053 = n3047 & ~n3052 ;
  assign n3058 = n3057 ^ n3053 ;
  assign n3059 = n3056 ^ x375 ;
  assign n3060 = n3059 ^ x503 ;
  assign n3061 = n3060 ^ n3056 ;
  assign n3062 = n1848 & n3061 ;
  assign n3063 = n3062 ^ n3059 ;
  assign n3064 = n3058 & ~n3063 ;
  assign n3066 = n3065 ^ n3064 ;
  assign n3067 = ~n1871 & n3066 ;
  assign n3069 = n3068 ^ n3067 ;
  assign n3070 = ~n1864 & n3069 ;
  assign n3074 = n3073 ^ n3070 ;
  assign n3076 = n1194 & n1848 ;
  assign n3075 = n3072 ^ x378 ;
  assign n3077 = n3076 ^ n3075 ;
  assign n3078 = n3074 & ~n3077 ;
  assign n3082 = n3081 ^ n3078 ;
  assign n3083 = n3080 ^ x123 ;
  assign n3084 = n3083 ^ x251 ;
  assign n3085 = n3084 ^ n3080 ;
  assign n3086 = n1180 & n3085 ;
  assign n3087 = n3086 ^ n3083 ;
  assign n3088 = ~n3082 & ~n3087 ;
  assign n3092 = n3091 ^ n3088 ;
  assign n3093 = n3090 ^ x124 ;
  assign n3094 = n3093 ^ x252 ;
  assign n3095 = n3094 ^ n3090 ;
  assign n3096 = n1180 & n3095 ;
  assign n3097 = n3096 ^ n3093 ;
  assign n3098 = n3092 & ~n3097 ;
  assign n3102 = n3101 ^ n3098 ;
  assign n3103 = n3100 ^ x381 ;
  assign n3104 = n3103 ^ x509 ;
  assign n3105 = n3104 ^ n3100 ;
  assign n3106 = n1848 & n3105 ;
  assign n3107 = n3106 ^ n3103 ;
  assign n3108 = ~n3102 & ~n3107 ;
  assign n3110 = n3109 ^ n3108 ;
  assign n3112 = n1186 & n1848 ;
  assign n3111 = n1856 ^ x382 ;
  assign n3113 = n3112 ^ n3111 ;
  assign n3114 = n3110 & ~n3113 ;
  assign n1857 = n1856 ^ n1853 ;
  assign n3115 = n3114 ^ n1857 ;
  assign n3116 = ~n1854 & n3115 ;
  assign n3117 = n3116 ^ n1853 ;
  assign n3118 = n1851 & n3117 ;
  assign n3119 = n3118 ^ n1850 ;
  assign n3120 = n2214 & ~n3117 ;
  assign n3121 = n3120 ^ n2213 ;
  assign n3122 = n2231 & ~n3117 ;
  assign n3123 = n3122 ^ n2224 ;
  assign n3124 = n2242 & ~n3117 ;
  assign n3125 = n3124 ^ n2235 ;
  assign n3126 = n2207 & ~n3117 ;
  assign n3127 = n3126 ^ n2206 ;
  assign n3128 = n2200 & ~n3117 ;
  assign n3129 = n3128 ^ n2199 ;
  assign n3130 = n2259 & ~n3117 ;
  assign n3131 = n3130 ^ n2252 ;
  assign n3132 = n2193 & ~n3117 ;
  assign n3133 = n3132 ^ n2192 ;
  assign n3134 = n2273 & ~n3117 ;
  assign n3135 = n3134 ^ n2266 ;
  assign n3136 = n2284 & ~n3117 ;
  assign n3137 = n3136 ^ n2277 ;
  assign n3138 = n2186 & ~n3117 ;
  assign n3139 = n3138 ^ n2185 ;
  assign n3140 = n2179 & ~n3117 ;
  assign n3141 = n3140 ^ n2178 ;
  assign n3142 = n2172 & ~n3117 ;
  assign n3143 = n3142 ^ n2171 ;
  assign n3144 = n2304 & ~n3117 ;
  assign n3145 = n3144 ^ n2297 ;
  assign n3146 = n2315 & ~n3117 ;
  assign n3147 = n3146 ^ n2308 ;
  assign n3148 = n2165 & ~n3117 ;
  assign n3149 = n3148 ^ n2164 ;
  assign n3150 = n2329 & ~n3117 ;
  assign n3151 = n3150 ^ n2322 ;
  assign n3152 = n2158 & ~n3117 ;
  assign n3153 = n3152 ^ n2157 ;
  assign n3154 = n2151 & ~n3117 ;
  assign n3155 = n3154 ^ n2150 ;
  assign n3156 = n2346 & ~n3117 ;
  assign n3157 = n3156 ^ n2339 ;
  assign n3158 = n2144 & ~n3117 ;
  assign n3159 = n3158 ^ n2143 ;
  assign n3160 = n2360 & ~n3117 ;
  assign n3161 = n3160 ^ n2353 ;
  assign n3162 = n2371 & ~n3117 ;
  assign n3163 = n3162 ^ n2364 ;
  assign n3164 = n2382 & ~n3117 ;
  assign n3165 = n3164 ^ n2375 ;
  assign n3166 = n2137 & ~n3117 ;
  assign n3167 = n3166 ^ n2136 ;
  assign n3168 = n2130 & ~n3117 ;
  assign n3169 = n3168 ^ n2129 ;
  assign n3170 = n2123 & ~n3117 ;
  assign n3171 = n3170 ^ n2122 ;
  assign n3172 = n2402 & ~n3117 ;
  assign n3173 = n3172 ^ n2395 ;
  assign n3174 = n2116 & ~n3117 ;
  assign n3175 = n3174 ^ n2115 ;
  assign n3176 = n2109 & ~n3117 ;
  assign n3177 = n3176 ^ n2108 ;
  assign n3178 = n2419 & ~n3117 ;
  assign n3179 = n3178 ^ n2412 ;
  assign n3180 = n2102 & ~n3117 ;
  assign n3181 = n3180 ^ n2101 ;
  assign n3182 = n2095 & ~n3117 ;
  assign n3183 = n3182 ^ n2094 ;
  assign n3184 = n2088 & ~n3117 ;
  assign n3185 = n3184 ^ n2087 ;
  assign n3186 = n2439 & ~n3117 ;
  assign n3187 = n3186 ^ n2432 ;
  assign n3188 = n2081 & ~n3117 ;
  assign n3189 = n3188 ^ n2080 ;
  assign n3190 = n2074 & ~n3117 ;
  assign n3191 = n3190 ^ n2073 ;
  assign n3192 = n2456 & ~n3117 ;
  assign n3193 = n3192 ^ n2449 ;
  assign n3194 = n2067 & ~n3117 ;
  assign n3195 = n3194 ^ n2066 ;
  assign n3196 = n2062 & ~n3117 ;
  assign n3197 = n3196 ^ n2061 ;
  assign n3198 = n2057 & ~n3117 ;
  assign n3199 = n3198 ^ n2056 ;
  assign n3200 = n2052 & ~n3117 ;
  assign n3201 = n3200 ^ n2051 ;
  assign n3202 = n2047 & ~n3117 ;
  assign n3203 = n3202 ^ n2046 ;
  assign n3204 = n2479 & ~n3117 ;
  assign n3205 = n3204 ^ n2474 ;
  assign n3206 = n2487 & ~n3117 ;
  assign n3207 = n3206 ^ n2482 ;
  assign n3208 = n2042 & ~n3117 ;
  assign n3209 = n3208 ^ n2041 ;
  assign n3210 = n2037 & ~n3117 ;
  assign n3211 = n3210 ^ n2036 ;
  assign n3212 = n2032 & ~n3117 ;
  assign n3213 = n3212 ^ n2031 ;
  assign n3214 = n2504 & ~n3117 ;
  assign n3215 = n3214 ^ n2499 ;
  assign n3216 = n2027 & ~n3117 ;
  assign n3217 = n3216 ^ n2026 ;
  assign n3218 = n2516 & ~n3117 ;
  assign n3219 = n3218 ^ n2511 ;
  assign n3220 = n2525 & ~n3117 ;
  assign n3221 = n3220 ^ n2520 ;
  assign n3222 = n2021 & ~n3117 ;
  assign n3223 = n3222 ^ n2020 ;
  assign n3224 = n2539 & ~n3117 ;
  assign n3225 = n3224 ^ n2532 ;
  assign n3226 = n2014 & ~n3117 ;
  assign n3227 = n3226 ^ n2013 ;
  assign n3228 = n2553 & ~n3117 ;
  assign n3229 = n3228 ^ n2546 ;
  assign n3230 = n2007 & ~n3117 ;
  assign n3231 = n3230 ^ n2006 ;
  assign n3232 = n2567 & ~n3117 ;
  assign n3233 = n3232 ^ n2560 ;
  assign n3234 = n2575 & ~n3117 ;
  assign n3235 = n3234 ^ n2570 ;
  assign n3236 = n2583 & ~n3117 ;
  assign n3237 = n3236 ^ n2578 ;
  assign n3238 = n2000 & ~n3117 ;
  assign n3239 = n3238 ^ n1999 ;
  assign n3240 = n2594 & ~n3117 ;
  assign n3241 = n3240 ^ n2589 ;
  assign n3242 = n1995 & ~n3117 ;
  assign n3243 = n3242 ^ n1994 ;
  assign n3244 = n1990 & ~n3117 ;
  assign n3245 = n3244 ^ n1989 ;
  assign n3246 = n1985 & ~n3117 ;
  assign n3247 = n3246 ^ n1984 ;
  assign n3248 = n1979 & ~n3117 ;
  assign n3249 = n3248 ^ n1978 ;
  assign n3250 = n1972 & ~n3117 ;
  assign n3251 = n3250 ^ n1971 ;
  assign n3252 = n1966 & ~n3117 ;
  assign n3253 = n3252 ^ n1965 ;
  assign n3254 = n2620 & ~n3117 ;
  assign n3255 = n3254 ^ n2615 ;
  assign n3256 = n1961 & ~n3117 ;
  assign n3257 = n3256 ^ n1960 ;
  assign n3258 = n1956 & ~n3117 ;
  assign n3259 = n3258 ^ n1955 ;
  assign n3260 = n1951 & ~n3117 ;
  assign n3261 = n3260 ^ n1950 ;
  assign n3262 = n1946 & ~n3117 ;
  assign n3263 = n3262 ^ n1945 ;
  assign n3264 = n2642 & ~n3117 ;
  assign n3265 = n3264 ^ n2635 ;
  assign n3266 = n2652 & ~n3117 ;
  assign n3267 = n3266 ^ n2645 ;
  assign n3268 = n2663 & n3117 ;
  assign n3269 = n3268 ^ n2656 ;
  assign n3270 = n2673 & ~n3117 ;
  assign n3271 = n3270 ^ n2666 ;
  assign n3272 = n2683 & ~n3117 ;
  assign n3273 = n3272 ^ n2676 ;
  assign n3274 = n2693 & ~n3117 ;
  assign n3275 = n3274 ^ n2686 ;
  assign n3276 = n2703 & ~n3117 ;
  assign n3277 = n3276 ^ n2696 ;
  assign n3278 = n1940 & ~n3117 ;
  assign n3279 = n3278 ^ n1939 ;
  assign n3280 = n1934 & ~n3117 ;
  assign n3281 = n3280 ^ n1933 ;
  assign n3282 = n2720 & n3117 ;
  assign n3283 = n3282 ^ n2713 ;
  assign n3284 = n2731 & ~n3117 ;
  assign n3285 = n3284 ^ n2724 ;
  assign n3286 = n2742 & ~n3117 ;
  assign n3287 = n3286 ^ n2735 ;
  assign n3288 = n2753 & ~n3117 ;
  assign n3289 = n3288 ^ n2746 ;
  assign n3290 = n2764 & ~n3117 ;
  assign n3291 = n3290 ^ n2757 ;
  assign n3292 = n2775 & ~n3117 ;
  assign n3293 = n3292 ^ n2768 ;
  assign n3294 = n2786 & n3117 ;
  assign n3295 = n3294 ^ n2779 ;
  assign n3296 = n2797 & n3117 ;
  assign n3297 = n3296 ^ n2790 ;
  assign n3298 = n2808 & n3117 ;
  assign n3299 = n3298 ^ n2801 ;
  assign n3300 = n2819 & ~n3117 ;
  assign n3301 = n3300 ^ n2812 ;
  assign n3302 = n2830 & ~n3117 ;
  assign n3303 = n3302 ^ n2823 ;
  assign n3304 = n2841 & ~n3117 ;
  assign n3305 = n3304 ^ n2834 ;
  assign n3306 = n2852 & n3117 ;
  assign n3307 = n3306 ^ n2845 ;
  assign n3308 = n2863 & n3117 ;
  assign n3309 = n3308 ^ n2856 ;
  assign n3310 = n1927 & ~n3117 ;
  assign n3311 = n3310 ^ n1926 ;
  assign n3312 = n1920 & ~n3117 ;
  assign n3313 = n3312 ^ n1919 ;
  assign n3314 = n2880 & n3117 ;
  assign n3315 = n3314 ^ n2873 ;
  assign n3316 = n2891 & n3117 ;
  assign n3317 = n3316 ^ n2884 ;
  assign n3318 = n1913 & ~n3117 ;
  assign n3319 = n3318 ^ n1912 ;
  assign n3320 = n1906 & ~n3117 ;
  assign n3321 = n3320 ^ n1905 ;
  assign n3322 = n2908 & n3117 ;
  assign n3323 = n3322 ^ n2901 ;
  assign n3324 = n2919 & ~n3117 ;
  assign n3325 = n3324 ^ n2912 ;
  assign n3326 = n1899 & ~n3117 ;
  assign n3327 = n3326 ^ n1898 ;
  assign n3328 = n2933 & n3117 ;
  assign n3329 = n3328 ^ n2926 ;
  assign n3330 = n2944 & ~n3117 ;
  assign n3331 = n3330 ^ n2937 ;
  assign n3332 = n2955 & ~n3117 ;
  assign n3333 = n3332 ^ n2948 ;
  assign n3334 = n1892 & ~n3117 ;
  assign n3335 = n3334 ^ n1891 ;
  assign n3336 = n1885 & ~n3117 ;
  assign n3337 = n3336 ^ n1884 ;
  assign n3338 = n1878 & ~n3117 ;
  assign n3339 = n3338 ^ n1877 ;
  assign n3340 = n2975 & n3117 ;
  assign n3341 = n3340 ^ n2968 ;
  assign n3342 = n2986 & n3117 ;
  assign n3343 = n3342 ^ n2979 ;
  assign n3344 = n2997 & ~n3117 ;
  assign n3345 = n3344 ^ n2990 ;
  assign n3346 = n3008 & n3117 ;
  assign n3347 = n3346 ^ n3001 ;
  assign n3348 = n3019 & n3117 ;
  assign n3349 = n3348 ^ n3012 ;
  assign n3350 = n3030 & ~n3117 ;
  assign n3351 = n3350 ^ n3023 ;
  assign n3352 = n3041 & ~n3117 ;
  assign n3353 = n3352 ^ n3034 ;
  assign n3354 = n3052 & ~n3117 ;
  assign n3355 = n3354 ^ n3045 ;
  assign n3356 = n3063 & ~n3117 ;
  assign n3357 = n3356 ^ n3056 ;
  assign n3358 = n1871 & ~n3117 ;
  assign n3359 = n3358 ^ n1870 ;
  assign n3360 = n1864 & ~n3117 ;
  assign n3361 = n3360 ^ n1863 ;
  assign n3362 = n3077 & ~n3117 ;
  assign n3363 = n3362 ^ n3072 ;
  assign n3364 = n3087 & n3117 ;
  assign n3365 = n3364 ^ n3080 ;
  assign n3366 = n3097 & n3117 ;
  assign n3367 = n3366 ^ n3090 ;
  assign n3368 = n3107 & ~n3117 ;
  assign n3369 = n3368 ^ n3100 ;
  assign n3370 = n3113 & ~n3117 ;
  assign n3371 = n3370 ^ n1856 ;
  assign n3372 = n1852 & n1853 ;
  assign n3373 = n1848 ^ n1180 ;
  assign n3374 = n3117 & n3373 ;
  assign n3375 = n3374 ^ n1848 ;
  assign y0 = n3119 ;
  assign y1 = n3121 ;
  assign y2 = n3123 ;
  assign y3 = n3125 ;
  assign y4 = n3127 ;
  assign y5 = n3129 ;
  assign y6 = n3131 ;
  assign y7 = n3133 ;
  assign y8 = n3135 ;
  assign y9 = n3137 ;
  assign y10 = n3139 ;
  assign y11 = n3141 ;
  assign y12 = n3143 ;
  assign y13 = n3145 ;
  assign y14 = n3147 ;
  assign y15 = n3149 ;
  assign y16 = n3151 ;
  assign y17 = n3153 ;
  assign y18 = n3155 ;
  assign y19 = n3157 ;
  assign y20 = n3159 ;
  assign y21 = n3161 ;
  assign y22 = n3163 ;
  assign y23 = n3165 ;
  assign y24 = n3167 ;
  assign y25 = n3169 ;
  assign y26 = n3171 ;
  assign y27 = n3173 ;
  assign y28 = n3175 ;
  assign y29 = n3177 ;
  assign y30 = n3179 ;
  assign y31 = n3181 ;
  assign y32 = n3183 ;
  assign y33 = n3185 ;
  assign y34 = n3187 ;
  assign y35 = n3189 ;
  assign y36 = n3191 ;
  assign y37 = n3193 ;
  assign y38 = n3195 ;
  assign y39 = n3197 ;
  assign y40 = n3199 ;
  assign y41 = n3201 ;
  assign y42 = n3203 ;
  assign y43 = n3205 ;
  assign y44 = n3207 ;
  assign y45 = n3209 ;
  assign y46 = n3211 ;
  assign y47 = n3213 ;
  assign y48 = n3215 ;
  assign y49 = n3217 ;
  assign y50 = n3219 ;
  assign y51 = n3221 ;
  assign y52 = n3223 ;
  assign y53 = n3225 ;
  assign y54 = n3227 ;
  assign y55 = n3229 ;
  assign y56 = n3231 ;
  assign y57 = n3233 ;
  assign y58 = n3235 ;
  assign y59 = n3237 ;
  assign y60 = n3239 ;
  assign y61 = n3241 ;
  assign y62 = n3243 ;
  assign y63 = n3245 ;
  assign y64 = n3247 ;
  assign y65 = n3249 ;
  assign y66 = n3251 ;
  assign y67 = n3253 ;
  assign y68 = n3255 ;
  assign y69 = n3257 ;
  assign y70 = n3259 ;
  assign y71 = n3261 ;
  assign y72 = n3263 ;
  assign y73 = n3265 ;
  assign y74 = n3267 ;
  assign y75 = n3269 ;
  assign y76 = n3271 ;
  assign y77 = n3273 ;
  assign y78 = n3275 ;
  assign y79 = n3277 ;
  assign y80 = n3279 ;
  assign y81 = n3281 ;
  assign y82 = n3283 ;
  assign y83 = n3285 ;
  assign y84 = n3287 ;
  assign y85 = n3289 ;
  assign y86 = n3291 ;
  assign y87 = n3293 ;
  assign y88 = n3295 ;
  assign y89 = n3297 ;
  assign y90 = n3299 ;
  assign y91 = n3301 ;
  assign y92 = n3303 ;
  assign y93 = n3305 ;
  assign y94 = n3307 ;
  assign y95 = n3309 ;
  assign y96 = n3311 ;
  assign y97 = n3313 ;
  assign y98 = n3315 ;
  assign y99 = n3317 ;
  assign y100 = n3319 ;
  assign y101 = n3321 ;
  assign y102 = n3323 ;
  assign y103 = n3325 ;
  assign y104 = n3327 ;
  assign y105 = n3329 ;
  assign y106 = n3331 ;
  assign y107 = n3333 ;
  assign y108 = n3335 ;
  assign y109 = n3337 ;
  assign y110 = n3339 ;
  assign y111 = n3341 ;
  assign y112 = n3343 ;
  assign y113 = n3345 ;
  assign y114 = n3347 ;
  assign y115 = n3349 ;
  assign y116 = n3351 ;
  assign y117 = n3353 ;
  assign y118 = n3355 ;
  assign y119 = n3357 ;
  assign y120 = n3359 ;
  assign y121 = n3361 ;
  assign y122 = n3363 ;
  assign y123 = n3365 ;
  assign y124 = n3367 ;
  assign y125 = n3369 ;
  assign y126 = n3371 ;
  assign y127 = n3372 ;
  assign y128 = n3375 ;
  assign y129 = ~n3117 ;
endmodule
