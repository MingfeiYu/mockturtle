module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, y0, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, y1, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, y2, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, y3, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152, y4, n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528, n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552, n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, y5, n_5612, n_5613, n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677, n_5678, n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705, n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713, n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743, n_5744, n_5745, n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772, n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789, n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907, n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, y6, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983, n_5984, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107, y7, n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208, n_6209, y8, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240, n_6241, n_6242, y9, n_6243, n_6244, n_6245, n_6246, y10, n_6247, n_6248, n_6249, n_6250, y11, n_6251, n_6252, n_6253, n_6254, y12, n_6255, n_6256, n_6257, n_6258, y13, n_6259, n_6260, n_6261, n_6262, y14, n_6263, n_6264, n_6265, n_6266, y15, n_6267, n_6268, n_6269, n_6270, y16, n_6271, n_6272, n_6273, n_6274, y17, n_6275, n_6276, n_6277, n_6278, y18, n_6279, n_6280, n_6281, n_6282, y19, n_6283, n_6284, n_6285, n_6286, y20, n_6287, n_6288, n_6289, n_6290, y21, n_6291, n_6292, n_6293, n_6294, y22, n_6295, n_6296, n_6297, n_6298, y23, n_6299, n_6300, n_6301, n_6302, y24, n_6303, n_6304, n_6305, n_6306, y25, n_6307, n_6308, n_6309, n_6310, y26, n_6311, n_6312, n_6313, n_6314, y27, n_6315, n_6316, n_6317, n_6318, y28, n_6319, n_6320, n_6321, n_6322, y29, n_6323, n_6324, n_6325, n_6326, y30, n_6327, n_6328, n_6329, n_6330, y31, n_6331, n_6332, n_6333, n_6334, y32, n_6335, n_6336, n_6337, n_6338, y33, n_6339, n_6340, n_6341, n_6342, y34, n_6343, n_6344, n_6345, n_6346, y35, n_6347, n_6348, n_6349, n_6350, y36, n_6351, n_6352, n_6353, n_6354, y37, n_6355, n_6356, n_6357, n_6358, y38, n_6359, n_6360, n_6361, n_6362, y39, n_6363, n_6364, n_6365, n_6366, y40, n_6367, n_6368, n_6369, n_6370, y41, n_6371, n_6372, n_6373, n_6374, y42, n_6375, n_6376, n_6377, n_6378, y43, n_6379, n_6380, n_6381, n_6382, y44, n_6383, n_6384, n_6385, n_6386, y45, n_6387, n_6388, n_6389, n_6390, y46, n_6391, n_6392, n_6393, n_6394, y47, n_6395, n_6396, n_6397, n_6398, y48, n_6399, n_6400, n_6401, n_6402, y49, n_6403, n_6404, n_6405, n_6406, y50, n_6407, n_6408, n_6409, n_6410, y51, n_6411, n_6412, n_6413, n_6414, y52, n_6415, n_6416, n_6417, n_6418, y53, n_6419, n_6420, n_6421, n_6422, y54, n_6423, n_6424, n_6425, n_6426, y55, n_6427, n_6428, n_6429, n_6430, y56, n_6431, n_6432, n_6433, n_6434, y57, n_6435, n_6436, n_6437, n_6438, y58, n_6439, n_6440, n_6441, n_6442, y59, n_6443, n_6444, n_6445, n_6446, y60, n_6447, n_6448, n_6449, n_6450, y61, n_6451, n_6452, n_6453, n_6454, y62, n_6455, n_6456, n_6457, y63;
assign n_0 = x0 & x32;
assign n_1 = x1 & x32;
assign n_2 = x2 & x32;
assign n_3 = x3 & x32;
assign n_4 = x4 & x32;
assign n_5 = x5 & x32;
assign n_6 = x6 & x32;
assign n_7 = x7 & x32;
assign n_8 = x8 & x32;
assign n_9 = x9 & x32;
assign n_10 = x10 & x32;
assign n_11 = x11 & x32;
assign n_12 = x12 & x32;
assign n_13 = x13 & x32;
assign n_14 = x14 & x32;
assign n_15 = x15 & x32;
assign n_16 = x16 & x32;
assign n_17 = x17 & x32;
assign n_18 = x18 & x32;
assign n_19 = x19 & x32;
assign n_20 = x20 & x32;
assign n_21 = x21 & x32;
assign n_22 = x22 & x32;
assign n_23 = x23 & x32;
assign n_24 = x24 & x32;
assign n_25 = x25 & x32;
assign n_26 = x26 & x32;
assign n_27 = x27 & x32;
assign n_28 = x28 & x32;
assign n_29 = x29 & x32;
assign n_30 = x30 & x32;
assign n_31 = x31 & x32;
assign n_32 = ~x32 & x33;
assign n_33 = x33 ^ x0;
assign n_34 = x34 ^ x33;
assign n_35 = x35 ^ x34;
assign n_36 = x35 ^ x0;
assign n_37 = x35 ^ x31;
assign n_38 = x36 ^ x35;
assign n_39 = x37 ^ x36;
assign n_40 = x37 ^ x0;
assign n_41 = x37 ^ x31;
assign n_42 = x38 ^ x37;
assign n_43 = x39 ^ x38;
assign n_44 = x39 ^ x0;
assign n_45 = x39 ^ x31;
assign n_46 = x40 ^ x39;
assign n_47 = x41 ^ x40;
assign n_48 = x41 ^ x0;
assign n_49 = x41 ^ x31;
assign n_50 = x42 ^ x41;
assign n_51 = x43 ^ x42;
assign n_52 = x43 ^ x0;
assign n_53 = x43 ^ x31;
assign n_54 = x44 ^ x43;
assign n_55 = x45 ^ x44;
assign n_56 = x45 ^ x0;
assign n_57 = x45 ^ x31;
assign n_58 = x46 ^ x45;
assign n_59 = x47 ^ x46;
assign n_60 = x47 ^ x0;
assign n_61 = x47 ^ x31;
assign n_62 = x48 ^ x47;
assign n_63 = x49 ^ x48;
assign n_64 = x49 ^ x0;
assign n_65 = x49 ^ x31;
assign n_66 = x50 ^ x49;
assign n_67 = x51 ^ x50;
assign n_68 = x51 ^ x0;
assign n_69 = x51 ^ x31;
assign n_70 = x52 ^ x51;
assign n_71 = x53 ^ x52;
assign n_72 = x53 ^ x0;
assign n_73 = x53 ^ x31;
assign n_74 = x54 ^ x53;
assign n_75 = x55 ^ x54;
assign n_76 = x55 ^ x0;
assign n_77 = x55 ^ x31;
assign n_78 = x56 ^ x55;
assign n_79 = x57 ^ x56;
assign n_80 = x57 ^ x0;
assign n_81 = x57 ^ x31;
assign n_82 = x58 ^ x57;
assign n_83 = x59 ^ x58;
assign n_84 = x59 ^ x0;
assign n_85 = x59 ^ x31;
assign n_86 = x60 ^ x59;
assign n_87 = x61 ^ x60;
assign n_88 = x61 ^ x0;
assign n_89 = x61 ^ x31;
assign n_90 = x62 ^ x61;
assign n_91 = x63 ^ x62;
assign n_92 = x0 & x63;
assign n_93 = x1 & x63;
assign n_94 = x2 & x63;
assign n_95 = x3 & x63;
assign n_96 = x4 & x63;
assign n_97 = x5 & x63;
assign n_98 = x6 & x63;
assign n_99 = x7 & x63;
assign n_100 = x8 & x63;
assign n_101 = x9 & x63;
assign n_102 = x10 & x63;
assign n_103 = x11 & x63;
assign n_104 = x12 & x63;
assign n_105 = x13 & x63;
assign n_106 = x14 & x63;
assign n_107 = x15 & x63;
assign n_108 = x16 & x63;
assign n_109 = x17 & x63;
assign n_110 = x18 & x63;
assign n_111 = x19 & x63;
assign n_112 = x20 & x63;
assign n_113 = x21 & x63;
assign n_114 = x22 & x63;
assign n_115 = x23 & x63;
assign n_116 = x24 & x63;
assign n_117 = x25 & x63;
assign n_118 = x26 & x63;
assign n_119 = x27 & x63;
assign n_120 = x28 & x63;
assign n_121 = x63 ^ x31;
assign n_122 = x29 & x63;
assign n_123 = x30 & x63;
assign n_124 = x33 & ~n_0;
assign y0 = n_0;
assign n_125 = n_32 ^ x33;
assign n_126 = ~x0 & n_32;
assign n_127 = ~x1 & n_32;
assign n_128 = ~x2 & n_32;
assign n_129 = ~x3 & n_32;
assign n_130 = ~x4 & n_32;
assign n_131 = ~x5 & n_32;
assign n_132 = ~x6 & n_32;
assign n_133 = ~x7 & n_32;
assign n_134 = ~x8 & n_32;
assign n_135 = ~x9 & n_32;
assign n_136 = ~x10 & n_32;
assign n_137 = ~x11 & n_32;
assign n_138 = ~x12 & n_32;
assign n_139 = ~x13 & n_32;
assign n_140 = ~x14 & n_32;
assign n_141 = ~x15 & n_32;
assign n_142 = ~x16 & n_32;
assign n_143 = ~x17 & n_32;
assign n_144 = ~x18 & n_32;
assign n_145 = ~x19 & n_32;
assign n_146 = ~x20 & n_32;
assign n_147 = ~x21 & n_32;
assign n_148 = ~x22 & n_32;
assign n_149 = ~x23 & n_32;
assign n_150 = ~x24 & n_32;
assign n_151 = ~x25 & n_32;
assign n_152 = ~x26 & n_32;
assign n_153 = ~x27 & n_32;
assign n_154 = ~x28 & n_32;
assign n_155 = ~x29 & n_32;
assign n_156 = ~x30 & n_32;
assign n_157 = x31 & n_32;
assign n_158 = x0 & n_34;
assign n_159 = ~n_34 & n_33;
assign n_160 = x35 & n_34;
assign n_161 = ~n_34 & n_35;
assign n_162 = n_34 & n_37;
assign n_163 = x0 & n_38;
assign n_164 = x37 & n_38;
assign n_165 = n_36 & ~n_38;
assign n_166 = ~n_38 & n_39;
assign n_167 = n_38 & n_41;
assign n_168 = x0 & n_42;
assign n_169 = n_40 & ~n_42;
assign n_170 = x39 & n_42;
assign n_171 = ~n_42 & n_43;
assign n_172 = n_42 & n_45;
assign n_173 = x0 & n_46;
assign n_174 = x41 & n_46;
assign n_175 = n_44 & ~n_46;
assign n_176 = ~n_46 & n_47;
assign n_177 = n_46 & n_49;
assign n_178 = x0 & n_50;
assign n_179 = ~x43 & n_50;
assign n_180 = n_48 & ~n_50;
assign n_181 = ~n_50 & n_51;
assign n_182 = n_50 & n_53;
assign n_183 = x0 & n_54;
assign n_184 = n_52 & ~n_54;
assign n_185 = x45 & n_54;
assign n_186 = ~n_54 & n_55;
assign n_187 = n_54 & n_57;
assign n_188 = x0 & n_58;
assign n_189 = ~x47 & n_58;
assign n_190 = n_56 & ~n_58;
assign n_191 = ~n_58 & n_59;
assign n_192 = n_58 & n_61;
assign n_193 = x0 & n_62;
assign n_194 = x49 & n_62;
assign n_195 = n_60 & ~n_62;
assign n_196 = ~n_62 & n_63;
assign n_197 = n_62 & n_65;
assign n_198 = x0 & n_66;
assign n_199 = ~x51 & n_66;
assign n_200 = n_64 & ~n_66;
assign n_201 = ~n_66 & n_67;
assign n_202 = n_66 & n_69;
assign n_203 = x0 & n_70;
assign n_204 = n_68 & ~n_70;
assign n_205 = x53 & n_70;
assign n_206 = ~n_70 & n_71;
assign n_207 = n_70 & n_73;
assign n_208 = x0 & n_74;
assign n_209 = n_72 & ~n_74;
assign n_210 = x55 & n_74;
assign n_211 = ~n_74 & n_75;
assign n_212 = n_74 & n_77;
assign n_213 = x0 & n_78;
assign n_214 = n_76 & ~n_78;
assign n_215 = x57 & n_78;
assign n_216 = ~n_78 & n_79;
assign n_217 = n_78 & n_81;
assign n_218 = x0 & n_82;
assign n_219 = ~x59 & n_82;
assign n_220 = n_80 & ~n_82;
assign n_221 = ~n_82 & n_83;
assign n_222 = n_82 & n_85;
assign n_223 = x0 & n_86;
assign n_224 = x61 & n_86;
assign n_225 = n_84 & ~n_86;
assign n_226 = ~n_86 & n_87;
assign n_227 = n_86 & n_89;
assign n_228 = x0 & n_90;
assign n_229 = x63 & n_90;
assign n_230 = n_88 & ~n_90;
assign n_231 = ~n_90 & n_91;
assign n_232 = n_90 & n_121;
assign n_233 = n_125 ^ n_126;
assign n_234 = n_127 ^ n_125;
assign n_235 = n_128 ^ n_125;
assign n_236 = n_129 ^ n_125;
assign n_237 = n_130 ^ n_125;
assign n_238 = n_131 ^ n_125;
assign n_239 = n_132 ^ n_125;
assign n_240 = n_133 ^ n_125;
assign n_241 = n_134 ^ n_125;
assign n_242 = n_135 ^ n_125;
assign n_243 = n_136 ^ n_125;
assign n_244 = n_137 ^ n_125;
assign n_245 = n_138 ^ n_125;
assign n_246 = n_139 ^ n_125;
assign n_247 = n_140 ^ n_125;
assign n_248 = n_141 ^ n_125;
assign n_249 = n_142 ^ n_125;
assign n_250 = n_143 ^ n_125;
assign n_251 = n_144 ^ n_125;
assign n_252 = n_145 ^ n_125;
assign n_253 = n_146 ^ n_125;
assign n_254 = n_147 ^ n_125;
assign n_255 = n_148 ^ n_125;
assign n_256 = n_149 ^ n_125;
assign n_257 = n_150 ^ n_125;
assign n_258 = n_151 ^ n_125;
assign n_259 = n_152 ^ n_125;
assign n_260 = n_153 ^ n_125;
assign n_261 = n_154 ^ n_125;
assign n_262 = n_155 ^ n_125;
assign n_263 = n_156 ^ n_125;
assign n_264 = n_157 ^ x33;
assign n_265 = n_159 ^ x0;
assign n_266 = ~x1 & ~n_160;
assign n_267 = n_160 ^ n_34;
assign n_268 = ~x2 & ~n_160;
assign n_269 = ~x3 & ~n_160;
assign n_270 = ~x4 & ~n_160;
assign n_271 = ~x5 & ~n_160;
assign n_272 = ~x6 & ~n_160;
assign n_273 = ~x7 & ~n_160;
assign n_274 = ~x8 & ~n_160;
assign n_275 = ~x9 & ~n_160;
assign n_276 = ~x10 & ~n_160;
assign n_277 = ~x11 & ~n_160;
assign n_278 = ~x12 & ~n_160;
assign n_279 = ~x13 & ~n_160;
assign n_280 = ~x14 & ~n_160;
assign n_281 = ~x15 & ~n_160;
assign n_282 = ~x16 & ~n_160;
assign n_283 = ~x17 & ~n_160;
assign n_284 = ~x18 & ~n_160;
assign n_285 = ~x19 & ~n_160;
assign n_286 = ~x20 & ~n_160;
assign n_287 = ~x21 & ~n_160;
assign n_288 = ~x22 & ~n_160;
assign n_289 = ~x23 & ~n_160;
assign n_290 = ~x24 & ~n_160;
assign n_291 = ~x25 & ~n_160;
assign n_292 = ~x26 & ~n_160;
assign n_293 = ~x27 & ~n_160;
assign n_294 = ~x28 & ~n_160;
assign n_295 = ~x29 & ~n_160;
assign n_296 = ~x30 & ~n_160;
assign n_297 = n_161 & n_36;
assign n_298 = x35 & n_161;
assign n_299 = n_161 & n_37;
assign n_300 = ~x1 & ~n_164;
assign n_301 = n_164 ^ n_38;
assign n_302 = ~x2 & ~n_164;
assign n_303 = ~x3 & ~n_164;
assign n_304 = ~x4 & ~n_164;
assign n_305 = ~x5 & ~n_164;
assign n_306 = ~x6 & ~n_164;
assign n_307 = ~x7 & ~n_164;
assign n_308 = ~x8 & ~n_164;
assign n_309 = ~x9 & ~n_164;
assign n_310 = ~x10 & ~n_164;
assign n_311 = ~x11 & ~n_164;
assign n_312 = ~x12 & ~n_164;
assign n_313 = ~x13 & ~n_164;
assign n_314 = ~x14 & ~n_164;
assign n_315 = ~x15 & ~n_164;
assign n_316 = ~x16 & ~n_164;
assign n_317 = ~x17 & ~n_164;
assign n_318 = ~x18 & ~n_164;
assign n_319 = ~x19 & ~n_164;
assign n_320 = ~x20 & ~n_164;
assign n_321 = ~x21 & ~n_164;
assign n_322 = ~x22 & ~n_164;
assign n_323 = ~x23 & ~n_164;
assign n_324 = ~x24 & ~n_164;
assign n_325 = ~x25 & ~n_164;
assign n_326 = ~x26 & ~n_164;
assign n_327 = ~x27 & ~n_164;
assign n_328 = ~x28 & ~n_164;
assign n_329 = ~x29 & ~n_164;
assign n_330 = ~x30 & ~n_164;
assign n_331 = n_165 ^ x0;
assign n_332 = n_166 & n_40;
assign n_333 = x37 & n_166;
assign n_334 = n_166 & n_41;
assign n_335 = n_169 ^ x0;
assign n_336 = ~x1 & ~n_170;
assign n_337 = n_170 ^ n_42;
assign n_338 = ~x2 & ~n_170;
assign n_339 = ~x3 & ~n_170;
assign n_340 = ~x4 & ~n_170;
assign n_341 = ~x5 & ~n_170;
assign n_342 = ~x6 & ~n_170;
assign n_343 = ~x7 & ~n_170;
assign n_344 = ~x8 & ~n_170;
assign n_345 = ~x9 & ~n_170;
assign n_346 = ~x10 & ~n_170;
assign n_347 = ~x11 & ~n_170;
assign n_348 = ~x12 & ~n_170;
assign n_349 = ~x13 & ~n_170;
assign n_350 = ~x14 & ~n_170;
assign n_351 = ~x15 & ~n_170;
assign n_352 = ~x16 & ~n_170;
assign n_353 = ~x17 & ~n_170;
assign n_354 = ~x18 & ~n_170;
assign n_355 = ~x19 & ~n_170;
assign n_356 = ~x20 & ~n_170;
assign n_357 = ~x21 & ~n_170;
assign n_358 = ~x22 & ~n_170;
assign n_359 = ~x23 & ~n_170;
assign n_360 = ~x24 & ~n_170;
assign n_361 = ~x25 & ~n_170;
assign n_362 = ~x26 & ~n_170;
assign n_363 = ~x27 & ~n_170;
assign n_364 = ~x28 & ~n_170;
assign n_365 = ~x29 & ~n_170;
assign n_366 = ~x30 & ~n_170;
assign n_367 = n_171 & n_44;
assign n_368 = x39 & n_171;
assign n_369 = n_171 & n_45;
assign n_370 = ~x1 & ~n_174;
assign n_371 = n_174 ^ n_46;
assign n_372 = ~x2 & ~n_174;
assign n_373 = ~x3 & ~n_174;
assign n_374 = ~x4 & ~n_174;
assign n_375 = ~x5 & ~n_174;
assign n_376 = ~x6 & ~n_174;
assign n_377 = ~x7 & ~n_174;
assign n_378 = ~x8 & ~n_174;
assign n_379 = ~x9 & ~n_174;
assign n_380 = ~x10 & ~n_174;
assign n_381 = ~x11 & ~n_174;
assign n_382 = ~x12 & ~n_174;
assign n_383 = ~x13 & ~n_174;
assign n_384 = ~x14 & ~n_174;
assign n_385 = ~x15 & ~n_174;
assign n_386 = ~x16 & ~n_174;
assign n_387 = ~x17 & ~n_174;
assign n_388 = ~x18 & ~n_174;
assign n_389 = ~x19 & ~n_174;
assign n_390 = ~x20 & ~n_174;
assign n_391 = ~x21 & ~n_174;
assign n_392 = ~x22 & ~n_174;
assign n_393 = ~x23 & ~n_174;
assign n_394 = ~x24 & ~n_174;
assign n_395 = ~x25 & ~n_174;
assign n_396 = ~x26 & ~n_174;
assign n_397 = ~x27 & ~n_174;
assign n_398 = ~x28 & ~n_174;
assign n_399 = ~x29 & ~n_174;
assign n_400 = ~x30 & ~n_174;
assign n_401 = n_175 ^ x0;
assign n_402 = n_176 & n_48;
assign n_403 = x41 & n_176;
assign n_404 = n_176 & n_49;
assign n_405 = x1 & ~n_179;
assign n_406 = n_179 ^ n_50;
assign n_407 = x2 & ~n_179;
assign n_408 = x3 & ~n_179;
assign n_409 = x4 & ~n_179;
assign n_410 = x5 & ~n_179;
assign n_411 = x6 & ~n_179;
assign n_412 = x7 & ~n_179;
assign n_413 = x8 & ~n_179;
assign n_414 = x9 & ~n_179;
assign n_415 = x10 & ~n_179;
assign n_416 = x11 & ~n_179;
assign n_417 = x12 & ~n_179;
assign n_418 = x13 & ~n_179;
assign n_419 = x14 & ~n_179;
assign n_420 = x15 & ~n_179;
assign n_421 = x16 & ~n_179;
assign n_422 = x17 & ~n_179;
assign n_423 = x18 & ~n_179;
assign n_424 = x19 & ~n_179;
assign n_425 = x20 & ~n_179;
assign n_426 = x21 & ~n_179;
assign n_427 = x22 & ~n_179;
assign n_428 = x23 & ~n_179;
assign n_429 = x24 & ~n_179;
assign n_430 = x25 & ~n_179;
assign n_431 = x26 & ~n_179;
assign n_432 = x27 & ~n_179;
assign n_433 = x28 & ~n_179;
assign n_434 = x29 & ~n_179;
assign n_435 = x30 & ~n_179;
assign n_436 = n_180 ^ x0;
assign n_437 = n_181 & n_52;
assign n_438 = ~x43 & n_181;
assign n_439 = n_181 & n_53;
assign n_440 = n_184 ^ x0;
assign n_441 = ~x1 & ~n_185;
assign n_442 = n_185 ^ n_54;
assign n_443 = ~x2 & ~n_185;
assign n_444 = ~x3 & ~n_185;
assign n_445 = ~x4 & ~n_185;
assign n_446 = ~x5 & ~n_185;
assign n_447 = ~x6 & ~n_185;
assign n_448 = ~x7 & ~n_185;
assign n_449 = ~x8 & ~n_185;
assign n_450 = ~x9 & ~n_185;
assign n_451 = ~x10 & ~n_185;
assign n_452 = ~x11 & ~n_185;
assign n_453 = ~x12 & ~n_185;
assign n_454 = ~x13 & ~n_185;
assign n_455 = ~x14 & ~n_185;
assign n_456 = ~x15 & ~n_185;
assign n_457 = ~x16 & ~n_185;
assign n_458 = ~x17 & ~n_185;
assign n_459 = ~x18 & ~n_185;
assign n_460 = ~x19 & ~n_185;
assign n_461 = ~x20 & ~n_185;
assign n_462 = ~x21 & ~n_185;
assign n_463 = ~x22 & ~n_185;
assign n_464 = ~x23 & ~n_185;
assign n_465 = ~x24 & ~n_185;
assign n_466 = ~x25 & ~n_185;
assign n_467 = ~x26 & ~n_185;
assign n_468 = ~x27 & ~n_185;
assign n_469 = ~x28 & ~n_185;
assign n_470 = ~x29 & ~n_185;
assign n_471 = ~x30 & ~n_185;
assign n_472 = n_186 & n_56;
assign n_473 = x45 & n_186;
assign n_474 = n_186 & n_57;
assign n_475 = x1 & ~n_189;
assign n_476 = n_189 ^ n_58;
assign n_477 = x2 & ~n_189;
assign n_478 = x3 & ~n_189;
assign n_479 = x4 & ~n_189;
assign n_480 = x5 & ~n_189;
assign n_481 = x6 & ~n_189;
assign n_482 = x7 & ~n_189;
assign n_483 = x8 & ~n_189;
assign n_484 = x9 & ~n_189;
assign n_485 = x10 & ~n_189;
assign n_486 = x11 & ~n_189;
assign n_487 = x12 & ~n_189;
assign n_488 = x13 & ~n_189;
assign n_489 = x14 & ~n_189;
assign n_490 = x15 & ~n_189;
assign n_491 = x16 & ~n_189;
assign n_492 = x17 & ~n_189;
assign n_493 = x18 & ~n_189;
assign n_494 = x19 & ~n_189;
assign n_495 = x20 & ~n_189;
assign n_496 = x21 & ~n_189;
assign n_497 = x22 & ~n_189;
assign n_498 = x23 & ~n_189;
assign n_499 = x24 & ~n_189;
assign n_500 = x25 & ~n_189;
assign n_501 = x26 & ~n_189;
assign n_502 = x27 & ~n_189;
assign n_503 = x28 & ~n_189;
assign n_504 = x29 & ~n_189;
assign n_505 = x30 & ~n_189;
assign n_506 = n_190 ^ x0;
assign n_507 = n_191 & n_60;
assign n_508 = ~x47 & n_191;
assign n_509 = n_191 & n_61;
assign n_510 = ~x1 & ~n_194;
assign n_511 = n_194 ^ n_62;
assign n_512 = ~x2 & ~n_194;
assign n_513 = ~x3 & ~n_194;
assign n_514 = ~x4 & ~n_194;
assign n_515 = ~x5 & ~n_194;
assign n_516 = ~x6 & ~n_194;
assign n_517 = ~x7 & ~n_194;
assign n_518 = ~x8 & ~n_194;
assign n_519 = ~x9 & ~n_194;
assign n_520 = ~x10 & ~n_194;
assign n_521 = ~x11 & ~n_194;
assign n_522 = ~x12 & ~n_194;
assign n_523 = ~x13 & ~n_194;
assign n_524 = ~x14 & ~n_194;
assign n_525 = ~x15 & ~n_194;
assign n_526 = ~x16 & ~n_194;
assign n_527 = ~x17 & ~n_194;
assign n_528 = ~x18 & ~n_194;
assign n_529 = ~x19 & ~n_194;
assign n_530 = ~x20 & ~n_194;
assign n_531 = ~x21 & ~n_194;
assign n_532 = ~x22 & ~n_194;
assign n_533 = ~x23 & ~n_194;
assign n_534 = ~x24 & ~n_194;
assign n_535 = ~x25 & ~n_194;
assign n_536 = ~x26 & ~n_194;
assign n_537 = ~x27 & ~n_194;
assign n_538 = ~x28 & ~n_194;
assign n_539 = ~x29 & ~n_194;
assign n_540 = ~x30 & ~n_194;
assign n_541 = n_195 ^ x0;
assign n_542 = n_196 & n_64;
assign n_543 = x49 & n_196;
assign n_544 = n_196 & n_65;
assign n_545 = x1 & ~n_199;
assign n_546 = n_199 ^ n_66;
assign n_547 = x2 & ~n_199;
assign n_548 = x3 & ~n_199;
assign n_549 = x4 & ~n_199;
assign n_550 = x5 & ~n_199;
assign n_551 = x6 & ~n_199;
assign n_552 = x7 & ~n_199;
assign n_553 = x8 & ~n_199;
assign n_554 = x9 & ~n_199;
assign n_555 = x10 & ~n_199;
assign n_556 = x11 & ~n_199;
assign n_557 = x12 & ~n_199;
assign n_558 = x13 & ~n_199;
assign n_559 = x14 & ~n_199;
assign n_560 = x15 & ~n_199;
assign n_561 = x16 & ~n_199;
assign n_562 = x17 & ~n_199;
assign n_563 = x18 & ~n_199;
assign n_564 = x19 & ~n_199;
assign n_565 = x20 & ~n_199;
assign n_566 = x21 & ~n_199;
assign n_567 = x22 & ~n_199;
assign n_568 = x23 & ~n_199;
assign n_569 = x24 & ~n_199;
assign n_570 = x25 & ~n_199;
assign n_571 = x26 & ~n_199;
assign n_572 = x27 & ~n_199;
assign n_573 = x28 & ~n_199;
assign n_574 = x29 & ~n_199;
assign n_575 = x30 & ~n_199;
assign n_576 = n_200 ^ x0;
assign n_577 = n_201 & n_68;
assign n_578 = ~x51 & n_201;
assign n_579 = n_201 & n_69;
assign n_580 = n_204 ^ x0;
assign n_581 = ~x1 & ~n_205;
assign n_582 = n_205 ^ n_70;
assign n_583 = ~x2 & ~n_205;
assign n_584 = ~x3 & ~n_205;
assign n_585 = ~x4 & ~n_205;
assign n_586 = ~x5 & ~n_205;
assign n_587 = ~x6 & ~n_205;
assign n_588 = ~x7 & ~n_205;
assign n_589 = ~x8 & ~n_205;
assign n_590 = ~x9 & ~n_205;
assign n_591 = ~x10 & ~n_205;
assign n_592 = ~x11 & ~n_205;
assign n_593 = ~x12 & ~n_205;
assign n_594 = ~x13 & ~n_205;
assign n_595 = ~x14 & ~n_205;
assign n_596 = ~x15 & ~n_205;
assign n_597 = ~x16 & ~n_205;
assign n_598 = ~x17 & ~n_205;
assign n_599 = ~x18 & ~n_205;
assign n_600 = ~x19 & ~n_205;
assign n_601 = ~x20 & ~n_205;
assign n_602 = ~x21 & ~n_205;
assign n_603 = ~x22 & ~n_205;
assign n_604 = ~x23 & ~n_205;
assign n_605 = ~x24 & ~n_205;
assign n_606 = ~x25 & ~n_205;
assign n_607 = ~x26 & ~n_205;
assign n_608 = ~x27 & ~n_205;
assign n_609 = ~x28 & ~n_205;
assign n_610 = ~x29 & ~n_205;
assign n_611 = ~x30 & ~n_205;
assign n_612 = n_206 & n_72;
assign n_613 = x53 & n_206;
assign n_614 = n_206 & n_73;
assign n_615 = n_209 ^ x0;
assign n_616 = ~x1 & ~n_210;
assign n_617 = n_210 ^ n_74;
assign n_618 = ~x2 & ~n_210;
assign n_619 = ~x3 & ~n_210;
assign n_620 = ~x4 & ~n_210;
assign n_621 = ~x5 & ~n_210;
assign n_622 = ~x6 & ~n_210;
assign n_623 = ~x7 & ~n_210;
assign n_624 = ~x8 & ~n_210;
assign n_625 = ~x9 & ~n_210;
assign n_626 = ~x10 & ~n_210;
assign n_627 = ~x11 & ~n_210;
assign n_628 = ~x12 & ~n_210;
assign n_629 = ~x13 & ~n_210;
assign n_630 = ~x14 & ~n_210;
assign n_631 = ~x15 & ~n_210;
assign n_632 = ~x16 & ~n_210;
assign n_633 = ~x17 & ~n_210;
assign n_634 = ~x18 & ~n_210;
assign n_635 = ~x19 & ~n_210;
assign n_636 = ~x20 & ~n_210;
assign n_637 = ~x21 & ~n_210;
assign n_638 = ~x22 & ~n_210;
assign n_639 = ~x23 & ~n_210;
assign n_640 = ~x24 & ~n_210;
assign n_641 = ~x25 & ~n_210;
assign n_642 = ~x26 & ~n_210;
assign n_643 = ~x27 & ~n_210;
assign n_644 = ~x28 & ~n_210;
assign n_645 = ~x29 & ~n_210;
assign n_646 = ~x30 & ~n_210;
assign n_647 = n_211 & n_76;
assign n_648 = x55 & n_211;
assign n_649 = n_211 & n_77;
assign n_650 = n_214 ^ x0;
assign n_651 = ~x1 & ~n_215;
assign n_652 = n_215 ^ n_78;
assign n_653 = ~x2 & ~n_215;
assign n_654 = ~x3 & ~n_215;
assign n_655 = ~x4 & ~n_215;
assign n_656 = ~x5 & ~n_215;
assign n_657 = ~x6 & ~n_215;
assign n_658 = ~x7 & ~n_215;
assign n_659 = ~x8 & ~n_215;
assign n_660 = ~x9 & ~n_215;
assign n_661 = ~x10 & ~n_215;
assign n_662 = ~x11 & ~n_215;
assign n_663 = ~x12 & ~n_215;
assign n_664 = ~x13 & ~n_215;
assign n_665 = ~x14 & ~n_215;
assign n_666 = ~x15 & ~n_215;
assign n_667 = ~x16 & ~n_215;
assign n_668 = ~x17 & ~n_215;
assign n_669 = ~x18 & ~n_215;
assign n_670 = ~x19 & ~n_215;
assign n_671 = ~x20 & ~n_215;
assign n_672 = ~x21 & ~n_215;
assign n_673 = ~x22 & ~n_215;
assign n_674 = ~x23 & ~n_215;
assign n_675 = ~x24 & ~n_215;
assign n_676 = ~x25 & ~n_215;
assign n_677 = ~x26 & ~n_215;
assign n_678 = ~x27 & ~n_215;
assign n_679 = ~x28 & ~n_215;
assign n_680 = ~x29 & ~n_215;
assign n_681 = ~x30 & ~n_215;
assign n_682 = n_216 & n_80;
assign n_683 = x57 & n_216;
assign n_684 = n_216 & n_81;
assign n_685 = x1 & ~n_219;
assign n_686 = n_219 ^ n_82;
assign n_687 = x2 & ~n_219;
assign n_688 = x3 & ~n_219;
assign n_689 = x4 & ~n_219;
assign n_690 = x5 & ~n_219;
assign n_691 = x6 & ~n_219;
assign n_692 = x7 & ~n_219;
assign n_693 = x8 & ~n_219;
assign n_694 = x9 & ~n_219;
assign n_695 = x10 & ~n_219;
assign n_696 = x11 & ~n_219;
assign n_697 = x12 & ~n_219;
assign n_698 = x13 & ~n_219;
assign n_699 = x14 & ~n_219;
assign n_700 = x15 & ~n_219;
assign n_701 = x16 & ~n_219;
assign n_702 = x17 & ~n_219;
assign n_703 = x18 & ~n_219;
assign n_704 = x19 & ~n_219;
assign n_705 = x20 & ~n_219;
assign n_706 = x21 & ~n_219;
assign n_707 = x22 & ~n_219;
assign n_708 = x23 & ~n_219;
assign n_709 = x24 & ~n_219;
assign n_710 = x25 & ~n_219;
assign n_711 = x26 & ~n_219;
assign n_712 = x27 & ~n_219;
assign n_713 = x28 & ~n_219;
assign n_714 = x29 & ~n_219;
assign n_715 = x30 & ~n_219;
assign n_716 = n_220 ^ x0;
assign n_717 = n_221 & n_84;
assign n_718 = ~x59 & n_221;
assign n_719 = n_221 & n_85;
assign n_720 = ~x1 & ~n_224;
assign n_721 = n_224 ^ n_86;
assign n_722 = ~x2 & ~n_224;
assign n_723 = ~x3 & ~n_224;
assign n_724 = ~x4 & ~n_224;
assign n_725 = ~x5 & ~n_224;
assign n_726 = ~x6 & ~n_224;
assign n_727 = ~x7 & ~n_224;
assign n_728 = ~x8 & ~n_224;
assign n_729 = ~x9 & ~n_224;
assign n_730 = ~x10 & ~n_224;
assign n_731 = ~x11 & ~n_224;
assign n_732 = ~x12 & ~n_224;
assign n_733 = ~x13 & ~n_224;
assign n_734 = ~x14 & ~n_224;
assign n_735 = ~x15 & ~n_224;
assign n_736 = ~x16 & ~n_224;
assign n_737 = ~x17 & ~n_224;
assign n_738 = ~x18 & ~n_224;
assign n_739 = ~x19 & ~n_224;
assign n_740 = ~x20 & ~n_224;
assign n_741 = ~x21 & ~n_224;
assign n_742 = ~x22 & ~n_224;
assign n_743 = ~x23 & ~n_224;
assign n_744 = ~x24 & ~n_224;
assign n_745 = ~x25 & ~n_224;
assign n_746 = ~x26 & ~n_224;
assign n_747 = ~x27 & ~n_224;
assign n_748 = ~x28 & ~n_224;
assign n_749 = ~x29 & ~n_224;
assign n_750 = ~x30 & ~n_224;
assign n_751 = n_225 ^ x0;
assign n_752 = n_226 & n_88;
assign n_753 = x61 & n_226;
assign n_754 = n_226 & n_89;
assign n_755 = ~x1 & ~n_229;
assign n_756 = n_229 ^ n_90;
assign n_757 = ~x2 & ~n_229;
assign n_758 = ~x3 & ~n_229;
assign n_759 = ~x4 & ~n_229;
assign n_760 = ~x5 & ~n_229;
assign n_761 = ~x6 & ~n_229;
assign n_762 = ~x7 & ~n_229;
assign n_763 = ~x8 & ~n_229;
assign n_764 = ~x9 & ~n_229;
assign n_765 = ~x10 & ~n_229;
assign n_766 = ~x11 & ~n_229;
assign n_767 = ~x12 & ~n_229;
assign n_768 = ~x13 & ~n_229;
assign n_769 = ~x14 & ~n_229;
assign n_770 = ~x15 & ~n_229;
assign n_771 = ~x16 & ~n_229;
assign n_772 = ~x17 & ~n_229;
assign n_773 = ~x18 & ~n_229;
assign n_774 = ~x19 & ~n_229;
assign n_775 = ~x20 & ~n_229;
assign n_776 = ~x21 & ~n_229;
assign n_777 = ~x22 & ~n_229;
assign n_778 = ~x23 & ~n_229;
assign n_779 = ~x24 & ~n_229;
assign n_780 = ~x25 & ~n_229;
assign n_781 = ~x26 & ~n_229;
assign n_782 = ~x27 & ~n_229;
assign n_783 = ~x28 & ~n_229;
assign n_784 = ~x29 & ~n_229;
assign n_785 = ~x30 & ~n_229;
assign n_786 = n_230 ^ x0;
assign n_787 = x63 & n_231;
assign n_788 = n_231 & n_121;
assign n_789 = n_231 ^ n_90;
assign n_790 = n_1 ^ n_233;
assign n_791 = n_2 ^ n_234;
assign n_792 = n_3 ^ n_235;
assign n_793 = n_4 ^ n_236;
assign n_794 = n_5 ^ n_237;
assign n_795 = n_6 ^ n_238;
assign n_796 = n_7 ^ n_239;
assign n_797 = n_8 ^ n_240;
assign n_798 = n_9 ^ n_241;
assign n_799 = n_10 ^ n_242;
assign n_800 = n_11 ^ n_243;
assign n_801 = n_12 ^ n_244;
assign n_802 = n_13 ^ n_245;
assign n_803 = n_14 ^ n_246;
assign n_804 = n_15 ^ n_247;
assign n_805 = n_16 ^ n_248;
assign n_806 = n_17 ^ n_249;
assign n_807 = n_18 ^ n_250;
assign n_808 = n_19 ^ n_251;
assign n_809 = n_20 ^ n_252;
assign n_810 = n_21 ^ n_253;
assign n_811 = n_22 ^ n_254;
assign n_812 = n_23 ^ n_255;
assign n_813 = n_24 ^ n_256;
assign n_814 = n_25 ^ n_257;
assign n_815 = n_26 ^ n_258;
assign n_816 = n_27 ^ n_259;
assign n_817 = n_28 ^ n_260;
assign n_818 = n_29 ^ n_261;
assign n_819 = n_30 ^ n_262;
assign n_820 = n_31 ^ n_263;
assign n_821 = n_264 ^ n_92;
assign n_822 = x35 & ~n_265;
assign n_823 = x1 & ~n_267;
assign n_824 = x2 & ~n_267;
assign n_825 = x3 & ~n_267;
assign n_826 = x4 & ~n_267;
assign n_827 = x5 & ~n_267;
assign n_828 = x6 & ~n_267;
assign n_829 = x7 & ~n_267;
assign n_830 = x8 & ~n_267;
assign n_831 = x9 & ~n_267;
assign n_832 = x10 & ~n_267;
assign n_833 = x11 & ~n_267;
assign n_834 = x12 & ~n_267;
assign n_835 = x13 & ~n_267;
assign n_836 = x14 & ~n_267;
assign n_837 = x15 & ~n_267;
assign n_838 = x16 & ~n_267;
assign n_839 = x17 & ~n_267;
assign n_840 = x18 & ~n_267;
assign n_841 = x19 & ~n_267;
assign n_842 = x20 & ~n_267;
assign n_843 = x21 & ~n_267;
assign n_844 = x22 & ~n_267;
assign n_845 = x23 & ~n_267;
assign n_846 = x24 & ~n_267;
assign n_847 = x25 & ~n_267;
assign n_848 = x26 & ~n_267;
assign n_849 = x27 & ~n_267;
assign n_850 = x28 & ~n_267;
assign n_851 = x29 & ~n_267;
assign n_852 = x30 & ~n_267;
assign n_853 = ~x1 & n_298;
assign n_854 = n_298 ^ n_161;
assign n_855 = ~x2 & n_298;
assign n_856 = ~x3 & n_298;
assign n_857 = ~x4 & n_298;
assign n_858 = ~x5 & n_298;
assign n_859 = ~x6 & n_298;
assign n_860 = ~x7 & n_298;
assign n_861 = ~x8 & n_298;
assign n_862 = ~x9 & n_298;
assign n_863 = ~x10 & n_298;
assign n_864 = ~x11 & n_298;
assign n_865 = ~x12 & n_298;
assign n_866 = ~x13 & n_298;
assign n_867 = ~x14 & n_298;
assign n_868 = ~x15 & n_298;
assign n_869 = ~x16 & n_298;
assign n_870 = ~x17 & n_298;
assign n_871 = ~x18 & n_298;
assign n_872 = ~x19 & n_298;
assign n_873 = ~x20 & n_298;
assign n_874 = ~x21 & n_298;
assign n_875 = ~x22 & n_298;
assign n_876 = ~x23 & n_298;
assign n_877 = ~x24 & n_298;
assign n_878 = ~x25 & n_298;
assign n_879 = ~x26 & n_298;
assign n_880 = ~x27 & n_298;
assign n_881 = ~x28 & n_298;
assign n_882 = ~x29 & n_298;
assign n_883 = ~x30 & n_298;
assign n_884 = n_298 ^ n_160;
assign n_885 = n_299 ^ n_160;
assign n_886 = x1 & ~n_301;
assign n_887 = x2 & ~n_301;
assign n_888 = x3 & ~n_301;
assign n_889 = x4 & ~n_301;
assign n_890 = x5 & ~n_301;
assign n_891 = x6 & ~n_301;
assign n_892 = x7 & ~n_301;
assign n_893 = x8 & ~n_301;
assign n_894 = x9 & ~n_301;
assign n_895 = x10 & ~n_301;
assign n_896 = x11 & ~n_301;
assign n_897 = x12 & ~n_301;
assign n_898 = x13 & ~n_301;
assign n_899 = x14 & ~n_301;
assign n_900 = x15 & ~n_301;
assign n_901 = x16 & ~n_301;
assign n_902 = x17 & ~n_301;
assign n_903 = x18 & ~n_301;
assign n_904 = x19 & ~n_301;
assign n_905 = x20 & ~n_301;
assign n_906 = x21 & ~n_301;
assign n_907 = x22 & ~n_301;
assign n_908 = x23 & ~n_301;
assign n_909 = x24 & ~n_301;
assign n_910 = x25 & ~n_301;
assign n_911 = x26 & ~n_301;
assign n_912 = x27 & ~n_301;
assign n_913 = x28 & ~n_301;
assign n_914 = x29 & ~n_301;
assign n_915 = x30 & ~n_301;
assign n_916 = x37 & ~n_331;
assign n_917 = ~x1 & n_333;
assign n_918 = n_333 ^ n_166;
assign n_919 = ~x2 & n_333;
assign n_920 = ~x3 & n_333;
assign n_921 = ~x4 & n_333;
assign n_922 = ~x5 & n_333;
assign n_923 = ~x6 & n_333;
assign n_924 = ~x7 & n_333;
assign n_925 = ~x8 & n_333;
assign n_926 = ~x9 & n_333;
assign n_927 = ~x10 & n_333;
assign n_928 = ~x11 & n_333;
assign n_929 = ~x12 & n_333;
assign n_930 = ~x13 & n_333;
assign n_931 = ~x14 & n_333;
assign n_932 = ~x15 & n_333;
assign n_933 = ~x16 & n_333;
assign n_934 = ~x17 & n_333;
assign n_935 = ~x18 & n_333;
assign n_936 = ~x19 & n_333;
assign n_937 = ~x20 & n_333;
assign n_938 = ~x21 & n_333;
assign n_939 = ~x22 & n_333;
assign n_940 = ~x23 & n_333;
assign n_941 = ~x24 & n_333;
assign n_942 = ~x25 & n_333;
assign n_943 = ~x26 & n_333;
assign n_944 = ~x27 & n_333;
assign n_945 = ~x28 & n_333;
assign n_946 = ~x29 & n_333;
assign n_947 = ~x30 & n_333;
assign n_948 = n_333 ^ n_164;
assign n_949 = n_334 ^ n_164;
assign n_950 = x39 & ~n_335;
assign n_951 = x1 & ~n_337;
assign n_952 = x2 & ~n_337;
assign n_953 = x3 & ~n_337;
assign n_954 = x4 & ~n_337;
assign n_955 = x5 & ~n_337;
assign n_956 = x6 & ~n_337;
assign n_957 = x7 & ~n_337;
assign n_958 = x8 & ~n_337;
assign n_959 = x9 & ~n_337;
assign n_960 = x10 & ~n_337;
assign n_961 = x11 & ~n_337;
assign n_962 = x12 & ~n_337;
assign n_963 = x13 & ~n_337;
assign n_964 = x14 & ~n_337;
assign n_965 = x15 & ~n_337;
assign n_966 = x16 & ~n_337;
assign n_967 = x17 & ~n_337;
assign n_968 = x18 & ~n_337;
assign n_969 = x19 & ~n_337;
assign n_970 = x20 & ~n_337;
assign n_971 = x21 & ~n_337;
assign n_972 = x22 & ~n_337;
assign n_973 = x23 & ~n_337;
assign n_974 = x24 & ~n_337;
assign n_975 = x25 & ~n_337;
assign n_976 = x26 & ~n_337;
assign n_977 = x27 & ~n_337;
assign n_978 = x28 & ~n_337;
assign n_979 = x29 & ~n_337;
assign n_980 = x30 & ~n_337;
assign n_981 = ~x1 & n_368;
assign n_982 = n_368 ^ n_171;
assign n_983 = ~x2 & n_368;
assign n_984 = ~x3 & n_368;
assign n_985 = ~x4 & n_368;
assign n_986 = ~x5 & n_368;
assign n_987 = ~x6 & n_368;
assign n_988 = ~x7 & n_368;
assign n_989 = ~x8 & n_368;
assign n_990 = ~x9 & n_368;
assign n_991 = ~x10 & n_368;
assign n_992 = ~x11 & n_368;
assign n_993 = ~x12 & n_368;
assign n_994 = ~x13 & n_368;
assign n_995 = ~x14 & n_368;
assign n_996 = ~x15 & n_368;
assign n_997 = ~x16 & n_368;
assign n_998 = ~x17 & n_368;
assign n_999 = ~x18 & n_368;
assign n_1000 = ~x19 & n_368;
assign n_1001 = ~x20 & n_368;
assign n_1002 = ~x21 & n_368;
assign n_1003 = ~x22 & n_368;
assign n_1004 = ~x23 & n_368;
assign n_1005 = ~x24 & n_368;
assign n_1006 = ~x25 & n_368;
assign n_1007 = ~x26 & n_368;
assign n_1008 = ~x27 & n_368;
assign n_1009 = ~x28 & n_368;
assign n_1010 = ~x29 & n_368;
assign n_1011 = ~x30 & n_368;
assign n_1012 = n_368 ^ n_170;
assign n_1013 = n_369 ^ n_170;
assign n_1014 = x1 & ~n_371;
assign n_1015 = x2 & ~n_371;
assign n_1016 = x3 & ~n_371;
assign n_1017 = x4 & ~n_371;
assign n_1018 = x5 & ~n_371;
assign n_1019 = x6 & ~n_371;
assign n_1020 = x7 & ~n_371;
assign n_1021 = x8 & ~n_371;
assign n_1022 = x9 & ~n_371;
assign n_1023 = x10 & ~n_371;
assign n_1024 = x11 & ~n_371;
assign n_1025 = x12 & ~n_371;
assign n_1026 = x13 & ~n_371;
assign n_1027 = x14 & ~n_371;
assign n_1028 = x15 & ~n_371;
assign n_1029 = x16 & ~n_371;
assign n_1030 = x17 & ~n_371;
assign n_1031 = x18 & ~n_371;
assign n_1032 = x19 & ~n_371;
assign n_1033 = x20 & ~n_371;
assign n_1034 = x21 & ~n_371;
assign n_1035 = x22 & ~n_371;
assign n_1036 = x23 & ~n_371;
assign n_1037 = x24 & ~n_371;
assign n_1038 = x25 & ~n_371;
assign n_1039 = x26 & ~n_371;
assign n_1040 = x27 & ~n_371;
assign n_1041 = x28 & ~n_371;
assign n_1042 = x29 & ~n_371;
assign n_1043 = x30 & ~n_371;
assign n_1044 = x41 & ~n_401;
assign n_1045 = ~x1 & n_403;
assign n_1046 = n_403 ^ n_176;
assign n_1047 = ~x2 & n_403;
assign n_1048 = ~x3 & n_403;
assign n_1049 = ~x4 & n_403;
assign n_1050 = ~x5 & n_403;
assign n_1051 = ~x6 & n_403;
assign n_1052 = ~x7 & n_403;
assign n_1053 = ~x8 & n_403;
assign n_1054 = ~x9 & n_403;
assign n_1055 = ~x10 & n_403;
assign n_1056 = ~x11 & n_403;
assign n_1057 = ~x12 & n_403;
assign n_1058 = ~x13 & n_403;
assign n_1059 = ~x14 & n_403;
assign n_1060 = ~x15 & n_403;
assign n_1061 = ~x16 & n_403;
assign n_1062 = ~x17 & n_403;
assign n_1063 = ~x18 & n_403;
assign n_1064 = ~x19 & n_403;
assign n_1065 = ~x20 & n_403;
assign n_1066 = ~x21 & n_403;
assign n_1067 = ~x22 & n_403;
assign n_1068 = ~x23 & n_403;
assign n_1069 = ~x24 & n_403;
assign n_1070 = ~x25 & n_403;
assign n_1071 = ~x26 & n_403;
assign n_1072 = ~x27 & n_403;
assign n_1073 = ~x28 & n_403;
assign n_1074 = ~x29 & n_403;
assign n_1075 = ~x30 & n_403;
assign n_1076 = n_403 ^ n_174;
assign n_1077 = n_404 ^ n_174;
assign n_1078 = ~x1 & ~n_406;
assign n_1079 = ~x2 & ~n_406;
assign n_1080 = ~x3 & ~n_406;
assign n_1081 = ~x4 & ~n_406;
assign n_1082 = ~x5 & ~n_406;
assign n_1083 = ~x6 & ~n_406;
assign n_1084 = ~x7 & ~n_406;
assign n_1085 = ~x8 & ~n_406;
assign n_1086 = ~x9 & ~n_406;
assign n_1087 = ~x10 & ~n_406;
assign n_1088 = ~x11 & ~n_406;
assign n_1089 = ~x12 & ~n_406;
assign n_1090 = ~x13 & ~n_406;
assign n_1091 = ~x14 & ~n_406;
assign n_1092 = ~x15 & ~n_406;
assign n_1093 = ~x16 & ~n_406;
assign n_1094 = ~x17 & ~n_406;
assign n_1095 = ~x18 & ~n_406;
assign n_1096 = ~x19 & ~n_406;
assign n_1097 = ~x20 & ~n_406;
assign n_1098 = ~x21 & ~n_406;
assign n_1099 = ~x22 & ~n_406;
assign n_1100 = ~x23 & ~n_406;
assign n_1101 = ~x24 & ~n_406;
assign n_1102 = ~x25 & ~n_406;
assign n_1103 = ~x26 & ~n_406;
assign n_1104 = ~x27 & ~n_406;
assign n_1105 = ~x28 & ~n_406;
assign n_1106 = ~x29 & ~n_406;
assign n_1107 = ~x30 & ~n_406;
assign n_1108 = x43 & ~n_436;
assign n_1109 = x1 & n_438;
assign n_1110 = n_438 ^ n_181;
assign n_1111 = x2 & n_438;
assign n_1112 = x3 & n_438;
assign n_1113 = x4 & n_438;
assign n_1114 = x5 & n_438;
assign n_1115 = x6 & n_438;
assign n_1116 = x7 & n_438;
assign n_1117 = x8 & n_438;
assign n_1118 = x9 & n_438;
assign n_1119 = x10 & n_438;
assign n_1120 = x11 & n_438;
assign n_1121 = x12 & n_438;
assign n_1122 = x13 & n_438;
assign n_1123 = x14 & n_438;
assign n_1124 = x15 & n_438;
assign n_1125 = x16 & n_438;
assign n_1126 = x17 & n_438;
assign n_1127 = x18 & n_438;
assign n_1128 = x19 & n_438;
assign n_1129 = x20 & n_438;
assign n_1130 = x21 & n_438;
assign n_1131 = x22 & n_438;
assign n_1132 = x23 & n_438;
assign n_1133 = x24 & n_438;
assign n_1134 = x25 & n_438;
assign n_1135 = x26 & n_438;
assign n_1136 = x27 & n_438;
assign n_1137 = x28 & n_438;
assign n_1138 = x29 & n_438;
assign n_1139 = x30 & n_438;
assign n_1140 = n_439 ^ n_406;
assign n_1141 = x45 & ~n_440;
assign n_1142 = x1 & ~n_442;
assign n_1143 = x2 & ~n_442;
assign n_1144 = x3 & ~n_442;
assign n_1145 = x4 & ~n_442;
assign n_1146 = x5 & ~n_442;
assign n_1147 = x6 & ~n_442;
assign n_1148 = x7 & ~n_442;
assign n_1149 = x8 & ~n_442;
assign n_1150 = x9 & ~n_442;
assign n_1151 = x10 & ~n_442;
assign n_1152 = x11 & ~n_442;
assign n_1153 = x12 & ~n_442;
assign n_1154 = x13 & ~n_442;
assign n_1155 = x14 & ~n_442;
assign n_1156 = x15 & ~n_442;
assign n_1157 = x16 & ~n_442;
assign n_1158 = x17 & ~n_442;
assign n_1159 = x18 & ~n_442;
assign n_1160 = x19 & ~n_442;
assign n_1161 = x20 & ~n_442;
assign n_1162 = x21 & ~n_442;
assign n_1163 = x22 & ~n_442;
assign n_1164 = x23 & ~n_442;
assign n_1165 = x24 & ~n_442;
assign n_1166 = x25 & ~n_442;
assign n_1167 = x26 & ~n_442;
assign n_1168 = x27 & ~n_442;
assign n_1169 = x28 & ~n_442;
assign n_1170 = x29 & ~n_442;
assign n_1171 = x30 & ~n_442;
assign n_1172 = ~x1 & n_473;
assign n_1173 = n_473 ^ n_186;
assign n_1174 = ~x2 & n_473;
assign n_1175 = ~x3 & n_473;
assign n_1176 = ~x4 & n_473;
assign n_1177 = ~x5 & n_473;
assign n_1178 = ~x6 & n_473;
assign n_1179 = ~x7 & n_473;
assign n_1180 = ~x8 & n_473;
assign n_1181 = ~x9 & n_473;
assign n_1182 = ~x10 & n_473;
assign n_1183 = ~x11 & n_473;
assign n_1184 = ~x12 & n_473;
assign n_1185 = ~x13 & n_473;
assign n_1186 = ~x14 & n_473;
assign n_1187 = ~x15 & n_473;
assign n_1188 = ~x16 & n_473;
assign n_1189 = ~x17 & n_473;
assign n_1190 = ~x18 & n_473;
assign n_1191 = ~x19 & n_473;
assign n_1192 = ~x20 & n_473;
assign n_1193 = ~x21 & n_473;
assign n_1194 = ~x22 & n_473;
assign n_1195 = ~x23 & n_473;
assign n_1196 = ~x24 & n_473;
assign n_1197 = ~x25 & n_473;
assign n_1198 = ~x26 & n_473;
assign n_1199 = ~x27 & n_473;
assign n_1200 = ~x28 & n_473;
assign n_1201 = ~x29 & n_473;
assign n_1202 = ~x30 & n_473;
assign n_1203 = n_473 ^ n_185;
assign n_1204 = n_474 ^ n_185;
assign n_1205 = ~x1 & ~n_476;
assign n_1206 = ~x2 & ~n_476;
assign n_1207 = ~x3 & ~n_476;
assign n_1208 = ~x4 & ~n_476;
assign n_1209 = ~x5 & ~n_476;
assign n_1210 = ~x6 & ~n_476;
assign n_1211 = ~x7 & ~n_476;
assign n_1212 = ~x8 & ~n_476;
assign n_1213 = ~x9 & ~n_476;
assign n_1214 = ~x10 & ~n_476;
assign n_1215 = ~x11 & ~n_476;
assign n_1216 = ~x12 & ~n_476;
assign n_1217 = ~x13 & ~n_476;
assign n_1218 = ~x14 & ~n_476;
assign n_1219 = ~x15 & ~n_476;
assign n_1220 = ~x16 & ~n_476;
assign n_1221 = ~x17 & ~n_476;
assign n_1222 = ~x18 & ~n_476;
assign n_1223 = ~x19 & ~n_476;
assign n_1224 = ~x20 & ~n_476;
assign n_1225 = ~x21 & ~n_476;
assign n_1226 = ~x22 & ~n_476;
assign n_1227 = ~x23 & ~n_476;
assign n_1228 = ~x24 & ~n_476;
assign n_1229 = ~x25 & ~n_476;
assign n_1230 = ~x26 & ~n_476;
assign n_1231 = ~x27 & ~n_476;
assign n_1232 = ~x28 & ~n_476;
assign n_1233 = ~x29 & ~n_476;
assign n_1234 = ~x30 & ~n_476;
assign n_1235 = x47 & ~n_506;
assign n_1236 = x1 & n_508;
assign n_1237 = n_508 ^ n_191;
assign n_1238 = x2 & n_508;
assign n_1239 = x3 & n_508;
assign n_1240 = x4 & n_508;
assign n_1241 = x5 & n_508;
assign n_1242 = x6 & n_508;
assign n_1243 = x7 & n_508;
assign n_1244 = x8 & n_508;
assign n_1245 = x9 & n_508;
assign n_1246 = x10 & n_508;
assign n_1247 = x11 & n_508;
assign n_1248 = x12 & n_508;
assign n_1249 = x13 & n_508;
assign n_1250 = x14 & n_508;
assign n_1251 = x15 & n_508;
assign n_1252 = x16 & n_508;
assign n_1253 = x17 & n_508;
assign n_1254 = x18 & n_508;
assign n_1255 = x19 & n_508;
assign n_1256 = x20 & n_508;
assign n_1257 = x21 & n_508;
assign n_1258 = x22 & n_508;
assign n_1259 = x23 & n_508;
assign n_1260 = x24 & n_508;
assign n_1261 = x25 & n_508;
assign n_1262 = x26 & n_508;
assign n_1263 = x27 & n_508;
assign n_1264 = x28 & n_508;
assign n_1265 = x29 & n_508;
assign n_1266 = x30 & n_508;
assign n_1267 = n_509 ^ n_476;
assign n_1268 = x1 & ~n_511;
assign n_1269 = x2 & ~n_511;
assign n_1270 = x3 & ~n_511;
assign n_1271 = x4 & ~n_511;
assign n_1272 = x5 & ~n_511;
assign n_1273 = x6 & ~n_511;
assign n_1274 = x7 & ~n_511;
assign n_1275 = x8 & ~n_511;
assign n_1276 = x9 & ~n_511;
assign n_1277 = x10 & ~n_511;
assign n_1278 = x11 & ~n_511;
assign n_1279 = x12 & ~n_511;
assign n_1280 = x13 & ~n_511;
assign n_1281 = x14 & ~n_511;
assign n_1282 = x15 & ~n_511;
assign n_1283 = x16 & ~n_511;
assign n_1284 = x17 & ~n_511;
assign n_1285 = x18 & ~n_511;
assign n_1286 = x19 & ~n_511;
assign n_1287 = x20 & ~n_511;
assign n_1288 = x21 & ~n_511;
assign n_1289 = x22 & ~n_511;
assign n_1290 = x23 & ~n_511;
assign n_1291 = x24 & ~n_511;
assign n_1292 = x25 & ~n_511;
assign n_1293 = x26 & ~n_511;
assign n_1294 = x27 & ~n_511;
assign n_1295 = x28 & ~n_511;
assign n_1296 = x29 & ~n_511;
assign n_1297 = x30 & ~n_511;
assign n_1298 = x49 & ~n_541;
assign n_1299 = ~x1 & n_543;
assign n_1300 = n_543 ^ n_196;
assign n_1301 = ~x2 & n_543;
assign n_1302 = ~x3 & n_543;
assign n_1303 = ~x4 & n_543;
assign n_1304 = ~x5 & n_543;
assign n_1305 = ~x6 & n_543;
assign n_1306 = ~x7 & n_543;
assign n_1307 = ~x8 & n_543;
assign n_1308 = ~x9 & n_543;
assign n_1309 = ~x10 & n_543;
assign n_1310 = ~x11 & n_543;
assign n_1311 = ~x12 & n_543;
assign n_1312 = ~x13 & n_543;
assign n_1313 = ~x14 & n_543;
assign n_1314 = ~x15 & n_543;
assign n_1315 = ~x16 & n_543;
assign n_1316 = ~x17 & n_543;
assign n_1317 = ~x18 & n_543;
assign n_1318 = ~x19 & n_543;
assign n_1319 = ~x20 & n_543;
assign n_1320 = ~x21 & n_543;
assign n_1321 = ~x22 & n_543;
assign n_1322 = ~x23 & n_543;
assign n_1323 = ~x24 & n_543;
assign n_1324 = ~x25 & n_543;
assign n_1325 = ~x26 & n_543;
assign n_1326 = ~x27 & n_543;
assign n_1327 = ~x28 & n_543;
assign n_1328 = ~x29 & n_543;
assign n_1329 = ~x30 & n_543;
assign n_1330 = n_543 ^ n_194;
assign n_1331 = n_544 ^ n_194;
assign n_1332 = ~x1 & ~n_546;
assign n_1333 = ~x2 & ~n_546;
assign n_1334 = ~x3 & ~n_546;
assign n_1335 = ~x4 & ~n_546;
assign n_1336 = ~x5 & ~n_546;
assign n_1337 = ~x6 & ~n_546;
assign n_1338 = ~x7 & ~n_546;
assign n_1339 = ~x8 & ~n_546;
assign n_1340 = ~x9 & ~n_546;
assign n_1341 = ~x10 & ~n_546;
assign n_1342 = ~x11 & ~n_546;
assign n_1343 = ~x12 & ~n_546;
assign n_1344 = ~x13 & ~n_546;
assign n_1345 = ~x14 & ~n_546;
assign n_1346 = ~x15 & ~n_546;
assign n_1347 = ~x16 & ~n_546;
assign n_1348 = ~x17 & ~n_546;
assign n_1349 = ~x18 & ~n_546;
assign n_1350 = ~x19 & ~n_546;
assign n_1351 = ~x20 & ~n_546;
assign n_1352 = ~x21 & ~n_546;
assign n_1353 = ~x22 & ~n_546;
assign n_1354 = ~x23 & ~n_546;
assign n_1355 = ~x24 & ~n_546;
assign n_1356 = ~x25 & ~n_546;
assign n_1357 = ~x26 & ~n_546;
assign n_1358 = ~x27 & ~n_546;
assign n_1359 = ~x28 & ~n_546;
assign n_1360 = ~x29 & ~n_546;
assign n_1361 = ~x30 & ~n_546;
assign n_1362 = x51 & ~n_576;
assign n_1363 = x1 & n_578;
assign n_1364 = n_578 ^ n_201;
assign n_1365 = x2 & n_578;
assign n_1366 = x3 & n_578;
assign n_1367 = x4 & n_578;
assign n_1368 = x5 & n_578;
assign n_1369 = x6 & n_578;
assign n_1370 = x7 & n_578;
assign n_1371 = x8 & n_578;
assign n_1372 = x9 & n_578;
assign n_1373 = x10 & n_578;
assign n_1374 = x11 & n_578;
assign n_1375 = x12 & n_578;
assign n_1376 = x13 & n_578;
assign n_1377 = x14 & n_578;
assign n_1378 = x15 & n_578;
assign n_1379 = x16 & n_578;
assign n_1380 = x17 & n_578;
assign n_1381 = x18 & n_578;
assign n_1382 = x19 & n_578;
assign n_1383 = x20 & n_578;
assign n_1384 = x21 & n_578;
assign n_1385 = x22 & n_578;
assign n_1386 = x23 & n_578;
assign n_1387 = x24 & n_578;
assign n_1388 = x25 & n_578;
assign n_1389 = x26 & n_578;
assign n_1390 = x27 & n_578;
assign n_1391 = x28 & n_578;
assign n_1392 = x29 & n_578;
assign n_1393 = x30 & n_578;
assign n_1394 = n_579 ^ n_546;
assign n_1395 = x53 & ~n_580;
assign n_1396 = x1 & ~n_582;
assign n_1397 = x2 & ~n_582;
assign n_1398 = x3 & ~n_582;
assign n_1399 = x4 & ~n_582;
assign n_1400 = x5 & ~n_582;
assign n_1401 = x6 & ~n_582;
assign n_1402 = x7 & ~n_582;
assign n_1403 = x8 & ~n_582;
assign n_1404 = x9 & ~n_582;
assign n_1405 = x10 & ~n_582;
assign n_1406 = x11 & ~n_582;
assign n_1407 = x12 & ~n_582;
assign n_1408 = x13 & ~n_582;
assign n_1409 = x14 & ~n_582;
assign n_1410 = x15 & ~n_582;
assign n_1411 = x16 & ~n_582;
assign n_1412 = x17 & ~n_582;
assign n_1413 = x18 & ~n_582;
assign n_1414 = x19 & ~n_582;
assign n_1415 = x20 & ~n_582;
assign n_1416 = x21 & ~n_582;
assign n_1417 = x22 & ~n_582;
assign n_1418 = x23 & ~n_582;
assign n_1419 = x24 & ~n_582;
assign n_1420 = x25 & ~n_582;
assign n_1421 = x26 & ~n_582;
assign n_1422 = x27 & ~n_582;
assign n_1423 = x28 & ~n_582;
assign n_1424 = x29 & ~n_582;
assign n_1425 = x30 & ~n_582;
assign n_1426 = ~x1 & n_613;
assign n_1427 = n_613 ^ n_206;
assign n_1428 = ~x2 & n_613;
assign n_1429 = ~x3 & n_613;
assign n_1430 = ~x4 & n_613;
assign n_1431 = ~x5 & n_613;
assign n_1432 = ~x6 & n_613;
assign n_1433 = ~x7 & n_613;
assign n_1434 = ~x8 & n_613;
assign n_1435 = ~x9 & n_613;
assign n_1436 = ~x10 & n_613;
assign n_1437 = ~x11 & n_613;
assign n_1438 = ~x12 & n_613;
assign n_1439 = ~x13 & n_613;
assign n_1440 = ~x14 & n_613;
assign n_1441 = ~x15 & n_613;
assign n_1442 = ~x16 & n_613;
assign n_1443 = ~x17 & n_613;
assign n_1444 = ~x18 & n_613;
assign n_1445 = ~x19 & n_613;
assign n_1446 = ~x20 & n_613;
assign n_1447 = ~x21 & n_613;
assign n_1448 = ~x22 & n_613;
assign n_1449 = ~x23 & n_613;
assign n_1450 = ~x24 & n_613;
assign n_1451 = ~x25 & n_613;
assign n_1452 = ~x26 & n_613;
assign n_1453 = ~x27 & n_613;
assign n_1454 = ~x28 & n_613;
assign n_1455 = ~x29 & n_613;
assign n_1456 = ~x30 & n_613;
assign n_1457 = n_613 ^ n_205;
assign n_1458 = n_614 ^ n_205;
assign n_1459 = x55 & ~n_615;
assign n_1460 = x1 & ~n_617;
assign n_1461 = x2 & ~n_617;
assign n_1462 = x3 & ~n_617;
assign n_1463 = x4 & ~n_617;
assign n_1464 = x5 & ~n_617;
assign n_1465 = x6 & ~n_617;
assign n_1466 = x7 & ~n_617;
assign n_1467 = x8 & ~n_617;
assign n_1468 = x9 & ~n_617;
assign n_1469 = x10 & ~n_617;
assign n_1470 = x11 & ~n_617;
assign n_1471 = x12 & ~n_617;
assign n_1472 = x13 & ~n_617;
assign n_1473 = x14 & ~n_617;
assign n_1474 = x15 & ~n_617;
assign n_1475 = x16 & ~n_617;
assign n_1476 = x17 & ~n_617;
assign n_1477 = x18 & ~n_617;
assign n_1478 = x19 & ~n_617;
assign n_1479 = x20 & ~n_617;
assign n_1480 = x21 & ~n_617;
assign n_1481 = x22 & ~n_617;
assign n_1482 = x23 & ~n_617;
assign n_1483 = x24 & ~n_617;
assign n_1484 = x25 & ~n_617;
assign n_1485 = x26 & ~n_617;
assign n_1486 = x27 & ~n_617;
assign n_1487 = x28 & ~n_617;
assign n_1488 = x29 & ~n_617;
assign n_1489 = x30 & ~n_617;
assign n_1490 = ~x1 & n_648;
assign n_1491 = n_648 ^ n_211;
assign n_1492 = ~x2 & n_648;
assign n_1493 = ~x3 & n_648;
assign n_1494 = ~x4 & n_648;
assign n_1495 = ~x5 & n_648;
assign n_1496 = ~x6 & n_648;
assign n_1497 = ~x7 & n_648;
assign n_1498 = ~x8 & n_648;
assign n_1499 = ~x9 & n_648;
assign n_1500 = ~x10 & n_648;
assign n_1501 = ~x11 & n_648;
assign n_1502 = ~x12 & n_648;
assign n_1503 = ~x13 & n_648;
assign n_1504 = ~x14 & n_648;
assign n_1505 = ~x15 & n_648;
assign n_1506 = ~x16 & n_648;
assign n_1507 = ~x17 & n_648;
assign n_1508 = ~x18 & n_648;
assign n_1509 = ~x19 & n_648;
assign n_1510 = ~x20 & n_648;
assign n_1511 = ~x21 & n_648;
assign n_1512 = ~x22 & n_648;
assign n_1513 = ~x23 & n_648;
assign n_1514 = ~x24 & n_648;
assign n_1515 = ~x25 & n_648;
assign n_1516 = ~x26 & n_648;
assign n_1517 = ~x27 & n_648;
assign n_1518 = ~x28 & n_648;
assign n_1519 = ~x29 & n_648;
assign n_1520 = ~x30 & n_648;
assign n_1521 = n_648 ^ n_210;
assign n_1522 = n_649 ^ n_210;
assign n_1523 = x57 & ~n_650;
assign n_1524 = x1 & ~n_652;
assign n_1525 = x2 & ~n_652;
assign n_1526 = x3 & ~n_652;
assign n_1527 = x4 & ~n_652;
assign n_1528 = x5 & ~n_652;
assign n_1529 = x6 & ~n_652;
assign n_1530 = x7 & ~n_652;
assign n_1531 = x8 & ~n_652;
assign n_1532 = x9 & ~n_652;
assign n_1533 = x10 & ~n_652;
assign n_1534 = x11 & ~n_652;
assign n_1535 = x12 & ~n_652;
assign n_1536 = x13 & ~n_652;
assign n_1537 = x14 & ~n_652;
assign n_1538 = x15 & ~n_652;
assign n_1539 = x16 & ~n_652;
assign n_1540 = x17 & ~n_652;
assign n_1541 = x18 & ~n_652;
assign n_1542 = x19 & ~n_652;
assign n_1543 = x20 & ~n_652;
assign n_1544 = x21 & ~n_652;
assign n_1545 = x22 & ~n_652;
assign n_1546 = x23 & ~n_652;
assign n_1547 = x24 & ~n_652;
assign n_1548 = x25 & ~n_652;
assign n_1549 = x26 & ~n_652;
assign n_1550 = x27 & ~n_652;
assign n_1551 = x28 & ~n_652;
assign n_1552 = x29 & ~n_652;
assign n_1553 = x30 & ~n_652;
assign n_1554 = ~x1 & n_683;
assign n_1555 = n_683 ^ n_216;
assign n_1556 = ~x2 & n_683;
assign n_1557 = ~x3 & n_683;
assign n_1558 = ~x4 & n_683;
assign n_1559 = ~x5 & n_683;
assign n_1560 = ~x6 & n_683;
assign n_1561 = ~x7 & n_683;
assign n_1562 = ~x8 & n_683;
assign n_1563 = ~x9 & n_683;
assign n_1564 = ~x10 & n_683;
assign n_1565 = ~x11 & n_683;
assign n_1566 = ~x12 & n_683;
assign n_1567 = ~x13 & n_683;
assign n_1568 = ~x14 & n_683;
assign n_1569 = ~x15 & n_683;
assign n_1570 = ~x16 & n_683;
assign n_1571 = ~x17 & n_683;
assign n_1572 = ~x18 & n_683;
assign n_1573 = ~x19 & n_683;
assign n_1574 = ~x20 & n_683;
assign n_1575 = ~x21 & n_683;
assign n_1576 = ~x22 & n_683;
assign n_1577 = ~x23 & n_683;
assign n_1578 = ~x24 & n_683;
assign n_1579 = ~x25 & n_683;
assign n_1580 = ~x26 & n_683;
assign n_1581 = ~x27 & n_683;
assign n_1582 = ~x28 & n_683;
assign n_1583 = ~x29 & n_683;
assign n_1584 = ~x30 & n_683;
assign n_1585 = n_683 ^ n_215;
assign n_1586 = n_684 ^ n_215;
assign n_1587 = ~x1 & ~n_686;
assign n_1588 = ~x2 & ~n_686;
assign n_1589 = ~x3 & ~n_686;
assign n_1590 = ~x4 & ~n_686;
assign n_1591 = ~x5 & ~n_686;
assign n_1592 = ~x6 & ~n_686;
assign n_1593 = ~x7 & ~n_686;
assign n_1594 = ~x8 & ~n_686;
assign n_1595 = ~x9 & ~n_686;
assign n_1596 = ~x10 & ~n_686;
assign n_1597 = ~x11 & ~n_686;
assign n_1598 = ~x12 & ~n_686;
assign n_1599 = ~x13 & ~n_686;
assign n_1600 = ~x14 & ~n_686;
assign n_1601 = ~x15 & ~n_686;
assign n_1602 = ~x16 & ~n_686;
assign n_1603 = ~x17 & ~n_686;
assign n_1604 = ~x18 & ~n_686;
assign n_1605 = ~x19 & ~n_686;
assign n_1606 = ~x20 & ~n_686;
assign n_1607 = ~x21 & ~n_686;
assign n_1608 = ~x22 & ~n_686;
assign n_1609 = ~x23 & ~n_686;
assign n_1610 = ~x24 & ~n_686;
assign n_1611 = ~x25 & ~n_686;
assign n_1612 = ~x26 & ~n_686;
assign n_1613 = ~x27 & ~n_686;
assign n_1614 = ~x28 & ~n_686;
assign n_1615 = ~x29 & ~n_686;
assign n_1616 = ~x30 & ~n_686;
assign n_1617 = x59 & ~n_716;
assign n_1618 = x1 & n_718;
assign n_1619 = n_718 ^ n_221;
assign n_1620 = x2 & n_718;
assign n_1621 = x3 & n_718;
assign n_1622 = x4 & n_718;
assign n_1623 = x5 & n_718;
assign n_1624 = x6 & n_718;
assign n_1625 = x7 & n_718;
assign n_1626 = x8 & n_718;
assign n_1627 = x9 & n_718;
assign n_1628 = x10 & n_718;
assign n_1629 = x11 & n_718;
assign n_1630 = x12 & n_718;
assign n_1631 = x13 & n_718;
assign n_1632 = x14 & n_718;
assign n_1633 = x15 & n_718;
assign n_1634 = x16 & n_718;
assign n_1635 = x17 & n_718;
assign n_1636 = x18 & n_718;
assign n_1637 = x19 & n_718;
assign n_1638 = x20 & n_718;
assign n_1639 = x21 & n_718;
assign n_1640 = x22 & n_718;
assign n_1641 = x23 & n_718;
assign n_1642 = x24 & n_718;
assign n_1643 = x25 & n_718;
assign n_1644 = x26 & n_718;
assign n_1645 = x27 & n_718;
assign n_1646 = x28 & n_718;
assign n_1647 = x29 & n_718;
assign n_1648 = x30 & n_718;
assign n_1649 = n_719 ^ n_686;
assign n_1650 = x1 & ~n_721;
assign n_1651 = x2 & ~n_721;
assign n_1652 = x3 & ~n_721;
assign n_1653 = x4 & ~n_721;
assign n_1654 = x5 & ~n_721;
assign n_1655 = x6 & ~n_721;
assign n_1656 = x7 & ~n_721;
assign n_1657 = x8 & ~n_721;
assign n_1658 = x9 & ~n_721;
assign n_1659 = x10 & ~n_721;
assign n_1660 = x11 & ~n_721;
assign n_1661 = x12 & ~n_721;
assign n_1662 = x13 & ~n_721;
assign n_1663 = x14 & ~n_721;
assign n_1664 = x15 & ~n_721;
assign n_1665 = x16 & ~n_721;
assign n_1666 = x17 & ~n_721;
assign n_1667 = x18 & ~n_721;
assign n_1668 = x19 & ~n_721;
assign n_1669 = x20 & ~n_721;
assign n_1670 = x21 & ~n_721;
assign n_1671 = x22 & ~n_721;
assign n_1672 = x23 & ~n_721;
assign n_1673 = x24 & ~n_721;
assign n_1674 = x25 & ~n_721;
assign n_1675 = x26 & ~n_721;
assign n_1676 = x27 & ~n_721;
assign n_1677 = x28 & ~n_721;
assign n_1678 = x29 & ~n_721;
assign n_1679 = x30 & ~n_721;
assign n_1680 = x61 & ~n_751;
assign n_1681 = ~x1 & n_753;
assign n_1682 = n_753 ^ n_226;
assign n_1683 = ~x2 & n_753;
assign n_1684 = ~x3 & n_753;
assign n_1685 = ~x4 & n_753;
assign n_1686 = ~x5 & n_753;
assign n_1687 = ~x6 & n_753;
assign n_1688 = ~x7 & n_753;
assign n_1689 = ~x8 & n_753;
assign n_1690 = ~x9 & n_753;
assign n_1691 = ~x10 & n_753;
assign n_1692 = ~x11 & n_753;
assign n_1693 = ~x12 & n_753;
assign n_1694 = ~x13 & n_753;
assign n_1695 = ~x14 & n_753;
assign n_1696 = ~x15 & n_753;
assign n_1697 = ~x16 & n_753;
assign n_1698 = ~x17 & n_753;
assign n_1699 = ~x18 & n_753;
assign n_1700 = ~x19 & n_753;
assign n_1701 = ~x20 & n_753;
assign n_1702 = ~x21 & n_753;
assign n_1703 = ~x22 & n_753;
assign n_1704 = ~x23 & n_753;
assign n_1705 = ~x24 & n_753;
assign n_1706 = ~x25 & n_753;
assign n_1707 = ~x26 & n_753;
assign n_1708 = ~x27 & n_753;
assign n_1709 = ~x28 & n_753;
assign n_1710 = ~x29 & n_753;
assign n_1711 = ~x30 & n_753;
assign n_1712 = n_753 ^ n_224;
assign n_1713 = n_754 ^ n_224;
assign n_1714 = x1 & ~n_756;
assign n_1715 = x2 & ~n_756;
assign n_1716 = x3 & ~n_756;
assign n_1717 = x4 & ~n_756;
assign n_1718 = x5 & ~n_756;
assign n_1719 = x6 & ~n_756;
assign n_1720 = x7 & ~n_756;
assign n_1721 = x8 & ~n_756;
assign n_1722 = x9 & ~n_756;
assign n_1723 = x10 & ~n_756;
assign n_1724 = x11 & ~n_756;
assign n_1725 = x12 & ~n_756;
assign n_1726 = x13 & ~n_756;
assign n_1727 = x14 & ~n_756;
assign n_1728 = x15 & ~n_756;
assign n_1729 = x16 & ~n_756;
assign n_1730 = x17 & ~n_756;
assign n_1731 = x18 & ~n_756;
assign n_1732 = x19 & ~n_756;
assign n_1733 = x20 & ~n_756;
assign n_1734 = x21 & ~n_756;
assign n_1735 = x22 & ~n_756;
assign n_1736 = x23 & ~n_756;
assign n_1737 = x24 & ~n_756;
assign n_1738 = x25 & ~n_756;
assign n_1739 = x26 & ~n_756;
assign n_1740 = x27 & ~n_756;
assign n_1741 = x28 & ~n_756;
assign n_1742 = x29 & ~n_756;
assign n_1743 = x30 & ~n_756;
assign n_1744 = x63 & ~n_786;
assign n_1745 = ~x0 & n_787;
assign n_1746 = n_787 ^ n_231;
assign n_1747 = ~x1 & n_787;
assign n_1748 = ~x2 & n_787;
assign n_1749 = ~x3 & n_787;
assign n_1750 = ~x4 & n_787;
assign n_1751 = ~x5 & n_787;
assign n_1752 = ~x6 & n_787;
assign n_1753 = ~x7 & n_787;
assign n_1754 = ~x8 & n_787;
assign n_1755 = ~x9 & n_787;
assign n_1756 = ~x10 & n_787;
assign n_1757 = ~x11 & n_787;
assign n_1758 = ~x12 & n_787;
assign n_1759 = ~x13 & n_787;
assign n_1760 = ~x14 & n_787;
assign n_1761 = ~x15 & n_787;
assign n_1762 = ~x16 & n_787;
assign n_1763 = ~x17 & n_787;
assign n_1764 = ~x18 & n_787;
assign n_1765 = ~x19 & n_787;
assign n_1766 = ~x20 & n_787;
assign n_1767 = ~x21 & n_787;
assign n_1768 = ~x22 & n_787;
assign n_1769 = ~x23 & n_787;
assign n_1770 = ~x24 & n_787;
assign n_1771 = ~x25 & n_787;
assign n_1772 = ~x26 & n_787;
assign n_1773 = ~x27 & n_787;
assign n_1774 = ~x28 & n_787;
assign n_1775 = ~x29 & n_787;
assign n_1776 = ~x30 & n_787;
assign n_1777 = n_788 ^ n_229;
assign n_1778 = n_789 ^ x31;
assign n_1779 = n_124 ^ n_790;
assign n_1780 = n_790 & n_124;
assign n_1781 = n_158 ^ n_791;
assign n_1782 = n_163 ^ n_793;
assign n_1783 = n_168 ^ n_795;
assign n_1784 = n_173 ^ n_797;
assign n_1785 = n_188 ^ n_803;
assign n_1786 = n_193 ^ n_805;
assign n_1787 = n_198 ^ n_807;
assign n_1788 = n_203 ^ n_809;
assign n_1789 = n_228 ^ n_819;
assign n_1790 = n_822 ^ n_792;
assign n_1791 = n_792 & n_822;
assign n_1792 = n_266 ^ n_823;
assign n_1793 = n_268 ^ n_824;
assign n_1794 = n_269 ^ n_825;
assign n_1795 = n_270 ^ n_826;
assign n_1796 = n_271 ^ n_827;
assign n_1797 = n_272 ^ n_828;
assign n_1798 = n_273 ^ n_829;
assign n_1799 = n_274 ^ n_830;
assign n_1800 = n_275 ^ n_831;
assign n_1801 = n_276 ^ n_832;
assign n_1802 = n_277 ^ n_833;
assign n_1803 = n_278 ^ n_834;
assign n_1804 = n_279 ^ n_835;
assign n_1805 = n_280 ^ n_836;
assign n_1806 = n_281 ^ n_837;
assign n_1807 = n_282 ^ n_838;
assign n_1808 = n_283 ^ n_839;
assign n_1809 = n_284 ^ n_840;
assign n_1810 = n_285 ^ n_841;
assign n_1811 = n_286 ^ n_842;
assign n_1812 = n_287 ^ n_843;
assign n_1813 = n_288 ^ n_844;
assign n_1814 = n_289 ^ n_845;
assign n_1815 = n_290 ^ n_846;
assign n_1816 = n_291 ^ n_847;
assign n_1817 = n_292 ^ n_848;
assign n_1818 = n_293 ^ n_849;
assign n_1819 = n_294 ^ n_850;
assign n_1820 = n_295 ^ n_851;
assign n_1821 = n_296 ^ n_852;
assign n_1822 = x1 & n_854;
assign n_1823 = x2 & n_854;
assign n_1824 = x3 & n_854;
assign n_1825 = x4 & n_854;
assign n_1826 = x5 & n_854;
assign n_1827 = x6 & n_854;
assign n_1828 = x7 & n_854;
assign n_1829 = x8 & n_854;
assign n_1830 = x9 & n_854;
assign n_1831 = x10 & n_854;
assign n_1832 = x11 & n_854;
assign n_1833 = x12 & n_854;
assign n_1834 = x13 & n_854;
assign n_1835 = x14 & n_854;
assign n_1836 = x15 & n_854;
assign n_1837 = x16 & n_854;
assign n_1838 = x17 & n_854;
assign n_1839 = x18 & n_854;
assign n_1840 = x19 & n_854;
assign n_1841 = x20 & n_854;
assign n_1842 = x21 & n_854;
assign n_1843 = x22 & n_854;
assign n_1844 = x23 & n_854;
assign n_1845 = x24 & n_854;
assign n_1846 = x25 & n_854;
assign n_1847 = x26 & n_854;
assign n_1848 = x27 & n_854;
assign n_1849 = x28 & n_854;
assign n_1850 = x29 & n_854;
assign n_1851 = x30 & n_854;
assign n_1852 = n_885 ^ x33;
assign n_1853 = n_300 ^ n_886;
assign n_1854 = n_302 ^ n_887;
assign n_1855 = n_303 ^ n_888;
assign n_1856 = n_304 ^ n_889;
assign n_1857 = n_305 ^ n_890;
assign n_1858 = n_306 ^ n_891;
assign n_1859 = n_307 ^ n_892;
assign n_1860 = n_308 ^ n_893;
assign n_1861 = n_309 ^ n_894;
assign n_1862 = n_310 ^ n_895;
assign n_1863 = n_311 ^ n_896;
assign n_1864 = n_312 ^ n_897;
assign n_1865 = n_313 ^ n_898;
assign n_1866 = n_314 ^ n_899;
assign n_1867 = n_315 ^ n_900;
assign n_1868 = n_316 ^ n_901;
assign n_1869 = n_317 ^ n_902;
assign n_1870 = n_318 ^ n_903;
assign n_1871 = n_319 ^ n_904;
assign n_1872 = n_320 ^ n_905;
assign n_1873 = n_321 ^ n_906;
assign n_1874 = n_322 ^ n_907;
assign n_1875 = n_323 ^ n_908;
assign n_1876 = n_324 ^ n_909;
assign n_1877 = n_325 ^ n_910;
assign n_1878 = n_326 ^ n_911;
assign n_1879 = n_327 ^ n_912;
assign n_1880 = n_328 ^ n_913;
assign n_1881 = n_329 ^ n_914;
assign n_1882 = n_330 ^ n_915;
assign n_1883 = n_916 ^ n_794;
assign n_1884 = n_794 & n_916;
assign n_1885 = x1 & n_918;
assign n_1886 = x2 & n_918;
assign n_1887 = x3 & n_918;
assign n_1888 = x4 & n_918;
assign n_1889 = x5 & n_918;
assign n_1890 = x6 & n_918;
assign n_1891 = x7 & n_918;
assign n_1892 = x8 & n_918;
assign n_1893 = x9 & n_918;
assign n_1894 = x10 & n_918;
assign n_1895 = x11 & n_918;
assign n_1896 = x12 & n_918;
assign n_1897 = x13 & n_918;
assign n_1898 = x14 & n_918;
assign n_1899 = x15 & n_918;
assign n_1900 = x16 & n_918;
assign n_1901 = x17 & n_918;
assign n_1902 = x18 & n_918;
assign n_1903 = x19 & n_918;
assign n_1904 = x20 & n_918;
assign n_1905 = x21 & n_918;
assign n_1906 = x22 & n_918;
assign n_1907 = x23 & n_918;
assign n_1908 = x24 & n_918;
assign n_1909 = x25 & n_918;
assign n_1910 = x26 & n_918;
assign n_1911 = x27 & n_918;
assign n_1912 = x28 & n_918;
assign n_1913 = x29 & n_918;
assign n_1914 = x30 & n_918;
assign n_1915 = n_96 ^ n_949;
assign n_1916 = n_950 ^ n_796;
assign n_1917 = n_796 & n_950;
assign n_1918 = n_336 ^ n_951;
assign n_1919 = n_338 ^ n_952;
assign n_1920 = n_339 ^ n_953;
assign n_1921 = n_340 ^ n_954;
assign n_1922 = n_341 ^ n_955;
assign n_1923 = n_342 ^ n_956;
assign n_1924 = n_343 ^ n_957;
assign n_1925 = n_344 ^ n_958;
assign n_1926 = n_345 ^ n_959;
assign n_1927 = n_346 ^ n_960;
assign n_1928 = n_347 ^ n_961;
assign n_1929 = n_348 ^ n_962;
assign n_1930 = n_349 ^ n_963;
assign n_1931 = n_350 ^ n_964;
assign n_1932 = n_351 ^ n_965;
assign n_1933 = n_352 ^ n_966;
assign n_1934 = n_353 ^ n_967;
assign n_1935 = n_354 ^ n_968;
assign n_1936 = n_355 ^ n_969;
assign n_1937 = n_356 ^ n_970;
assign n_1938 = n_357 ^ n_971;
assign n_1939 = n_358 ^ n_972;
assign n_1940 = n_359 ^ n_973;
assign n_1941 = n_360 ^ n_974;
assign n_1942 = n_361 ^ n_975;
assign n_1943 = n_362 ^ n_976;
assign n_1944 = n_363 ^ n_977;
assign n_1945 = n_364 ^ n_978;
assign n_1946 = n_365 ^ n_979;
assign n_1947 = n_366 ^ n_980;
assign n_1948 = x1 & n_982;
assign n_1949 = x2 & n_982;
assign n_1950 = x3 & n_982;
assign n_1951 = x4 & n_982;
assign n_1952 = x5 & n_982;
assign n_1953 = x6 & n_982;
assign n_1954 = x7 & n_982;
assign n_1955 = x8 & n_982;
assign n_1956 = x9 & n_982;
assign n_1957 = x10 & n_982;
assign n_1958 = x11 & n_982;
assign n_1959 = x12 & n_982;
assign n_1960 = x13 & n_982;
assign n_1961 = x14 & n_982;
assign n_1962 = x15 & n_982;
assign n_1963 = x16 & n_982;
assign n_1964 = x17 & n_982;
assign n_1965 = x18 & n_982;
assign n_1966 = x19 & n_982;
assign n_1967 = x20 & n_982;
assign n_1968 = x21 & n_982;
assign n_1969 = x22 & n_982;
assign n_1970 = x23 & n_982;
assign n_1971 = x24 & n_982;
assign n_1972 = x25 & n_982;
assign n_1973 = x26 & n_982;
assign n_1974 = x27 & n_982;
assign n_1975 = x28 & n_982;
assign n_1976 = x29 & n_982;
assign n_1977 = x30 & n_982;
assign n_1978 = n_370 ^ n_1014;
assign n_1979 = n_372 ^ n_1015;
assign n_1980 = n_373 ^ n_1016;
assign n_1981 = n_374 ^ n_1017;
assign n_1982 = n_375 ^ n_1018;
assign n_1983 = n_376 ^ n_1019;
assign n_1984 = n_377 ^ n_1020;
assign n_1985 = n_378 ^ n_1021;
assign n_1986 = n_379 ^ n_1022;
assign n_1987 = n_380 ^ n_1023;
assign n_1988 = n_381 ^ n_1024;
assign n_1989 = n_382 ^ n_1025;
assign n_1990 = n_383 ^ n_1026;
assign n_1991 = n_384 ^ n_1027;
assign n_1992 = n_385 ^ n_1028;
assign n_1993 = n_386 ^ n_1029;
assign n_1994 = n_387 ^ n_1030;
assign n_1995 = n_388 ^ n_1031;
assign n_1996 = n_389 ^ n_1032;
assign n_1997 = n_390 ^ n_1033;
assign n_1998 = n_391 ^ n_1034;
assign n_1999 = n_392 ^ n_1035;
assign n_2000 = n_393 ^ n_1036;
assign n_2001 = n_394 ^ n_1037;
assign n_2002 = n_395 ^ n_1038;
assign n_2003 = n_396 ^ n_1039;
assign n_2004 = n_397 ^ n_1040;
assign n_2005 = n_398 ^ n_1041;
assign n_2006 = n_399 ^ n_1042;
assign n_2007 = n_400 ^ n_1043;
assign n_2008 = x1 & n_1046;
assign n_2009 = x2 & n_1046;
assign n_2010 = x3 & n_1046;
assign n_2011 = x4 & n_1046;
assign n_2012 = x5 & n_1046;
assign n_2013 = x6 & n_1046;
assign n_2014 = x7 & n_1046;
assign n_2015 = x8 & n_1046;
assign n_2016 = x9 & n_1046;
assign n_2017 = x10 & n_1046;
assign n_2018 = x11 & n_1046;
assign n_2019 = x12 & n_1046;
assign n_2020 = x13 & n_1046;
assign n_2021 = x14 & n_1046;
assign n_2022 = x15 & n_1046;
assign n_2023 = x16 & n_1046;
assign n_2024 = x17 & n_1046;
assign n_2025 = x18 & n_1046;
assign n_2026 = x19 & n_1046;
assign n_2027 = x20 & n_1046;
assign n_2028 = x21 & n_1046;
assign n_2029 = x22 & n_1046;
assign n_2030 = x23 & n_1046;
assign n_2031 = x24 & n_1046;
assign n_2032 = x25 & n_1046;
assign n_2033 = x26 & n_1046;
assign n_2034 = x27 & n_1046;
assign n_2035 = x28 & n_1046;
assign n_2036 = x29 & n_1046;
assign n_2037 = x30 & n_1046;
assign n_2038 = n_405 ^ n_1078;
assign n_2039 = n_407 ^ n_1079;
assign n_2040 = n_408 ^ n_1080;
assign n_2041 = n_409 ^ n_1081;
assign n_2042 = n_410 ^ n_1082;
assign n_2043 = n_411 ^ n_1083;
assign n_2044 = n_412 ^ n_1084;
assign n_2045 = n_413 ^ n_1085;
assign n_2046 = n_414 ^ n_1086;
assign n_2047 = n_415 ^ n_1087;
assign n_2048 = n_416 ^ n_1088;
assign n_2049 = n_417 ^ n_1089;
assign n_2050 = n_418 ^ n_1090;
assign n_2051 = n_419 ^ n_1091;
assign n_2052 = n_420 ^ n_1092;
assign n_2053 = n_421 ^ n_1093;
assign n_2054 = n_422 ^ n_1094;
assign n_2055 = n_423 ^ n_1095;
assign n_2056 = n_424 ^ n_1096;
assign n_2057 = n_425 ^ n_1097;
assign n_2058 = n_426 ^ n_1098;
assign n_2059 = n_427 ^ n_1099;
assign n_2060 = n_428 ^ n_1100;
assign n_2061 = n_429 ^ n_1101;
assign n_2062 = n_430 ^ n_1102;
assign n_2063 = n_431 ^ n_1103;
assign n_2064 = n_432 ^ n_1104;
assign n_2065 = n_433 ^ n_1105;
assign n_2066 = n_434 ^ n_1106;
assign n_2067 = n_435 ^ n_1107;
assign n_2068 = ~x1 & n_1110;
assign n_2069 = ~x2 & n_1110;
assign n_2070 = ~x3 & n_1110;
assign n_2071 = ~x4 & n_1110;
assign n_2072 = ~x5 & n_1110;
assign n_2073 = ~x6 & n_1110;
assign n_2074 = ~x7 & n_1110;
assign n_2075 = ~x8 & n_1110;
assign n_2076 = ~x9 & n_1110;
assign n_2077 = ~x10 & n_1110;
assign n_2078 = ~x11 & n_1110;
assign n_2079 = ~x12 & n_1110;
assign n_2080 = ~x13 & n_1110;
assign n_2081 = ~x14 & n_1110;
assign n_2082 = ~x15 & n_1110;
assign n_2083 = ~x16 & n_1110;
assign n_2084 = ~x17 & n_1110;
assign n_2085 = ~x18 & n_1110;
assign n_2086 = ~x19 & n_1110;
assign n_2087 = ~x20 & n_1110;
assign n_2088 = ~x21 & n_1110;
assign n_2089 = ~x22 & n_1110;
assign n_2090 = ~x23 & n_1110;
assign n_2091 = ~x24 & n_1110;
assign n_2092 = ~x25 & n_1110;
assign n_2093 = ~x26 & n_1110;
assign n_2094 = ~x27 & n_1110;
assign n_2095 = ~x28 & n_1110;
assign n_2096 = ~x29 & n_1110;
assign n_2097 = ~x30 & n_1110;
assign n_2098 = n_1110 ^ n_406;
assign n_2099 = n_1140 ^ n_102;
assign n_2100 = n_1141 ^ n_802;
assign n_2101 = n_802 & n_1141;
assign n_2102 = n_441 ^ n_1142;
assign n_2103 = n_443 ^ n_1143;
assign n_2104 = n_444 ^ n_1144;
assign n_2105 = n_445 ^ n_1145;
assign n_2106 = n_446 ^ n_1146;
assign n_2107 = n_447 ^ n_1147;
assign n_2108 = n_448 ^ n_1148;
assign n_2109 = n_449 ^ n_1149;
assign n_2110 = n_450 ^ n_1150;
assign n_2111 = n_451 ^ n_1151;
assign n_2112 = n_452 ^ n_1152;
assign n_2113 = n_453 ^ n_1153;
assign n_2114 = n_454 ^ n_1154;
assign n_2115 = n_455 ^ n_1155;
assign n_2116 = n_456 ^ n_1156;
assign n_2117 = n_457 ^ n_1157;
assign n_2118 = n_458 ^ n_1158;
assign n_2119 = n_459 ^ n_1159;
assign n_2120 = n_460 ^ n_1160;
assign n_2121 = n_461 ^ n_1161;
assign n_2122 = n_462 ^ n_1162;
assign n_2123 = n_463 ^ n_1163;
assign n_2124 = n_464 ^ n_1164;
assign n_2125 = n_465 ^ n_1165;
assign n_2126 = n_466 ^ n_1166;
assign n_2127 = n_467 ^ n_1167;
assign n_2128 = n_468 ^ n_1168;
assign n_2129 = n_469 ^ n_1169;
assign n_2130 = n_470 ^ n_1170;
assign n_2131 = n_471 ^ n_1171;
assign n_2132 = x1 & n_1173;
assign n_2133 = x2 & n_1173;
assign n_2134 = x3 & n_1173;
assign n_2135 = x4 & n_1173;
assign n_2136 = x5 & n_1173;
assign n_2137 = x6 & n_1173;
assign n_2138 = x7 & n_1173;
assign n_2139 = x8 & n_1173;
assign n_2140 = x9 & n_1173;
assign n_2141 = x10 & n_1173;
assign n_2142 = x11 & n_1173;
assign n_2143 = x12 & n_1173;
assign n_2144 = x13 & n_1173;
assign n_2145 = x14 & n_1173;
assign n_2146 = x15 & n_1173;
assign n_2147 = x16 & n_1173;
assign n_2148 = x17 & n_1173;
assign n_2149 = x18 & n_1173;
assign n_2150 = x19 & n_1173;
assign n_2151 = x20 & n_1173;
assign n_2152 = x21 & n_1173;
assign n_2153 = x22 & n_1173;
assign n_2154 = x23 & n_1173;
assign n_2155 = x24 & n_1173;
assign n_2156 = x25 & n_1173;
assign n_2157 = x26 & n_1173;
assign n_2158 = x27 & n_1173;
assign n_2159 = x28 & n_1173;
assign n_2160 = x29 & n_1173;
assign n_2161 = x30 & n_1173;
assign n_2162 = n_475 ^ n_1205;
assign n_2163 = n_477 ^ n_1206;
assign n_2164 = n_478 ^ n_1207;
assign n_2165 = n_479 ^ n_1208;
assign n_2166 = n_480 ^ n_1209;
assign n_2167 = n_481 ^ n_1210;
assign n_2168 = n_482 ^ n_1211;
assign n_2169 = n_483 ^ n_1212;
assign n_2170 = n_484 ^ n_1213;
assign n_2171 = n_485 ^ n_1214;
assign n_2172 = n_486 ^ n_1215;
assign n_2173 = n_487 ^ n_1216;
assign n_2174 = n_488 ^ n_1217;
assign n_2175 = n_489 ^ n_1218;
assign n_2176 = n_490 ^ n_1219;
assign n_2177 = n_491 ^ n_1220;
assign n_2178 = n_492 ^ n_1221;
assign n_2179 = n_493 ^ n_1222;
assign n_2180 = n_494 ^ n_1223;
assign n_2181 = n_495 ^ n_1224;
assign n_2182 = n_496 ^ n_1225;
assign n_2183 = n_497 ^ n_1226;
assign n_2184 = n_498 ^ n_1227;
assign n_2185 = n_499 ^ n_1228;
assign n_2186 = n_500 ^ n_1229;
assign n_2187 = n_501 ^ n_1230;
assign n_2188 = n_502 ^ n_1231;
assign n_2189 = n_503 ^ n_1232;
assign n_2190 = n_504 ^ n_1233;
assign n_2191 = n_505 ^ n_1234;
assign n_2192 = n_1235 ^ n_804;
assign n_2193 = n_804 & n_1235;
assign n_2194 = ~x1 & n_1237;
assign n_2195 = ~x2 & n_1237;
assign n_2196 = ~x3 & n_1237;
assign n_2197 = ~x4 & n_1237;
assign n_2198 = ~x5 & n_1237;
assign n_2199 = ~x6 & n_1237;
assign n_2200 = ~x7 & n_1237;
assign n_2201 = ~x8 & n_1237;
assign n_2202 = ~x9 & n_1237;
assign n_2203 = ~x10 & n_1237;
assign n_2204 = ~x11 & n_1237;
assign n_2205 = ~x12 & n_1237;
assign n_2206 = ~x13 & n_1237;
assign n_2207 = ~x14 & n_1237;
assign n_2208 = ~x15 & n_1237;
assign n_2209 = ~x16 & n_1237;
assign n_2210 = ~x17 & n_1237;
assign n_2211 = ~x18 & n_1237;
assign n_2212 = ~x19 & n_1237;
assign n_2213 = ~x20 & n_1237;
assign n_2214 = ~x21 & n_1237;
assign n_2215 = ~x22 & n_1237;
assign n_2216 = ~x23 & n_1237;
assign n_2217 = ~x24 & n_1237;
assign n_2218 = ~x25 & n_1237;
assign n_2219 = ~x26 & n_1237;
assign n_2220 = ~x27 & n_1237;
assign n_2221 = ~x28 & n_1237;
assign n_2222 = ~x29 & n_1237;
assign n_2223 = ~x30 & n_1237;
assign n_2224 = n_1237 ^ n_476;
assign n_2225 = n_510 ^ n_1268;
assign n_2226 = n_512 ^ n_1269;
assign n_2227 = n_513 ^ n_1270;
assign n_2228 = n_514 ^ n_1271;
assign n_2229 = n_515 ^ n_1272;
assign n_2230 = n_516 ^ n_1273;
assign n_2231 = n_517 ^ n_1274;
assign n_2232 = n_518 ^ n_1275;
assign n_2233 = n_519 ^ n_1276;
assign n_2234 = n_520 ^ n_1277;
assign n_2235 = n_521 ^ n_1278;
assign n_2236 = n_522 ^ n_1279;
assign n_2237 = n_523 ^ n_1280;
assign n_2238 = n_524 ^ n_1281;
assign n_2239 = n_525 ^ n_1282;
assign n_2240 = n_526 ^ n_1283;
assign n_2241 = n_527 ^ n_1284;
assign n_2242 = n_528 ^ n_1285;
assign n_2243 = n_529 ^ n_1286;
assign n_2244 = n_530 ^ n_1287;
assign n_2245 = n_531 ^ n_1288;
assign n_2246 = n_532 ^ n_1289;
assign n_2247 = n_533 ^ n_1290;
assign n_2248 = n_534 ^ n_1291;
assign n_2249 = n_535 ^ n_1292;
assign n_2250 = n_536 ^ n_1293;
assign n_2251 = n_537 ^ n_1294;
assign n_2252 = n_538 ^ n_1295;
assign n_2253 = n_539 ^ n_1296;
assign n_2254 = n_540 ^ n_1297;
assign n_2255 = n_1298 ^ n_806;
assign n_2256 = n_806 & n_1298;
assign n_2257 = x1 & n_1300;
assign n_2258 = x2 & n_1300;
assign n_2259 = x3 & n_1300;
assign n_2260 = x4 & n_1300;
assign n_2261 = x5 & n_1300;
assign n_2262 = x6 & n_1300;
assign n_2263 = x7 & n_1300;
assign n_2264 = x8 & n_1300;
assign n_2265 = x9 & n_1300;
assign n_2266 = x10 & n_1300;
assign n_2267 = x11 & n_1300;
assign n_2268 = x12 & n_1300;
assign n_2269 = x13 & n_1300;
assign n_2270 = x14 & n_1300;
assign n_2271 = x15 & n_1300;
assign n_2272 = x16 & n_1300;
assign n_2273 = x17 & n_1300;
assign n_2274 = x18 & n_1300;
assign n_2275 = x19 & n_1300;
assign n_2276 = x20 & n_1300;
assign n_2277 = x21 & n_1300;
assign n_2278 = x22 & n_1300;
assign n_2279 = x23 & n_1300;
assign n_2280 = x24 & n_1300;
assign n_2281 = x25 & n_1300;
assign n_2282 = x26 & n_1300;
assign n_2283 = x27 & n_1300;
assign n_2284 = x28 & n_1300;
assign n_2285 = x29 & n_1300;
assign n_2286 = x30 & n_1300;
assign n_2287 = n_545 ^ n_1332;
assign n_2288 = n_547 ^ n_1333;
assign n_2289 = n_548 ^ n_1334;
assign n_2290 = n_549 ^ n_1335;
assign n_2291 = n_550 ^ n_1336;
assign n_2292 = n_551 ^ n_1337;
assign n_2293 = n_552 ^ n_1338;
assign n_2294 = n_553 ^ n_1339;
assign n_2295 = n_554 ^ n_1340;
assign n_2296 = n_555 ^ n_1341;
assign n_2297 = n_556 ^ n_1342;
assign n_2298 = n_557 ^ n_1343;
assign n_2299 = n_558 ^ n_1344;
assign n_2300 = n_559 ^ n_1345;
assign n_2301 = n_560 ^ n_1346;
assign n_2302 = n_561 ^ n_1347;
assign n_2303 = n_562 ^ n_1348;
assign n_2304 = n_563 ^ n_1349;
assign n_2305 = n_564 ^ n_1350;
assign n_2306 = n_565 ^ n_1351;
assign n_2307 = n_566 ^ n_1352;
assign n_2308 = n_567 ^ n_1353;
assign n_2309 = n_568 ^ n_1354;
assign n_2310 = n_569 ^ n_1355;
assign n_2311 = n_570 ^ n_1356;
assign n_2312 = n_571 ^ n_1357;
assign n_2313 = n_572 ^ n_1358;
assign n_2314 = n_573 ^ n_1359;
assign n_2315 = n_574 ^ n_1360;
assign n_2316 = n_575 ^ n_1361;
assign n_2317 = n_1362 ^ n_808;
assign n_2318 = n_808 & n_1362;
assign n_2319 = ~x1 & n_1364;
assign n_2320 = ~x2 & n_1364;
assign n_2321 = ~x3 & n_1364;
assign n_2322 = ~x4 & n_1364;
assign n_2323 = ~x5 & n_1364;
assign n_2324 = ~x6 & n_1364;
assign n_2325 = ~x7 & n_1364;
assign n_2326 = ~x8 & n_1364;
assign n_2327 = ~x9 & n_1364;
assign n_2328 = ~x10 & n_1364;
assign n_2329 = ~x11 & n_1364;
assign n_2330 = ~x12 & n_1364;
assign n_2331 = ~x13 & n_1364;
assign n_2332 = ~x14 & n_1364;
assign n_2333 = ~x15 & n_1364;
assign n_2334 = ~x16 & n_1364;
assign n_2335 = ~x17 & n_1364;
assign n_2336 = ~x18 & n_1364;
assign n_2337 = ~x19 & n_1364;
assign n_2338 = ~x20 & n_1364;
assign n_2339 = ~x21 & n_1364;
assign n_2340 = ~x22 & n_1364;
assign n_2341 = ~x23 & n_1364;
assign n_2342 = ~x24 & n_1364;
assign n_2343 = ~x25 & n_1364;
assign n_2344 = ~x26 & n_1364;
assign n_2345 = ~x27 & n_1364;
assign n_2346 = ~x28 & n_1364;
assign n_2347 = ~x29 & n_1364;
assign n_2348 = ~x30 & n_1364;
assign n_2349 = n_1364 ^ n_546;
assign n_2350 = n_581 ^ n_1396;
assign n_2351 = n_583 ^ n_1397;
assign n_2352 = n_584 ^ n_1398;
assign n_2353 = n_585 ^ n_1399;
assign n_2354 = n_586 ^ n_1400;
assign n_2355 = n_587 ^ n_1401;
assign n_2356 = n_588 ^ n_1402;
assign n_2357 = n_589 ^ n_1403;
assign n_2358 = n_590 ^ n_1404;
assign n_2359 = n_591 ^ n_1405;
assign n_2360 = n_592 ^ n_1406;
assign n_2361 = n_593 ^ n_1407;
assign n_2362 = n_594 ^ n_1408;
assign n_2363 = n_595 ^ n_1409;
assign n_2364 = n_596 ^ n_1410;
assign n_2365 = n_597 ^ n_1411;
assign n_2366 = n_598 ^ n_1412;
assign n_2367 = n_599 ^ n_1413;
assign n_2368 = n_600 ^ n_1414;
assign n_2369 = n_601 ^ n_1415;
assign n_2370 = n_602 ^ n_1416;
assign n_2371 = n_603 ^ n_1417;
assign n_2372 = n_604 ^ n_1418;
assign n_2373 = n_605 ^ n_1419;
assign n_2374 = n_606 ^ n_1420;
assign n_2375 = n_607 ^ n_1421;
assign n_2376 = n_608 ^ n_1422;
assign n_2377 = n_609 ^ n_1423;
assign n_2378 = n_610 ^ n_1424;
assign n_2379 = n_611 ^ n_1425;
assign n_2380 = x1 & n_1427;
assign n_2381 = x2 & n_1427;
assign n_2382 = x3 & n_1427;
assign n_2383 = x4 & n_1427;
assign n_2384 = x5 & n_1427;
assign n_2385 = x6 & n_1427;
assign n_2386 = x7 & n_1427;
assign n_2387 = x8 & n_1427;
assign n_2388 = x9 & n_1427;
assign n_2389 = x10 & n_1427;
assign n_2390 = x11 & n_1427;
assign n_2391 = x12 & n_1427;
assign n_2392 = x13 & n_1427;
assign n_2393 = x14 & n_1427;
assign n_2394 = x15 & n_1427;
assign n_2395 = x16 & n_1427;
assign n_2396 = x17 & n_1427;
assign n_2397 = x18 & n_1427;
assign n_2398 = x19 & n_1427;
assign n_2399 = x20 & n_1427;
assign n_2400 = x21 & n_1427;
assign n_2401 = x22 & n_1427;
assign n_2402 = x23 & n_1427;
assign n_2403 = x24 & n_1427;
assign n_2404 = x25 & n_1427;
assign n_2405 = x26 & n_1427;
assign n_2406 = x27 & n_1427;
assign n_2407 = x28 & n_1427;
assign n_2408 = x29 & n_1427;
assign n_2409 = x30 & n_1427;
assign n_2410 = n_113 ^ n_1458;
assign n_2411 = n_616 ^ n_1460;
assign n_2412 = n_618 ^ n_1461;
assign n_2413 = n_619 ^ n_1462;
assign n_2414 = n_620 ^ n_1463;
assign n_2415 = n_621 ^ n_1464;
assign n_2416 = n_622 ^ n_1465;
assign n_2417 = n_623 ^ n_1466;
assign n_2418 = n_624 ^ n_1467;
assign n_2419 = n_625 ^ n_1468;
assign n_2420 = n_626 ^ n_1469;
assign n_2421 = n_627 ^ n_1470;
assign n_2422 = n_628 ^ n_1471;
assign n_2423 = n_629 ^ n_1472;
assign n_2424 = n_630 ^ n_1473;
assign n_2425 = n_631 ^ n_1474;
assign n_2426 = n_632 ^ n_1475;
assign n_2427 = n_633 ^ n_1476;
assign n_2428 = n_634 ^ n_1477;
assign n_2429 = n_635 ^ n_1478;
assign n_2430 = n_636 ^ n_1479;
assign n_2431 = n_637 ^ n_1480;
assign n_2432 = n_638 ^ n_1481;
assign n_2433 = n_639 ^ n_1482;
assign n_2434 = n_640 ^ n_1483;
assign n_2435 = n_641 ^ n_1484;
assign n_2436 = n_642 ^ n_1485;
assign n_2437 = n_643 ^ n_1486;
assign n_2438 = n_644 ^ n_1487;
assign n_2439 = n_645 ^ n_1488;
assign n_2440 = n_646 ^ n_1489;
assign n_2441 = x1 & n_1491;
assign n_2442 = x2 & n_1491;
assign n_2443 = x3 & n_1491;
assign n_2444 = x4 & n_1491;
assign n_2445 = x5 & n_1491;
assign n_2446 = x6 & n_1491;
assign n_2447 = x7 & n_1491;
assign n_2448 = x8 & n_1491;
assign n_2449 = x9 & n_1491;
assign n_2450 = x10 & n_1491;
assign n_2451 = x11 & n_1491;
assign n_2452 = x12 & n_1491;
assign n_2453 = x13 & n_1491;
assign n_2454 = x14 & n_1491;
assign n_2455 = x15 & n_1491;
assign n_2456 = x16 & n_1491;
assign n_2457 = x17 & n_1491;
assign n_2458 = x18 & n_1491;
assign n_2459 = x19 & n_1491;
assign n_2460 = x20 & n_1491;
assign n_2461 = x21 & n_1491;
assign n_2462 = x22 & n_1491;
assign n_2463 = x23 & n_1491;
assign n_2464 = x24 & n_1491;
assign n_2465 = x25 & n_1491;
assign n_2466 = x26 & n_1491;
assign n_2467 = x27 & n_1491;
assign n_2468 = x28 & n_1491;
assign n_2469 = x29 & n_1491;
assign n_2470 = x30 & n_1491;
assign n_2471 = n_651 ^ n_1524;
assign n_2472 = n_653 ^ n_1525;
assign n_2473 = n_654 ^ n_1526;
assign n_2474 = n_655 ^ n_1527;
assign n_2475 = n_656 ^ n_1528;
assign n_2476 = n_657 ^ n_1529;
assign n_2477 = n_658 ^ n_1530;
assign n_2478 = n_659 ^ n_1531;
assign n_2479 = n_660 ^ n_1532;
assign n_2480 = n_661 ^ n_1533;
assign n_2481 = n_662 ^ n_1534;
assign n_2482 = n_663 ^ n_1535;
assign n_2483 = n_664 ^ n_1536;
assign n_2484 = n_665 ^ n_1537;
assign n_2485 = n_666 ^ n_1538;
assign n_2486 = n_667 ^ n_1539;
assign n_2487 = n_668 ^ n_1540;
assign n_2488 = n_669 ^ n_1541;
assign n_2489 = n_670 ^ n_1542;
assign n_2490 = n_671 ^ n_1543;
assign n_2491 = n_672 ^ n_1544;
assign n_2492 = n_673 ^ n_1545;
assign n_2493 = n_674 ^ n_1546;
assign n_2494 = n_675 ^ n_1547;
assign n_2495 = n_676 ^ n_1548;
assign n_2496 = n_677 ^ n_1549;
assign n_2497 = n_678 ^ n_1550;
assign n_2498 = n_679 ^ n_1551;
assign n_2499 = n_680 ^ n_1552;
assign n_2500 = n_681 ^ n_1553;
assign n_2501 = x1 & n_1555;
assign n_2502 = x2 & n_1555;
assign n_2503 = x3 & n_1555;
assign n_2504 = x4 & n_1555;
assign n_2505 = x5 & n_1555;
assign n_2506 = x6 & n_1555;
assign n_2507 = x7 & n_1555;
assign n_2508 = x8 & n_1555;
assign n_2509 = x9 & n_1555;
assign n_2510 = x10 & n_1555;
assign n_2511 = x11 & n_1555;
assign n_2512 = x12 & n_1555;
assign n_2513 = x13 & n_1555;
assign n_2514 = x14 & n_1555;
assign n_2515 = x15 & n_1555;
assign n_2516 = x16 & n_1555;
assign n_2517 = x17 & n_1555;
assign n_2518 = x18 & n_1555;
assign n_2519 = x19 & n_1555;
assign n_2520 = x20 & n_1555;
assign n_2521 = x21 & n_1555;
assign n_2522 = x22 & n_1555;
assign n_2523 = x23 & n_1555;
assign n_2524 = x24 & n_1555;
assign n_2525 = x25 & n_1555;
assign n_2526 = x26 & n_1555;
assign n_2527 = x27 & n_1555;
assign n_2528 = x28 & n_1555;
assign n_2529 = x29 & n_1555;
assign n_2530 = x30 & n_1555;
assign n_2531 = n_116 ^ n_1586;
assign n_2532 = n_685 ^ n_1587;
assign n_2533 = n_687 ^ n_1588;
assign n_2534 = n_688 ^ n_1589;
assign n_2535 = n_689 ^ n_1590;
assign n_2536 = n_690 ^ n_1591;
assign n_2537 = n_691 ^ n_1592;
assign n_2538 = n_692 ^ n_1593;
assign n_2539 = n_693 ^ n_1594;
assign n_2540 = n_694 ^ n_1595;
assign n_2541 = n_695 ^ n_1596;
assign n_2542 = n_696 ^ n_1597;
assign n_2543 = n_697 ^ n_1598;
assign n_2544 = n_698 ^ n_1599;
assign n_2545 = n_699 ^ n_1600;
assign n_2546 = n_700 ^ n_1601;
assign n_2547 = n_701 ^ n_1602;
assign n_2548 = n_702 ^ n_1603;
assign n_2549 = n_703 ^ n_1604;
assign n_2550 = n_704 ^ n_1605;
assign n_2551 = n_705 ^ n_1606;
assign n_2552 = n_706 ^ n_1607;
assign n_2553 = n_707 ^ n_1608;
assign n_2554 = n_708 ^ n_1609;
assign n_2555 = n_709 ^ n_1610;
assign n_2556 = n_710 ^ n_1611;
assign n_2557 = n_711 ^ n_1612;
assign n_2558 = n_712 ^ n_1613;
assign n_2559 = n_713 ^ n_1614;
assign n_2560 = n_714 ^ n_1615;
assign n_2561 = n_715 ^ n_1616;
assign n_2562 = ~x1 & n_1619;
assign n_2563 = ~x2 & n_1619;
assign n_2564 = ~x3 & n_1619;
assign n_2565 = ~x4 & n_1619;
assign n_2566 = ~x5 & n_1619;
assign n_2567 = ~x6 & n_1619;
assign n_2568 = ~x7 & n_1619;
assign n_2569 = ~x8 & n_1619;
assign n_2570 = ~x9 & n_1619;
assign n_2571 = ~x10 & n_1619;
assign n_2572 = ~x11 & n_1619;
assign n_2573 = ~x12 & n_1619;
assign n_2574 = ~x13 & n_1619;
assign n_2575 = ~x14 & n_1619;
assign n_2576 = ~x15 & n_1619;
assign n_2577 = ~x16 & n_1619;
assign n_2578 = ~x17 & n_1619;
assign n_2579 = ~x18 & n_1619;
assign n_2580 = ~x19 & n_1619;
assign n_2581 = ~x20 & n_1619;
assign n_2582 = ~x21 & n_1619;
assign n_2583 = ~x22 & n_1619;
assign n_2584 = ~x23 & n_1619;
assign n_2585 = ~x24 & n_1619;
assign n_2586 = ~x25 & n_1619;
assign n_2587 = ~x26 & n_1619;
assign n_2588 = ~x27 & n_1619;
assign n_2589 = ~x28 & n_1619;
assign n_2590 = ~x29 & n_1619;
assign n_2591 = ~x30 & n_1619;
assign n_2592 = n_1619 ^ n_686;
assign n_2593 = n_720 ^ n_1650;
assign n_2594 = n_722 ^ n_1651;
assign n_2595 = n_723 ^ n_1652;
assign n_2596 = n_724 ^ n_1653;
assign n_2597 = n_725 ^ n_1654;
assign n_2598 = n_726 ^ n_1655;
assign n_2599 = n_727 ^ n_1656;
assign n_2600 = n_728 ^ n_1657;
assign n_2601 = n_729 ^ n_1658;
assign n_2602 = n_730 ^ n_1659;
assign n_2603 = n_731 ^ n_1660;
assign n_2604 = n_732 ^ n_1661;
assign n_2605 = n_733 ^ n_1662;
assign n_2606 = n_734 ^ n_1663;
assign n_2607 = n_735 ^ n_1664;
assign n_2608 = n_736 ^ n_1665;
assign n_2609 = n_737 ^ n_1666;
assign n_2610 = n_738 ^ n_1667;
assign n_2611 = n_739 ^ n_1668;
assign n_2612 = n_740 ^ n_1669;
assign n_2613 = n_741 ^ n_1670;
assign n_2614 = n_742 ^ n_1671;
assign n_2615 = n_743 ^ n_1672;
assign n_2616 = n_744 ^ n_1673;
assign n_2617 = n_745 ^ n_1674;
assign n_2618 = n_746 ^ n_1675;
assign n_2619 = n_747 ^ n_1676;
assign n_2620 = n_748 ^ n_1677;
assign n_2621 = n_749 ^ n_1678;
assign n_2622 = n_750 ^ n_1679;
assign n_2623 = n_1680 ^ n_818;
assign n_2624 = n_818 & n_1680;
assign n_2625 = x1 & n_1682;
assign n_2626 = x2 & n_1682;
assign n_2627 = x3 & n_1682;
assign n_2628 = x4 & n_1682;
assign n_2629 = x5 & n_1682;
assign n_2630 = x6 & n_1682;
assign n_2631 = x7 & n_1682;
assign n_2632 = x8 & n_1682;
assign n_2633 = x9 & n_1682;
assign n_2634 = x10 & n_1682;
assign n_2635 = x11 & n_1682;
assign n_2636 = x12 & n_1682;
assign n_2637 = x13 & n_1682;
assign n_2638 = x14 & n_1682;
assign n_2639 = x15 & n_1682;
assign n_2640 = x16 & n_1682;
assign n_2641 = x17 & n_1682;
assign n_2642 = x18 & n_1682;
assign n_2643 = x19 & n_1682;
assign n_2644 = x20 & n_1682;
assign n_2645 = x21 & n_1682;
assign n_2646 = x22 & n_1682;
assign n_2647 = x23 & n_1682;
assign n_2648 = x24 & n_1682;
assign n_2649 = x25 & n_1682;
assign n_2650 = x26 & n_1682;
assign n_2651 = x27 & n_1682;
assign n_2652 = x28 & n_1682;
assign n_2653 = x29 & n_1682;
assign n_2654 = x30 & n_1682;
assign n_2655 = n_1712 ^ n_122;
assign n_2656 = n_120 ^ n_1713;
assign n_2657 = n_755 ^ n_1714;
assign n_2658 = n_757 ^ n_1715;
assign n_2659 = n_758 ^ n_1716;
assign n_2660 = n_759 ^ n_1717;
assign n_2661 = n_760 ^ n_1718;
assign n_2662 = n_761 ^ n_1719;
assign n_2663 = n_762 ^ n_1720;
assign n_2664 = n_763 ^ n_1721;
assign n_2665 = n_764 ^ n_1722;
assign n_2666 = n_765 ^ n_1723;
assign n_2667 = n_766 ^ n_1724;
assign n_2668 = n_767 ^ n_1725;
assign n_2669 = n_768 ^ n_1726;
assign n_2670 = n_769 ^ n_1727;
assign n_2671 = n_770 ^ n_1728;
assign n_2672 = n_771 ^ n_1729;
assign n_2673 = n_772 ^ n_1730;
assign n_2674 = n_773 ^ n_1731;
assign n_2675 = n_774 ^ n_1732;
assign n_2676 = n_775 ^ n_1733;
assign n_2677 = n_776 ^ n_1734;
assign n_2678 = n_777 ^ n_1735;
assign n_2679 = n_778 ^ n_1736;
assign n_2680 = n_779 ^ n_1737;
assign n_2681 = n_780 ^ n_1738;
assign n_2682 = n_781 ^ n_1739;
assign n_2683 = n_782 ^ n_1740;
assign n_2684 = n_783 ^ n_1741;
assign n_2685 = n_784 ^ n_1742;
assign n_2686 = n_785 ^ n_1743;
assign n_2687 = n_1744 ^ n_820;
assign n_2688 = n_820 & n_1744;
assign n_2689 = x0 & n_1746;
assign n_2690 = x1 & n_1746;
assign n_2691 = x2 & n_1746;
assign n_2692 = x3 & n_1746;
assign n_2693 = x4 & n_1746;
assign n_2694 = x5 & n_1746;
assign n_2695 = x6 & n_1746;
assign n_2696 = x7 & n_1746;
assign n_2697 = x8 & n_1746;
assign n_2698 = x9 & n_1746;
assign n_2699 = x10 & n_1746;
assign n_2700 = x11 & n_1746;
assign n_2701 = x12 & n_1746;
assign n_2702 = x13 & n_1746;
assign n_2703 = x14 & n_1746;
assign n_2704 = x15 & n_1746;
assign n_2705 = x16 & n_1746;
assign n_2706 = x17 & n_1746;
assign n_2707 = x18 & n_1746;
assign n_2708 = x19 & n_1746;
assign n_2709 = x20 & n_1746;
assign n_2710 = x21 & n_1746;
assign n_2711 = x22 & n_1746;
assign n_2712 = x23 & n_1746;
assign n_2713 = x24 & n_1746;
assign n_2714 = x25 & n_1746;
assign n_2715 = x26 & n_1746;
assign n_2716 = x27 & n_1746;
assign n_2717 = x28 & n_1746;
assign n_2718 = x29 & n_1746;
assign n_2719 = x30 & n_1746;
assign n_2720 = n_1777 ^ n_123;
assign n_2721 = x63 & n_1778;
assign y1 = n_1779;
assign n_2722 = n_158 ^ n_1780;
assign n_2723 = n_1781 ^ n_1780;
assign n_2724 = n_297 ^ n_1792;
assign n_2725 = n_853 ^ n_1822;
assign n_2726 = n_855 ^ n_1823;
assign n_2727 = n_856 ^ n_1824;
assign n_2728 = n_857 ^ n_1825;
assign n_2729 = n_858 ^ n_1826;
assign n_2730 = n_859 ^ n_1827;
assign n_2731 = n_860 ^ n_1828;
assign n_2732 = n_861 ^ n_1829;
assign n_2733 = n_862 ^ n_1830;
assign n_2734 = n_863 ^ n_1831;
assign n_2735 = n_864 ^ n_1832;
assign n_2736 = n_865 ^ n_1833;
assign n_2737 = n_866 ^ n_1834;
assign n_2738 = n_867 ^ n_1835;
assign n_2739 = n_868 ^ n_1836;
assign n_2740 = n_869 ^ n_1837;
assign n_2741 = n_870 ^ n_1838;
assign n_2742 = n_871 ^ n_1839;
assign n_2743 = n_872 ^ n_1840;
assign n_2744 = n_873 ^ n_1841;
assign n_2745 = n_874 ^ n_1842;
assign n_2746 = n_875 ^ n_1843;
assign n_2747 = n_876 ^ n_1844;
assign n_2748 = n_877 ^ n_1845;
assign n_2749 = n_878 ^ n_1846;
assign n_2750 = n_879 ^ n_1847;
assign n_2751 = n_880 ^ n_1848;
assign n_2752 = n_881 ^ n_1849;
assign n_2753 = n_882 ^ n_1850;
assign n_2754 = n_883 ^ n_1851;
assign n_2755 = n_332 ^ n_1853;
assign n_2756 = n_917 ^ n_1885;
assign n_2757 = n_919 ^ n_1886;
assign n_2758 = n_920 ^ n_1887;
assign n_2759 = n_921 ^ n_1888;
assign n_2760 = n_922 ^ n_1889;
assign n_2761 = n_923 ^ n_1890;
assign n_2762 = n_924 ^ n_1891;
assign n_2763 = n_925 ^ n_1892;
assign n_2764 = n_926 ^ n_1893;
assign n_2765 = n_927 ^ n_1894;
assign n_2766 = n_928 ^ n_1895;
assign n_2767 = n_929 ^ n_1896;
assign n_2768 = n_930 ^ n_1897;
assign n_2769 = n_931 ^ n_1898;
assign n_2770 = n_932 ^ n_1899;
assign n_2771 = n_933 ^ n_1900;
assign n_2772 = n_934 ^ n_1901;
assign n_2773 = n_935 ^ n_1902;
assign n_2774 = n_936 ^ n_1903;
assign n_2775 = n_937 ^ n_1904;
assign n_2776 = n_938 ^ n_1905;
assign n_2777 = n_939 ^ n_1906;
assign n_2778 = n_940 ^ n_1907;
assign n_2779 = n_941 ^ n_1908;
assign n_2780 = n_942 ^ n_1909;
assign n_2781 = n_943 ^ n_1910;
assign n_2782 = n_944 ^ n_1911;
assign n_2783 = n_945 ^ n_1912;
assign n_2784 = n_946 ^ n_1913;
assign n_2785 = n_947 ^ n_1914;
assign n_2786 = n_367 ^ n_1918;
assign n_2787 = n_981 ^ n_1948;
assign n_2788 = n_983 ^ n_1949;
assign n_2789 = n_984 ^ n_1950;
assign n_2790 = n_985 ^ n_1951;
assign n_2791 = n_986 ^ n_1952;
assign n_2792 = n_987 ^ n_1953;
assign n_2793 = n_988 ^ n_1954;
assign n_2794 = n_989 ^ n_1955;
assign n_2795 = n_990 ^ n_1956;
assign n_2796 = n_991 ^ n_1957;
assign n_2797 = n_992 ^ n_1958;
assign n_2798 = n_993 ^ n_1959;
assign n_2799 = n_994 ^ n_1960;
assign n_2800 = n_995 ^ n_1961;
assign n_2801 = n_996 ^ n_1962;
assign n_2802 = n_997 ^ n_1963;
assign n_2803 = n_998 ^ n_1964;
assign n_2804 = n_999 ^ n_1965;
assign n_2805 = n_1000 ^ n_1966;
assign n_2806 = n_1001 ^ n_1967;
assign n_2807 = n_1002 ^ n_1968;
assign n_2808 = n_1003 ^ n_1969;
assign n_2809 = n_1004 ^ n_1970;
assign n_2810 = n_1005 ^ n_1971;
assign n_2811 = n_1006 ^ n_1972;
assign n_2812 = n_1007 ^ n_1973;
assign n_2813 = n_1008 ^ n_1974;
assign n_2814 = n_1009 ^ n_1975;
assign n_2815 = n_1010 ^ n_1976;
assign n_2816 = n_1011 ^ n_1977;
assign n_2817 = n_402 ^ n_1978;
assign n_2818 = n_1045 ^ n_2008;
assign n_2819 = n_1047 ^ n_2009;
assign n_2820 = n_1048 ^ n_2010;
assign n_2821 = n_1049 ^ n_2011;
assign n_2822 = n_1050 ^ n_2012;
assign n_2823 = n_1051 ^ n_2013;
assign n_2824 = n_1052 ^ n_2014;
assign n_2825 = n_1053 ^ n_2015;
assign n_2826 = n_1054 ^ n_2016;
assign n_2827 = n_1055 ^ n_2017;
assign n_2828 = n_1056 ^ n_2018;
assign n_2829 = n_1057 ^ n_2019;
assign n_2830 = n_1058 ^ n_2020;
assign n_2831 = n_1059 ^ n_2021;
assign n_2832 = n_1060 ^ n_2022;
assign n_2833 = n_1061 ^ n_2023;
assign n_2834 = n_1062 ^ n_2024;
assign n_2835 = n_1063 ^ n_2025;
assign n_2836 = n_1064 ^ n_2026;
assign n_2837 = n_1065 ^ n_2027;
assign n_2838 = n_1066 ^ n_2028;
assign n_2839 = n_1067 ^ n_2029;
assign n_2840 = n_1068 ^ n_2030;
assign n_2841 = n_1069 ^ n_2031;
assign n_2842 = n_1070 ^ n_2032;
assign n_2843 = n_1071 ^ n_2033;
assign n_2844 = n_1072 ^ n_2034;
assign n_2845 = n_1073 ^ n_2035;
assign n_2846 = n_1074 ^ n_2036;
assign n_2847 = n_1075 ^ n_2037;
assign n_2848 = n_437 ^ n_2038;
assign n_2849 = n_1109 ^ n_2068;
assign n_2850 = n_1111 ^ n_2069;
assign n_2851 = n_1112 ^ n_2070;
assign n_2852 = n_1113 ^ n_2071;
assign n_2853 = n_1114 ^ n_2072;
assign n_2854 = n_1115 ^ n_2073;
assign n_2855 = n_1116 ^ n_2074;
assign n_2856 = n_1117 ^ n_2075;
assign n_2857 = n_1118 ^ n_2076;
assign n_2858 = n_1119 ^ n_2077;
assign n_2859 = n_1120 ^ n_2078;
assign n_2860 = n_1121 ^ n_2079;
assign n_2861 = n_1122 ^ n_2080;
assign n_2862 = n_1123 ^ n_2081;
assign n_2863 = n_1124 ^ n_2082;
assign n_2864 = n_1125 ^ n_2083;
assign n_2865 = n_1126 ^ n_2084;
assign n_2866 = n_1127 ^ n_2085;
assign n_2867 = n_1128 ^ n_2086;
assign n_2868 = n_1129 ^ n_2087;
assign n_2869 = n_1130 ^ n_2088;
assign n_2870 = n_1131 ^ n_2089;
assign n_2871 = n_1132 ^ n_2090;
assign n_2872 = n_1133 ^ n_2091;
assign n_2873 = n_1134 ^ n_2092;
assign n_2874 = n_1135 ^ n_2093;
assign n_2875 = n_1136 ^ n_2094;
assign n_2876 = n_1137 ^ n_2095;
assign n_2877 = n_1138 ^ n_2096;
assign n_2878 = n_1139 ^ n_2097;
assign n_2879 = n_472 ^ n_2102;
assign n_2880 = n_1172 ^ n_2132;
assign n_2881 = n_1174 ^ n_2133;
assign n_2882 = n_1175 ^ n_2134;
assign n_2883 = n_1176 ^ n_2135;
assign n_2884 = n_1177 ^ n_2136;
assign n_2885 = n_1178 ^ n_2137;
assign n_2886 = n_1179 ^ n_2138;
assign n_2887 = n_1180 ^ n_2139;
assign n_2888 = n_1181 ^ n_2140;
assign n_2889 = n_1182 ^ n_2141;
assign n_2890 = n_1183 ^ n_2142;
assign n_2891 = n_1184 ^ n_2143;
assign n_2892 = n_1185 ^ n_2144;
assign n_2893 = n_1186 ^ n_2145;
assign n_2894 = n_1187 ^ n_2146;
assign n_2895 = n_1188 ^ n_2147;
assign n_2896 = n_1189 ^ n_2148;
assign n_2897 = n_1190 ^ n_2149;
assign n_2898 = n_1191 ^ n_2150;
assign n_2899 = n_1192 ^ n_2151;
assign n_2900 = n_1193 ^ n_2152;
assign n_2901 = n_1194 ^ n_2153;
assign n_2902 = n_1195 ^ n_2154;
assign n_2903 = n_1196 ^ n_2155;
assign n_2904 = n_1197 ^ n_2156;
assign n_2905 = n_1198 ^ n_2157;
assign n_2906 = n_1199 ^ n_2158;
assign n_2907 = n_1200 ^ n_2159;
assign n_2908 = n_1201 ^ n_2160;
assign n_2909 = n_1202 ^ n_2161;
assign n_2910 = n_507 ^ n_2162;
assign n_2911 = n_1236 ^ n_2194;
assign n_2912 = n_1238 ^ n_2195;
assign n_2913 = n_1239 ^ n_2196;
assign n_2914 = n_1240 ^ n_2197;
assign n_2915 = n_1241 ^ n_2198;
assign n_2916 = n_1242 ^ n_2199;
assign n_2917 = n_1243 ^ n_2200;
assign n_2918 = n_1244 ^ n_2201;
assign n_2919 = n_1245 ^ n_2202;
assign n_2920 = n_1246 ^ n_2203;
assign n_2921 = n_1247 ^ n_2204;
assign n_2922 = n_1248 ^ n_2205;
assign n_2923 = n_1249 ^ n_2206;
assign n_2924 = n_1250 ^ n_2207;
assign n_2925 = n_1251 ^ n_2208;
assign n_2926 = n_1252 ^ n_2209;
assign n_2927 = n_1253 ^ n_2210;
assign n_2928 = n_1254 ^ n_2211;
assign n_2929 = n_1255 ^ n_2212;
assign n_2930 = n_1256 ^ n_2213;
assign n_2931 = n_1257 ^ n_2214;
assign n_2932 = n_1258 ^ n_2215;
assign n_2933 = n_1259 ^ n_2216;
assign n_2934 = n_1260 ^ n_2217;
assign n_2935 = n_1261 ^ n_2218;
assign n_2936 = n_1262 ^ n_2219;
assign n_2937 = n_1263 ^ n_2220;
assign n_2938 = n_1264 ^ n_2221;
assign n_2939 = n_1265 ^ n_2222;
assign n_2940 = n_1266 ^ n_2223;
assign n_2941 = n_542 ^ n_2225;
assign n_2942 = n_1299 ^ n_2257;
assign n_2943 = n_1301 ^ n_2258;
assign n_2944 = n_1302 ^ n_2259;
assign n_2945 = n_1303 ^ n_2260;
assign n_2946 = n_1304 ^ n_2261;
assign n_2947 = n_1305 ^ n_2262;
assign n_2948 = n_1306 ^ n_2263;
assign n_2949 = n_1307 ^ n_2264;
assign n_2950 = n_1308 ^ n_2265;
assign n_2951 = n_1309 ^ n_2266;
assign n_2952 = n_1310 ^ n_2267;
assign n_2953 = n_1311 ^ n_2268;
assign n_2954 = n_1312 ^ n_2269;
assign n_2955 = n_1313 ^ n_2270;
assign n_2956 = n_1314 ^ n_2271;
assign n_2957 = n_1315 ^ n_2272;
assign n_2958 = n_1316 ^ n_2273;
assign n_2959 = n_1317 ^ n_2274;
assign n_2960 = n_1318 ^ n_2275;
assign n_2961 = n_1319 ^ n_2276;
assign n_2962 = n_1320 ^ n_2277;
assign n_2963 = n_1321 ^ n_2278;
assign n_2964 = n_1322 ^ n_2279;
assign n_2965 = n_1323 ^ n_2280;
assign n_2966 = n_1324 ^ n_2281;
assign n_2967 = n_1325 ^ n_2282;
assign n_2968 = n_1326 ^ n_2283;
assign n_2969 = n_1327 ^ n_2284;
assign n_2970 = n_1328 ^ n_2285;
assign n_2971 = n_1329 ^ n_2286;
assign n_2972 = n_577 ^ n_2287;
assign n_2973 = n_1363 ^ n_2319;
assign n_2974 = n_1365 ^ n_2320;
assign n_2975 = n_1366 ^ n_2321;
assign n_2976 = n_1367 ^ n_2322;
assign n_2977 = n_1368 ^ n_2323;
assign n_2978 = n_1369 ^ n_2324;
assign n_2979 = n_1370 ^ n_2325;
assign n_2980 = n_1371 ^ n_2326;
assign n_2981 = n_1372 ^ n_2327;
assign n_2982 = n_1373 ^ n_2328;
assign n_2983 = n_1374 ^ n_2329;
assign n_2984 = n_1375 ^ n_2330;
assign n_2985 = n_1376 ^ n_2331;
assign n_2986 = n_1377 ^ n_2332;
assign n_2987 = n_1378 ^ n_2333;
assign n_2988 = n_1379 ^ n_2334;
assign n_2989 = n_1380 ^ n_2335;
assign n_2990 = n_1381 ^ n_2336;
assign n_2991 = n_1382 ^ n_2337;
assign n_2992 = n_1383 ^ n_2338;
assign n_2993 = n_1384 ^ n_2339;
assign n_2994 = n_1385 ^ n_2340;
assign n_2995 = n_1386 ^ n_2341;
assign n_2996 = n_1387 ^ n_2342;
assign n_2997 = n_1388 ^ n_2343;
assign n_2998 = n_1389 ^ n_2344;
assign n_2999 = n_1390 ^ n_2345;
assign n_3000 = n_1391 ^ n_2346;
assign n_3001 = n_1392 ^ n_2347;
assign n_3002 = n_1393 ^ n_2348;
assign n_3003 = n_612 ^ n_2350;
assign n_3004 = n_1426 ^ n_2380;
assign n_3005 = n_1428 ^ n_2381;
assign n_3006 = n_1429 ^ n_2382;
assign n_3007 = n_1430 ^ n_2383;
assign n_3008 = n_1431 ^ n_2384;
assign n_3009 = n_1432 ^ n_2385;
assign n_3010 = n_1433 ^ n_2386;
assign n_3011 = n_1434 ^ n_2387;
assign n_3012 = n_1435 ^ n_2388;
assign n_3013 = n_1436 ^ n_2389;
assign n_3014 = n_1437 ^ n_2390;
assign n_3015 = n_1438 ^ n_2391;
assign n_3016 = n_1439 ^ n_2392;
assign n_3017 = n_1440 ^ n_2393;
assign n_3018 = n_1441 ^ n_2394;
assign n_3019 = n_1442 ^ n_2395;
assign n_3020 = n_1443 ^ n_2396;
assign n_3021 = n_1444 ^ n_2397;
assign n_3022 = n_1445 ^ n_2398;
assign n_3023 = n_1446 ^ n_2399;
assign n_3024 = n_1447 ^ n_2400;
assign n_3025 = n_1448 ^ n_2401;
assign n_3026 = n_1449 ^ n_2402;
assign n_3027 = n_1450 ^ n_2403;
assign n_3028 = n_1451 ^ n_2404;
assign n_3029 = n_1452 ^ n_2405;
assign n_3030 = n_1453 ^ n_2406;
assign n_3031 = n_1454 ^ n_2407;
assign n_3032 = n_1455 ^ n_2408;
assign n_3033 = n_1456 ^ n_2409;
assign n_3034 = n_647 ^ n_2411;
assign n_3035 = n_1490 ^ n_2441;
assign n_3036 = n_1492 ^ n_2442;
assign n_3037 = n_1493 ^ n_2443;
assign n_3038 = n_1494 ^ n_2444;
assign n_3039 = n_1495 ^ n_2445;
assign n_3040 = n_1496 ^ n_2446;
assign n_3041 = n_1497 ^ n_2447;
assign n_3042 = n_1498 ^ n_2448;
assign n_3043 = n_1499 ^ n_2449;
assign n_3044 = n_1500 ^ n_2450;
assign n_3045 = n_1501 ^ n_2451;
assign n_3046 = n_1502 ^ n_2452;
assign n_3047 = n_1503 ^ n_2453;
assign n_3048 = n_1504 ^ n_2454;
assign n_3049 = n_1505 ^ n_2455;
assign n_3050 = n_1506 ^ n_2456;
assign n_3051 = n_1507 ^ n_2457;
assign n_3052 = n_1508 ^ n_2458;
assign n_3053 = n_1509 ^ n_2459;
assign n_3054 = n_1510 ^ n_2460;
assign n_3055 = n_1511 ^ n_2461;
assign n_3056 = n_1512 ^ n_2462;
assign n_3057 = n_1513 ^ n_2463;
assign n_3058 = n_1514 ^ n_2464;
assign n_3059 = n_1515 ^ n_2465;
assign n_3060 = n_1516 ^ n_2466;
assign n_3061 = n_1517 ^ n_2467;
assign n_3062 = n_1518 ^ n_2468;
assign n_3063 = n_1519 ^ n_2469;
assign n_3064 = n_1520 ^ n_2470;
assign n_3065 = n_682 ^ n_2471;
assign n_3066 = n_1554 ^ n_2501;
assign n_3067 = n_1556 ^ n_2502;
assign n_3068 = n_1557 ^ n_2503;
assign n_3069 = n_1558 ^ n_2504;
assign n_3070 = n_1559 ^ n_2505;
assign n_3071 = n_1560 ^ n_2506;
assign n_3072 = n_1561 ^ n_2507;
assign n_3073 = n_1562 ^ n_2508;
assign n_3074 = n_1563 ^ n_2509;
assign n_3075 = n_1564 ^ n_2510;
assign n_3076 = n_1565 ^ n_2511;
assign n_3077 = n_1566 ^ n_2512;
assign n_3078 = n_1567 ^ n_2513;
assign n_3079 = n_1568 ^ n_2514;
assign n_3080 = n_1569 ^ n_2515;
assign n_3081 = n_1570 ^ n_2516;
assign n_3082 = n_1571 ^ n_2517;
assign n_3083 = n_1572 ^ n_2518;
assign n_3084 = n_1573 ^ n_2519;
assign n_3085 = n_1574 ^ n_2520;
assign n_3086 = n_1575 ^ n_2521;
assign n_3087 = n_1576 ^ n_2522;
assign n_3088 = n_1577 ^ n_2523;
assign n_3089 = n_1578 ^ n_2524;
assign n_3090 = n_1579 ^ n_2525;
assign n_3091 = n_1580 ^ n_2526;
assign n_3092 = n_1581 ^ n_2527;
assign n_3093 = n_1582 ^ n_2528;
assign n_3094 = n_1583 ^ n_2529;
assign n_3095 = n_1584 ^ n_2530;
assign n_3096 = n_717 ^ n_2532;
assign n_3097 = n_1618 ^ n_2562;
assign n_3098 = n_1620 ^ n_2563;
assign n_3099 = n_1621 ^ n_2564;
assign n_3100 = n_1622 ^ n_2565;
assign n_3101 = n_1623 ^ n_2566;
assign n_3102 = n_1624 ^ n_2567;
assign n_3103 = n_1625 ^ n_2568;
assign n_3104 = n_1626 ^ n_2569;
assign n_3105 = n_1627 ^ n_2570;
assign n_3106 = n_1628 ^ n_2571;
assign n_3107 = n_1629 ^ n_2572;
assign n_3108 = n_1630 ^ n_2573;
assign n_3109 = n_1631 ^ n_2574;
assign n_3110 = n_1632 ^ n_2575;
assign n_3111 = n_1633 ^ n_2576;
assign n_3112 = n_1634 ^ n_2577;
assign n_3113 = n_1635 ^ n_2578;
assign n_3114 = n_1636 ^ n_2579;
assign n_3115 = n_1637 ^ n_2580;
assign n_3116 = n_1638 ^ n_2581;
assign n_3117 = n_1639 ^ n_2582;
assign n_3118 = n_1640 ^ n_2583;
assign n_3119 = n_1641 ^ n_2584;
assign n_3120 = n_1642 ^ n_2585;
assign n_3121 = n_1643 ^ n_2586;
assign n_3122 = n_1644 ^ n_2587;
assign n_3123 = n_1645 ^ n_2588;
assign n_3124 = n_1646 ^ n_2589;
assign n_3125 = n_1647 ^ n_2590;
assign n_3126 = n_1648 ^ n_2591;
assign n_3127 = n_2592 ^ n_119;
assign n_3128 = n_752 ^ n_2593;
assign n_3129 = n_1681 ^ n_2625;
assign n_3130 = n_1683 ^ n_2626;
assign n_3131 = n_1684 ^ n_2627;
assign n_3132 = n_1685 ^ n_2628;
assign n_3133 = n_1686 ^ n_2629;
assign n_3134 = n_1687 ^ n_2630;
assign n_3135 = n_1688 ^ n_2631;
assign n_3136 = n_1689 ^ n_2632;
assign n_3137 = n_1690 ^ n_2633;
assign n_3138 = n_1691 ^ n_2634;
assign n_3139 = n_1692 ^ n_2635;
assign n_3140 = n_1693 ^ n_2636;
assign n_3141 = n_1694 ^ n_2637;
assign n_3142 = n_1695 ^ n_2638;
assign n_3143 = n_1696 ^ n_2639;
assign n_3144 = n_1697 ^ n_2640;
assign n_3145 = n_1698 ^ n_2641;
assign n_3146 = n_1699 ^ n_2642;
assign n_3147 = n_1700 ^ n_2643;
assign n_3148 = n_1701 ^ n_2644;
assign n_3149 = n_1702 ^ n_2645;
assign n_3150 = n_1703 ^ n_2646;
assign n_3151 = n_1704 ^ n_2647;
assign n_3152 = n_1705 ^ n_2648;
assign n_3153 = n_1706 ^ n_2649;
assign n_3154 = n_1707 ^ n_2650;
assign n_3155 = n_1708 ^ n_2651;
assign n_3156 = n_1709 ^ n_2652;
assign n_3157 = n_1710 ^ n_2653;
assign n_3158 = n_1711 ^ n_2654;
assign n_3159 = n_1745 ^ n_2689;
assign n_3160 = n_1747 ^ n_2690;
assign n_3161 = n_1748 ^ n_2691;
assign n_3162 = n_1749 ^ n_2692;
assign n_3163 = n_1750 ^ n_2693;
assign n_3164 = n_1751 ^ n_2694;
assign n_3165 = n_1752 ^ n_2695;
assign n_3166 = n_1753 ^ n_2696;
assign n_3167 = n_1754 ^ n_2697;
assign n_3168 = n_1755 ^ n_2698;
assign n_3169 = n_1756 ^ n_2699;
assign n_3170 = n_1757 ^ n_2700;
assign n_3171 = n_1758 ^ n_2701;
assign n_3172 = n_1759 ^ n_2702;
assign n_3173 = n_1760 ^ n_2703;
assign n_3174 = n_1761 ^ n_2704;
assign n_3175 = n_1762 ^ n_2705;
assign n_3176 = n_1763 ^ n_2706;
assign n_3177 = n_1764 ^ n_2707;
assign n_3178 = n_1765 ^ n_2708;
assign n_3179 = n_1766 ^ n_2709;
assign n_3180 = n_1767 ^ n_2710;
assign n_3181 = n_1768 ^ n_2711;
assign n_3182 = n_1769 ^ n_2712;
assign n_3183 = n_1770 ^ n_2713;
assign n_3184 = n_1771 ^ n_2714;
assign n_3185 = n_1772 ^ n_2715;
assign n_3186 = n_1773 ^ n_2716;
assign n_3187 = n_1774 ^ n_2717;
assign n_3188 = n_1775 ^ n_2718;
assign n_3189 = n_1776 ^ n_2719;
assign n_3190 = n_2721 ^ n_123;
assign n_3191 = ~n_1781 & n_2722;
assign y2 = n_2723;
assign n_3192 = n_1790 ^ n_2724;
assign n_3193 = n_2725 ^ n_1793;
assign n_3194 = n_2726 ^ n_1794;
assign n_3195 = n_2727 ^ n_1795;
assign n_3196 = n_2728 ^ n_1796;
assign n_3197 = n_2729 ^ n_1797;
assign n_3198 = n_2730 ^ n_1798;
assign n_3199 = n_2731 ^ n_1799;
assign n_3200 = n_2732 ^ n_1800;
assign n_3201 = n_2733 ^ n_1801;
assign n_3202 = n_2734 ^ n_1802;
assign n_3203 = n_2735 ^ n_1803;
assign n_3204 = n_2736 ^ n_1804;
assign n_3205 = n_2737 ^ n_1805;
assign n_3206 = n_2738 ^ n_1806;
assign n_3207 = n_2739 ^ n_1807;
assign n_3208 = n_2740 ^ n_1808;
assign n_3209 = n_2741 ^ n_1809;
assign n_3210 = n_2742 ^ n_1810;
assign n_3211 = n_2743 ^ n_1811;
assign n_3212 = n_2744 ^ n_1812;
assign n_3213 = n_2745 ^ n_1813;
assign n_3214 = n_2746 ^ n_1814;
assign n_3215 = n_2747 ^ n_1815;
assign n_3216 = n_2748 ^ n_1816;
assign n_3217 = n_2749 ^ n_1817;
assign n_3218 = n_2750 ^ n_1818;
assign n_3219 = n_2751 ^ n_1819;
assign n_3220 = n_2752 ^ n_1820;
assign n_3221 = n_2753 ^ n_1821;
assign n_3222 = n_162 ^ n_2754;
assign n_3223 = n_2755 ^ n_1883;
assign n_3224 = n_2756 ^ n_1854;
assign n_3225 = n_2757 ^ n_1855;
assign n_3226 = n_2758 ^ n_1856;
assign n_3227 = n_2759 ^ n_1857;
assign n_3228 = n_2760 ^ n_1858;
assign n_3229 = n_2761 ^ n_1859;
assign n_3230 = n_2762 ^ n_1860;
assign n_3231 = n_2763 ^ n_1861;
assign n_3232 = n_2764 ^ n_1862;
assign n_3233 = n_2765 ^ n_1863;
assign n_3234 = n_2766 ^ n_1864;
assign n_3235 = n_2767 ^ n_1865;
assign n_3236 = n_2768 ^ n_1866;
assign n_3237 = n_2769 ^ n_1867;
assign n_3238 = n_2770 ^ n_1868;
assign n_3239 = n_2771 ^ n_1869;
assign n_3240 = n_2772 ^ n_1870;
assign n_3241 = n_2773 ^ n_1871;
assign n_3242 = n_2774 ^ n_1872;
assign n_3243 = n_2775 ^ n_1873;
assign n_3244 = n_2776 ^ n_1874;
assign n_3245 = n_2777 ^ n_1875;
assign n_3246 = n_2778 ^ n_1876;
assign n_3247 = n_2779 ^ n_1877;
assign n_3248 = n_2780 ^ n_1878;
assign n_3249 = n_2781 ^ n_1879;
assign n_3250 = n_2782 ^ n_1880;
assign n_3251 = n_2783 ^ n_1881;
assign n_3252 = n_2784 ^ n_1882;
assign n_3253 = n_167 ^ n_2785;
assign n_3254 = n_2787 ^ n_1919;
assign n_3255 = n_2788 ^ n_1920;
assign n_3256 = n_2789 ^ n_1921;
assign n_3257 = n_2790 ^ n_1922;
assign n_3258 = n_2791 ^ n_1923;
assign n_3259 = n_2792 ^ n_1924;
assign n_3260 = n_2793 ^ n_1925;
assign n_3261 = n_2794 ^ n_1926;
assign n_3262 = n_2795 ^ n_1927;
assign n_3263 = n_2796 ^ n_1928;
assign n_3264 = n_2797 ^ n_1929;
assign n_3265 = n_2798 ^ n_1930;
assign n_3266 = n_2799 ^ n_1931;
assign n_3267 = n_2800 ^ n_1932;
assign n_3268 = n_2801 ^ n_1933;
assign n_3269 = n_2802 ^ n_1934;
assign n_3270 = n_2803 ^ n_1935;
assign n_3271 = n_2804 ^ n_1936;
assign n_3272 = n_2805 ^ n_1937;
assign n_3273 = n_2806 ^ n_1938;
assign n_3274 = n_2807 ^ n_1939;
assign n_3275 = n_2808 ^ n_1940;
assign n_3276 = n_2809 ^ n_1941;
assign n_3277 = n_2810 ^ n_1942;
assign n_3278 = n_2811 ^ n_1943;
assign n_3279 = n_2812 ^ n_1944;
assign n_3280 = n_2813 ^ n_1945;
assign n_3281 = n_2814 ^ n_1946;
assign n_3282 = n_2815 ^ n_1947;
assign n_3283 = n_172 ^ n_2816;
assign n_3284 = n_2817 ^ n_798;
assign n_3285 = n_2818 ^ n_1979;
assign n_3286 = n_2819 ^ n_1980;
assign n_3287 = n_2820 ^ n_1981;
assign n_3288 = n_2821 ^ n_1982;
assign n_3289 = n_2822 ^ n_1983;
assign n_3290 = n_2823 ^ n_1984;
assign n_3291 = n_2824 ^ n_1985;
assign n_3292 = n_2825 ^ n_1986;
assign n_3293 = n_2826 ^ n_1987;
assign n_3294 = n_2827 ^ n_1988;
assign n_3295 = n_2828 ^ n_1989;
assign n_3296 = n_2829 ^ n_1990;
assign n_3297 = n_2830 ^ n_1991;
assign n_3298 = n_2831 ^ n_1992;
assign n_3299 = n_2832 ^ n_1993;
assign n_3300 = n_2833 ^ n_1994;
assign n_3301 = n_2834 ^ n_1995;
assign n_3302 = n_2835 ^ n_1996;
assign n_3303 = n_2836 ^ n_1997;
assign n_3304 = n_2837 ^ n_1998;
assign n_3305 = n_2838 ^ n_1999;
assign n_3306 = n_2839 ^ n_2000;
assign n_3307 = n_2840 ^ n_2001;
assign n_3308 = n_2841 ^ n_2002;
assign n_3309 = n_2842 ^ n_2003;
assign n_3310 = n_2843 ^ n_2004;
assign n_3311 = n_2844 ^ n_2005;
assign n_3312 = n_2845 ^ n_2006;
assign n_3313 = n_2846 ^ n_2007;
assign n_3314 = n_177 ^ n_2847;
assign n_3315 = n_2849 ^ n_2039;
assign n_3316 = n_2850 ^ n_2040;
assign n_3317 = n_2851 ^ n_2041;
assign n_3318 = n_2852 ^ n_2042;
assign n_3319 = n_2853 ^ n_2043;
assign n_3320 = n_2854 ^ n_2044;
assign n_3321 = n_2855 ^ n_2045;
assign n_3322 = n_2856 ^ n_2046;
assign n_3323 = n_2857 ^ n_2047;
assign n_3324 = n_2858 ^ n_2048;
assign n_3325 = n_2859 ^ n_2049;
assign n_3326 = n_2860 ^ n_2050;
assign n_3327 = n_2861 ^ n_2051;
assign n_3328 = n_2862 ^ n_2052;
assign n_3329 = n_2863 ^ n_2053;
assign n_3330 = n_2864 ^ n_2054;
assign n_3331 = n_2865 ^ n_2055;
assign n_3332 = n_2866 ^ n_2056;
assign n_3333 = n_2867 ^ n_2057;
assign n_3334 = n_2868 ^ n_2058;
assign n_3335 = n_2869 ^ n_2059;
assign n_3336 = n_2870 ^ n_2060;
assign n_3337 = n_2871 ^ n_2061;
assign n_3338 = n_2872 ^ n_2062;
assign n_3339 = n_2873 ^ n_2063;
assign n_3340 = n_2874 ^ n_2064;
assign n_3341 = n_2875 ^ n_2065;
assign n_3342 = n_2876 ^ n_2066;
assign n_3343 = n_2877 ^ n_2067;
assign n_3344 = n_182 ^ n_2878;
assign n_3345 = n_2880 ^ n_2103;
assign n_3346 = n_2881 ^ n_2104;
assign n_3347 = n_2882 ^ n_2105;
assign n_3348 = n_2883 ^ n_2106;
assign n_3349 = n_2884 ^ n_2107;
assign n_3350 = n_2885 ^ n_2108;
assign n_3351 = n_2886 ^ n_2109;
assign n_3352 = n_2887 ^ n_2110;
assign n_3353 = n_2888 ^ n_2111;
assign n_3354 = n_2889 ^ n_2112;
assign n_3355 = n_2890 ^ n_2113;
assign n_3356 = n_2891 ^ n_2114;
assign n_3357 = n_2892 ^ n_2115;
assign n_3358 = n_2893 ^ n_2116;
assign n_3359 = n_2894 ^ n_2117;
assign n_3360 = n_2895 ^ n_2118;
assign n_3361 = n_2896 ^ n_2119;
assign n_3362 = n_2897 ^ n_2120;
assign n_3363 = n_2898 ^ n_2121;
assign n_3364 = n_2899 ^ n_2122;
assign n_3365 = n_2900 ^ n_2123;
assign n_3366 = n_2901 ^ n_2124;
assign n_3367 = n_2902 ^ n_2125;
assign n_3368 = n_2903 ^ n_2126;
assign n_3369 = n_2904 ^ n_2127;
assign n_3370 = n_2905 ^ n_2128;
assign n_3371 = n_2906 ^ n_2129;
assign n_3372 = n_2907 ^ n_2130;
assign n_3373 = n_2908 ^ n_2131;
assign n_3374 = n_187 ^ n_2909;
assign n_3375 = n_2911 ^ n_2163;
assign n_3376 = n_2912 ^ n_2164;
assign n_3377 = n_2913 ^ n_2165;
assign n_3378 = n_2914 ^ n_2166;
assign n_3379 = n_2915 ^ n_2167;
assign n_3380 = n_2916 ^ n_2168;
assign n_3381 = n_2917 ^ n_2169;
assign n_3382 = n_2918 ^ n_2170;
assign n_3383 = n_2919 ^ n_2171;
assign n_3384 = n_2920 ^ n_2172;
assign n_3385 = n_2921 ^ n_2173;
assign n_3386 = n_2922 ^ n_2174;
assign n_3387 = n_2923 ^ n_2175;
assign n_3388 = n_2924 ^ n_2176;
assign n_3389 = n_2925 ^ n_2177;
assign n_3390 = n_2926 ^ n_2178;
assign n_3391 = n_2927 ^ n_2179;
assign n_3392 = n_2928 ^ n_2180;
assign n_3393 = n_2929 ^ n_2181;
assign n_3394 = n_2930 ^ n_2182;
assign n_3395 = n_2931 ^ n_2183;
assign n_3396 = n_2932 ^ n_2184;
assign n_3397 = n_2933 ^ n_2185;
assign n_3398 = n_2934 ^ n_2186;
assign n_3399 = n_2935 ^ n_2187;
assign n_3400 = n_2936 ^ n_2188;
assign n_3401 = n_2937 ^ n_2189;
assign n_3402 = n_2938 ^ n_2190;
assign n_3403 = n_2939 ^ n_2191;
assign n_3404 = n_192 ^ n_2940;
assign n_3405 = n_2942 ^ n_2226;
assign n_3406 = n_2943 ^ n_2227;
assign n_3407 = n_2944 ^ n_2228;
assign n_3408 = n_2945 ^ n_2229;
assign n_3409 = n_2946 ^ n_2230;
assign n_3410 = n_2947 ^ n_2231;
assign n_3411 = n_2948 ^ n_2232;
assign n_3412 = n_2949 ^ n_2233;
assign n_3413 = n_2950 ^ n_2234;
assign n_3414 = n_2951 ^ n_2235;
assign n_3415 = n_2952 ^ n_2236;
assign n_3416 = n_2953 ^ n_2237;
assign n_3417 = n_2954 ^ n_2238;
assign n_3418 = n_2955 ^ n_2239;
assign n_3419 = n_2956 ^ n_2240;
assign n_3420 = n_2957 ^ n_2241;
assign n_3421 = n_2958 ^ n_2242;
assign n_3422 = n_2959 ^ n_2243;
assign n_3423 = n_2960 ^ n_2244;
assign n_3424 = n_2961 ^ n_2245;
assign n_3425 = n_2962 ^ n_2246;
assign n_3426 = n_2963 ^ n_2247;
assign n_3427 = n_2964 ^ n_2248;
assign n_3428 = n_2965 ^ n_2249;
assign n_3429 = n_2966 ^ n_2250;
assign n_3430 = n_2967 ^ n_2251;
assign n_3431 = n_2968 ^ n_2252;
assign n_3432 = n_2969 ^ n_2253;
assign n_3433 = n_2970 ^ n_2254;
assign n_3434 = n_197 ^ n_2971;
assign n_3435 = n_2973 ^ n_2288;
assign n_3436 = n_2974 ^ n_2289;
assign n_3437 = n_2975 ^ n_2290;
assign n_3438 = n_2976 ^ n_2291;
assign n_3439 = n_2977 ^ n_2292;
assign n_3440 = n_2978 ^ n_2293;
assign n_3441 = n_2979 ^ n_2294;
assign n_3442 = n_2980 ^ n_2295;
assign n_3443 = n_2981 ^ n_2296;
assign n_3444 = n_2982 ^ n_2297;
assign n_3445 = n_2983 ^ n_2298;
assign n_3446 = n_2984 ^ n_2299;
assign n_3447 = n_2985 ^ n_2300;
assign n_3448 = n_2986 ^ n_2301;
assign n_3449 = n_2987 ^ n_2302;
assign n_3450 = n_2988 ^ n_2303;
assign n_3451 = n_2989 ^ n_2304;
assign n_3452 = n_2990 ^ n_2305;
assign n_3453 = n_2991 ^ n_2306;
assign n_3454 = n_2992 ^ n_2307;
assign n_3455 = n_2993 ^ n_2308;
assign n_3456 = n_2994 ^ n_2309;
assign n_3457 = n_2995 ^ n_2310;
assign n_3458 = n_2996 ^ n_2311;
assign n_3459 = n_2997 ^ n_2312;
assign n_3460 = n_2998 ^ n_2313;
assign n_3461 = n_2999 ^ n_2314;
assign n_3462 = n_3000 ^ n_2315;
assign n_3463 = n_3001 ^ n_2316;
assign n_3464 = n_202 ^ n_3002;
assign n_3465 = n_3004 ^ n_2351;
assign n_3466 = n_3005 ^ n_2352;
assign n_3467 = n_3006 ^ n_2353;
assign n_3468 = n_3007 ^ n_2354;
assign n_3469 = n_3008 ^ n_2355;
assign n_3470 = n_3009 ^ n_2356;
assign n_3471 = n_3010 ^ n_2357;
assign n_3472 = n_3011 ^ n_2358;
assign n_3473 = n_3012 ^ n_2359;
assign n_3474 = n_3013 ^ n_2360;
assign n_3475 = n_3014 ^ n_2361;
assign n_3476 = n_3015 ^ n_2362;
assign n_3477 = n_3016 ^ n_2363;
assign n_3478 = n_3017 ^ n_2364;
assign n_3479 = n_3018 ^ n_2365;
assign n_3480 = n_3019 ^ n_2366;
assign n_3481 = n_3020 ^ n_2367;
assign n_3482 = n_3021 ^ n_2368;
assign n_3483 = n_3022 ^ n_2369;
assign n_3484 = n_3023 ^ n_2370;
assign n_3485 = n_3024 ^ n_2371;
assign n_3486 = n_3025 ^ n_2372;
assign n_3487 = n_3026 ^ n_2373;
assign n_3488 = n_3027 ^ n_2374;
assign n_3489 = n_3028 ^ n_2375;
assign n_3490 = n_3029 ^ n_2376;
assign n_3491 = n_3030 ^ n_2377;
assign n_3492 = n_3031 ^ n_2378;
assign n_3493 = n_3032 ^ n_2379;
assign n_3494 = n_207 ^ n_3033;
assign n_3495 = n_3035 ^ n_2412;
assign n_3496 = n_3036 ^ n_2413;
assign n_3497 = n_3037 ^ n_2414;
assign n_3498 = n_3038 ^ n_2415;
assign n_3499 = n_3039 ^ n_2416;
assign n_3500 = n_3040 ^ n_2417;
assign n_3501 = n_3041 ^ n_2418;
assign n_3502 = n_3042 ^ n_2419;
assign n_3503 = n_3043 ^ n_2420;
assign n_3504 = n_3044 ^ n_2421;
assign n_3505 = n_3045 ^ n_2422;
assign n_3506 = n_3046 ^ n_2423;
assign n_3507 = n_3047 ^ n_2424;
assign n_3508 = n_3048 ^ n_2425;
assign n_3509 = n_3049 ^ n_2426;
assign n_3510 = n_3050 ^ n_2427;
assign n_3511 = n_3051 ^ n_2428;
assign n_3512 = n_3052 ^ n_2429;
assign n_3513 = n_3053 ^ n_2430;
assign n_3514 = n_3054 ^ n_2431;
assign n_3515 = n_3055 ^ n_2432;
assign n_3516 = n_3056 ^ n_2433;
assign n_3517 = n_3057 ^ n_2434;
assign n_3518 = n_3058 ^ n_2435;
assign n_3519 = n_3059 ^ n_2436;
assign n_3520 = n_3060 ^ n_2437;
assign n_3521 = n_3061 ^ n_2438;
assign n_3522 = n_3062 ^ n_2439;
assign n_3523 = n_3063 ^ n_2440;
assign n_3524 = n_212 ^ n_3064;
assign n_3525 = n_3066 ^ n_2472;
assign n_3526 = n_3067 ^ n_2473;
assign n_3527 = n_3068 ^ n_2474;
assign n_3528 = n_3069 ^ n_2475;
assign n_3529 = n_3070 ^ n_2476;
assign n_3530 = n_3071 ^ n_2477;
assign n_3531 = n_3072 ^ n_2478;
assign n_3532 = n_3073 ^ n_2479;
assign n_3533 = n_3074 ^ n_2480;
assign n_3534 = n_3075 ^ n_2481;
assign n_3535 = n_3076 ^ n_2482;
assign n_3536 = n_3077 ^ n_2483;
assign n_3537 = n_3078 ^ n_2484;
assign n_3538 = n_3079 ^ n_2485;
assign n_3539 = n_3080 ^ n_2486;
assign n_3540 = n_3081 ^ n_2487;
assign n_3541 = n_3082 ^ n_2488;
assign n_3542 = n_3083 ^ n_2489;
assign n_3543 = n_3084 ^ n_2490;
assign n_3544 = n_3085 ^ n_2491;
assign n_3545 = n_3086 ^ n_2492;
assign n_3546 = n_3087 ^ n_2493;
assign n_3547 = n_3088 ^ n_2494;
assign n_3548 = n_3089 ^ n_2495;
assign n_3549 = n_3090 ^ n_2496;
assign n_3550 = n_3091 ^ n_2497;
assign n_3551 = n_3092 ^ n_2498;
assign n_3552 = n_3093 ^ n_2499;
assign n_3553 = n_3094 ^ n_2500;
assign n_3554 = n_217 ^ n_3095;
assign n_3555 = n_3097 ^ n_2533;
assign n_3556 = n_3098 ^ n_2534;
assign n_3557 = n_3099 ^ n_2535;
assign n_3558 = n_3100 ^ n_2536;
assign n_3559 = n_3101 ^ n_2537;
assign n_3560 = n_3102 ^ n_2538;
assign n_3561 = n_3103 ^ n_2539;
assign n_3562 = n_3104 ^ n_2540;
assign n_3563 = n_3105 ^ n_2541;
assign n_3564 = n_3106 ^ n_2542;
assign n_3565 = n_3107 ^ n_2543;
assign n_3566 = n_3108 ^ n_2544;
assign n_3567 = n_3109 ^ n_2545;
assign n_3568 = n_3110 ^ n_2546;
assign n_3569 = n_3111 ^ n_2547;
assign n_3570 = n_3112 ^ n_2548;
assign n_3571 = n_3113 ^ n_2549;
assign n_3572 = n_3114 ^ n_2550;
assign n_3573 = n_3115 ^ n_2551;
assign n_3574 = n_3116 ^ n_2552;
assign n_3575 = n_3117 ^ n_2553;
assign n_3576 = n_3118 ^ n_2554;
assign n_3577 = n_3119 ^ n_2555;
assign n_3578 = n_3120 ^ n_2556;
assign n_3579 = n_3121 ^ n_2557;
assign n_3580 = n_3122 ^ n_2558;
assign n_3581 = n_3123 ^ n_2559;
assign n_3582 = n_3124 ^ n_2560;
assign n_3583 = n_3125 ^ n_2561;
assign n_3584 = n_222 ^ n_3126;
assign n_3585 = n_3128 ^ n_2623;
assign n_3586 = n_3129 ^ n_2594;
assign n_3587 = n_3130 ^ n_2595;
assign n_3588 = n_3131 ^ n_2596;
assign n_3589 = n_3132 ^ n_2597;
assign n_3590 = n_3133 ^ n_2598;
assign n_3591 = n_3134 ^ n_2599;
assign n_3592 = n_3135 ^ n_2600;
assign n_3593 = n_3136 ^ n_2601;
assign n_3594 = n_3137 ^ n_2602;
assign n_3595 = n_3138 ^ n_2603;
assign n_3596 = n_3139 ^ n_2604;
assign n_3597 = n_3140 ^ n_2605;
assign n_3598 = n_3141 ^ n_2606;
assign n_3599 = n_3142 ^ n_2607;
assign n_3600 = n_3143 ^ n_2608;
assign n_3601 = n_3144 ^ n_2609;
assign n_3602 = n_3145 ^ n_2610;
assign n_3603 = n_3146 ^ n_2611;
assign n_3604 = n_3147 ^ n_2612;
assign n_3605 = n_3148 ^ n_2613;
assign n_3606 = n_3149 ^ n_2614;
assign n_3607 = n_3150 ^ n_2615;
assign n_3608 = n_3151 ^ n_2616;
assign n_3609 = n_3152 ^ n_2617;
assign n_3610 = n_3153 ^ n_2618;
assign n_3611 = n_3154 ^ n_2619;
assign n_3612 = n_3155 ^ n_2620;
assign n_3613 = n_3156 ^ n_2621;
assign n_3614 = n_3157 ^ n_2622;
assign n_3615 = n_227 ^ n_3158;
assign n_3616 = n_3159 ^ n_2657;
assign n_3617 = n_3160 ^ n_2658;
assign n_3618 = n_3161 ^ n_2659;
assign n_3619 = n_3162 ^ n_2660;
assign n_3620 = n_3163 ^ n_2661;
assign n_3621 = n_3164 ^ n_2662;
assign n_3622 = n_3165 ^ n_2663;
assign n_3623 = n_3166 ^ n_2664;
assign n_3624 = n_3167 ^ n_2665;
assign n_3625 = n_3168 ^ n_2666;
assign n_3626 = n_3169 ^ n_2667;
assign n_3627 = n_3170 ^ n_2668;
assign n_3628 = n_3171 ^ n_2669;
assign n_3629 = n_3172 ^ n_2670;
assign n_3630 = n_3173 ^ n_2671;
assign n_3631 = n_3174 ^ n_2672;
assign n_3632 = n_3175 ^ n_2673;
assign n_3633 = n_3176 ^ n_2674;
assign n_3634 = n_3177 ^ n_2675;
assign n_3635 = n_3178 ^ n_2676;
assign n_3636 = n_3179 ^ n_2677;
assign n_3637 = n_3180 ^ n_2678;
assign n_3638 = n_3181 ^ n_2679;
assign n_3639 = n_3182 ^ n_2680;
assign n_3640 = n_3183 ^ n_2681;
assign n_3641 = n_3184 ^ n_2682;
assign n_3642 = n_3185 ^ n_2683;
assign n_3643 = n_3186 ^ n_2684;
assign n_3644 = n_3187 ^ n_2685;
assign n_3645 = n_3188 ^ n_2686;
assign n_3646 = n_232 ^ n_3189;
assign n_3647 = n_3191 ^ n_1780;
assign n_3648 = n_163 ^ n_3193;
assign n_3649 = n_3193 ^ n_793;
assign n_3650 = n_2755 ^ n_3194;
assign n_3651 = n_1783 ^ n_3195;
assign n_3652 = n_795 ^ n_3195;
assign n_3653 = n_2786 ^ n_3196;
assign n_3654 = n_1044 ^ n_3198;
assign n_3655 = ~n_3198 & n_1044;
assign n_3656 = n_178 ^ n_3199;
assign n_3657 = n_1108 ^ n_3200;
assign n_3658 = ~n_3200 & n_1108;
assign n_3659 = n_183 ^ n_3201;
assign n_3660 = n_1785 ^ n_3203;
assign n_3661 = n_803 ^ n_3203;
assign n_3662 = n_2910 ^ n_3204;
assign n_3663 = n_1786 ^ n_3205;
assign n_3664 = n_805 ^ n_3205;
assign n_3665 = n_2972 ^ n_3208;
assign n_3666 = n_1395 ^ n_3210;
assign n_3667 = ~n_3210 & n_1395;
assign n_3668 = n_208 ^ n_3211;
assign n_3669 = n_1459 ^ n_3212;
assign n_3670 = ~n_3212 & n_1459;
assign n_3671 = n_213 ^ n_3213;
assign n_3672 = n_1523 ^ n_3214;
assign n_3673 = ~n_3214 & n_1523;
assign n_3674 = n_218 ^ n_3215;
assign n_3675 = n_1617 ^ n_3216;
assign n_3676 = ~n_3216 & n_1617;
assign n_3677 = n_223 ^ n_3217;
assign n_3678 = n_1789 ^ n_3219;
assign n_3679 = n_819 ^ n_3219;
assign n_3680 = n_821 ^ n_3221;
assign n_3681 = n_264 ^ n_3221;
assign n_3682 = n_1884 ^ n_3224;
assign n_3683 = n_3196 ^ n_3225;
assign n_3684 = n_2786 ^ n_3225;
assign n_3685 = n_3226 ^ n_3197;
assign n_3686 = n_3226 ^ n_1917;
assign n_3687 = n_2848 ^ n_3229;
assign n_3688 = n_3239 ^ n_810;
assign n_3689 = n_3241 ^ n_812;
assign n_3690 = n_3241 ^ n_3034;
assign n_3691 = n_3065 ^ n_3243;
assign n_3692 = n_3245 ^ n_3096;
assign n_3693 = n_884 ^ n_3253;
assign n_3694 = n_1784 ^ n_3254;
assign n_3695 = n_797 ^ n_3254;
assign n_3696 = n_2817 ^ n_3255;
assign n_3697 = n_3199 ^ n_3256;
assign n_3698 = n_3257 ^ n_800;
assign n_3699 = n_183 ^ n_3258;
assign n_3700 = n_3201 ^ n_3258;
assign n_3701 = n_3259 ^ n_3202;
assign n_3702 = n_3260 ^ n_3232;
assign n_3703 = n_2910 ^ n_3261;
assign n_3704 = n_1787 ^ n_3264;
assign n_3705 = n_807 ^ n_3264;
assign n_3706 = n_1788 ^ n_3266;
assign n_3707 = n_809 ^ n_3266;
assign n_3708 = n_208 ^ n_3268;
assign n_3709 = n_3211 ^ n_3268;
assign n_3710 = n_3213 ^ n_3270;
assign n_3711 = n_3215 ^ n_3272;
assign n_3712 = n_223 ^ n_3274;
assign n_3713 = n_3217 ^ n_3274;
assign n_3714 = n_3275 ^ n_3218;
assign n_3715 = n_3277 ^ n_3220;
assign n_3716 = n_3222 ^ n_3279;
assign n_3717 = n_948 ^ n_3283;
assign n_3718 = n_3285 ^ n_799;
assign n_3719 = n_3285 ^ n_3228;
assign n_3720 = n_3286 ^ n_3257;
assign n_3721 = n_3287 ^ n_801;
assign n_3722 = n_3202 ^ n_3288;
assign n_3723 = n_3289 ^ n_3260;
assign n_3724 = n_3289 ^ n_3232;
assign n_3725 = n_3290 ^ n_3233;
assign n_3726 = n_3262 ^ n_3291;
assign n_3727 = n_3292 ^ n_3206;
assign n_3728 = n_3292 ^ n_3235;
assign n_3729 = n_3293 ^ n_3236;
assign n_3730 = n_2972 ^ n_3294;
assign n_3731 = n_3295 ^ n_3238;
assign n_3732 = n_3296 ^ n_3003;
assign n_3733 = n_3309 ^ n_3252;
assign n_3734 = n_3309 ^ n_94;
assign n_3735 = n_884 ^ n_3310;
assign n_3736 = n_3253 ^ n_3310;
assign n_3737 = n_1012 ^ n_3314;
assign n_3738 = n_3287 ^ n_3315;
assign n_3739 = n_3316 ^ n_3231;
assign n_3740 = n_3316 ^ n_2879;
assign n_3741 = n_3290 ^ n_3318;
assign n_3742 = n_3233 ^ n_3318;
assign n_3743 = n_3319 ^ n_3234;
assign n_3744 = n_3320 ^ n_2255;
assign n_3745 = n_3293 ^ n_3321;
assign n_3746 = n_3322 ^ n_3237;
assign n_3747 = n_3239 ^ n_3324;
assign n_3748 = n_3325 ^ n_3240;
assign n_3749 = n_3242 ^ n_3327;
assign n_3750 = n_3328 ^ n_814;
assign n_3751 = n_3330 ^ n_816;
assign n_3752 = n_3247 ^ n_3332;
assign n_3753 = n_3333 ^ n_3248;
assign n_3754 = n_3250 ^ n_3335;
assign n_3755 = n_3336 ^ n_3251;
assign n_3756 = n_3339 ^ n_3282;
assign n_3757 = n_948 ^ n_3340;
assign n_3758 = n_3283 ^ n_3340;
assign n_3759 = n_3341 ^ n_98;
assign n_3760 = n_1076 ^ n_3344;
assign n_3761 = n_3345 ^ n_3317;
assign n_3762 = n_3345 ^ n_2101;
assign n_3763 = n_2192 ^ n_3346;
assign n_3764 = n_3234 ^ n_3347;
assign n_3765 = n_3348 ^ n_3320;
assign n_3766 = n_2256 ^ n_3349;
assign n_3767 = n_3322 ^ n_3350;
assign n_3768 = n_3351 ^ n_3323;
assign n_3769 = n_3351 ^ n_2318;
assign n_3770 = n_3325 ^ n_3353;
assign n_3771 = n_3354 ^ n_3326;
assign n_3772 = n_3243 ^ n_3356;
assign n_3773 = n_3357 ^ n_3244;
assign n_3774 = n_3246 ^ n_3359;
assign n_3775 = n_3366 ^ n_3281;
assign n_3776 = n_1012 ^ n_3370;
assign n_3777 = n_3314 ^ n_3370;
assign n_3778 = n_100 ^ n_3371;
assign n_3779 = n_2098 ^ n_3374;
assign n_3780 = n_3375 ^ n_3262;
assign n_3781 = n_3376 ^ n_3263;
assign n_3782 = n_3376 ^ n_2941;
assign n_3783 = n_3377 ^ n_3207;
assign n_3784 = n_3378 ^ n_3265;
assign n_3785 = n_3379 ^ n_3209;
assign n_3786 = n_3380 ^ n_3267;
assign n_3787 = n_3381 ^ n_3297;
assign n_3788 = n_3382 ^ n_3269;
assign n_3789 = n_3383 ^ n_3299;
assign n_3790 = n_3384 ^ n_3271;
assign n_3791 = n_3385 ^ n_3301;
assign n_3792 = n_3386 ^ n_3273;
assign n_3793 = n_3275 ^ n_3388;
assign n_3794 = n_3389 ^ n_3276;
assign n_3795 = n_3278 ^ n_3391;
assign n_3796 = n_3392 ^ n_93;
assign n_3797 = n_3311 ^ n_3395;
assign n_3798 = n_3344 ^ n_3400;
assign n_3799 = n_1140 ^ n_3401;
assign n_3800 = n_1203 ^ n_3404;
assign n_3801 = n_3405 ^ n_3377;
assign n_3802 = n_3378 ^ n_3406;
assign n_3803 = n_3407 ^ n_3379;
assign n_3804 = n_3407 ^ n_3209;
assign n_3805 = n_3267 ^ n_3408;
assign n_3806 = n_3409 ^ n_3381;
assign n_3807 = n_3269 ^ n_3410;
assign n_3808 = n_3411 ^ n_3383;
assign n_3809 = n_3411 ^ n_3299;
assign n_3810 = n_3384 ^ n_3412;
assign n_3811 = n_3413 ^ n_3385;
assign n_3812 = n_3413 ^ n_3301;
assign n_3813 = n_3386 ^ n_3414;
assign n_3814 = n_3415 ^ n_3387;
assign n_3815 = n_3415 ^ n_3303;
assign n_3816 = n_3416 ^ n_3304;
assign n_3817 = n_3389 ^ n_3417;
assign n_3818 = n_3418 ^ n_3390;
assign n_3819 = n_3418 ^ n_3306;
assign n_3820 = n_3419 ^ n_3307;
assign n_3821 = n_3420 ^ n_3222;
assign n_3822 = n_95 ^ n_3422;
assign n_3823 = n_3424 ^ n_97;
assign n_3824 = n_1013 ^ n_3425;
assign n_3825 = n_3374 ^ n_3430;
assign n_3826 = n_1204 ^ n_3431;
assign n_3827 = n_105 ^ n_3432;
assign n_3828 = n_106 ^ n_3433;
assign n_3829 = n_2224 ^ n_3434;
assign n_3830 = n_3435 ^ n_3295;
assign n_3831 = n_3436 ^ n_3296;
assign n_3832 = n_3437 ^ n_811;
assign n_3833 = n_3438 ^ n_3298;
assign n_3834 = n_3439 ^ n_813;
assign n_3835 = n_3440 ^ n_3300;
assign n_3836 = n_3442 ^ n_3302;
assign n_3837 = n_3443 ^ n_817;
assign n_3838 = n_3304 ^ n_3444;
assign n_3839 = n_3445 ^ n_3305;
assign n_3840 = n_3446 ^ n_3249;
assign n_3841 = n_3419 ^ n_3447;
assign n_3842 = n_3448 ^ n_3308;
assign n_3843 = n_3449 ^ n_3421;
assign n_3844 = n_3449 ^ n_3337;
assign n_3845 = n_95 ^ n_3450;
assign n_3846 = n_3422 ^ n_3450;
assign n_3847 = n_3282 ^ n_3451;
assign n_3848 = n_3452 ^ n_3368;
assign n_3849 = n_3453 ^ n_3313;
assign n_3850 = n_99 ^ n_3454;
assign n_3851 = n_3454 ^ n_3313;
assign n_3852 = n_1077 ^ n_3455;
assign n_3853 = n_3456 ^ n_101;
assign n_3854 = n_3404 ^ n_3460;
assign n_3855 = n_107 ^ n_3462;
assign n_3856 = n_1330 ^ n_3464;
assign n_3857 = n_3465 ^ n_3437;
assign n_3858 = n_3298 ^ n_3466;
assign n_3859 = n_3467 ^ n_3439;
assign n_3860 = n_3300 ^ n_3468;
assign n_3861 = n_3440 ^ n_3468;
assign n_3862 = n_3469 ^ n_3441;
assign n_3863 = n_3469 ^ n_815;
assign n_3864 = n_3442 ^ n_3470;
assign n_3865 = n_3471 ^ n_3443;
assign n_3866 = n_3472 ^ n_3247;
assign n_3867 = n_3445 ^ n_3473;
assign n_3868 = n_3474 ^ n_3446;
assign n_3869 = n_3474 ^ n_3249;
assign n_3870 = n_3475 ^ n_3250;
assign n_3871 = n_3475 ^ n_3335;
assign n_3872 = n_3308 ^ n_3476;
assign n_3873 = n_3478 ^ n_3338;
assign n_3874 = n_3479 ^ n_3367;
assign n_3875 = n_3480 ^ n_3452;
assign n_3876 = n_3481 ^ n_3369;
assign n_3877 = n_3482 ^ n_3398;
assign n_3878 = n_3371 ^ n_3483;
assign n_3879 = n_3484 ^ n_3343;
assign n_3880 = n_3485 ^ n_3373;
assign n_3881 = n_103 ^ n_3486;
assign n_3882 = n_3487 ^ n_104;
assign n_3883 = n_3434 ^ n_3490;
assign n_3884 = n_3463 ^ n_3491;
assign n_3885 = n_110 ^ n_3493;
assign n_3886 = n_2349 ^ n_3494;
assign n_3887 = n_3495 ^ n_3242;
assign n_3888 = n_3495 ^ n_3327;
assign n_3889 = n_814 ^ n_3496;
assign n_3890 = n_3328 ^ n_3496;
assign n_3891 = n_3497 ^ n_3329;
assign n_3892 = n_3330 ^ n_3498;
assign n_3893 = n_3499 ^ n_3331;
assign n_3894 = n_3333 ^ n_3501;
assign n_3895 = n_3502 ^ n_3334;
assign n_3896 = n_3503 ^ n_3363;
assign n_3897 = n_3251 ^ n_3504;
assign n_3898 = n_3505 ^ n_3477;
assign n_3899 = n_3505 ^ n_3280;
assign n_3900 = n_3338 ^ n_3506;
assign n_3901 = n_3478 ^ n_3506;
assign n_3902 = n_3367 ^ n_3507;
assign n_3903 = n_3369 ^ n_3509;
assign n_3904 = n_3510 ^ n_3482;
assign n_3905 = n_3511 ^ n_3399;
assign n_3906 = n_3513 ^ n_3485;
assign n_3907 = n_3513 ^ n_3373;
assign n_3908 = n_3486 ^ n_3514;
assign n_3909 = n_1204 ^ n_3515;
assign n_3910 = n_3431 ^ n_3515;
assign n_3911 = n_3516 ^ n_3403;
assign n_3912 = n_3433 ^ n_3517;
assign n_3913 = n_1330 ^ n_3520;
assign n_3914 = n_3464 ^ n_3520;
assign n_3915 = n_1457 ^ n_3524;
assign n_3916 = n_3329 ^ n_3525;
assign n_3917 = n_3526 ^ n_3245;
assign n_3918 = n_3331 ^ n_3527;
assign n_3919 = n_3528 ^ n_3500;
assign n_3920 = n_3528 ^ n_3360;
assign n_3921 = n_3529 ^ n_3361;
assign n_3922 = n_3502 ^ n_3530;
assign n_3923 = n_3531 ^ n_3503;
assign n_3924 = n_3531 ^ n_3363;
assign n_3925 = n_3532 ^ n_3364;
assign n_3926 = n_3533 ^ n_3365;
assign n_3927 = n_3366 ^ n_3534;
assign n_3928 = n_3535 ^ n_3311;
assign n_3929 = n_3535 ^ n_3395;
assign n_3930 = n_3536 ^ n_3508;
assign n_3931 = n_3536 ^ n_3312;
assign n_3932 = n_3537 ^ n_3397;
assign n_3933 = n_3538 ^ n_3342;
assign n_3934 = n_3511 ^ n_3539;
assign n_3935 = n_3399 ^ n_3539;
assign n_3936 = n_3540 ^ n_3512;
assign n_3937 = n_3540 ^ n_3428;
assign n_3938 = n_3541 ^ n_3429;
assign n_3939 = n_3543 ^ n_3403;
assign n_3940 = n_3544 ^ n_3516;
assign n_3941 = n_3544 ^ n_3403;
assign n_3942 = n_3545 ^ n_3461;
assign n_3943 = n_3462 ^ n_3546;
assign n_3944 = n_3547 ^ n_3463;
assign n_3945 = n_109 ^ n_3548;
assign n_3946 = n_3493 ^ n_3549;
assign n_3947 = n_3494 ^ n_3550;
assign n_3948 = n_3551 ^ n_112;
assign n_3949 = n_114 ^ n_3553;
assign n_3950 = n_1521 ^ n_3554;
assign n_3951 = n_3555 ^ n_3246;
assign n_3952 = n_3128 ^ n_3556;
assign n_3953 = n_3361 ^ n_3557;
assign n_3954 = n_3558 ^ n_3362;
assign n_3955 = n_3364 ^ n_3560;
assign n_3956 = n_3532 ^ n_3560;
assign n_3957 = n_3533 ^ n_3561;
assign n_3958 = n_3562 ^ n_3394;
assign n_3959 = n_3563 ^ n_3423;
assign n_3960 = n_3564 ^ n_3396;
assign n_3961 = n_3397 ^ n_3565;
assign n_3962 = n_3566 ^ n_3538;
assign n_3963 = n_3567 ^ n_3427;
assign n_3964 = n_3568 ^ n_3372;
assign n_3965 = n_3429 ^ n_3569;
assign n_3966 = n_3570 ^ n_3542;
assign n_3967 = n_3570 ^ n_3458;
assign n_3968 = n_3571 ^ n_3459;
assign n_3969 = n_3572 ^ n_3488;
assign n_3970 = n_3545 ^ n_3573;
assign n_3971 = n_3461 ^ n_3573;
assign n_3972 = n_3574 ^ n_1267;
assign n_3973 = n_3576 ^ n_3492;
assign n_3974 = n_3577 ^ n_3521;
assign n_3975 = n_111 ^ n_3578;
assign n_3976 = n_3578 ^ n_3522;
assign n_3977 = n_3579 ^ n_3523;
assign n_3978 = n_3524 ^ n_3580;
assign n_3979 = n_114 ^ n_3581;
assign n_3980 = n_3581 ^ n_3553;
assign n_3981 = n_3582 ^ n_115;
assign n_3982 = n_117 ^ n_3583;
assign n_3983 = n_1585 ^ n_3584;
assign n_3984 = n_2624 ^ n_3586;
assign n_3985 = n_3558 ^ n_3587;
assign n_3986 = n_3588 ^ n_3559;
assign n_3987 = n_3588 ^ n_2688;
assign n_3988 = n_3589 ^ x33;
assign n_3989 = n_3590 ^ n_3393;
assign n_3990 = n_3394 ^ n_3591;
assign n_3991 = n_3562 ^ n_3591;
assign n_3992 = n_3592 ^ n_3563;
assign n_3993 = n_3396 ^ n_3593;
assign n_3994 = n_3425 ^ n_3594;
assign n_3995 = n_3595 ^ n_3426;
assign n_3996 = n_3427 ^ n_3596;
assign n_3997 = n_3597 ^ n_3568;
assign n_3998 = n_3598 ^ n_3457;
assign n_3999 = n_3599 ^ n_3402;
assign n_4000 = n_3571 ^ n_3600;
assign n_4001 = n_3459 ^ n_3600;
assign n_4002 = n_3601 ^ n_3572;
assign n_4003 = n_3602 ^ n_3489;
assign n_4004 = n_3604 ^ n_3575;
assign n_4005 = n_3604 ^ n_1331;
assign n_4006 = n_3576 ^ n_3605;
assign n_4007 = n_3577 ^ n_3606;
assign n_4008 = n_3607 ^ n_1394;
assign n_4009 = n_3579 ^ n_3608;
assign n_4010 = n_3609 ^ n_3552;
assign n_4011 = n_3554 ^ n_3611;
assign n_4012 = n_3612 ^ n_3583;
assign n_4013 = n_117 ^ n_3613;
assign n_4014 = n_3613 ^ n_3583;
assign n_4015 = n_118 ^ n_3614;
assign n_4016 = n_2592 ^ n_3615;
assign n_4017 = n_3277 ^ n_3616;
assign n_4018 = n_3617 ^ n_3278;
assign n_4019 = n_3617 ^ n_3391;
assign n_4020 = n_3618 ^ n_3392;
assign n_4021 = n_3590 ^ n_3619;
assign n_4022 = n_3620 ^ n_885;
assign n_4023 = n_96 ^ n_3621;
assign n_4024 = n_3621 ^ n_949;
assign n_4025 = n_3622 ^ n_3424;
assign n_4026 = n_3623 ^ n_3341;
assign n_4027 = n_3595 ^ n_3624;
assign n_4028 = n_1077 ^ n_3625;
assign n_4029 = n_3455 ^ n_3625;
assign n_4030 = n_3626 ^ n_3456;
assign n_4031 = n_3598 ^ n_3627;
assign n_4032 = n_3457 ^ n_3627;
assign n_4033 = n_3628 ^ n_3599;
assign n_4034 = n_3628 ^ n_3402;
assign n_4035 = n_3629 ^ n_3487;
assign n_4036 = n_105 ^ n_3630;
assign n_4037 = n_3630 ^ n_3432;
assign n_4038 = n_3602 ^ n_3631;
assign n_4039 = n_3632 ^ n_3603;
assign n_4040 = n_3632 ^ n_3518;
assign n_4041 = n_3633 ^ n_3519;
assign n_4042 = n_3633 ^ n_108;
assign n_4043 = n_109 ^ n_3634;
assign n_4044 = n_3634 ^ n_3548;
assign n_4045 = n_1394 ^ n_3635;
assign n_4046 = n_3636 ^ n_3607;
assign n_4047 = n_3637 ^ n_3551;
assign n_4048 = n_3609 ^ n_3638;
assign n_4049 = n_3552 ^ n_3638;
assign n_4050 = n_3639 ^ n_3610;
assign n_4051 = n_3639 ^ n_1522;
assign n_4052 = n_3640 ^ n_3582;
assign n_4053 = n_116 ^ n_3641;
assign n_4054 = n_3641 ^ n_1586;
assign n_4055 = n_1585 ^ n_3642;
assign n_4056 = n_3584 ^ n_3642;
assign n_4057 = n_3614 ^ n_3643;
assign n_4058 = n_3644 ^ n_1649;
assign n_4059 = n_120 ^ n_3645;
assign n_4060 = n_3645 ^ n_1713;
assign n_4061 = n_1712 ^ n_3646;
assign n_4062 = n_3647 ^ n_3192;
assign n_4063 = n_3647 ^ n_2724;
assign n_4064 = n_3648 ^ n_793;
assign n_4065 = n_1782 & n_3649;
assign n_4066 = n_3650 ^ n_1883;
assign n_4067 = n_3650 & n_3223;
assign n_4068 = n_3651 ^ n_1884;
assign n_4069 = n_1783 & n_3652;
assign n_4070 = n_3653 ^ n_3225;
assign n_4071 = n_3654 ^ n_3227;
assign n_4072 = n_3656 ^ n_3256;
assign n_4073 = n_2848 ^ n_3657;
assign n_4074 = n_3658 ^ n_3230;
assign n_4075 = n_3659 ^ n_3258;
assign n_4076 = n_1785 & n_3661;
assign n_4077 = n_3662 ^ n_3261;
assign n_4078 = n_1786 & n_3664;
assign n_4079 = n_3665 ^ n_3294;
assign n_4080 = n_3666 ^ n_3352;
assign n_4081 = n_3668 ^ n_3268;
assign n_4082 = n_3354 ^ n_3669;
assign n_4083 = n_3670 ^ n_3355;
assign n_4084 = n_3671 ^ n_3270;
assign n_4085 = n_3357 ^ n_3673;
assign n_4086 = n_3674 ^ n_3272;
assign n_4087 = n_3675 ^ n_3358;
assign n_4088 = n_3677 ^ n_3274;
assign n_4089 = n_1789 & n_3679;
assign n_4090 = n_821 & n_3681;
assign n_4091 = n_3651 ^ n_3682;
assign n_4092 = ~n_3683 & n_3684;
assign n_4093 = n_3685 ^ n_1917;
assign n_4094 = n_3685 & n_3686;
assign n_4095 = n_3687 ^ n_3657;
assign n_4096 = n_3688 ^ n_3324;
assign n_4097 = n_3689 ^ n_3034;
assign n_4098 = ~n_3689 & ~n_3690;
assign n_4099 = n_3691 ^ n_3356;
assign n_4100 = n_3693 ^ n_3310;
assign n_4101 = n_1784 & n_3695;
assign n_4102 = n_3696 ^ n_798;
assign n_4103 = ~n_3696 & ~n_3284;
assign n_4104 = ~n_3656 & ~n_3697;
assign n_4105 = ~n_3699 & ~n_3700;
assign n_4106 = n_3701 ^ n_3288;
assign n_4107 = n_3662 & ~n_3703;
assign n_4108 = n_1787 & n_3705;
assign n_4109 = n_1788 & n_3707;
assign n_4110 = ~n_3708 & ~n_3709;
assign n_4111 = ~n_3671 & ~n_3710;
assign n_4112 = ~n_3674 & ~n_3711;
assign n_4113 = ~n_3712 & ~n_3713;
assign n_4114 = n_3714 ^ n_3388;
assign n_4115 = n_3715 ^ n_3616;
assign n_4116 = n_3717 ^ n_3340;
assign n_4117 = n_3718 ^ n_3228;
assign n_4118 = ~n_3718 & ~n_3719;
assign n_4119 = n_3720 ^ n_800;
assign n_4120 = ~n_3720 & ~n_3698;
assign n_4121 = n_3721 ^ n_3315;
assign n_4122 = n_3701 & ~n_3722;
assign n_4123 = n_3723 ^ n_3232;
assign n_4124 = n_3702 & ~n_3724;
assign n_4125 = n_3725 ^ n_3318;
assign n_4126 = n_3727 ^ n_3235;
assign n_4127 = n_3727 & ~n_3728;
assign n_4128 = n_3729 ^ n_3321;
assign n_4129 = ~n_3665 & n_3730;
assign n_4130 = n_3733 ^ n_94;
assign n_4131 = ~n_3733 & ~n_3734;
assign n_4132 = n_3735 & n_3736;
assign n_4133 = n_3737 ^ n_3370;
assign n_4134 = ~n_3721 & ~n_3738;
assign n_4135 = n_3739 ^ n_2879;
assign n_4136 = n_3739 & ~n_3740;
assign n_4137 = n_3741 & ~n_3742;
assign n_4138 = n_3743 ^ n_3347;
assign n_4139 = ~n_3729 & n_3745;
assign n_4140 = n_3746 ^ n_3350;
assign n_4141 = ~n_3688 & ~n_3747;
assign n_4142 = n_3748 ^ n_3353;
assign n_4143 = n_3750 ^ n_3496;
assign n_4144 = n_3751 ^ n_3498;
assign n_4145 = n_3753 ^ n_3501;
assign n_4146 = n_3755 ^ n_3504;
assign n_4147 = n_3756 ^ n_3451;
assign n_4148 = n_3757 & n_3758;
assign n_4149 = n_3760 ^ n_3400;
assign n_4150 = n_3761 ^ n_2101;
assign n_4151 = n_3761 & n_3762;
assign n_4152 = ~n_3743 & n_3764;
assign n_4153 = n_3765 ^ n_2255;
assign n_4154 = n_3765 & n_3744;
assign n_4155 = n_3746 & ~n_3767;
assign n_4156 = n_3768 ^ n_2318;
assign n_4157 = n_3768 & n_3769;
assign n_4158 = n_3748 & ~n_3770;
assign n_4159 = n_3771 ^ n_3669;
assign n_4160 = n_3691 & ~n_3772;
assign n_4161 = n_3773 ^ n_3673;
assign n_4162 = n_3775 ^ n_3534;
assign n_4163 = n_3776 & n_3777;
assign n_4164 = n_3778 ^ n_3483;
assign n_4165 = n_3779 ^ n_3430;
assign n_4166 = n_3780 ^ n_3291;
assign n_4167 = n_3780 & ~n_3726;
assign n_4168 = n_3781 ^ n_2941;
assign n_4169 = ~n_3781 & n_3782;
assign n_4170 = n_3784 ^ n_3406;
assign n_4171 = n_3786 ^ n_3408;
assign n_4172 = n_3788 ^ n_3410;
assign n_4173 = n_3790 ^ n_3412;
assign n_4174 = n_3792 ^ n_3414;
assign n_4175 = n_3714 & ~n_3793;
assign n_4176 = n_3794 ^ n_3417;
assign n_4177 = ~n_3760 & n_3798;
assign n_4178 = n_3799 ^ n_102;
assign n_4179 = n_3799 & n_2099;
assign n_4180 = n_3800 ^ n_3460;
assign n_4181 = n_3801 ^ n_3207;
assign n_4182 = ~n_3801 & n_3783;
assign n_4183 = n_3784 & ~n_3802;
assign n_4184 = n_3803 ^ n_3209;
assign n_4185 = ~n_3785 & n_3804;
assign n_4186 = n_3786 & ~n_3805;
assign n_4187 = n_3806 ^ n_3297;
assign n_4188 = ~n_3806 & n_3787;
assign n_4189 = ~n_3788 & n_3807;
assign n_4190 = n_3808 ^ n_3299;
assign n_4191 = ~n_3789 & n_3809;
assign n_4192 = n_3790 & ~n_3810;
assign n_4193 = n_3811 ^ n_3301;
assign n_4194 = ~n_3791 & n_3812;
assign n_4195 = n_3792 & ~n_3813;
assign n_4196 = n_3814 ^ n_3303;
assign n_4197 = n_3814 & ~n_3815;
assign n_4198 = n_3816 ^ n_3444;
assign n_4199 = n_3794 & ~n_3817;
assign n_4200 = n_3818 ^ n_3306;
assign n_4201 = ~n_3818 & n_3819;
assign n_4202 = n_3820 ^ n_3447;
assign n_4203 = n_3821 ^ n_3279;
assign n_4204 = n_3821 & ~n_3716;
assign n_4205 = n_3822 ^ n_3450;
assign n_4206 = n_3824 ^ n_3594;
assign n_4207 = ~n_3779 & n_3825;
assign n_4208 = n_3826 ^ n_3515;
assign n_4209 = n_3828 ^ n_3517;
assign n_4210 = n_3829 ^ n_3490;
assign n_4211 = n_3830 ^ n_3238;
assign n_4212 = n_3830 & ~n_3731;
assign n_4213 = n_3831 ^ n_3003;
assign n_4214 = ~n_3831 & n_3732;
assign n_4215 = n_3833 ^ n_3466;
assign n_4216 = n_3835 ^ n_3468;
assign n_4217 = n_3836 ^ n_3470;
assign n_4218 = n_3816 & ~n_3838;
assign n_4219 = n_3839 ^ n_3473;
assign n_4220 = n_3820 & ~n_3841;
assign n_4221 = n_3842 ^ n_3476;
assign n_4222 = n_3843 ^ n_3337;
assign n_4223 = n_3843 & ~n_3844;
assign n_4224 = ~n_3845 & ~n_3846;
assign n_4225 = n_3756 & ~n_3847;
assign n_4226 = n_3850 ^ n_3313;
assign n_4227 = ~n_3850 & ~n_3851;
assign n_4228 = n_3852 ^ n_3625;
assign n_4229 = ~n_3800 & n_3854;
assign n_4230 = n_3855 ^ n_3546;
assign n_4231 = n_3856 ^ n_3520;
assign n_4232 = n_3857 ^ n_811;
assign n_4233 = ~n_3857 & ~n_3832;
assign n_4234 = ~n_3833 & n_3858;
assign n_4235 = n_3859 ^ n_813;
assign n_4236 = ~n_3859 & ~n_3834;
assign n_4237 = n_3860 & ~n_3861;
assign n_4238 = n_3862 ^ n_815;
assign n_4239 = ~n_3862 & ~n_3863;
assign n_4240 = n_3836 & ~n_3864;
assign n_4241 = n_3865 ^ n_817;
assign n_4242 = ~n_3865 & ~n_3837;
assign n_4243 = n_3866 ^ n_3332;
assign n_4244 = n_3866 & ~n_3752;
assign n_4245 = n_3839 & ~n_3867;
assign n_4246 = n_3868 ^ n_3249;
assign n_4247 = n_3840 & ~n_3869;
assign n_4248 = n_3870 ^ n_3335;
assign n_4249 = n_3754 & ~n_3871;
assign n_4250 = n_3842 & ~n_3872;
assign n_4251 = n_3873 ^ n_3506;
assign n_4252 = n_3874 ^ n_3507;
assign n_4253 = n_3875 ^ n_3368;
assign n_4254 = ~n_3875 & n_3848;
assign n_4255 = n_3876 ^ n_3509;
assign n_4256 = ~n_3778 & ~n_3878;
assign n_4257 = n_3881 ^ n_3514;
assign n_4258 = ~n_3829 & n_3883;
assign n_4259 = n_3885 ^ n_3549;
assign n_4260 = n_3886 ^ n_3550;
assign n_4261 = n_3887 ^ n_3327;
assign n_4262 = ~n_3749 & n_3888;
assign n_4263 = ~n_3889 & ~n_3890;
assign n_4264 = n_3891 ^ n_3525;
assign n_4265 = ~n_3751 & ~n_3892;
assign n_4266 = n_3893 ^ n_3527;
assign n_4267 = n_3753 & ~n_3894;
assign n_4268 = n_3895 ^ n_3530;
assign n_4269 = ~n_3755 & n_3897;
assign n_4270 = n_3898 ^ n_3280;
assign n_4271 = ~n_3898 & n_3899;
assign n_4272 = n_3900 & ~n_3901;
assign n_4273 = n_3874 & ~n_3902;
assign n_4274 = ~n_3876 & n_3903;
assign n_4275 = n_3904 ^ n_3398;
assign n_4276 = ~n_3904 & n_3877;
assign n_4277 = n_3905 ^ n_3539;
assign n_4278 = n_3906 ^ n_3373;
assign n_4279 = n_3880 & ~n_3907;
assign n_4280 = ~n_3881 & ~n_3908;
assign n_4281 = ~n_3909 & ~n_3910;
assign n_4282 = ~n_3828 & ~n_3912;
assign n_4283 = n_3913 & n_3914;
assign n_4284 = n_3915 ^ n_3580;
assign n_4285 = n_3891 & ~n_3916;
assign n_4286 = n_3917 ^ n_3096;
assign n_4287 = n_3917 & ~n_3692;
assign n_4288 = ~n_3893 & n_3918;
assign n_4289 = n_3919 ^ n_3360;
assign n_4290 = n_3919 & ~n_3920;
assign n_4291 = n_3921 ^ n_3557;
assign n_4292 = ~n_3895 & n_3922;
assign n_4293 = n_3923 ^ n_3363;
assign n_4294 = n_3896 & ~n_3924;
assign n_4295 = n_3925 ^ n_3560;
assign n_4296 = n_3926 ^ n_3561;
assign n_4297 = n_3775 & ~n_3927;
assign n_4298 = n_3928 ^ n_3395;
assign n_4299 = n_3797 & ~n_3929;
assign n_4300 = n_3930 ^ n_3312;
assign n_4301 = n_3930 & ~n_3931;
assign n_4302 = n_3932 ^ n_3565;
assign n_4303 = n_3934 & ~n_3935;
assign n_4304 = n_3936 ^ n_3428;
assign n_4305 = n_3936 & ~n_3937;
assign n_4306 = n_3938 ^ n_3569;
assign n_4307 = n_3940 ^ n_3403;
assign n_4308 = ~n_3911 & n_3941;
assign n_4309 = n_3942 ^ n_3573;
assign n_4310 = ~n_3855 & ~n_3943;
assign n_4311 = n_3944 ^ n_3491;
assign n_4312 = n_3944 & ~n_3884;
assign n_4313 = ~n_3885 & ~n_3946;
assign n_4314 = ~n_3886 & n_3947;
assign n_4315 = n_3950 ^ n_3611;
assign n_4316 = n_3951 ^ n_3359;
assign n_4317 = ~n_3951 & n_3774;
assign n_4318 = n_3952 ^ n_2623;
assign n_4319 = n_3952 & n_3585;
assign n_4320 = n_3921 & ~n_3953;
assign n_4321 = n_3954 ^ n_3587;
assign n_4322 = n_3955 & ~n_3956;
assign n_4323 = n_3926 & ~n_3957;
assign n_4324 = n_3958 ^ n_3591;
assign n_4325 = n_3960 ^ n_3593;
assign n_4326 = ~n_3932 & n_3961;
assign n_4327 = n_3962 ^ n_3342;
assign n_4328 = ~n_3962 & n_3933;
assign n_4329 = n_3963 ^ n_3596;
assign n_4330 = n_3938 & ~n_3965;
assign n_4331 = n_3966 ^ n_3458;
assign n_4332 = n_3966 & ~n_3967;
assign n_4333 = n_3968 ^ n_3600;
assign n_4334 = n_3970 & ~n_3971;
assign n_4335 = n_3973 ^ n_3605;
assign n_4336 = n_3974 ^ n_3606;
assign n_4337 = n_3975 ^ n_3522;
assign n_4338 = ~n_3975 & ~n_3976;
assign n_4339 = n_3977 ^ n_3608;
assign n_4340 = ~n_3915 & n_3978;
assign n_4341 = n_3979 ^ n_3553;
assign n_4342 = n_3949 & n_3980;
assign n_4343 = n_3983 ^ n_3642;
assign n_4344 = ~n_3954 & n_3985;
assign n_4345 = n_3986 ^ n_2688;
assign n_4346 = n_3986 & n_3987;
assign n_4347 = n_3989 ^ n_3619;
assign n_4348 = n_3990 & ~n_3991;
assign n_4349 = n_3992 ^ n_3423;
assign n_4350 = ~n_3992 & n_3959;
assign n_4351 = ~n_3960 & n_3993;
assign n_4352 = ~n_3824 & ~n_3994;
assign n_4353 = n_3995 ^ n_3624;
assign n_4354 = ~n_3963 & n_3996;
assign n_4355 = n_3997 ^ n_3372;
assign n_4356 = ~n_3997 & n_3964;
assign n_4357 = n_3998 ^ n_3627;
assign n_4358 = n_4000 & ~n_4001;
assign n_4359 = n_4002 ^ n_3488;
assign n_4360 = ~n_4002 & n_3969;
assign n_4361 = n_4003 ^ n_3631;
assign n_4362 = n_4004 ^ n_1331;
assign n_4363 = ~n_4004 & n_4005;
assign n_4364 = n_3973 & ~n_4006;
assign n_4365 = ~n_3974 & n_4007;
assign n_4366 = n_3977 & ~n_4009;
assign n_4367 = n_4010 ^ n_3638;
assign n_4368 = ~n_3950 & n_4011;
assign n_4369 = n_4013 ^ n_3583;
assign n_4370 = ~n_3982 & ~n_4014;
assign n_4371 = n_4015 ^ n_3643;
assign n_4372 = n_4016 ^ n_119;
assign n_4373 = n_4016 & ~n_3127;
assign n_4374 = n_3715 & ~n_4017;
assign n_4375 = n_4018 ^ n_3391;
assign n_4376 = ~n_3795 & n_4019;
assign n_4377 = n_4020 ^ n_93;
assign n_4378 = ~n_4020 & ~n_3796;
assign n_4379 = ~n_3989 & n_4021;
assign n_4380 = n_4023 ^ n_949;
assign n_4381 = ~n_1915 & ~n_4024;
assign n_4382 = n_4025 ^ n_97;
assign n_4383 = ~n_4025 & ~n_3823;
assign n_4384 = n_4026 ^ n_98;
assign n_4385 = ~n_4026 & ~n_3759;
assign n_4386 = n_3995 & ~n_4027;
assign n_4387 = ~n_4028 & ~n_4029;
assign n_4388 = n_4030 ^ n_101;
assign n_4389 = ~n_4030 & ~n_3853;
assign n_4390 = n_4031 & ~n_4032;
assign n_4391 = n_4033 ^ n_3402;
assign n_4392 = n_3999 & ~n_4034;
assign n_4393 = n_4035 ^ n_104;
assign n_4394 = ~n_4035 & ~n_3882;
assign n_4395 = n_4036 ^ n_3432;
assign n_4396 = ~n_3827 & ~n_4037;
assign n_4397 = n_4003 & ~n_4038;
assign n_4398 = n_4039 ^ n_3518;
assign n_4399 = n_4039 & ~n_4040;
assign n_4400 = n_4041 ^ n_108;
assign n_4401 = ~n_4041 & ~n_4042;
assign n_4402 = n_4043 ^ n_3548;
assign n_4403 = ~n_3945 & ~n_4044;
assign n_4404 = n_4046 ^ n_1394;
assign n_4405 = ~n_4046 & ~n_4008;
assign n_4406 = n_4047 ^ n_112;
assign n_4407 = ~n_4047 & ~n_3948;
assign n_4408 = n_4048 & ~n_4049;
assign n_4409 = n_4050 ^ n_1522;
assign n_4410 = ~n_4050 & ~n_4051;
assign n_4411 = n_4052 ^ n_115;
assign n_4412 = ~n_4052 & ~n_3981;
assign n_4413 = n_4053 ^ n_1586;
assign n_4414 = n_2531 & n_4054;
assign n_4415 = n_4055 & n_4056;
assign n_4416 = ~n_4015 & ~n_4057;
assign n_4417 = n_4059 ^ n_1713;
assign n_4418 = ~n_2656 & ~n_4060;
assign n_4419 = n_4061 ^ n_122;
assign n_4420 = n_4061 & ~n_2655;
assign y3 = ~n_4062;
assign n_4421 = n_3192 & ~n_4063;
assign n_4422 = n_4064 ^ n_1791;
assign n_4423 = n_4065 ^ n_163;
assign n_4424 = n_4067 ^ n_3194;
assign n_4425 = ~n_3682 & n_4068;
assign n_4426 = n_4069 ^ n_168;
assign n_4427 = n_1916 ^ n_4070;
assign n_4428 = n_3655 ^ n_4072;
assign n_4429 = n_3687 & ~n_4073;
assign n_4430 = n_4076 ^ n_188;
assign n_4431 = n_4078 ^ n_193;
assign n_4432 = n_3771 & ~n_4082;
assign n_4433 = n_3773 & n_4085;
assign n_4434 = n_4089 ^ n_228;
assign n_4435 = n_4090 ^ n_92;
assign n_4436 = n_4092 ^ n_2786;
assign n_4437 = n_3694 ^ n_4093;
assign n_4438 = n_4094 ^ n_3197;
assign n_4439 = n_4098 ^ n_812;
assign n_4440 = n_4101 ^ n_173;
assign n_4441 = n_4103 ^ n_798;
assign n_4442 = n_4104 ^ n_178;
assign n_4443 = n_4105 ^ n_183;
assign n_4444 = n_4107 ^ n_3204;
assign n_4445 = n_4108 ^ n_198;
assign n_4446 = n_4109 ^ n_203;
assign n_4447 = n_4110 ^ n_208;
assign n_4448 = n_4111 ^ n_213;
assign n_4449 = n_4112 ^ n_218;
assign n_4450 = n_4113 ^ n_223;
assign n_4451 = n_4118 ^ n_799;
assign n_4452 = n_4120 ^ n_800;
assign n_4453 = n_4121 ^ n_4075;
assign n_4454 = n_4122 ^ n_3259;
assign n_4455 = n_4124 ^ n_3260;
assign n_4456 = n_4125 ^ n_4077;
assign n_4457 = n_4127 ^ n_3206;
assign n_4458 = n_4128 ^ n_3704;
assign n_4459 = n_4129 ^ n_3294;
assign n_4460 = n_4131 ^ n_94;
assign n_4461 = n_4132 ^ n_884;
assign n_4462 = n_4134 ^ n_801;
assign n_4463 = n_4135 ^ n_4106;
assign n_4464 = n_4136 ^ n_3231;
assign n_4465 = n_4137 ^ n_3290;
assign n_4466 = n_4138 ^ n_3663;
assign n_4467 = n_4139 ^ n_3321;
assign n_4468 = n_4141 ^ n_810;
assign n_4469 = n_3678 ^ n_4145;
assign n_4470 = n_4148 ^ n_948;
assign n_4471 = n_4150 ^ n_4123;
assign n_4472 = n_4151 ^ n_3317;
assign n_4473 = n_4152 ^ n_3347;
assign n_4474 = n_4126 ^ n_4153;
assign n_4475 = n_4154 ^ n_3348;
assign n_4476 = n_4155 ^ n_3237;
assign n_4477 = n_4157 ^ n_3323;
assign n_4478 = n_4158 ^ n_3240;
assign n_4479 = n_4160 ^ n_3065;
assign n_4480 = n_4163 ^ n_1012;
assign n_4481 = n_4138 ^ n_4166;
assign n_4482 = n_4167 ^ n_3375;
assign n_4483 = n_4168 ^ n_4126;
assign n_4484 = n_4169 ^ n_2941;
assign n_4485 = n_4140 ^ n_4170;
assign n_4486 = n_4172 ^ n_4159;
assign n_4487 = n_4174 ^ n_4144;
assign n_4488 = n_4175 ^ n_3218;
assign n_4489 = n_4177 ^ n_1076;
assign n_4490 = n_4179 ^ n_102;
assign n_4491 = n_4182 ^ n_3207;
assign n_4492 = n_4183 ^ n_3265;
assign n_4493 = n_4184 ^ n_3706;
assign n_4494 = n_4185 ^ n_3407;
assign n_4495 = n_4186 ^ n_3380;
assign n_4496 = n_4142 ^ n_4187;
assign n_4497 = n_4188 ^ n_3297;
assign n_4498 = n_4189 ^ n_3410;
assign n_4499 = n_4084 ^ n_4190;
assign n_4500 = n_4191 ^ n_3411;
assign n_4501 = n_4192 ^ n_3271;
assign n_4502 = n_4194 ^ n_3413;
assign n_4503 = n_4195 ^ n_3273;
assign n_4504 = n_4197 ^ n_3387;
assign n_4505 = n_4199 ^ n_3276;
assign n_4506 = n_4115 ^ n_4200;
assign n_4507 = n_4201 ^ n_3306;
assign n_4508 = n_4203 ^ n_4146;
assign n_4509 = n_4204 ^ n_3279;
assign n_4510 = n_4205 ^ n_4100;
assign n_4511 = n_4207 ^ n_2098;
assign n_4512 = n_4184 ^ n_4211;
assign n_4513 = n_4212 ^ n_3435;
assign n_4514 = n_4213 ^ n_4171;
assign n_4515 = n_4214 ^ n_3003;
assign n_4516 = n_4097 ^ n_4215;
assign n_4517 = n_4216 ^ n_4173;
assign n_4518 = n_4216 ^ n_4143;
assign n_4519 = n_4218 ^ n_3416;
assign n_4520 = n_4219 ^ n_4176;
assign n_4521 = n_4220 ^ n_3307;
assign n_4522 = n_4146 ^ n_4221;
assign n_4523 = n_4203 ^ n_4221;
assign n_4524 = n_4223 ^ n_3421;
assign n_4525 = n_4224 ^ n_95;
assign n_4526 = n_4225 ^ n_3339;
assign n_4527 = n_4227 ^ n_99;
assign n_4528 = n_4229 ^ n_1203;
assign n_4529 = n_4232 ^ n_4081;
assign n_4530 = n_4233 ^ n_811;
assign n_4531 = n_4234 ^ n_3466;
assign n_4532 = n_4235 ^ n_4084;
assign n_4533 = n_4235 ^ n_4190;
assign n_4534 = n_4236 ^ n_813;
assign n_4535 = n_4237 ^ n_3300;
assign n_4536 = n_4086 ^ n_4238;
assign n_4537 = n_4239 ^ n_815;
assign n_4538 = n_4240 ^ n_3302;
assign n_4539 = n_4088 ^ n_4241;
assign n_4540 = n_4242 ^ n_817;
assign n_4541 = n_4244 ^ n_3472;
assign n_4542 = n_4245 ^ n_3305;
assign n_4543 = n_4247 ^ n_3446;
assign n_4544 = n_4248 ^ n_4202;
assign n_4545 = n_4249 ^ n_3250;
assign n_4546 = n_4250 ^ n_3448;
assign n_4547 = n_4254 ^ n_3368;
assign n_4548 = n_4256 ^ n_100;
assign n_4549 = n_4258 ^ n_2224;
assign n_4550 = n_4262 ^ n_3495;
assign n_4551 = n_4263 ^ n_814;
assign n_4552 = n_4264 ^ n_4193;
assign n_4553 = n_4264 ^ n_4161;
assign n_4554 = n_4265 ^ n_816;
assign n_4555 = n_4267 ^ n_3248;
assign n_4556 = n_4268 ^ n_4246;
assign n_4557 = n_4269 ^ n_3504;
assign n_4558 = n_4270 ^ n_4130;
assign n_4559 = n_4271 ^ n_3280;
assign n_4560 = n_4272 ^ n_3338;
assign n_4561 = n_4273 ^ n_3479;
assign n_4562 = n_4274 ^ n_3509;
assign n_4563 = n_4275 ^ n_4133;
assign n_4564 = n_4276 ^ n_3398;
assign n_4565 = n_4277 ^ n_4228;
assign n_4566 = n_4279 ^ n_3513;
assign n_4567 = n_4280 ^ n_103;
assign n_4568 = n_4281 ^ n_1204;
assign n_4569 = n_4282 ^ n_106;
assign n_4570 = n_4283 ^ n_1330;
assign n_4571 = n_4285 ^ n_3497;
assign n_4572 = n_4286 ^ n_4174;
assign n_4573 = n_4287 ^ n_3526;
assign n_4574 = n_4288 ^ n_3527;
assign n_4575 = n_4289 ^ n_4198;
assign n_4576 = n_4289 ^ n_4243;
assign n_4577 = n_4290 ^ n_3500;
assign n_4578 = n_4291 ^ n_3678;
assign n_4579 = n_4291 ^ n_4145;
assign n_4580 = n_4292 ^ n_3530;
assign n_4581 = n_4248 ^ n_4293;
assign n_4582 = n_4294 ^ n_3503;
assign n_4583 = n_4130 ^ n_4296;
assign n_4584 = n_4270 ^ n_4296;
assign n_4585 = n_4297 ^ n_3281;
assign n_4586 = n_4252 ^ n_4298;
assign n_4587 = n_4299 ^ n_3311;
assign n_4588 = n_4301 ^ n_3508;
assign n_4589 = n_4302 ^ n_4206;
assign n_4590 = n_4303 ^ n_3511;
assign n_4591 = n_4305 ^ n_3512;
assign n_4592 = n_4178 ^ n_4306;
assign n_4593 = n_4308 ^ n_3544;
assign n_4594 = n_4310 ^ n_107;
assign n_4595 = n_4312 ^ n_3547;
assign n_4596 = n_4313 ^ n_110;
assign n_4597 = n_4314 ^ n_2349;
assign n_4598 = n_4316 ^ n_4088;
assign n_4599 = n_4316 ^ n_4241;
assign n_4600 = n_4317 ^ n_3359;
assign n_4601 = n_4319 ^ n_3556;
assign n_4602 = n_4320 ^ n_3529;
assign n_4603 = n_4321 ^ n_4115;
assign n_4604 = n_4322 ^ n_3364;
assign n_4605 = n_4323 ^ n_3365;
assign n_4606 = n_4324 ^ n_4251;
assign n_4607 = n_4324 ^ n_4162;
assign n_4608 = n_4116 ^ n_4325;
assign n_4609 = n_4326 ^ n_3565;
assign n_4610 = n_4328 ^ n_3342;
assign n_4611 = n_4277 ^ n_4329;
assign n_4612 = n_4228 ^ n_4329;
assign n_4613 = n_4330 ^ n_3541;
assign n_4614 = n_4331 ^ n_4165;
assign n_4615 = n_4332 ^ n_3542;
assign n_4616 = n_4208 ^ n_4333;
assign n_4617 = n_4334 ^ n_3545;
assign n_4618 = n_4335 ^ n_4231;
assign n_4619 = n_4338 ^ n_111;
assign n_4620 = n_4340 ^ n_1457;
assign n_4621 = n_4342 ^ n_114;
assign n_4622 = n_4344 ^ n_3587;
assign n_4623 = n_4346 ^ n_3559;
assign n_4624 = n_4347 ^ n_4222;
assign n_4625 = n_4348 ^ n_3394;
assign n_4626 = n_4349 ^ n_4252;
assign n_4627 = n_4349 ^ n_4298;
assign n_4628 = n_4350 ^ n_3423;
assign n_4629 = n_4351 ^ n_3593;
assign n_4630 = n_4352 ^ n_1013;
assign n_4631 = n_4353 ^ n_4327;
assign n_4632 = n_4353 ^ n_4226;
assign n_4633 = n_4354 ^ n_3596;
assign n_4634 = n_4355 ^ n_4149;
assign n_4635 = n_4355 ^ n_4304;
assign n_4636 = n_4356 ^ n_3372;
assign n_4637 = n_4357 ^ n_4278;
assign n_4638 = n_4358 ^ n_3571;
assign n_4639 = n_4359 ^ n_4180;
assign n_4640 = n_4360 ^ n_3488;
assign n_4641 = n_4361 ^ n_4209;
assign n_4642 = n_4311 ^ n_4362;
assign n_4643 = n_4363 ^ n_1331;
assign n_4644 = n_4364 ^ n_3492;
assign n_4645 = n_4365 ^ n_3606;
assign n_4646 = n_4366 ^ n_3523;
assign n_4647 = n_4367 ^ n_4284;
assign n_4648 = n_4368 ^ n_1521;
assign n_4649 = n_4343 ^ n_4369;
assign n_4650 = n_4370 ^ n_117;
assign n_4651 = n_1649 ^ n_4371;
assign n_4652 = n_4373 ^ n_119;
assign n_4653 = n_4374 ^ n_3220;
assign n_4654 = n_4375 ^ n_4345;
assign n_4655 = n_4376 ^ n_3617;
assign n_4656 = n_4377 ^ n_4295;
assign n_4657 = n_4378 ^ n_93;
assign n_4658 = n_4379 ^ n_3619;
assign n_4659 = n_4381 ^ n_96;
assign n_4660 = n_4382 ^ n_4116;
assign n_4661 = n_4382 ^ n_4325;
assign n_4662 = n_4383 ^ n_97;
assign n_4663 = n_4384 ^ n_4255;
assign n_4664 = n_4385 ^ n_98;
assign n_4665 = n_4386 ^ n_3426;
assign n_4666 = n_4387 ^ n_1077;
assign n_4667 = n_4389 ^ n_101;
assign n_4668 = n_4390 ^ n_3598;
assign n_4669 = n_4391 ^ n_4257;
assign n_4670 = n_4392 ^ n_3599;
assign n_4671 = n_4393 ^ n_4208;
assign n_4672 = n_4393 ^ n_4333;
assign n_4673 = n_4394 ^ n_104;
assign n_4674 = n_4395 ^ n_4359;
assign n_4675 = n_4396 ^ n_105;
assign n_4676 = n_4397 ^ n_3489;
assign n_4677 = n_4398 ^ n_4210;
assign n_4678 = n_4399 ^ n_3603;
assign n_4679 = n_4400 ^ n_4311;
assign n_4680 = n_4401 ^ n_108;
assign n_4681 = n_4231 ^ n_4402;
assign n_4682 = n_4403 ^ n_109;
assign n_4683 = n_4404 ^ n_4337;
assign n_4684 = n_4405 ^ n_1394;
assign n_4685 = n_4406 ^ n_4339;
assign n_4686 = n_4407 ^ n_112;
assign n_4687 = n_4408 ^ n_3609;
assign n_4688 = n_4410 ^ n_1522;
assign n_4689 = n_4411 ^ n_3553;
assign n_4690 = n_4412 ^ n_115;
assign n_4691 = n_4414 ^ n_116;
assign n_4692 = n_4415 ^ n_1585;
assign n_4693 = n_4416 ^ n_118;
assign n_4694 = n_4418 ^ n_120;
assign n_4695 = n_4419 ^ n_1713;
assign n_4696 = n_4420 ^ n_122;
assign n_4697 = n_4421 ^ n_3647;
assign n_4698 = n_4423 ^ n_4066;
assign n_4699 = n_4424 ^ n_4091;
assign n_4700 = n_4425 ^ n_3224;
assign n_4701 = n_4426 ^ n_1916;
assign n_4702 = n_4426 ^ n_4070;
assign n_4703 = n_4429 ^ n_3229;
assign n_4704 = n_4430 ^ n_3763;
assign n_4705 = n_4430 ^ n_2192;
assign n_4706 = n_4432 ^ n_3326;
assign n_4707 = n_4433 ^ n_3244;
assign n_4708 = n_4434 ^ n_2687;
assign n_4709 = n_4435 ^ n_3988;
assign n_4710 = n_4435 ^ n_3589;
assign n_4711 = n_4436 ^ n_3694;
assign n_4712 = n_4436 ^ n_4093;
assign n_4713 = n_4438 ^ n_4102;
assign n_4714 = n_4439 ^ n_4261;
assign n_4715 = n_4440 ^ n_4071;
assign n_4716 = n_4440 ^ n_3654;
assign n_4717 = n_4441 ^ n_3655;
assign n_4718 = n_4443 ^ n_2100;
assign n_4719 = n_4444 ^ n_2193;
assign n_4720 = n_4445 ^ n_2317;
assign n_4721 = n_4446 ^ n_4096;
assign n_4722 = n_4448 ^ n_4099;
assign n_4723 = n_4449 ^ n_4087;
assign n_4724 = n_4449 ^ n_3675;
assign n_4725 = n_4451 ^ n_4442;
assign n_4726 = n_4451 ^ n_4119;
assign n_4727 = n_4452 ^ n_4074;
assign n_4728 = n_4452 ^ n_3658;
assign n_4729 = n_4454 ^ n_3660;
assign n_4730 = n_4455 ^ n_4125;
assign n_4731 = n_4455 ^ n_4077;
assign n_4732 = n_4457 ^ n_4128;
assign n_4733 = n_4460 ^ n_4022;
assign n_4734 = n_4460 ^ n_3620;
assign n_4735 = n_4443 ^ n_4462;
assign n_4736 = n_4464 ^ n_4454;
assign n_4737 = n_4444 ^ n_4465;
assign n_4738 = n_4466 ^ n_4166;
assign n_4739 = n_4467 ^ n_4140;
assign n_4740 = n_4467 ^ n_4170;
assign n_4741 = n_4468 ^ n_3667;
assign n_4742 = n_4473 ^ n_4431;
assign n_4743 = n_4475 ^ n_4181;
assign n_4744 = n_4477 ^ n_4171;
assign n_4745 = n_4478 ^ n_4447;
assign n_4746 = n_4479 ^ n_4086;
assign n_4747 = n_4480 ^ n_4164;
assign n_4748 = n_4466 & ~n_4481;
assign n_4749 = n_4473 ^ n_4482;
assign n_4750 = n_4483 ^ n_4153;
assign n_4751 = ~n_4483 & ~n_4474;
assign n_4752 = n_4484 ^ n_3766;
assign n_4753 = n_4484 ^ n_2256;
assign n_4754 = n_4488 ^ n_3984;
assign n_4755 = n_4488 ^ n_2624;
assign n_4756 = n_4490 ^ n_3373;
assign n_4757 = n_4445 ^ n_4491;
assign n_4758 = n_4492 ^ n_4476;
assign n_4759 = n_4492 ^ n_4459;
assign n_4760 = n_4493 ^ n_4211;
assign n_4761 = n_4494 ^ n_4080;
assign n_4762 = n_4494 ^ n_3666;
assign n_4763 = n_4495 ^ n_4142;
assign n_4764 = n_4495 ^ n_4187;
assign n_4765 = n_4497 ^ n_4097;
assign n_4766 = n_4439 ^ n_4498;
assign n_4767 = n_4500 ^ n_3672;
assign n_4768 = n_4503 ^ n_3676;
assign n_4769 = n_4450 ^ n_4504;
assign n_4770 = n_4434 ^ n_4505;
assign n_4771 = n_4508 ^ n_4221;
assign n_4772 = n_4493 & ~n_4512;
assign n_4773 = n_4513 ^ n_4446;
assign n_4774 = n_4477 ^ n_4514;
assign n_4775 = n_4468 ^ n_4515;
assign n_4776 = n_4517 ^ n_4143;
assign n_4777 = n_4517 & n_4518;
assign n_4778 = n_4522 & n_4523;
assign n_4779 = n_4525 ^ n_4461;
assign n_4780 = n_4526 ^ n_949;
assign n_4781 = n_4528 ^ n_1267;
assign n_4782 = n_4530 ^ n_4478;
assign n_4783 = n_4531 ^ n_4083;
assign n_4784 = n_4531 ^ n_3670;
assign n_4785 = n_4532 ^ n_4190;
assign n_4786 = ~n_4499 & n_4533;
assign n_4787 = n_4500 ^ n_4534;
assign n_4788 = n_4535 ^ n_4501;
assign n_4789 = n_4537 ^ n_4502;
assign n_4790 = n_4503 ^ n_4538;
assign n_4791 = n_4540 ^ n_4450;
assign n_4792 = n_4541 ^ n_4519;
assign n_4793 = n_4544 ^ n_4293;
assign n_4794 = n_4545 ^ n_4377;
assign n_4795 = n_4546 ^ n_4509;
assign n_4796 = n_4547 ^ n_4470;
assign n_4797 = n_4550 ^ n_4448;
assign n_4798 = n_4535 ^ n_4551;
assign n_4799 = n_4552 ^ n_4161;
assign n_4800 = n_4552 & n_4553;
assign n_4801 = n_4554 ^ n_4196;
assign n_4802 = n_4555 ^ n_4542;
assign n_4803 = n_4509 ^ n_4557;
assign n_4804 = n_4558 ^ n_4296;
assign n_4805 = n_4559 ^ n_4524;
assign n_4806 = n_4461 ^ n_4560;
assign n_4807 = n_4525 ^ n_4560;
assign n_4808 = n_4526 ^ n_4561;
assign n_4809 = n_4564 ^ n_3343;
assign n_4810 = n_4565 ^ n_4329;
assign n_4811 = n_4331 ^ n_4566;
assign n_4812 = n_4567 ^ n_4511;
assign n_4813 = n_4569 ^ n_4230;
assign n_4814 = n_4570 ^ n_4045;
assign n_4815 = n_4570 ^ n_3635;
assign n_4816 = n_4502 ^ n_4571;
assign n_4817 = n_4572 ^ n_4144;
assign n_4818 = ~n_4572 & ~n_4487;
assign n_4819 = n_4573 ^ n_4554;
assign n_4820 = n_4574 ^ n_4114;
assign n_4821 = n_4575 ^ n_4243;
assign n_4822 = ~n_4575 & n_4576;
assign n_4823 = n_4541 ^ n_4577;
assign n_4824 = n_4578 ^ n_4145;
assign n_4825 = n_4469 & ~n_4579;
assign n_4826 = n_4580 ^ n_3680;
assign n_4827 = n_4544 & ~n_4581;
assign n_4828 = ~n_4583 & ~n_4584;
assign n_4829 = n_4585 ^ n_4147;
assign n_4830 = n_4547 ^ n_4588;
assign n_4831 = n_4548 ^ n_4590;
assign n_4832 = n_4591 ^ n_4178;
assign n_4833 = n_4591 ^ n_4306;
assign n_4834 = n_4593 ^ n_4309;
assign n_4835 = n_4549 ^ n_4594;
assign n_4836 = n_4596 ^ n_4260;
assign n_4837 = n_4597 ^ n_1458;
assign n_4838 = n_4598 ^ n_4241;
assign n_4839 = n_4539 & n_4599;
assign n_4840 = n_4600 ^ n_4574;
assign n_4841 = n_4601 ^ n_4520;
assign n_4842 = n_4601 ^ n_4219;
assign n_4843 = n_4555 ^ n_4602;
assign n_4844 = n_4603 ^ n_4200;
assign n_4845 = ~n_4603 & n_4506;
assign n_4846 = n_4604 ^ n_4347;
assign n_4847 = n_4604 ^ n_4222;
assign n_4848 = n_4559 ^ n_4605;
assign n_4849 = n_4524 ^ n_4605;
assign n_4850 = n_4606 ^ n_4162;
assign n_4851 = ~n_4606 & n_4607;
assign n_4852 = n_4609 ^ n_4562;
assign n_4853 = n_4564 ^ n_4610;
assign n_4854 = n_4611 & n_4612;
assign n_4855 = n_4490 ^ n_4613;
assign n_4856 = n_4614 ^ n_4566;
assign n_4857 = n_4567 ^ n_4615;
assign n_4858 = n_4511 ^ n_4615;
assign n_4859 = n_4617 ^ n_4569;
assign n_4860 = n_4618 ^ n_4402;
assign n_4861 = n_1458 ^ n_4619;
assign n_4862 = n_4597 ^ n_4619;
assign n_4863 = n_4620 ^ n_4409;
assign n_4864 = n_4621 ^ n_4315;
assign n_4865 = n_4622 ^ n_4580;
assign n_4866 = n_4625 ^ n_4585;
assign n_4867 = n_4626 ^ n_4298;
assign n_4868 = ~n_4586 & n_4627;
assign n_4869 = n_4628 ^ n_4587;
assign n_4870 = n_4628 ^ n_4253;
assign n_4871 = n_4629 ^ n_3849;
assign n_4872 = n_4629 ^ n_3453;
assign n_4873 = n_4562 ^ n_4630;
assign n_4874 = n_4631 ^ n_4226;
assign n_4875 = ~n_4631 & ~n_4632;
assign n_4876 = n_4633 ^ n_3879;
assign n_4877 = n_4633 ^ n_3484;
assign n_4878 = n_4634 ^ n_4304;
assign n_4879 = ~n_4634 & ~n_4635;
assign n_4880 = n_4636 ^ n_4489;
assign n_4881 = n_4638 ^ n_4568;
assign n_4882 = n_1267 ^ n_4640;
assign n_4883 = n_4528 ^ n_4640;
assign n_4884 = n_4645 ^ n_4596;
assign n_4885 = n_4646 ^ n_2410;
assign n_4886 = n_4646 ^ n_1458;
assign n_4887 = n_4648 ^ n_4413;
assign n_4888 = n_4652 ^ n_4417;
assign n_4889 = n_4653 ^ n_4507;
assign n_4890 = n_4653 ^ n_4543;
assign n_4891 = n_4655 ^ n_4521;
assign n_4892 = n_4655 ^ n_4582;
assign n_4893 = n_4657 ^ n_1852;
assign n_4894 = n_4657 ^ n_885;
assign n_4895 = n_4658 ^ n_4205;
assign n_4896 = n_4658 ^ n_4100;
assign n_4897 = n_4659 ^ n_4300;
assign n_4898 = n_4660 ^ n_4325;
assign n_4899 = ~n_4608 & n_4661;
assign n_4900 = n_4662 ^ n_4384;
assign n_4901 = n_4664 ^ n_4275;
assign n_4902 = n_4665 ^ n_4480;
assign n_4903 = n_4666 ^ n_4548;
assign n_4904 = n_4666 ^ n_4590;
assign n_4905 = n_4667 ^ n_4636;
assign n_4906 = n_4667 ^ n_4489;
assign n_4907 = n_4668 ^ n_4391;
assign n_4908 = n_4670 ^ n_3939;
assign n_4909 = n_4670 ^ n_3543;
assign n_4910 = n_4671 ^ n_4333;
assign n_4911 = ~n_4616 & n_4672;
assign n_4912 = n_4638 ^ n_4673;
assign n_4913 = n_4674 ^ n_4180;
assign n_4914 = n_4674 & ~n_4639;
assign n_4915 = n_4675 ^ n_4361;
assign n_4916 = n_4676 ^ n_3972;
assign n_4917 = n_4676 ^ n_3574;
assign n_4918 = n_4678 ^ n_4549;
assign n_4919 = n_4679 ^ n_4362;
assign n_4920 = n_4679 & n_4642;
assign n_4921 = n_4680 ^ n_1331;
assign n_4922 = n_4680 ^ n_4595;
assign n_4923 = ~n_4618 & ~n_4681;
assign n_4924 = n_4682 ^ n_4644;
assign n_4925 = n_4682 ^ n_4336;
assign n_4926 = n_4339 ^ n_4684;
assign n_4927 = n_4685 ^ n_4684;
assign n_4928 = n_4686 ^ n_4367;
assign n_4929 = n_4686 ^ n_4284;
assign n_4930 = n_4687 ^ n_4620;
assign n_4931 = n_4688 ^ n_3553;
assign n_4932 = n_4688 ^ n_4411;
assign n_4933 = n_4690 ^ n_4012;
assign n_4934 = n_4690 ^ n_3612;
assign n_4935 = n_4691 ^ n_4343;
assign n_4936 = n_4692 ^ n_1649;
assign n_4937 = n_4692 ^ n_4371;
assign n_4938 = n_4693 ^ n_4058;
assign n_4939 = n_4693 ^ n_3644;
assign n_4940 = n_4419 ^ n_4694;
assign n_4941 = n_4695 ^ n_4694;
assign n_4942 = n_4696 ^ n_2720;
assign n_4943 = n_4696 ^ n_1777;
assign n_4944 = n_4697 ^ n_4422;
assign n_4945 = n_4697 ^ n_1791;
assign n_4946 = n_4701 ^ n_4070;
assign n_4947 = ~n_4427 & n_4702;
assign n_4948 = n_4703 ^ n_4453;
assign n_4949 = n_4703 ^ n_4121;
assign n_4950 = n_4704 ^ n_4472;
assign n_4951 = ~n_3763 & ~n_4705;
assign n_4952 = n_4707 ^ n_4217;
assign n_4953 = n_4708 ^ n_4505;
assign n_4954 = ~n_3988 & n_4710;
assign n_4955 = n_4711 ^ n_4093;
assign n_4956 = ~n_4437 & n_4712;
assign n_4957 = n_4713 ^ n_4715;
assign n_4958 = n_4102 ^ n_4715;
assign n_4959 = n_4438 ^ n_4715;
assign n_4960 = n_4071 & n_4716;
assign n_4961 = n_4717 ^ n_4072;
assign n_4962 = ~n_4717 & n_4428;
assign n_4963 = n_4718 ^ n_4462;
assign n_4964 = n_4719 ^ n_4465;
assign n_4965 = n_4720 ^ n_4491;
assign n_4966 = n_4707 ^ n_4723;
assign n_4967 = n_4087 & n_4724;
assign n_4968 = n_4725 ^ n_4119;
assign n_4969 = ~n_4725 & n_4726;
assign n_4970 = ~n_4074 & ~n_4728;
assign n_4971 = n_4730 ^ n_4077;
assign n_4972 = n_4456 & ~n_4731;
assign n_4973 = n_4732 ^ n_3704;
assign n_4974 = ~n_4732 & n_4458;
assign n_4975 = ~n_4022 & n_4734;
assign n_4976 = n_4718 & ~n_4735;
assign n_4977 = n_4736 ^ n_3660;
assign n_4978 = ~n_4736 & n_4729;
assign n_4979 = ~n_4719 & ~n_4737;
assign n_4980 = n_4739 ^ n_4170;
assign n_4981 = n_4485 & ~n_4740;
assign n_4982 = n_4741 ^ n_4515;
assign n_4983 = n_4742 ^ n_4482;
assign n_4984 = n_4514 & ~n_4744;
assign n_4985 = n_4746 ^ n_4238;
assign n_4986 = n_4746 & n_4536;
assign n_4987 = n_4748 ^ n_3663;
assign n_4988 = ~n_4742 & ~n_4749;
assign n_4989 = n_4751 ^ n_4153;
assign n_4990 = n_4743 ^ n_4752;
assign n_4991 = n_4475 ^ n_4752;
assign n_4992 = ~n_3766 & n_4753;
assign n_4993 = ~n_3984 & n_4755;
assign n_4994 = n_4756 ^ n_4613;
assign n_4995 = n_4720 & n_4757;
assign n_4996 = n_4758 ^ n_4459;
assign n_4997 = n_4758 & ~n_4759;
assign n_4998 = n_4080 & ~n_4762;
assign n_4999 = n_4763 ^ n_4187;
assign n_5000 = n_4496 & ~n_4764;
assign n_5001 = n_4765 ^ n_4215;
assign n_5002 = n_4765 & ~n_4516;
assign n_5003 = n_4766 ^ n_4261;
assign n_5004 = n_4766 & ~n_4714;
assign n_5005 = n_4767 ^ n_4534;
assign n_5006 = n_4768 ^ n_4538;
assign n_5007 = n_4708 & n_4770;
assign n_5008 = n_4772 ^ n_3706;
assign n_5009 = n_4773 ^ n_4096;
assign n_5010 = n_4773 & n_4721;
assign n_5011 = n_4741 & n_4775;
assign n_5012 = n_4777 ^ n_4173;
assign n_5013 = n_4778 ^ n_4146;
assign n_5014 = n_4779 ^ n_4560;
assign n_5015 = n_4780 ^ n_4561;
assign n_5016 = n_4781 ^ n_4640;
assign n_5017 = n_4782 ^ n_4447;
assign n_5018 = n_4782 & ~n_4745;
assign n_5019 = n_4706 ^ n_4783;
assign n_5020 = ~n_4083 & n_4784;
assign n_5021 = n_4786 ^ n_4084;
assign n_5022 = n_4767 & n_4787;
assign n_5023 = n_4788 ^ n_4551;
assign n_5024 = n_4789 ^ n_4571;
assign n_5025 = ~n_4768 & ~n_4790;
assign n_5026 = n_4791 ^ n_4504;
assign n_5027 = ~n_4791 & ~n_4769;
assign n_5028 = n_4792 ^ n_4577;
assign n_5029 = n_4794 ^ n_4295;
assign n_5030 = n_4794 & ~n_4656;
assign n_5031 = n_4795 ^ n_4557;
assign n_5032 = n_4796 ^ n_4588;
assign n_5033 = n_4797 ^ n_4099;
assign n_5034 = n_4797 & ~n_4722;
assign n_5035 = n_4788 & n_4798;
assign n_5036 = n_4800 ^ n_4193;
assign n_5037 = n_4802 ^ n_4602;
assign n_5038 = n_4795 & ~n_4803;
assign n_5039 = n_4805 ^ n_4605;
assign n_5040 = n_4806 & n_4807;
assign n_5041 = ~n_4780 & ~n_4808;
assign n_5042 = n_4809 ^ n_4610;
assign n_5043 = ~n_4614 & ~n_4811;
assign n_5044 = n_4812 ^ n_4615;
assign n_5045 = n_4814 ^ n_4259;
assign n_5046 = n_4045 & ~n_4815;
assign n_5047 = n_4789 & n_4816;
assign n_5048 = n_4818 ^ n_4144;
assign n_5049 = n_4819 ^ n_4196;
assign n_5050 = n_4819 & ~n_4801;
assign n_5051 = n_4822 ^ n_4243;
assign n_5052 = ~n_4792 & n_4823;
assign n_5053 = n_4825 ^ n_3678;
assign n_5054 = n_4827 ^ n_4202;
assign n_5055 = n_4828 ^ n_4130;
assign n_5056 = n_4796 & ~n_4830;
assign n_5057 = n_4832 ^ n_4306;
assign n_5058 = n_4592 & ~n_4833;
assign n_5059 = n_4837 ^ n_4619;
assign n_5060 = n_4839 ^ n_4088;
assign n_5061 = n_4840 ^ n_4114;
assign n_5062 = ~n_4840 & n_4820;
assign n_5063 = n_4520 & ~n_4842;
assign n_5064 = n_4802 & ~n_4843;
assign n_5065 = n_4845 ^ n_4200;
assign n_5066 = n_4846 ^ n_4222;
assign n_5067 = n_4624 & ~n_4847;
assign n_5068 = n_4848 & ~n_4849;
assign n_5069 = n_4851 ^ n_4162;
assign n_5070 = n_4852 ^ n_4630;
assign n_5071 = ~n_4809 & ~n_4853;
assign n_5072 = n_4854 ^ n_4277;
assign n_5073 = ~n_4756 & n_4855;
assign n_5074 = ~n_4857 & ~n_4858;
assign n_5075 = n_4859 ^ n_4230;
assign n_5076 = n_4859 & n_4813;
assign n_5077 = ~n_4861 & n_4862;
assign n_5078 = n_4865 ^ n_3680;
assign n_5079 = ~n_4865 & n_4826;
assign n_5080 = n_4866 ^ n_4147;
assign n_5081 = ~n_4866 & n_4829;
assign n_5082 = n_4868 ^ n_4349;
assign n_5083 = n_4869 ^ n_4253;
assign n_5084 = ~n_4869 & n_4870;
assign n_5085 = n_4871 ^ n_4589;
assign n_5086 = n_4871 ^ n_4302;
assign n_5087 = ~n_3849 & ~n_4872;
assign n_5088 = n_4852 & n_4873;
assign n_5089 = n_4875 ^ n_4226;
assign n_5090 = n_4876 ^ n_4388;
assign n_5091 = n_3879 & ~n_4877;
assign n_5092 = n_4879 ^ n_4149;
assign n_5093 = n_4881 ^ n_4673;
assign n_5094 = n_4882 & ~n_4883;
assign n_5095 = n_4884 ^ n_4260;
assign n_5096 = n_4884 & n_4836;
assign n_5097 = n_2410 & n_4886;
assign n_5098 = n_4889 ^ n_4543;
assign n_5099 = n_4889 & ~n_4890;
assign n_5100 = n_4891 ^ n_4582;
assign n_5101 = ~n_4891 & n_4892;
assign n_5102 = n_1852 & n_4894;
assign n_5103 = n_4895 ^ n_4100;
assign n_5104 = n_4510 & n_4896;
assign n_5105 = n_4899 ^ n_4116;
assign n_5106 = n_4900 ^ n_4255;
assign n_5107 = ~n_4900 & ~n_4663;
assign n_5108 = n_4901 ^ n_4133;
assign n_5109 = n_4901 & ~n_4563;
assign n_5110 = n_4902 ^ n_4164;
assign n_5111 = ~n_4902 & ~n_4747;
assign n_5112 = n_4903 ^ n_4590;
assign n_5113 = ~n_4831 & n_4904;
assign n_5114 = n_4905 ^ n_4489;
assign n_5115 = n_4880 & n_4906;
assign n_5116 = n_4907 ^ n_4257;
assign n_5117 = ~n_4907 & ~n_4669;
assign n_5118 = ~n_3939 & ~n_4909;
assign n_5119 = n_4911 ^ n_4208;
assign n_5120 = ~n_4881 & n_4912;
assign n_5121 = n_4914 ^ n_4180;
assign n_5122 = n_4915 ^ n_4209;
assign n_5123 = n_4915 & ~n_4641;
assign n_5124 = n_4916 ^ n_4677;
assign n_5125 = n_4916 ^ n_4398;
assign n_5126 = ~n_3972 & ~n_4917;
assign n_5127 = n_4918 ^ n_4594;
assign n_5128 = ~n_4918 & ~n_4835;
assign n_5129 = n_4920 ^ n_4362;
assign n_5130 = n_4921 ^ n_4595;
assign n_5131 = n_4921 & n_4922;
assign n_5132 = n_4923 ^ n_4335;
assign n_5133 = n_4924 ^ n_4336;
assign n_5134 = n_4924 & ~n_4925;
assign n_5135 = ~n_4685 & n_4926;
assign n_5136 = n_4928 ^ n_4284;
assign n_5137 = ~n_4647 & ~n_4929;
assign n_5138 = n_4930 ^ n_4409;
assign n_5139 = ~n_4930 & ~n_4863;
assign n_5140 = n_4931 ^ n_4411;
assign n_5141 = ~n_4689 & ~n_4932;
assign n_5142 = n_4933 ^ n_4887;
assign n_5143 = n_4933 ^ n_4648;
assign n_5144 = ~n_4012 & n_4934;
assign n_5145 = n_4935 ^ n_4369;
assign n_5146 = ~n_4935 & n_4649;
assign n_5147 = n_4936 ^ n_4371;
assign n_5148 = ~n_4651 & n_4937;
assign n_5149 = n_4938 ^ n_4372;
assign n_5150 = ~n_4058 & n_4939;
assign n_5151 = ~n_4695 & n_4940;
assign n_5152 = ~n_2720 & ~n_4943;
assign y4 = ~n_4944;
assign n_5153 = n_4422 & n_4945;
assign n_5154 = n_4946 ^ n_4700;
assign n_5155 = n_4947 ^ n_1916;
assign n_5156 = n_4727 ^ n_4948;
assign n_5157 = n_4453 & n_4949;
assign n_5158 = n_4951 ^ n_3346;
assign n_5159 = n_4952 ^ n_4723;
assign n_5160 = n_4954 ^ x33;
assign n_5161 = n_4956 ^ n_3694;
assign n_5162 = n_4958 & n_4959;
assign n_5163 = n_4960 ^ n_3227;
assign n_5164 = n_4117 ^ n_4961;
assign n_5165 = n_4962 ^ n_4072;
assign n_5166 = n_4079 ^ n_4965;
assign n_5167 = n_4952 & n_4966;
assign n_5168 = n_4967 ^ n_3358;
assign n_5169 = n_4968 ^ n_4095;
assign n_5170 = n_4969 ^ n_4119;
assign n_5171 = n_4970 ^ n_3230;
assign n_5172 = n_4972 ^ n_4125;
assign n_5173 = n_4974 ^ n_3704;
assign n_5174 = n_4975 ^ n_885;
assign n_5175 = n_4976 ^ n_2100;
assign n_5176 = n_4978 ^ n_3660;
assign n_5177 = n_4979 ^ n_2193;
assign n_5178 = n_4981 ^ n_4140;
assign n_5179 = n_4984 ^ n_4213;
assign n_5180 = n_4799 ^ n_4985;
assign n_5181 = n_4986 ^ n_4238;
assign n_5182 = n_4983 ^ n_4987;
assign n_5183 = n_4988 ^ n_4431;
assign n_5184 = n_4989 ^ n_4973;
assign n_5185 = n_4743 & n_4991;
assign n_5186 = n_4992 ^ n_3349;
assign n_5187 = n_4993 ^ n_3586;
assign n_5188 = n_4995 ^ n_2317;
assign n_5189 = n_4996 ^ n_4760;
assign n_5190 = n_4997 ^ n_4476;
assign n_5191 = n_4998 ^ n_3352;
assign n_5192 = n_5000 ^ n_4142;
assign n_5193 = n_5002 ^ n_4215;
assign n_5194 = n_5003 ^ n_4785;
assign n_5195 = n_5004 ^ n_4261;
assign n_5196 = n_5005 ^ n_4776;
assign n_5197 = n_5007 ^ n_2687;
assign n_5198 = n_5008 ^ n_4774;
assign n_5199 = n_4761 ^ n_5009;
assign n_5200 = n_5010 ^ n_4096;
assign n_5201 = n_5011 ^ n_3667;
assign n_5202 = n_4893 ^ n_5013;
assign n_5203 = n_5017 ^ n_5001;
assign n_5204 = n_5018 ^ n_4447;
assign n_5205 = n_5020 ^ n_3355;
assign n_5206 = n_5022 ^ n_3672;
assign n_5207 = n_5023 ^ n_4799;
assign n_5208 = n_5023 ^ n_4985;
assign n_5209 = n_5025 ^ n_3676;
assign n_5210 = n_5027 ^ n_4504;
assign n_5211 = n_5028 ^ n_4841;
assign n_5212 = n_5029 ^ n_4771;
assign n_5213 = n_5030 ^ n_4295;
assign n_5214 = n_5033 ^ n_5021;
assign n_5215 = n_5034 ^ n_4099;
assign n_5216 = n_5035 ^ n_4501;
assign n_5217 = n_5036 ^ n_4817;
assign n_5218 = n_5037 ^ n_4953;
assign n_5219 = n_5038 ^ n_4546;
assign n_5220 = n_5040 ^ n_4461;
assign n_5221 = n_5041 ^ n_949;
assign n_5222 = n_4527 ^ n_5042;
assign n_5223 = n_5043 ^ n_4165;
assign n_5224 = n_4908 ^ n_5044;
assign n_5225 = n_5046 ^ n_1394;
assign n_5226 = n_5047 ^ n_4571;
assign n_5227 = n_5049 ^ n_5006;
assign n_5228 = n_5049 ^ n_5048;
assign n_5229 = n_5050 ^ n_4196;
assign n_5230 = n_4754 ^ n_5051;
assign n_5231 = n_5052 ^ n_4577;
assign n_5232 = n_5053 ^ n_4844;
assign n_5233 = n_4709 ^ n_5054;
assign n_5234 = n_5055 ^ n_5039;
assign n_5235 = n_5056 ^ n_4470;
assign n_5236 = n_5058 ^ n_4178;
assign n_5237 = n_5059 ^ n_4927;
assign n_5238 = n_4318 ^ n_5060;
assign n_5239 = n_5026 ^ n_5061;
assign n_5240 = n_5062 ^ n_4114;
assign n_5241 = n_5063 ^ n_4176;
assign n_5242 = n_5064 ^ n_4542;
assign n_5243 = n_5066 ^ n_4804;
assign n_5244 = n_5067 ^ n_4347;
assign n_5245 = n_5068 ^ n_4559;
assign n_5246 = n_5069 ^ n_4867;
assign n_5247 = n_5071 ^ n_3343;
assign n_5248 = n_5073 ^ n_3373;
assign n_5249 = n_5074 ^ n_4567;
assign n_5250 = n_5076 ^ n_4230;
assign n_5251 = n_5077 ^ n_1458;
assign n_5252 = n_5065 ^ n_5078;
assign n_5253 = n_5079 ^ n_3680;
assign n_5254 = n_5014 ^ n_5080;
assign n_5255 = n_5081 ^ n_4147;
assign n_5256 = n_5082 ^ n_4898;
assign n_5257 = n_5083 ^ n_5015;
assign n_5258 = n_5084 ^ n_4253;
assign n_5259 = ~n_4589 & n_5086;
assign n_5260 = n_5087 ^ n_3313;
assign n_5261 = n_5088 ^ n_4609;
assign n_5262 = n_5091 ^ n_3343;
assign n_5263 = n_5094 ^ n_1267;
assign n_5264 = n_5096 ^ n_4260;
assign n_5265 = n_5097 ^ n_113;
assign n_5266 = n_5098 ^ n_4793;
assign n_5267 = n_5099 ^ n_4507;
assign n_5268 = n_5100 ^ n_4709;
assign n_5269 = n_5100 ^ n_5054;
assign n_5270 = n_5101 ^ n_4582;
assign n_5271 = n_5102 ^ x33;
assign n_5272 = n_5103 ^ n_4850;
assign n_5273 = n_5104 ^ n_4205;
assign n_5274 = n_5106 ^ n_5105;
assign n_5275 = n_5107 ^ n_4255;
assign n_5276 = n_5108 ^ n_4874;
assign n_5277 = n_5109 ^ n_4133;
assign n_5278 = n_5110 ^ n_5089;
assign n_5279 = n_5111 ^ n_4164;
assign n_5280 = n_5112 ^ n_5072;
assign n_5281 = n_5113 ^ n_4548;
assign n_5282 = n_5114 ^ n_5092;
assign n_5283 = n_5115 ^ n_4636;
assign n_5284 = n_5116 ^ n_4856;
assign n_5285 = n_5117 ^ n_4257;
assign n_5286 = n_5118 ^ n_3403;
assign n_5287 = n_5119 ^ n_5093;
assign n_5288 = n_5119 ^ n_4913;
assign n_5289 = n_5120 ^ n_4568;
assign n_5290 = n_5121 ^ n_5016;
assign n_5291 = n_5016 ^ n_5122;
assign n_5292 = n_5123 ^ n_4209;
assign n_5293 = ~n_4677 & n_5125;
assign n_5294 = n_5126 ^ n_1267;
assign n_5295 = n_5128 ^ n_4594;
assign n_5296 = n_5129 ^ n_4860;
assign n_5297 = n_4643 ^ n_5130;
assign n_5298 = n_5131 ^ n_1331;
assign n_5299 = n_5133 ^ n_5132;
assign n_5300 = n_5134 ^ n_4336;
assign n_5301 = n_5135 ^ n_4406;
assign n_5302 = n_5137 ^ n_4367;
assign n_5303 = n_5139 ^ n_4409;
assign n_5304 = n_5140 ^ n_4864;
assign n_5305 = n_5140 ^ n_4621;
assign n_5306 = n_5141 ^ n_3553;
assign n_5307 = n_4887 & ~n_5143;
assign n_5308 = n_5144 ^ n_3583;
assign n_5309 = n_5146 ^ n_4369;
assign n_5310 = n_5147 ^ n_4650;
assign n_5311 = n_5148 ^ n_1649;
assign n_5312 = n_5150 ^ n_1649;
assign n_5313 = n_5151 ^ n_1713;
assign n_5314 = n_5152 ^ n_123;
assign n_5315 = n_5153 ^ n_4697;
assign n_5316 = n_5155 ^ n_4955;
assign n_5317 = n_5157 ^ n_4075;
assign n_5318 = n_5158 ^ n_4964;
assign n_5319 = n_4817 ^ n_5159;
assign n_5320 = n_5036 ^ n_5159;
assign n_5321 = n_5160 ^ n_5031;
assign n_5322 = n_5161 ^ n_4957;
assign n_5323 = n_5162 ^ n_4102;
assign n_5324 = n_5163 ^ n_4117;
assign n_5325 = n_5163 ^ n_4961;
assign n_5326 = n_4968 ^ n_5165;
assign n_5327 = n_5167 ^ n_4217;
assign n_5328 = n_4266 ^ n_5168;
assign n_5329 = n_5169 ^ n_5165;
assign n_5330 = n_5170 ^ n_4727;
assign n_5331 = n_5171 ^ n_4463;
assign n_5332 = n_5171 ^ n_4135;
assign n_5333 = n_5158 ^ n_5172;
assign n_5334 = n_5173 ^ n_4980;
assign n_5335 = n_4380 ^ n_5174;
assign n_5336 = n_5175 ^ n_4471;
assign n_5337 = n_5175 ^ n_4150;
assign n_5338 = n_5176 ^ n_4950;
assign n_5339 = n_5176 ^ n_4472;
assign n_5340 = n_5177 ^ n_4983;
assign n_5341 = n_4156 ^ n_5178;
assign n_5342 = n_5181 ^ n_5024;
assign n_5343 = n_5183 ^ n_4989;
assign n_5344 = n_5185 ^ n_4181;
assign n_5345 = n_5186 ^ n_4079;
assign n_5346 = n_5186 ^ n_4965;
assign n_5347 = n_5187 ^ n_5037;
assign n_5348 = n_5188 ^ n_4156;
assign n_5349 = n_5188 ^ n_5178;
assign n_5350 = n_5190 ^ n_4761;
assign n_5351 = n_5190 ^ n_5009;
assign n_5352 = n_5191 ^ n_4529;
assign n_5353 = n_5191 ^ n_4232;
assign n_5354 = n_5192 ^ n_5017;
assign n_5355 = n_5193 ^ n_5003;
assign n_5356 = n_5195 ^ n_5005;
assign n_5357 = n_5197 ^ n_5065;
assign n_5358 = n_5197 ^ n_5078;
assign n_5359 = n_5200 ^ n_4982;
assign n_5360 = n_5200 ^ n_5179;
assign n_5361 = n_5201 ^ n_4486;
assign n_5362 = n_5201 ^ n_4172;
assign n_5363 = n_5204 ^ n_4706;
assign n_5364 = n_5204 ^ n_4783;
assign n_5365 = n_5205 ^ n_5033;
assign n_5366 = n_5205 ^ n_5021;
assign n_5367 = n_5206 ^ n_5012;
assign n_5368 = n_5207 ^ n_4985;
assign n_5369 = ~n_5180 & n_5208;
assign n_5370 = n_5209 ^ n_4318;
assign n_5371 = n_5209 ^ n_5060;
assign n_5372 = n_5210 ^ n_4754;
assign n_5373 = n_5210 ^ n_5051;
assign n_5374 = n_5213 ^ n_4893;
assign n_5375 = n_5213 ^ n_5013;
assign n_5376 = n_5215 ^ n_5206;
assign n_5377 = n_5181 ^ n_5216;
assign n_5378 = n_5217 ^ n_5159;
assign n_5379 = n_5219 ^ n_4733;
assign n_5380 = n_5220 ^ n_4897;
assign n_5381 = n_5220 ^ n_4659;
assign n_5382 = n_5221 ^ n_5032;
assign n_5383 = n_5225 ^ n_4683;
assign n_5384 = n_5225 ^ n_4337;
assign n_5385 = n_5226 ^ n_4266;
assign n_5386 = n_5226 ^ n_5168;
assign n_5387 = n_5227 ^ n_5048;
assign n_5388 = ~n_5227 & n_5228;
assign n_5389 = n_5229 ^ n_5026;
assign n_5390 = n_5231 ^ n_4556;
assign n_5391 = n_5231 ^ n_4246;
assign n_5392 = n_5236 ^ n_4994;
assign n_5393 = n_5240 ^ n_5028;
assign n_5394 = n_5241 ^ n_5053;
assign n_5395 = n_5242 ^ n_4654;
assign n_5396 = n_5242 ^ n_4375;
assign n_5397 = n_5244 ^ n_5234;
assign n_5398 = n_5244 ^ n_5055;
assign n_5399 = n_5245 ^ n_4380;
assign n_5400 = n_5245 ^ n_5174;
assign n_5401 = n_5247 ^ n_5090;
assign n_5402 = n_5247 ^ n_4876;
assign n_5403 = n_5248 ^ n_4908;
assign n_5404 = n_5248 ^ n_5044;
assign n_5405 = n_5249 ^ n_4307;
assign n_5406 = n_5251 ^ n_4885;
assign n_5407 = n_4623 ^ n_5253;
assign n_5408 = n_5015 ^ n_5255;
assign n_5409 = n_5257 ^ n_5255;
assign n_5410 = n_5032 ^ n_5258;
assign n_5411 = n_5221 ^ n_5258;
assign n_5412 = n_5259 ^ n_4206;
assign n_5413 = n_5260 ^ n_5235;
assign n_5414 = n_5260 ^ n_5070;
assign n_5415 = n_5261 ^ n_4527;
assign n_5416 = n_5261 ^ n_5042;
assign n_5417 = n_5262 ^ n_5114;
assign n_5418 = n_5262 ^ n_5092;
assign n_5419 = n_5264 ^ n_5059;
assign n_5420 = n_5265 ^ n_4341;
assign n_5421 = n_5267 ^ n_4623;
assign n_5422 = n_5267 ^ n_5253;
assign n_5423 = n_5268 ^ n_5054;
assign n_5424 = n_5233 & ~n_5269;
assign n_5425 = n_5270 ^ n_5160;
assign n_5426 = n_4733 ^ n_5271;
assign n_5427 = n_5219 ^ n_5271;
assign n_5428 = n_5273 ^ n_5014;
assign n_5429 = n_5275 ^ n_5108;
assign n_5430 = n_5277 ^ n_5110;
assign n_5431 = n_5277 ^ n_5089;
assign n_5432 = n_5279 ^ n_5112;
assign n_5433 = n_5281 ^ n_4637;
assign n_5434 = n_5281 ^ n_4357;
assign n_5435 = n_5283 ^ n_5236;
assign n_5436 = n_5285 ^ n_5223;
assign n_5437 = n_5285 ^ n_4910;
assign n_5438 = n_4307 ^ n_5286;
assign n_5439 = n_5249 ^ n_5286;
assign n_5440 = n_5287 ^ n_4913;
assign n_5441 = n_5287 & ~n_5288;
assign n_5442 = n_5289 ^ n_4834;
assign n_5443 = n_5289 ^ n_4593;
assign n_5444 = n_5290 ^ n_5122;
assign n_5445 = n_5290 & n_5291;
assign n_5446 = n_5292 ^ n_5263;
assign n_5447 = n_5292 ^ n_5075;
assign n_5448 = n_5293 ^ n_4210;
assign n_5449 = n_5294 ^ n_5250;
assign n_5450 = n_5294 ^ n_5127;
assign n_5451 = n_5295 ^ n_4643;
assign n_5452 = n_5295 ^ n_5130;
assign n_5453 = n_5298 ^ n_5045;
assign n_5454 = n_5298 ^ n_4814;
assign n_5455 = n_5300 ^ n_5095;
assign n_5456 = n_4885 ^ n_5301;
assign n_5457 = n_5251 ^ n_5301;
assign n_5458 = n_5265 ^ n_5302;
assign n_5459 = n_5304 ^ n_5303;
assign n_5460 = n_4864 & n_5305;
assign n_5461 = n_5306 ^ n_5142;
assign n_5462 = n_5307 ^ n_4413;
assign n_5463 = n_5308 ^ n_5145;
assign n_5464 = n_5147 ^ n_5309;
assign n_5465 = n_5310 ^ n_5309;
assign n_5466 = n_5311 ^ n_5149;
assign n_5467 = n_5311 ^ n_4938;
assign n_5468 = n_5312 ^ n_4888;
assign n_5469 = n_5312 ^ n_4652;
assign n_5470 = n_5313 ^ n_4942;
assign n_5471 = n_5314 ^ n_3190;
assign n_5472 = n_5315 ^ n_4698;
assign n_5473 = n_5315 ^ n_4066;
assign n_5474 = n_5317 ^ n_4963;
assign n_5475 = n_5318 ^ n_5172;
assign n_5476 = n_5319 & n_5320;
assign n_5477 = n_5324 ^ n_4961;
assign n_5478 = n_5164 & n_5325;
assign n_5479 = ~n_5169 & ~n_5326;
assign n_5480 = n_5327 ^ n_4838;
assign n_5481 = n_5330 ^ n_4948;
assign n_5482 = n_5330 & n_5156;
assign n_5483 = n_5317 ^ n_5331;
assign n_5484 = n_4463 & ~n_5332;
assign n_5485 = ~n_5318 & ~n_5333;
assign n_5486 = n_5336 ^ n_4977;
assign n_5487 = ~n_4471 & ~n_5337;
assign n_5488 = n_4971 ^ n_5338;
assign n_5489 = n_4950 & ~n_5339;
assign n_5490 = n_5340 ^ n_4987;
assign n_5491 = ~n_5340 & ~n_5182;
assign n_5492 = n_5343 ^ n_4973;
assign n_5493 = ~n_5343 & ~n_5184;
assign n_5494 = n_5344 ^ n_5334;
assign n_5495 = n_5344 ^ n_4980;
assign n_5496 = n_5344 ^ n_5173;
assign n_5497 = n_5345 ^ n_4965;
assign n_5498 = n_5166 & ~n_5346;
assign n_5499 = n_5347 ^ n_4953;
assign n_5500 = ~n_5347 & n_5218;
assign n_5501 = n_5348 ^ n_5178;
assign n_5502 = ~n_5341 & n_5349;
assign n_5503 = n_5350 ^ n_5009;
assign n_5504 = n_5199 & ~n_5351;
assign n_5505 = n_5352 ^ n_4999;
assign n_5506 = n_4529 & n_5353;
assign n_5507 = n_5354 ^ n_5001;
assign n_5508 = ~n_5354 & ~n_5203;
assign n_5509 = n_5355 ^ n_4785;
assign n_5510 = n_5355 & ~n_5194;
assign n_5511 = n_5356 ^ n_4776;
assign n_5512 = n_5356 & n_5196;
assign n_5513 = n_5357 ^ n_5078;
assign n_5514 = n_5252 & n_5358;
assign n_5515 = n_5359 ^ n_5179;
assign n_5516 = ~n_5359 & n_5360;
assign n_5517 = n_4486 & n_5362;
assign n_5518 = n_5363 ^ n_4783;
assign n_5519 = ~n_5019 & ~n_5364;
assign n_5520 = n_5365 ^ n_5021;
assign n_5521 = n_5214 & n_5366;
assign n_5522 = n_5369 ^ n_4799;
assign n_5523 = n_5370 ^ n_5060;
assign n_5524 = n_5238 & ~n_5371;
assign n_5525 = n_5372 ^ n_5051;
assign n_5526 = ~n_5230 & ~n_5373;
assign n_5527 = n_5374 ^ n_5013;
assign n_5528 = ~n_5202 & ~n_5375;
assign n_5529 = n_5376 ^ n_5012;
assign n_5530 = ~n_5376 & n_5367;
assign n_5531 = n_5377 ^ n_5024;
assign n_5532 = n_5377 & n_5342;
assign n_5533 = n_5379 ^ n_5271;
assign n_5534 = n_5380 ^ n_5256;
assign n_5535 = n_5380 ^ n_5082;
assign n_5536 = ~n_4897 & n_5381;
assign n_5537 = n_5382 ^ n_5258;
assign n_5538 = n_4683 & n_5384;
assign n_5539 = n_5385 ^ n_5168;
assign n_5540 = n_5328 & ~n_5386;
assign n_5541 = n_5388 ^ n_5048;
assign n_5542 = n_5389 ^ n_5061;
assign n_5543 = ~n_5389 & n_5239;
assign n_5544 = n_4556 & ~n_5391;
assign n_5545 = n_5393 ^ n_4841;
assign n_5546 = ~n_5393 & n_5211;
assign n_5547 = n_5394 ^ n_4844;
assign n_5548 = ~n_5394 & n_5232;
assign n_5549 = ~n_4654 & ~n_5396;
assign n_5550 = ~n_5234 & n_5398;
assign n_5551 = n_5399 ^ n_5174;
assign n_5552 = n_5335 & n_5400;
assign n_5553 = n_4878 ^ n_5401;
assign n_5554 = ~n_5090 & n_5402;
assign n_5555 = n_5403 ^ n_5044;
assign n_5556 = n_5224 & n_5404;
assign n_5557 = n_5405 ^ n_5286;
assign n_5558 = n_5406 ^ n_5301;
assign n_5559 = ~n_5257 & n_5408;
assign n_5560 = n_5410 & n_5411;
assign n_5561 = n_5413 ^ n_5070;
assign n_5562 = n_5413 & n_5414;
assign n_5563 = n_5415 ^ n_5042;
assign n_5564 = n_5222 & n_5416;
assign n_5565 = n_5417 ^ n_5092;
assign n_5566 = n_5282 & n_5418;
assign n_5567 = n_5419 ^ n_4927;
assign n_5568 = ~n_5419 & ~n_5237;
assign n_5569 = n_5420 ^ n_5302;
assign n_5570 = n_5421 ^ n_5253;
assign n_5571 = n_5407 & ~n_5422;
assign n_5572 = n_5424 ^ n_4709;
assign n_5573 = n_5425 ^ n_5031;
assign n_5574 = n_5425 & ~n_5321;
assign n_5575 = n_5426 & ~n_5427;
assign n_5576 = n_5428 ^ n_5080;
assign n_5577 = ~n_5428 & ~n_5254;
assign n_5578 = n_5429 ^ n_4874;
assign n_5579 = ~n_5429 & ~n_5276;
assign n_5580 = n_5430 ^ n_5089;
assign n_5581 = n_5278 & ~n_5431;
assign n_5582 = n_5432 ^ n_5072;
assign n_5583 = n_5432 & n_5280;
assign n_5584 = n_5057 ^ n_5433;
assign n_5585 = ~n_4637 & n_5434;
assign n_5586 = n_5435 ^ n_4994;
assign n_5587 = ~n_5435 & ~n_5392;
assign n_5588 = n_5436 ^ n_4910;
assign n_5589 = ~n_5436 & ~n_5437;
assign n_5590 = ~n_5438 & ~n_5439;
assign n_5591 = n_5441 ^ n_4913;
assign n_5592 = n_4834 & n_5443;
assign n_5593 = n_5445 ^ n_5122;
assign n_5594 = n_5446 ^ n_5075;
assign n_5595 = n_5446 & ~n_5447;
assign n_5596 = n_5448 ^ n_4919;
assign n_5597 = n_5449 ^ n_5127;
assign n_5598 = ~n_5449 & n_5450;
assign n_5599 = n_5451 ^ n_5130;
assign n_5600 = n_5297 & n_5452;
assign n_5601 = n_5453 ^ n_5299;
assign n_5602 = n_5453 ^ n_5132;
assign n_5603 = ~n_5045 & n_5454;
assign n_5604 = ~n_5456 & n_5457;
assign n_5605 = ~n_5420 & n_5458;
assign n_5606 = n_5460 ^ n_4315;
assign n_5607 = n_5308 ^ n_5462;
assign n_5608 = n_5463 ^ n_5462;
assign n_5609 = n_5310 & ~n_5464;
assign n_5610 = n_5149 & ~n_5467;
assign n_5611 = n_4888 & ~n_5469;
assign y5 = n_5472;
assign n_5612 = ~n_4698 & n_5473;
assign n_5613 = n_5474 ^ n_5331;
assign n_5614 = n_4738 ^ n_5475;
assign n_5615 = n_5476 ^ n_4817;
assign n_5616 = n_5477 ^ n_5323;
assign n_5617 = n_5478 ^ n_4117;
assign n_5618 = n_5479 ^ n_4095;
assign n_5619 = n_5482 ^ n_4948;
assign n_5620 = n_5474 & n_5483;
assign n_5621 = n_5484 ^ n_4106;
assign n_5622 = n_5485 ^ n_4964;
assign n_5623 = n_5487 ^ n_4123;
assign n_5624 = n_5489 ^ n_4704;
assign n_5625 = n_4750 ^ n_5490;
assign n_5626 = n_5491 ^ n_4987;
assign n_5627 = n_4990 ^ n_5492;
assign n_5628 = n_5493 ^ n_4973;
assign n_5629 = n_5495 & ~n_5496;
assign n_5630 = n_5497 ^ n_5494;
assign n_5631 = n_5498 ^ n_4079;
assign n_5632 = n_5500 ^ n_4953;
assign n_5633 = n_5501 ^ n_5189;
assign n_5634 = n_5501 ^ n_4996;
assign n_5635 = n_5502 ^ n_4156;
assign n_5636 = n_5503 ^ n_5198;
assign n_5637 = n_5503 ^ n_4774;
assign n_5638 = n_5504 ^ n_4761;
assign n_5639 = n_5506 ^ n_4081;
assign n_5640 = n_5361 ^ n_5507;
assign n_5641 = n_5508 ^ n_5001;
assign n_5642 = n_5510 ^ n_4785;
assign n_5643 = n_5512 ^ n_4776;
assign n_5644 = n_5514 ^ n_5065;
assign n_5645 = n_5516 ^ n_4982;
assign n_5646 = n_5517 ^ n_4159;
assign n_5647 = n_5519 ^ n_4706;
assign n_5648 = n_5521 ^ n_5033;
assign n_5649 = n_5524 ^ n_4318;
assign n_5650 = n_5526 ^ n_4754;
assign n_5651 = n_5528 ^ n_4893;
assign n_5652 = n_5530 ^ n_5012;
assign n_5653 = n_5522 ^ n_5531;
assign n_5654 = n_5532 ^ n_5024;
assign n_5655 = n_5533 ^ n_5272;
assign n_5656 = n_5533 ^ n_5103;
assign n_5657 = n_5256 & n_5535;
assign n_5658 = n_5536 ^ n_4300;
assign n_5659 = n_5085 ^ n_5537;
assign n_5660 = n_5538 ^ n_4404;
assign n_5661 = n_5539 ^ n_5387;
assign n_5662 = n_5540 ^ n_4266;
assign n_5663 = n_4821 ^ n_5541;
assign n_5664 = n_5542 ^ n_5523;
assign n_5665 = n_5543 ^ n_5061;
assign n_5666 = n_5544 ^ n_4268;
assign n_5667 = n_5545 ^ n_5525;
assign n_5668 = n_5546 ^ n_4841;
assign n_5669 = n_5547 ^ n_5499;
assign n_5670 = n_5548 ^ n_4844;
assign n_5671 = n_5549 ^ n_4345;
assign n_5672 = n_5550 ^ n_5039;
assign n_5673 = n_5552 ^ n_4380;
assign n_5674 = n_5554 ^ n_4388;
assign n_5675 = n_5556 ^ n_4908;
assign n_5676 = n_5557 ^ n_5440;
assign n_5677 = n_5558 ^ n_5136;
assign n_5678 = n_5559 ^ n_5083;
assign n_5679 = n_5560 ^ n_5032;
assign n_5680 = n_5561 ^ n_5412;
assign n_5681 = n_5562 ^ n_5070;
assign n_5682 = n_4810 ^ n_5563;
assign n_5683 = n_5564 ^ n_4527;
assign n_5684 = n_5566 ^ n_5114;
assign n_5685 = n_5568 ^ n_4927;
assign n_5686 = n_5569 ^ n_5138;
assign n_5687 = n_5570 ^ n_5423;
assign n_5688 = n_5571 ^ n_4623;
assign n_5689 = n_5572 ^ n_5243;
assign n_5690 = n_5572 ^ n_5066;
assign n_5691 = n_5573 ^ n_5527;
assign n_5692 = n_5574 ^ n_5031;
assign n_5693 = n_5575 ^ n_4733;
assign n_5694 = n_5551 ^ n_5576;
assign n_5695 = n_5577 ^ n_5080;
assign n_5696 = n_5579 ^ n_4874;
assign n_5697 = n_5581 ^ n_5110;
assign n_5698 = n_5583 ^ n_5072;
assign n_5699 = n_5585 ^ n_4278;
assign n_5700 = n_5587 ^ n_4994;
assign n_5701 = n_5589 ^ n_4910;
assign n_5702 = n_5590 ^ n_4307;
assign n_5703 = n_5442 ^ n_5591;
assign n_5704 = n_5592 ^ n_4309;
assign n_5705 = n_5124 ^ n_5593;
assign n_5706 = n_5595 ^ n_5075;
assign n_5707 = n_5598 ^ n_5127;
assign n_5708 = n_5600 ^ n_4643;
assign n_5709 = ~n_5299 & ~n_5602;
assign n_5710 = n_5603 ^ n_4259;
assign n_5711 = n_5604 ^ n_4885;
assign n_5712 = n_5605 ^ n_4341;
assign n_5713 = n_5606 ^ n_5461;
assign n_5714 = n_5606 ^ n_5306;
assign n_5715 = n_5463 & n_5607;
assign n_5716 = n_5609 ^ n_4650;
assign n_5717 = n_5610 ^ n_4372;
assign n_5718 = n_5611 ^ n_4417;
assign n_5719 = n_5612 ^ n_5315;
assign n_5720 = n_5539 ^ n_5615;
assign n_5721 = n_5617 ^ n_5329;
assign n_5722 = n_5618 ^ n_5481;
assign n_5723 = n_5619 ^ n_5613;
assign n_5724 = n_5620 ^ n_4963;
assign n_5725 = n_5621 ^ n_5486;
assign n_5726 = n_5621 ^ n_5336;
assign n_5727 = n_5622 ^ n_4750;
assign n_5728 = n_5622 ^ n_5490;
assign n_5729 = n_5623 ^ n_4971;
assign n_5730 = n_5623 ^ n_5338;
assign n_5731 = n_5624 ^ n_4738;
assign n_5732 = n_5624 ^ n_5475;
assign n_5733 = n_5626 ^ n_4990;
assign n_5734 = n_5626 ^ n_5492;
assign n_5735 = n_5628 ^ n_5497;
assign n_5736 = n_5628 ^ n_5494;
assign n_5737 = n_5629 ^ n_4980;
assign n_5738 = n_5632 ^ n_5395;
assign n_5739 = n_5631 ^ n_5633;
assign n_5740 = n_5189 & ~n_5634;
assign n_5741 = n_5636 ^ n_5635;
assign n_5742 = n_5198 & ~n_5637;
assign n_5743 = n_5638 ^ n_5505;
assign n_5744 = n_5638 ^ n_5352;
assign n_5745 = n_5639 ^ n_5361;
assign n_5746 = n_5639 ^ n_5507;
assign n_5747 = n_5642 ^ n_5520;
assign n_5748 = n_5644 ^ n_5570;
assign n_5749 = n_5646 ^ n_5518;
assign n_5750 = n_5646 ^ n_5641;
assign n_5751 = n_5647 ^ n_5642;
assign n_5752 = n_5648 ^ n_5529;
assign n_5753 = n_5648 ^ n_5643;
assign n_5754 = n_5650 ^ n_5390;
assign n_5755 = n_5651 ^ n_5397;
assign n_5756 = n_5652 ^ n_5522;
assign n_5757 = n_5652 ^ n_5531;
assign n_5758 = n_5654 ^ n_5480;
assign n_5759 = n_5654 ^ n_5327;
assign n_5760 = n_5272 & ~n_5656;
assign n_5761 = n_5657 ^ n_4898;
assign n_5762 = n_5658 ^ n_5274;
assign n_5763 = n_5658 ^ n_5105;
assign n_5764 = n_5660 ^ n_5567;
assign n_5765 = n_5661 ^ n_5615;
assign n_5766 = n_5662 ^ n_4821;
assign n_5767 = n_5662 ^ n_5541;
assign n_5768 = n_5665 ^ n_4824;
assign n_5769 = n_5665 ^ n_5649;
assign n_5770 = n_5666 ^ n_5266;
assign n_5771 = n_5666 ^ n_5098;
assign n_5772 = n_5650 ^ n_5668;
assign n_5773 = n_5632 ^ n_5670;
assign n_5774 = n_5671 ^ n_5212;
assign n_5775 = n_5671 ^ n_5029;
assign n_5776 = n_5672 ^ n_5551;
assign n_5777 = n_5672 ^ n_5576;
assign n_5778 = n_5673 ^ n_5409;
assign n_5779 = n_5674 ^ n_5057;
assign n_5780 = n_5674 ^ n_5433;
assign n_5781 = n_5675 ^ n_5557;
assign n_5782 = n_5678 ^ n_5085;
assign n_5783 = n_5678 ^ n_5537;
assign n_5784 = n_5561 ^ n_5679;
assign n_5785 = n_5680 ^ n_5679;
assign n_5786 = n_5681 ^ n_4810;
assign n_5787 = n_5681 ^ n_5563;
assign n_5788 = n_5683 ^ n_4878;
assign n_5789 = n_5683 ^ n_5401;
assign n_5790 = n_5684 ^ n_5586;
assign n_5791 = n_5685 ^ n_5677;
assign n_5792 = n_5685 ^ n_5558;
assign n_5793 = n_5688 ^ n_5573;
assign n_5794 = ~n_5243 & ~n_5690;
assign n_5795 = n_5692 ^ n_5651;
assign n_5796 = n_5693 ^ n_5246;
assign n_5797 = n_5693 ^ n_5069;
assign n_5798 = n_5695 ^ n_5673;
assign n_5799 = n_5696 ^ n_5580;
assign n_5800 = n_5697 ^ n_5582;
assign n_5801 = n_5698 ^ n_5565;
assign n_5802 = n_5699 ^ n_5284;
assign n_5803 = n_5699 ^ n_4856;
assign n_5804 = n_5700 ^ n_5555;
assign n_5805 = n_5702 ^ n_5442;
assign n_5806 = n_5702 ^ n_5591;
assign n_5807 = n_5704 ^ n_5124;
assign n_5808 = n_5704 ^ n_5593;
assign n_5809 = n_5706 ^ n_5596;
assign n_5810 = n_5706 ^ n_5448;
assign n_5811 = n_5707 ^ n_5296;
assign n_5812 = n_5707 ^ n_5129;
assign n_5813 = n_5708 ^ n_5601;
assign n_5814 = n_5709 ^ n_5133;
assign n_5815 = n_5710 ^ n_5455;
assign n_5816 = n_5710 ^ n_5300;
assign n_5817 = n_5711 ^ n_5686;
assign n_5818 = n_5711 ^ n_5569;
assign n_5819 = n_5712 ^ n_5459;
assign n_5820 = n_5712 ^ n_5303;
assign n_5821 = n_5461 & n_5714;
assign n_5822 = n_5715 ^ n_5145;
assign n_5823 = n_5716 ^ n_5466;
assign n_5824 = n_5717 ^ n_5468;
assign n_5825 = n_5718 ^ n_4941;
assign n_5826 = n_5719 ^ n_4699;
assign n_5827 = n_5719 ^ n_4091;
assign n_5828 = ~n_5661 & n_5720;
assign n_5829 = n_5725 ^ n_5724;
assign n_5830 = n_5486 & ~n_5726;
assign n_5831 = n_5727 ^ n_5490;
assign n_5832 = ~n_5625 & n_5728;
assign n_5833 = n_5729 ^ n_5338;
assign n_5834 = n_5488 & ~n_5730;
assign n_5835 = n_5731 ^ n_5475;
assign n_5836 = ~n_5614 & n_5732;
assign n_5837 = n_5733 ^ n_5492;
assign n_5838 = ~n_5627 & ~n_5734;
assign n_5839 = n_5735 ^ n_5494;
assign n_5840 = n_5630 & ~n_5736;
assign n_5841 = n_5737 ^ n_5631;
assign n_5842 = n_5738 ^ n_5670;
assign n_5843 = n_5740 ^ n_4760;
assign n_5844 = n_5742 ^ n_5008;
assign n_5845 = n_5743 ^ n_5515;
assign n_5846 = n_5505 & ~n_5744;
assign n_5847 = n_5745 ^ n_5507;
assign n_5848 = n_5640 & ~n_5746;
assign n_5849 = n_5748 ^ n_5423;
assign n_5850 = ~n_5748 & n_5687;
assign n_5851 = n_5749 ^ n_5641;
assign n_5852 = n_5749 & n_5750;
assign n_5853 = n_5751 ^ n_5520;
assign n_5854 = ~n_5751 & n_5747;
assign n_5855 = n_5752 ^ n_5643;
assign n_5856 = ~n_5752 & ~n_5753;
assign n_5857 = n_5754 ^ n_5668;
assign n_5858 = n_5756 ^ n_5531;
assign n_5859 = ~n_5653 & ~n_5757;
assign n_5860 = n_5480 & n_5759;
assign n_5861 = n_5760 ^ n_4850;
assign n_5862 = n_5762 ^ n_5761;
assign n_5863 = ~n_5274 & n_5763;
assign n_5864 = n_5758 ^ n_5765;
assign n_5865 = n_5766 ^ n_5541;
assign n_5866 = ~n_5663 & n_5767;
assign n_5867 = n_5768 ^ n_5649;
assign n_5868 = n_5768 & n_5769;
assign n_5869 = n_5770 ^ n_5513;
assign n_5870 = n_5266 & ~n_5771;
assign n_5871 = ~n_5754 & n_5772;
assign n_5872 = ~n_5738 & ~n_5773;
assign n_5873 = n_5212 & ~n_5775;
assign n_5874 = n_5776 ^ n_5576;
assign n_5875 = n_5694 & ~n_5777;
assign n_5876 = n_5779 ^ n_5433;
assign n_5877 = n_5584 & n_5780;
assign n_5878 = n_5781 ^ n_5440;
assign n_5879 = n_5781 & ~n_5676;
assign n_5880 = n_5782 ^ n_5537;
assign n_5881 = ~n_5659 & n_5783;
assign n_5882 = ~n_5680 & ~n_5784;
assign n_5883 = n_5578 ^ n_5785;
assign n_5884 = n_5786 ^ n_5563;
assign n_5885 = ~n_5682 & n_5787;
assign n_5886 = n_5788 ^ n_5401;
assign n_5887 = ~n_5553 & n_5789;
assign n_5888 = ~n_5677 & n_5792;
assign n_5889 = n_5793 ^ n_5527;
assign n_5890 = n_5793 & n_5691;
assign n_5891 = n_5794 ^ n_4804;
assign n_5892 = n_5795 ^ n_5397;
assign n_5893 = n_5795 & n_5755;
assign n_5894 = n_5246 & ~n_5797;
assign n_5895 = n_5798 ^ n_5409;
assign n_5896 = n_5798 & n_5778;
assign n_5897 = n_5284 & ~n_5803;
assign n_5898 = n_5805 ^ n_5591;
assign n_5899 = ~n_5703 & ~n_5806;
assign n_5900 = n_5807 ^ n_5593;
assign n_5901 = n_5705 & ~n_5808;
assign n_5902 = n_5809 ^ n_5597;
assign n_5903 = n_5596 & n_5810;
assign n_5904 = n_5811 ^ n_5599;
assign n_5905 = n_5296 & n_5812;
assign n_5906 = n_5383 ^ n_5814;
assign n_5907 = n_5815 ^ n_5383;
assign n_5908 = n_5815 ^ n_5814;
assign n_5909 = n_5455 & n_5816;
assign n_5910 = n_5686 & n_5818;
assign n_5911 = ~n_5459 & n_5820;
assign n_5912 = n_5821 ^ n_5142;
assign n_5913 = n_5822 ^ n_5465;
assign y6 = ~n_5826;
assign n_5914 = n_4699 & n_5827;
assign n_5915 = n_5828 ^ n_5387;
assign n_5916 = n_5830 ^ n_4977;
assign n_5917 = n_5832 ^ n_4750;
assign n_5918 = n_5834 ^ n_4971;
assign n_5919 = n_5836 ^ n_4738;
assign n_5920 = n_5838 ^ n_4990;
assign n_5921 = n_5840 ^ n_5497;
assign n_5922 = n_5841 ^ n_5633;
assign n_5923 = ~n_5841 & n_5739;
assign n_5924 = n_5770 ^ n_5842;
assign n_5925 = n_5843 ^ n_5741;
assign n_5926 = n_5843 ^ n_5636;
assign n_5927 = n_5843 ^ n_5635;
assign n_5928 = n_5743 ^ n_5844;
assign n_5929 = n_5845 ^ n_5844;
assign n_5930 = n_5846 ^ n_4999;
assign n_5931 = n_5645 ^ n_5847;
assign n_5932 = n_5848 ^ n_5361;
assign n_5933 = n_5850 ^ n_5423;
assign n_5934 = n_5851 ^ n_5509;
assign n_5935 = n_5852 ^ n_5518;
assign n_5936 = n_5511 ^ n_5853;
assign n_5937 = n_5854 ^ n_5520;
assign n_5938 = n_5368 ^ n_5855;
assign n_5939 = n_5856 ^ n_5529;
assign n_5940 = n_5378 ^ n_5858;
assign n_5941 = n_5859 ^ n_5522;
assign n_5942 = n_5860 ^ n_4838;
assign n_5943 = n_5861 ^ n_5796;
assign n_5944 = n_5863 ^ n_5106;
assign n_5945 = n_5865 ^ n_5664;
assign n_5946 = n_5865 ^ n_5523;
assign n_5947 = n_5866 ^ n_4821;
assign n_5948 = n_5868 ^ n_4824;
assign n_5949 = n_5869 ^ n_5842;
assign n_5950 = n_5870 ^ n_4793;
assign n_5951 = n_5871 ^ n_5390;
assign n_5952 = n_5872 ^ n_5395;
assign n_5953 = n_5873 ^ n_4771;
assign n_5954 = n_5875 ^ n_5551;
assign n_5955 = n_5877 ^ n_5057;
assign n_5956 = n_5878 ^ n_5701;
assign n_5957 = n_5879 ^ n_5440;
assign n_5958 = n_5880 ^ n_5862;
assign n_5959 = n_5880 ^ n_5762;
assign n_5960 = n_5880 ^ n_5761;
assign n_5961 = n_5881 ^ n_5085;
assign n_5962 = n_5882 ^ n_5412;
assign n_5963 = n_5885 ^ n_4810;
assign n_5964 = n_5887 ^ n_4878;
assign n_5965 = n_5888 ^ n_5136;
assign n_5966 = n_5890 ^ n_5527;
assign n_5967 = n_5891 ^ n_5655;
assign n_5968 = n_5893 ^ n_5397;
assign n_5969 = n_5894 ^ n_4867;
assign n_5970 = n_5896 ^ n_5409;
assign n_5971 = n_5897 ^ n_5116;
assign n_5972 = n_5898 ^ n_5444;
assign n_5973 = n_5899 ^ n_5442;
assign n_5974 = n_5900 ^ n_5594;
assign n_5975 = n_5901 ^ n_5124;
assign n_5976 = n_5903 ^ n_4919;
assign n_5977 = n_5905 ^ n_4860;
assign n_5978 = n_5907 ^ n_5814;
assign n_5979 = ~n_5906 & ~n_5908;
assign n_5980 = n_5909 ^ n_5095;
assign n_5981 = n_5910 ^ n_5138;
assign n_5982 = n_5911 ^ n_5304;
assign n_5983 = n_5912 ^ n_5608;
assign n_5984 = n_5914 ^ n_5719;
assign n_5985 = n_5916 ^ n_5833;
assign n_5986 = n_5917 ^ n_5837;
assign n_5987 = n_5918 ^ n_5835;
assign n_5988 = n_5919 ^ n_5831;
assign n_5989 = n_5920 ^ n_5839;
assign n_5990 = n_5922 ^ n_5921;
assign n_5991 = n_5923 ^ n_5633;
assign n_5992 = ~n_5869 & n_5924;
assign n_5993 = n_5926 & n_5927;
assign n_5994 = ~n_5845 & ~n_5928;
assign n_5995 = n_5930 ^ n_5645;
assign n_5996 = n_5851 ^ n_5932;
assign n_5997 = n_5689 ^ n_5933;
assign n_5998 = n_5934 ^ n_5932;
assign n_5999 = n_5935 ^ n_5511;
assign n_6000 = n_5935 ^ n_5853;
assign n_6001 = n_5937 ^ n_5368;
assign n_6002 = n_5937 ^ n_5855;
assign n_6003 = n_5939 ^ n_5378;
assign n_6004 = n_5939 ^ n_5858;
assign n_6005 = n_5941 ^ n_5758;
assign n_6006 = n_5942 ^ n_5915;
assign n_6007 = n_5944 ^ n_5578;
assign n_6008 = n_5944 ^ n_5785;
assign n_6009 = n_5915 ^ n_5945;
assign n_6010 = ~n_5664 & ~n_5946;
assign n_6011 = n_5947 ^ n_5667;
assign n_6012 = n_5947 ^ n_5525;
assign n_6013 = n_5948 ^ n_5669;
assign n_6014 = n_5948 ^ n_5547;
assign n_6015 = n_5950 ^ n_5774;
assign n_6016 = n_5951 ^ n_5949;
assign n_6017 = n_5950 ^ n_5952;
assign n_6018 = n_5953 ^ n_5689;
assign n_6019 = n_5953 ^ n_5933;
assign n_6020 = n_5955 ^ n_5790;
assign n_6021 = n_5955 ^ n_5684;
assign n_6022 = n_5898 ^ n_5957;
assign n_6023 = n_5959 & n_5960;
assign n_6024 = n_5962 ^ n_5799;
assign n_6025 = n_5962 ^ n_5696;
assign n_6026 = n_5963 ^ n_5800;
assign n_6027 = n_5963 ^ n_5697;
assign n_6028 = n_5964 ^ n_5801;
assign n_6029 = n_5964 ^ n_5698;
assign n_6030 = n_5965 ^ n_5817;
assign n_6031 = n_5891 ^ n_5966;
assign n_6032 = n_5967 ^ n_5966;
assign n_6033 = n_5968 ^ n_5943;
assign n_6034 = n_5968 ^ n_5861;
assign n_6035 = n_5969 ^ n_5534;
assign n_6036 = n_5969 ^ n_5954;
assign n_6037 = n_5970 ^ n_5958;
assign n_6038 = n_5971 ^ n_5804;
assign n_6039 = n_5971 ^ n_5700;
assign n_6040 = n_5972 ^ n_5957;
assign n_6041 = n_5900 ^ n_5973;
assign n_6042 = n_5974 ^ n_5973;
assign n_6043 = n_5975 ^ n_5902;
assign n_6044 = n_5975 ^ n_5809;
assign n_6045 = n_5976 ^ n_5904;
assign n_6046 = n_5976 ^ n_5811;
assign n_6047 = n_5977 ^ n_5813;
assign n_6048 = n_5977 ^ n_5708;
assign n_6049 = n_5979 ^ n_5383;
assign n_6050 = n_5980 ^ n_5764;
assign n_6051 = n_5980 ^ n_5660;
assign n_6052 = n_5981 ^ n_5819;
assign n_6053 = n_5982 ^ n_5713;
assign n_6054 = n_5984 ^ n_5154;
assign n_6055 = n_5984 ^ n_4946;
assign n_6056 = n_5991 ^ n_5925;
assign n_6057 = n_5992 ^ n_5513;
assign n_6058 = n_5993 ^ n_5636;
assign n_6059 = n_5994 ^ n_5515;
assign n_6060 = n_5995 ^ n_5847;
assign n_6061 = ~n_5995 & ~n_5931;
assign n_6062 = n_5934 & ~n_5996;
assign n_6063 = n_5999 ^ n_5853;
assign n_6064 = n_5936 & ~n_6000;
assign n_6065 = n_6001 ^ n_5855;
assign n_6066 = n_5938 & ~n_6002;
assign n_6067 = n_6003 ^ n_5858;
assign n_6068 = ~n_5940 & n_6004;
assign n_6069 = n_6005 ^ n_5765;
assign n_6070 = ~n_6005 & ~n_5864;
assign n_6071 = n_6006 ^ n_5945;
assign n_6072 = n_6007 ^ n_5785;
assign n_6073 = n_5883 & n_6008;
assign n_6074 = n_6006 & ~n_6009;
assign n_6075 = n_6010 ^ n_5542;
assign n_6076 = n_6011 ^ n_5867;
assign n_6077 = ~n_5667 & n_6012;
assign n_6078 = n_6013 ^ n_5857;
assign n_6079 = n_5669 & ~n_6014;
assign n_6080 = n_6015 ^ n_5952;
assign n_6081 = ~n_6015 & n_6017;
assign n_6082 = n_6018 ^ n_5933;
assign n_6083 = ~n_5997 & n_6019;
assign n_6084 = n_6020 ^ n_5802;
assign n_6085 = n_5790 & n_6021;
assign n_6086 = n_5972 & ~n_6022;
assign n_6087 = n_6023 ^ n_5762;
assign n_6088 = n_6024 ^ n_5884;
assign n_6089 = n_5799 & ~n_6025;
assign n_6090 = n_6026 ^ n_5886;
assign n_6091 = n_5800 & ~n_6027;
assign n_6092 = n_6028 ^ n_5876;
assign n_6093 = n_5801 & n_6029;
assign n_6094 = ~n_5967 & ~n_6031;
assign n_6095 = n_6032 ^ n_5892;
assign n_6096 = n_6033 ^ n_5874;
assign n_6097 = n_5943 & n_6034;
assign n_6098 = n_6035 ^ n_5954;
assign n_6099 = ~n_6035 & ~n_6036;
assign n_6100 = n_6038 ^ n_5588;
assign n_6101 = ~n_5804 & ~n_6039;
assign n_6102 = ~n_5974 & n_6041;
assign n_6103 = ~n_5902 & ~n_6044;
assign n_6104 = n_5904 & ~n_6046;
assign n_6105 = ~n_5813 & ~n_6048;
assign n_6106 = n_6050 ^ n_6049;
assign n_6107 = ~n_5764 & n_6051;
assign y7 = n_6054;
assign n_6108 = ~n_5154 & ~n_6055;
assign n_6109 = n_6058 ^ n_5929;
assign n_6110 = n_6060 ^ n_6059;
assign n_6111 = n_6061 ^ n_5847;
assign n_6112 = n_6062 ^ n_5509;
assign n_6113 = n_6064 ^ n_5511;
assign n_6114 = n_6066 ^ n_5368;
assign n_6115 = n_6068 ^ n_5378;
assign n_6116 = n_6070 ^ n_5765;
assign n_6117 = n_6072 ^ n_5961;
assign n_6118 = n_6073 ^ n_5578;
assign n_6119 = n_6074 ^ n_5945;
assign n_6120 = n_5867 ^ n_6075;
assign n_6121 = n_6011 ^ n_6075;
assign n_6122 = n_6076 ^ n_6075;
assign n_6123 = n_6077 ^ n_5545;
assign n_6124 = n_6079 ^ n_5499;
assign n_6125 = n_6080 ^ n_5849;
assign n_6126 = n_6080 ^ n_6057;
assign n_6127 = n_6081 ^ n_5774;
assign n_6128 = n_6082 ^ n_5889;
assign n_6129 = n_6083 ^ n_5689;
assign n_6130 = n_6085 ^ n_5586;
assign n_6131 = n_6086 ^ n_5444;
assign n_6132 = n_5961 ^ n_6087;
assign n_6133 = n_6072 ^ n_6087;
assign n_6134 = n_6089 ^ n_5580;
assign n_6135 = n_6091 ^ n_5582;
assign n_6136 = n_6093 ^ n_5565;
assign n_6137 = n_6094 ^ n_5655;
assign n_6138 = n_6097 ^ n_5796;
assign n_6139 = n_6098 ^ n_5895;
assign n_6140 = n_6099 ^ n_5534;
assign n_6141 = n_6101 ^ n_5555;
assign n_6142 = n_6102 ^ n_5594;
assign n_6143 = n_6103 ^ n_5597;
assign n_6144 = n_6104 ^ n_5599;
assign n_6145 = n_6105 ^ n_5601;
assign n_6146 = n_6107 ^ n_5567;
assign n_6147 = n_6108 ^ n_5984;
assign n_6148 = n_6111 ^ n_5998;
assign n_6149 = n_6112 ^ n_6063;
assign n_6150 = n_6113 ^ n_6065;
assign n_6151 = n_6114 ^ n_6067;
assign n_6152 = n_6115 ^ n_6069;
assign n_6153 = n_6116 ^ n_6071;
assign n_6154 = n_6117 ^ n_6087;
assign n_6155 = n_6118 ^ n_6088;
assign n_6156 = n_6118 ^ n_6024;
assign n_6157 = ~n_6120 & n_6121;
assign n_6158 = n_6122 ^ n_6119;
assign n_6159 = n_6123 ^ n_6078;
assign n_6160 = n_6123 ^ n_6013;
assign n_6161 = n_6124 ^ n_5951;
assign n_6162 = n_6125 ^ n_6057;
assign n_6163 = n_6125 & n_6126;
assign n_6164 = n_6127 ^ n_6082;
assign n_6165 = n_6127 ^ n_6128;
assign n_6166 = n_6129 ^ n_6095;
assign n_6167 = n_6129 ^ n_6032;
assign n_6168 = n_6130 ^ n_6100;
assign n_6169 = n_6130 ^ n_6038;
assign n_6170 = n_6131 ^ n_6042;
assign n_6171 = ~n_6132 & n_6133;
assign n_6172 = n_6134 ^ n_6090;
assign n_6173 = n_6134 ^ n_6026;
assign n_6174 = n_6135 ^ n_6092;
assign n_6175 = n_6135 ^ n_6028;
assign n_6176 = n_6136 ^ n_6084;
assign n_6177 = n_6136 ^ n_6020;
assign n_6178 = n_6137 ^ n_6096;
assign n_6179 = n_6137 ^ n_6033;
assign n_6180 = n_6098 ^ n_6138;
assign n_6181 = n_6139 ^ n_6138;
assign n_6182 = n_6140 ^ n_6037;
assign n_6183 = n_6140 ^ n_5970;
assign n_6184 = n_6141 ^ n_5956;
assign n_6185 = n_6141 ^ n_5701;
assign n_6186 = n_6142 ^ n_6043;
assign n_6187 = n_6143 ^ n_6045;
assign n_6188 = n_6144 ^ n_6047;
assign n_6189 = n_6145 ^ n_5978;
assign n_6190 = n_6146 ^ n_5791;
assign n_6191 = n_6147 ^ n_5316;
assign n_6192 = n_6147 ^ n_4955;
assign n_6193 = ~n_6088 & ~n_6156;
assign n_6194 = n_6157 ^ n_5867;
assign n_6195 = ~n_6078 & ~n_6160;
assign n_6196 = n_6161 ^ n_5949;
assign n_6197 = ~n_6161 & n_6016;
assign n_6198 = n_6163 ^ n_5849;
assign n_6199 = n_6128 & n_6164;
assign n_6200 = n_6095 & n_6167;
assign n_6201 = n_6100 & n_6169;
assign n_6202 = n_6171 ^ n_5961;
assign n_6203 = ~n_6090 & ~n_6173;
assign n_6204 = n_6092 & ~n_6175;
assign n_6205 = ~n_6084 & ~n_6177;
assign n_6206 = ~n_6096 & n_6179;
assign n_6207 = ~n_6139 & n_6180;
assign n_6208 = ~n_6037 & ~n_6183;
assign n_6209 = n_5956 & ~n_6185;
assign y8 = n_6191;
assign n_6210 = ~n_5316 & n_6192;
assign n_6211 = n_6193 ^ n_5884;
assign n_6212 = n_6194 ^ n_6159;
assign n_6213 = n_6195 ^ n_5857;
assign n_6214 = n_6197 ^ n_5949;
assign n_6215 = n_6198 ^ n_6165;
assign n_6216 = n_6199 ^ n_5889;
assign n_6217 = n_6200 ^ n_5892;
assign n_6218 = n_6201 ^ n_5588;
assign n_6219 = n_6202 ^ n_6155;
assign n_6220 = n_6203 ^ n_5886;
assign n_6221 = n_6204 ^ n_5876;
assign n_6222 = n_6205 ^ n_5802;
assign n_6223 = n_6206 ^ n_5874;
assign n_6224 = n_6207 ^ n_5895;
assign n_6225 = n_6208 ^ n_5958;
assign n_6226 = n_6209 ^ n_5878;
assign n_6227 = n_6210 ^ n_6147;
assign n_6228 = n_6211 ^ n_6172;
assign n_6229 = n_6213 ^ n_6196;
assign n_6230 = n_6214 ^ n_6162;
assign n_6231 = n_6216 ^ n_6166;
assign n_6232 = n_6217 ^ n_6178;
assign n_6233 = n_6218 ^ n_6184;
assign n_6234 = n_6220 ^ n_6174;
assign n_6235 = n_6221 ^ n_6176;
assign n_6236 = n_6222 ^ n_6168;
assign n_6237 = n_6223 ^ n_6181;
assign n_6238 = n_6224 ^ n_6182;
assign n_6239 = n_6225 ^ n_6154;
assign n_6240 = n_6226 ^ n_6040;
assign n_6241 = n_6227 ^ n_5322;
assign n_6242 = n_6227 ^ n_4957;
assign y9 = n_6241;
assign n_6243 = ~n_5322 & ~n_6242;
assign n_6244 = n_6243 ^ n_6227;
assign n_6245 = n_6244 ^ n_5616;
assign n_6246 = n_6244 ^ n_5477;
assign y10 = ~n_6245;
assign n_6247 = n_5616 & ~n_6246;
assign n_6248 = n_6247 ^ n_6244;
assign n_6249 = n_6248 ^ n_5721;
assign n_6250 = n_6248 ^ n_5329;
assign y11 = ~n_6249;
assign n_6251 = n_5721 & ~n_6250;
assign n_6252 = n_6251 ^ n_6248;
assign n_6253 = n_6252 ^ n_5722;
assign n_6254 = n_6252 ^ n_5481;
assign y12 = ~n_6253;
assign n_6255 = n_5722 & n_6254;
assign n_6256 = n_6255 ^ n_6252;
assign n_6257 = n_6256 ^ n_5723;
assign n_6258 = n_6256 ^ n_5613;
assign y13 = n_6257;
assign n_6259 = ~n_5723 & ~n_6258;
assign n_6260 = n_6259 ^ n_6256;
assign n_6261 = n_6260 ^ n_5829;
assign n_6262 = n_6260 ^ n_5725;
assign y14 = ~n_6261;
assign n_6263 = n_5829 & ~n_6262;
assign n_6264 = n_6263 ^ n_6260;
assign n_6265 = n_6264 ^ n_5985;
assign n_6266 = n_6264 ^ n_5833;
assign y15 = n_6265;
assign n_6267 = ~n_5985 & ~n_6266;
assign n_6268 = n_6267 ^ n_6264;
assign n_6269 = n_6268 ^ n_5987;
assign n_6270 = n_6268 ^ n_5835;
assign y16 = ~n_6269;
assign n_6271 = n_5987 & n_6270;
assign n_6272 = n_6271 ^ n_6268;
assign n_6273 = n_6272 ^ n_5988;
assign n_6274 = n_6272 ^ n_5831;
assign y17 = n_6273;
assign n_6275 = ~n_5988 & ~n_6274;
assign n_6276 = n_6275 ^ n_6272;
assign n_6277 = n_6276 ^ n_5986;
assign n_6278 = n_6276 ^ n_5837;
assign y18 = n_6277;
assign n_6279 = ~n_5986 & n_6278;
assign n_6280 = n_6279 ^ n_6276;
assign n_6281 = n_6280 ^ n_5989;
assign n_6282 = n_6280 ^ n_5839;
assign y19 = ~n_6281;
assign n_6283 = n_5989 & ~n_6282;
assign n_6284 = n_6283 ^ n_6280;
assign n_6285 = n_6284 ^ n_5990;
assign n_6286 = n_6284 ^ n_5922;
assign y20 = n_6285;
assign n_6287 = ~n_5990 & ~n_6286;
assign n_6288 = n_6287 ^ n_6284;
assign n_6289 = n_6288 ^ n_6056;
assign n_6290 = n_6288 ^ n_5925;
assign y21 = ~n_6289;
assign n_6291 = n_6056 & n_6290;
assign n_6292 = n_6291 ^ n_6288;
assign n_6293 = n_6292 ^ n_6109;
assign n_6294 = n_6292 ^ n_5929;
assign y22 = ~n_6293;
assign n_6295 = n_6109 & n_6294;
assign n_6296 = n_6295 ^ n_6292;
assign n_6297 = n_6296 ^ n_6110;
assign n_6298 = n_6296 ^ n_6060;
assign y23 = n_6297;
assign n_6299 = ~n_6110 & n_6298;
assign n_6300 = n_6299 ^ n_6296;
assign n_6301 = n_6300 ^ n_6148;
assign n_6302 = n_6300 ^ n_5998;
assign y24 = n_6301;
assign n_6303 = ~n_6148 & n_6302;
assign n_6304 = n_6303 ^ n_6300;
assign n_6305 = n_6304 ^ n_6149;
assign n_6306 = n_6304 ^ n_6063;
assign y25 = ~n_6305;
assign n_6307 = n_6149 & ~n_6306;
assign n_6308 = n_6307 ^ n_6304;
assign n_6309 = n_6308 ^ n_6150;
assign n_6310 = n_6308 ^ n_6065;
assign y26 = n_6309;
assign n_6311 = ~n_6150 & ~n_6310;
assign n_6312 = n_6311 ^ n_6308;
assign n_6313 = n_6312 ^ n_6151;
assign n_6314 = n_6312 ^ n_6067;
assign y27 = ~n_6313;
assign n_6315 = n_6151 & n_6314;
assign n_6316 = n_6315 ^ n_6312;
assign n_6317 = n_6316 ^ n_6152;
assign n_6318 = n_6316 ^ n_6069;
assign y28 = n_6317;
assign n_6319 = ~n_6152 & ~n_6318;
assign n_6320 = n_6319 ^ n_6316;
assign n_6321 = n_6320 ^ n_6153;
assign n_6322 = n_6320 ^ n_6071;
assign y29 = ~n_6321;
assign n_6323 = n_6153 & n_6322;
assign n_6324 = n_6323 ^ n_6320;
assign n_6325 = n_6324 ^ n_6158;
assign n_6326 = n_6324 ^ n_6122;
assign y30 = n_6325;
assign n_6327 = ~n_6158 & ~n_6326;
assign n_6328 = n_6327 ^ n_6324;
assign n_6329 = n_6328 ^ n_6212;
assign n_6330 = n_6328 ^ n_6159;
assign y31 = n_6329;
assign n_6331 = ~n_6212 & n_6330;
assign n_6332 = n_6331 ^ n_6328;
assign n_6333 = n_6332 ^ n_6229;
assign n_6334 = n_6332 ^ n_6196;
assign y32 = ~n_6333;
assign n_6335 = n_6229 & ~n_6334;
assign n_6336 = n_6335 ^ n_6332;
assign n_6337 = n_6336 ^ n_6230;
assign n_6338 = n_6336 ^ n_6162;
assign y33 = ~n_6337;
assign n_6339 = n_6230 & n_6338;
assign n_6340 = n_6339 ^ n_6336;
assign n_6341 = n_6340 ^ n_6215;
assign n_6342 = n_6340 ^ n_6165;
assign y34 = ~n_6341;
assign n_6343 = n_6215 & n_6342;
assign n_6344 = n_6343 ^ n_6340;
assign n_6345 = n_6344 ^ n_6231;
assign n_6346 = n_6344 ^ n_6166;
assign y35 = ~n_6345;
assign n_6347 = n_6231 & n_6346;
assign n_6348 = n_6347 ^ n_6344;
assign n_6349 = n_6348 ^ n_6232;
assign n_6350 = n_6348 ^ n_6178;
assign y36 = ~n_6349;
assign n_6351 = n_6232 & n_6350;
assign n_6352 = n_6351 ^ n_6348;
assign n_6353 = n_6352 ^ n_6237;
assign n_6354 = n_6352 ^ n_6181;
assign y37 = ~n_6353;
assign n_6355 = n_6237 & n_6354;
assign n_6356 = n_6355 ^ n_6352;
assign n_6357 = n_6356 ^ n_6238;
assign n_6358 = n_6356 ^ n_6182;
assign y38 = n_6357;
assign n_6359 = ~n_6238 & ~n_6358;
assign n_6360 = n_6359 ^ n_6356;
assign n_6361 = n_6360 ^ n_6239;
assign n_6362 = n_6360 ^ n_6154;
assign y39 = ~n_6361;
assign n_6363 = n_6239 & n_6362;
assign n_6364 = n_6363 ^ n_6360;
assign n_6365 = n_6364 ^ n_6219;
assign n_6366 = n_6364 ^ n_6155;
assign y40 = n_6365;
assign n_6367 = ~n_6219 & ~n_6366;
assign n_6368 = n_6367 ^ n_6364;
assign n_6369 = n_6368 ^ n_6228;
assign n_6370 = n_6368 ^ n_6172;
assign y41 = n_6369;
assign n_6371 = ~n_6228 & ~n_6370;
assign n_6372 = n_6371 ^ n_6368;
assign n_6373 = n_6372 ^ n_6234;
assign n_6374 = n_6372 ^ n_6174;
assign y42 = ~n_6373;
assign n_6375 = n_6234 & n_6374;
assign n_6376 = n_6375 ^ n_6372;
assign n_6377 = n_6376 ^ n_6235;
assign n_6378 = n_6376 ^ n_6176;
assign y43 = n_6377;
assign n_6379 = ~n_6235 & n_6378;
assign n_6380 = n_6379 ^ n_6376;
assign n_6381 = n_6380 ^ n_6236;
assign n_6382 = n_6380 ^ n_6168;
assign y44 = n_6381;
assign n_6383 = ~n_6236 & n_6382;
assign n_6384 = n_6383 ^ n_6380;
assign n_6385 = n_6384 ^ n_6233;
assign n_6386 = n_6384 ^ n_6184;
assign y45 = n_6385;
assign n_6387 = ~n_6233 & ~n_6386;
assign n_6388 = n_6387 ^ n_6384;
assign n_6389 = n_6388 ^ n_6240;
assign n_6390 = n_6388 ^ n_6040;
assign y46 = ~n_6389;
assign n_6391 = n_6240 & n_6390;
assign n_6392 = n_6391 ^ n_6388;
assign n_6393 = n_6392 ^ n_6170;
assign n_6394 = n_6392 ^ n_6042;
assign y47 = ~n_6393;
assign n_6395 = n_6170 & ~n_6394;
assign n_6396 = n_6395 ^ n_6392;
assign n_6397 = n_6396 ^ n_6186;
assign n_6398 = n_6396 ^ n_6043;
assign y48 = n_6397;
assign n_6399 = ~n_6186 & n_6398;
assign n_6400 = n_6399 ^ n_6396;
assign n_6401 = n_6400 ^ n_6187;
assign n_6402 = n_6400 ^ n_6045;
assign y49 = n_6401;
assign n_6403 = ~n_6187 & n_6402;
assign n_6404 = n_6403 ^ n_6400;
assign n_6405 = n_6404 ^ n_6188;
assign n_6406 = n_6404 ^ n_6047;
assign y50 = n_6405;
assign n_6407 = ~n_6188 & n_6406;
assign n_6408 = n_6407 ^ n_6404;
assign n_6409 = n_6408 ^ n_6189;
assign n_6410 = n_6408 ^ n_5978;
assign y51 = ~n_6409;
assign n_6411 = n_6189 & ~n_6410;
assign n_6412 = n_6411 ^ n_6408;
assign n_6413 = n_6412 ^ n_6106;
assign n_6414 = n_6412 ^ n_6050;
assign y52 = ~n_6413;
assign n_6415 = n_6106 & n_6414;
assign n_6416 = n_6415 ^ n_6412;
assign n_6417 = n_6416 ^ n_6190;
assign n_6418 = n_6416 ^ n_5791;
assign y53 = ~n_6417;
assign n_6419 = n_6190 & n_6418;
assign n_6420 = n_6419 ^ n_6416;
assign n_6421 = n_6420 ^ n_6030;
assign n_6422 = n_6420 ^ n_5817;
assign y54 = n_6421;
assign n_6423 = ~n_6030 & ~n_6422;
assign n_6424 = n_6423 ^ n_6420;
assign n_6425 = n_6424 ^ n_6052;
assign n_6426 = n_6424 ^ n_5819;
assign y55 = n_6425;
assign n_6427 = ~n_6052 & n_6426;
assign n_6428 = n_6427 ^ n_6424;
assign n_6429 = n_6428 ^ n_6053;
assign n_6430 = n_6428 ^ n_5713;
assign y56 = ~n_6429;
assign n_6431 = n_6053 & n_6430;
assign n_6432 = n_6431 ^ n_6428;
assign n_6433 = n_6432 ^ n_5983;
assign n_6434 = n_6432 ^ n_5608;
assign y57 = n_6433;
assign n_6435 = ~n_5983 & ~n_6434;
assign n_6436 = n_6435 ^ n_6432;
assign n_6437 = n_6436 ^ n_5913;
assign n_6438 = n_6436 ^ n_5465;
assign y58 = n_6437;
assign n_6439 = ~n_5913 & n_6438;
assign n_6440 = n_6439 ^ n_6436;
assign n_6441 = n_6440 ^ n_5823;
assign n_6442 = n_6440 ^ n_5466;
assign y59 = ~n_6441;
assign n_6443 = n_5823 & ~n_6442;
assign n_6444 = n_6443 ^ n_6440;
assign n_6445 = n_6444 ^ n_5824;
assign n_6446 = n_6444 ^ n_5468;
assign y60 = ~n_6445;
assign n_6447 = n_5824 & n_6446;
assign n_6448 = n_6447 ^ n_6444;
assign n_6449 = n_6448 ^ n_5825;
assign n_6450 = n_6448 ^ n_4941;
assign y61 = ~n_6449;
assign n_6451 = n_5825 & ~n_6450;
assign n_6452 = n_6451 ^ n_6448;
assign n_6453 = n_6452 ^ n_5470;
assign n_6454 = n_6452 ^ n_4942;
assign y62 = ~n_6453;
assign n_6455 = n_5470 & ~n_6454;
assign n_6456 = n_6455 ^ n_6452;
assign n_6457 = n_6456 ^ n_5471;
assign y63 = n_6457;
endmodule