module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n211 , n212 , n213 , n214 , n217 , n218 , n219 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n273 , n274 , n275 , n276 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n295 , n296 , n297 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n449 , n450 , n451 , n452 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n539 , n540 , n541 , n542 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n639 , n640 , n641 , n642 , n647 , n648 , n649 , n650 , n651 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n786 , n787 , n788 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n872 , n873 , n874 , n875 , n876 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n913 , n914 , n915 , n920 , n921 , n922 , n923 , n924 , n925 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1110 , n1111 , n1112 , n1113 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1138 , n1139 , n1140 , n1141 , n1142 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1200 , n1201 , n1202 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1260 , n1261 , n1262 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1326 , n1327 , n1328 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1380 , n1381 , n1382 , n1383 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1489 , n1490 , n1491 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1521 , n1522 , n1523 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1604 , n1605 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1682 , n1683 , n1684 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1847 , n1848 , n1849 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1911 , n1912 , n1913 , n1914 , n1915 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2114 , n2116 , n2117 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2264 , n2265 , n2266 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2401 , n2402 , n2403 , n2404 , n2405 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2617 , n2618 , n2619 , n2620 , n2621 , n2624 , n2625 , n2626 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2814 , n2815 , n2816 , n2817 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3035 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3177 , n3178 , n3179 , n3180 , n3183 , n3184 , n3185 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3379 , n3380 , n3381 , n3382 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3448 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4757 , n4758 , n4759 , n4760 , n4761 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6741 , n6742 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7447 , n7448 , n7449 , n7450 , n7451 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8473 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9556 , n9557 , n9558 , n9559 , n9560 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10577 , n10578 , n10579 , n10580 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12627 , n12628 , n12629 , n12630 , n12631 , n12633 , n12634 , n12635 , n12636 , n12637 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14739 , n14740 , n14741 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14761 , n14762 , n14763 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15354 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15706 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15914 , n15915 , n15916 , n15917 , n15918 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16134 , n16135 , n16136 , n16137 , n16138 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16776 , n16777 , n16778 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17294 , n17295 , n17296 , n17297 , n17298 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17547 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18990 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19583 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19814 , n19815 , n19816 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20700 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23986 , n23987 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24825 , n24826 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24845 , n24846 , n24847 , n24848 , n24849 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 ;
  assign n129 = x122 ^ x34 ;
  assign n135 = x64 ^ x26 ;
  assign n136 = x81 ^ x2 ;
  assign n137 = n135 & n136 ;
  assign n138 = n137 ^ n135 ;
  assign n132 = x99 ^ x18 ;
  assign n133 = x90 ^ x10 ;
  assign n134 = n132 & ~n133 ;
  assign n143 = n134 ^ n132 ;
  assign n144 = n143 ^ n133 ;
  assign n151 = n144 ^ n132 ;
  assign n152 = n138 & ~n151 ;
  assign n202 = n152 ^ n151 ;
  assign n158 = n136 & ~n151 ;
  assign n203 = n202 ^ n158 ;
  assign n145 = n137 ^ n136 ;
  assign n146 = n144 & n145 ;
  assign n147 = n146 ^ n137 ;
  assign n142 = ~n133 & n137 ;
  assign n148 = n147 ^ n142 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n134 & ~n139 ;
  assign n199 = n148 ^ n140 ;
  assign n197 = n136 ^ n135 ;
  assign n198 = n197 ^ n132 ;
  assign n200 = n199 ^ n198 ;
  assign n204 = n203 ^ n200 ;
  assign n154 = n132 & n135 ;
  assign n155 = n154 ^ n143 ;
  assign n141 = n133 & n136 ;
  assign n149 = n148 ^ n141 ;
  assign n163 = n155 ^ n149 ;
  assign n156 = ~n136 & n155 ;
  assign n164 = n163 ^ n156 ;
  assign n160 = n133 ^ n132 ;
  assign n161 = n145 ^ n141 ;
  assign n162 = ~n160 & n161 ;
  assign n165 = n164 ^ n162 ;
  assign n166 = n165 ^ n146 ;
  assign n159 = n158 ^ n147 ;
  assign n167 = n166 ^ n159 ;
  assign n168 = n167 ^ n162 ;
  assign n186 = n168 ^ n161 ;
  assign n205 = n204 ^ n186 ;
  assign n188 = n138 & n143 ;
  assign n196 = n188 ^ n140 ;
  assign n201 = n200 ^ n196 ;
  assign n206 = n205 ^ n201 ;
  assign n1286 = ~n129 & n206 ;
  assign n1287 = n1286 ^ n205 ;
  assign n130 = x104 ^ x60 ;
  assign n214 = n167 ^ n149 ;
  assign n217 = n129 & n214 ;
  assign n218 = n217 ^ n149 ;
  assign n219 = n130 & n218 ;
  assign n1291 = n1287 ^ n219 ;
  assign n179 = n135 ^ n133 ;
  assign n195 = n179 ^ n168 ;
  assign n207 = n206 ^ n195 ;
  assign n208 = n207 ^ n203 ;
  assign n211 = ~n129 & ~n208 ;
  assign n212 = n211 ^ n203 ;
  assign n213 = n130 & ~n212 ;
  assign n1292 = n1291 ^ n213 ;
  assign n1293 = n1292 ^ x51 ;
  assign n1285 = n196 ^ n166 ;
  assign n1288 = n1287 ^ n1285 ;
  assign n182 = ~n139 & n144 ;
  assign n1282 = n182 ^ n166 ;
  assign n323 = n186 ^ n142 ;
  assign n1283 = n1282 ^ n323 ;
  assign n1284 = ~n129 & n1283 ;
  assign n1289 = n1288 ^ n1284 ;
  assign n1290 = n130 & ~n1289 ;
  assign n1294 = n1293 ^ n1290 ;
  assign n1295 = n1294 ^ x81 ;
  assign n1351 = x114 ^ x56 ;
  assign n1352 = x123 ^ x40 ;
  assign n1353 = n1351 & n1352 ;
  assign n1354 = x97 ^ x48 ;
  assign n1355 = x112 ^ x32 ;
  assign n1356 = n1354 & ~n1355 ;
  assign n1357 = n1353 & n1356 ;
  assign n1358 = x80 ^ x24 ;
  assign n1391 = x73 ^ x6 ;
  assign n1420 = ~n1358 & n1391 ;
  assign n1380 = n1354 ^ n1351 ;
  assign n1381 = n1355 ^ n1352 ;
  assign n1359 = n1355 ^ n1354 ;
  assign n1361 = n1352 & n1359 ;
  assign n1382 = n1381 ^ n1361 ;
  assign n1383 = ~n1380 & n1382 ;
  assign n1387 = n1383 ^ n1380 ;
  assign n1373 = n1354 ^ n1352 ;
  assign n1374 = ~n1355 & n1373 ;
  assign n1375 = n1374 ^ n1352 ;
  assign n1376 = ~n1351 & n1375 ;
  assign n1386 = n1376 ^ n1375 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1360 = n1353 & n1359 ;
  assign n1385 = n1360 ^ n1357 ;
  assign n1389 = n1388 ^ n1385 ;
  assign n1363 = n1353 ^ n1351 ;
  assign n1364 = n1363 ^ n1352 ;
  assign n1368 = n1356 ^ n1355 ;
  assign n1369 = n1368 ^ n1354 ;
  assign n1370 = ~n1364 & n1369 ;
  assign n1454 = n1389 ^ n1370 ;
  assign n1455 = n1420 & ~n1454 ;
  assign n1429 = n1356 ^ n1354 ;
  assign n1409 = n1363 & ~n1368 ;
  assign n1365 = n1364 ^ n1351 ;
  assign n1366 = n1356 & n1365 ;
  assign n1362 = n1361 ^ n1360 ;
  assign n1367 = n1366 ^ n1362 ;
  assign n1397 = n1383 ^ n1367 ;
  assign n1371 = n1356 & ~n1364 ;
  assign n1372 = n1371 ^ n1365 ;
  assign n1377 = n1376 ^ n1372 ;
  assign n1378 = n1377 ^ n1370 ;
  assign n1398 = n1397 ^ n1378 ;
  assign n1410 = n1409 ^ n1398 ;
  assign n1407 = n1363 & n1369 ;
  assign n1408 = n1407 ^ n1363 ;
  assign n1411 = n1410 ^ n1408 ;
  assign n1424 = n1411 ^ n1360 ;
  assign n1430 = n1429 ^ n1424 ;
  assign n1426 = n1424 ^ n1398 ;
  assign n1405 = n1365 ^ n1362 ;
  assign n1406 = n1405 ^ n1377 ;
  assign n1427 = n1426 ^ n1406 ;
  assign n1425 = n1424 ^ n1386 ;
  assign n1428 = n1427 ^ n1425 ;
  assign n1431 = n1430 ^ n1428 ;
  assign n1436 = n1431 ^ n1366 ;
  assign n1432 = n1431 ^ n1377 ;
  assign n1433 = n1432 ^ n1367 ;
  assign n1434 = n1433 ^ n1407 ;
  assign n1435 = n1434 ^ n1386 ;
  assign n1437 = n1436 ^ n1435 ;
  assign n1438 = n1391 & n1437 ;
  assign n1439 = n1438 ^ n1434 ;
  assign n1456 = n1455 ^ n1439 ;
  assign n1448 = n1420 ^ n1358 ;
  assign n1451 = n1409 ^ n1370 ;
  assign n1412 = n1411 ^ n1353 ;
  assign n1413 = n1412 ^ n1386 ;
  assign n1449 = n1413 ^ n1411 ;
  assign n1450 = n1449 ^ n1425 ;
  assign n1452 = n1451 ^ n1450 ;
  assign n1453 = ~n1448 & n1452 ;
  assign n1457 = n1456 ^ n1453 ;
  assign n1441 = n1439 ^ n1376 ;
  assign n1440 = n1439 ^ n1371 ;
  assign n1442 = n1441 ^ n1440 ;
  assign n1445 = ~n1391 & n1442 ;
  assign n1446 = n1445 ^ n1441 ;
  assign n1421 = n1420 ^ n1391 ;
  assign n1714 = n1448 ^ n1421 ;
  assign n1447 = n1446 & ~n1714 ;
  assign n1458 = n1457 ^ n1447 ;
  assign n1422 = n1409 & n1421 ;
  assign n1459 = n1458 ^ n1422 ;
  assign n1414 = n1413 ^ n1406 ;
  assign n1417 = ~n1391 & n1414 ;
  assign n1418 = n1417 ^ n1413 ;
  assign n1419 = n1358 & n1418 ;
  assign n1460 = n1459 ^ n1419 ;
  assign n1399 = n1398 ^ n1367 ;
  assign n1402 = n1358 & n1399 ;
  assign n1403 = n1402 ^ n1367 ;
  assign n1404 = ~n1391 & n1403 ;
  assign n1461 = n1460 ^ n1404 ;
  assign n1390 = n1398 ^ n1389 ;
  assign n1394 = ~n1390 & n1391 ;
  assign n1395 = n1394 ^ n1389 ;
  assign n1396 = n1358 & ~n1395 ;
  assign n1462 = n1461 ^ n1396 ;
  assign n1463 = ~n1357 & ~n1462 ;
  assign n1464 = n1463 ^ x59 ;
  assign n1465 = n1464 ^ x90 ;
  assign n1471 = ~n1295 & n1465 ;
  assign n1472 = n1471 ^ n1295 ;
  assign n227 = x78 ^ x38 ;
  assign n228 = x84 ^ x62 ;
  assign n229 = n227 & ~n228 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = x101 ^ x54 ;
  assign n232 = x126 ^ x46 ;
  assign n233 = ~n231 & n232 ;
  assign n234 = n233 ^ n231 ;
  assign n240 = n234 ^ n232 ;
  assign n251 = ~n230 & n240 ;
  assign n243 = n233 ^ n232 ;
  assign n244 = n229 & n243 ;
  assign n241 = n229 & n240 ;
  assign n237 = ~n230 & n233 ;
  assign n242 = n241 ^ n237 ;
  assign n245 = n244 ^ n242 ;
  assign n236 = n229 & n233 ;
  assign n238 = n237 ^ n236 ;
  assign n239 = n238 ^ n229 ;
  assign n246 = n245 ^ n239 ;
  assign n252 = n251 ^ n246 ;
  assign n273 = n252 ^ n236 ;
  assign n285 = n273 ^ n228 ;
  assign n255 = n230 ^ n227 ;
  assign n256 = n255 ^ n228 ;
  assign n257 = n243 & n256 ;
  assign n258 = n257 ^ n244 ;
  assign n259 = n258 ^ n243 ;
  assign n253 = n252 ^ n244 ;
  assign n235 = ~n230 & ~n234 ;
  assign n248 = n241 ^ n235 ;
  assign n249 = n248 ^ n238 ;
  assign n250 = n249 ^ n228 ;
  assign n254 = n253 ^ n250 ;
  assign n260 = n259 ^ n254 ;
  assign n284 = n260 ^ n239 ;
  assign n286 = n285 ^ n284 ;
  assign n282 = n232 ^ n228 ;
  assign n283 = n282 ^ n227 ;
  assign n287 = n286 ^ n283 ;
  assign n226 = x83 ^ x30 ;
  assign n276 = x124 ^ x4 ;
  assign n288 = n226 & n276 ;
  assign n289 = n288 ^ n276 ;
  assign n1316 = n287 & n289 ;
  assign n311 = n240 & n256 ;
  assign n1304 = n311 ^ n242 ;
  assign n1305 = n1304 ^ n284 ;
  assign n264 = n233 & n256 ;
  assign n263 = n238 ^ n233 ;
  assign n265 = n264 ^ n263 ;
  assign n262 = n240 & n255 ;
  assign n266 = n265 ^ n262 ;
  assign n261 = n260 ^ n255 ;
  assign n267 = n266 ^ n261 ;
  assign n1302 = n267 ^ n257 ;
  assign n1303 = n1302 ^ n265 ;
  assign n1306 = n1305 ^ n1303 ;
  assign n1307 = ~n226 & n1306 ;
  assign n1308 = n1307 ^ n284 ;
  assign n305 = n288 ^ n226 ;
  assign n268 = n267 ^ n234 ;
  assign n247 = n246 ^ n235 ;
  assign n269 = n268 ^ n247 ;
  assign n306 = n269 ^ n262 ;
  assign n307 = n305 & n306 ;
  assign n1311 = n1308 ^ n307 ;
  assign n292 = n254 ^ n251 ;
  assign n295 = ~n276 & ~n292 ;
  assign n296 = n295 ^ n251 ;
  assign n297 = n226 & n296 ;
  assign n1312 = n1311 ^ n297 ;
  assign n1313 = n1312 ^ x35 ;
  assign n1298 = n262 ^ n236 ;
  assign n1299 = n1298 ^ n255 ;
  assign n1300 = n1299 ^ n311 ;
  assign n1301 = n226 & n1300 ;
  assign n1309 = n1308 ^ n1301 ;
  assign n1310 = n276 & ~n1309 ;
  assign n1314 = n1313 ^ n1310 ;
  assign n315 = n254 ^ n246 ;
  assign n1296 = n276 ^ n226 ;
  assign n1297 = ~n315 & ~n1296 ;
  assign n1315 = n1314 ^ n1297 ;
  assign n1317 = n1316 ^ n1315 ;
  assign n1318 = n1317 ^ x99 ;
  assign n583 = x110 ^ x36 ;
  assign n582 = x92 ^ x62 ;
  assign n584 = n583 ^ n582 ;
  assign n585 = x68 ^ x20 ;
  assign n586 = x86 ^ x4 ;
  assign n587 = n585 & ~n586 ;
  assign n588 = n587 ^ n586 ;
  assign n589 = n588 ^ n585 ;
  assign n590 = n589 ^ n586 ;
  assign n591 = x93 ^ x28 ;
  assign n596 = n590 & n591 ;
  assign n592 = x116 ^ x12 ;
  assign n1342 = n596 ^ n592 ;
  assign n601 = n586 ^ n585 ;
  assign n602 = n601 ^ n591 ;
  assign n1343 = n1342 ^ n602 ;
  assign n1344 = ~n582 & n1343 ;
  assign n593 = n591 & n592 ;
  assign n619 = n593 ^ n592 ;
  assign n620 = n587 & n619 ;
  assign n1345 = n1344 ^ n620 ;
  assign n1346 = n584 & n1345 ;
  assign n626 = n590 & n619 ;
  assign n627 = n626 ^ n590 ;
  assign n628 = n627 ^ n596 ;
  assign n604 = ~n588 & ~n591 ;
  assign n629 = n628 ^ n604 ;
  assign n622 = n592 ^ n586 ;
  assign n630 = n629 ^ n622 ;
  assign n623 = ~n592 & ~n622 ;
  assign n624 = n623 ^ n591 ;
  assign n625 = ~n585 & n624 ;
  assign n631 = n630 ^ n625 ;
  assign n606 = n589 & n593 ;
  assign n632 = n631 ^ n606 ;
  assign n607 = n606 ^ n593 ;
  assign n605 = n604 ^ n588 ;
  assign n608 = n607 ^ n605 ;
  assign n603 = ~n585 & n602 ;
  assign n609 = n608 ^ n603 ;
  assign n610 = n609 ^ n591 ;
  assign n611 = n610 ^ n601 ;
  assign n594 = n593 ^ n591 ;
  assign n598 = n585 & ~n594 ;
  assign n599 = n598 ^ n585 ;
  assign n600 = n599 ^ n587 ;
  assign n612 = n611 ^ n600 ;
  assign n613 = n612 ^ n606 ;
  assign n614 = n613 ^ n593 ;
  assign n615 = n614 ^ n608 ;
  assign n595 = n590 & n594 ;
  assign n597 = n596 ^ n595 ;
  assign n616 = n615 ^ n597 ;
  assign n617 = n616 ^ n607 ;
  assign n618 = n617 ^ n595 ;
  assign n621 = n620 ^ n618 ;
  assign n633 = n632 ^ n621 ;
  assign n896 = n633 ^ n589 ;
  assign n858 = n604 ^ n585 ;
  assign n859 = n858 ^ n603 ;
  assign n897 = n896 ^ n859 ;
  assign n875 = n606 ^ n600 ;
  assign n876 = n875 ^ n631 ;
  assign n898 = n897 ^ n876 ;
  assign n1333 = ~n582 & ~n898 ;
  assign n1334 = n1333 ^ n876 ;
  assign n1335 = ~n583 & n1334 ;
  assign n1336 = n1335 ^ n620 ;
  assign n853 = n619 ^ n591 ;
  assign n884 = n876 ^ n853 ;
  assign n885 = n884 ^ n629 ;
  assign n663 = n582 & ~n583 ;
  assign n886 = n663 ^ n626 ;
  assign n887 = n886 ^ n583 ;
  assign n888 = ~n885 & n887 ;
  assign n889 = n888 ^ n626 ;
  assign n890 = n885 ^ n663 ;
  assign n891 = n890 ^ n582 ;
  assign n892 = n889 & ~n891 ;
  assign n893 = n892 ^ n885 ;
  assign n1337 = n1336 ^ n893 ;
  assign n895 = n853 ^ n618 ;
  assign n899 = n898 ^ n895 ;
  assign n900 = n582 & n899 ;
  assign n901 = n900 ^ n628 ;
  assign n902 = ~n583 & n901 ;
  assign n1338 = n1337 ^ n902 ;
  assign n1339 = n1338 ^ x43 ;
  assign n860 = n859 ^ n606 ;
  assign n654 = n599 ^ n595 ;
  assign n861 = n860 ^ n654 ;
  assign n1322 = n861 ^ n633 ;
  assign n1320 = n616 ^ n595 ;
  assign n1321 = n1320 ^ n654 ;
  assign n1323 = n1322 ^ n1321 ;
  assign n1326 = n583 & ~n1323 ;
  assign n1327 = n1326 ^ n1321 ;
  assign n1328 = ~n584 & n1327 ;
  assign n1340 = n1339 ^ n1328 ;
  assign n1319 = n582 & ~n613 ;
  assign n1341 = n1340 ^ n1319 ;
  assign n1347 = n1346 ^ n1341 ;
  assign n1348 = n1347 ^ x80 ;
  assign n1468 = n1318 & n1348 ;
  assign n1469 = n1468 ^ n1318 ;
  assign n1470 = n1469 ^ n1348 ;
  assign n1475 = n1470 ^ n1318 ;
  assign n1489 = ~n1472 & n1475 ;
  assign n474 = x85 ^ x2 ;
  assign n477 = x91 ^ x60 ;
  assign n476 = x100 ^ x36 ;
  assign n475 = x117 ^ x44 ;
  assign n483 = x102 ^ x52 ;
  assign n490 = n475 & ~n483 ;
  assign n495 = n476 & n490 ;
  assign n514 = ~n477 & n495 ;
  assign n484 = ~n477 & n483 ;
  assign n487 = n476 & n484 ;
  assign n481 = n475 & ~n476 ;
  assign n485 = n481 & n484 ;
  assign n486 = n485 ^ n484 ;
  assign n488 = n487 ^ n486 ;
  assign n575 = n514 ^ n488 ;
  assign n501 = n476 & n477 ;
  assign n502 = ~n475 & n501 ;
  assign n524 = n502 ^ n501 ;
  assign n517 = n514 ^ n495 ;
  assign n525 = n524 ^ n517 ;
  assign n1511 = n575 ^ n525 ;
  assign n496 = n495 ^ n490 ;
  assign n512 = ~n477 & n496 ;
  assign n532 = n512 ^ n496 ;
  assign n506 = n475 & n487 ;
  assign n507 = n506 ^ n487 ;
  assign n503 = n483 & n502 ;
  assign n504 = n503 ^ n502 ;
  assign n497 = n496 ^ n481 ;
  assign n492 = n476 ^ n475 ;
  assign n493 = n483 ^ n475 ;
  assign n494 = n492 & ~n493 ;
  assign n498 = n497 ^ n494 ;
  assign n505 = n504 ^ n498 ;
  assign n508 = n507 ^ n505 ;
  assign n491 = n490 ^ n483 ;
  assign n499 = n498 ^ n491 ;
  assign n482 = n481 ^ n476 ;
  assign n489 = n488 ^ n482 ;
  assign n500 = n499 ^ n489 ;
  assign n509 = n508 ^ n500 ;
  assign n478 = n477 ^ n476 ;
  assign n479 = n478 ^ n475 ;
  assign n480 = ~n475 & n479 ;
  assign n510 = n509 ^ n480 ;
  assign n511 = n510 ^ n507 ;
  assign n533 = n532 ^ n511 ;
  assign n534 = n533 ^ n506 ;
  assign n1512 = n1511 ^ n534 ;
  assign n548 = n497 ^ n485 ;
  assign n1510 = n548 ^ n511 ;
  assign n1513 = n1512 ^ n1510 ;
  assign n1514 = n474 & n1513 ;
  assign n1515 = n1514 ^ n1510 ;
  assign n473 = x67 ^ x28 ;
  assign n549 = ~n473 & n474 ;
  assign n550 = n549 ^ n473 ;
  assign n551 = n550 ^ n474 ;
  assign n552 = n551 ^ n473 ;
  assign n972 = n512 ^ n505 ;
  assign n973 = n552 & n972 ;
  assign n572 = n485 & n551 ;
  assign n974 = n973 ^ n572 ;
  assign n1531 = n1515 ^ n974 ;
  assign n554 = n474 ^ n473 ;
  assign n1528 = ~n473 & n508 ;
  assign n1529 = n1528 ^ n507 ;
  assign n1530 = ~n554 & n1529 ;
  assign n1532 = n1531 ^ n1530 ;
  assign n563 = n474 & n504 ;
  assign n555 = n525 ^ n500 ;
  assign n556 = n555 ^ n517 ;
  assign n557 = ~n473 & n556 ;
  assign n558 = n557 ^ n517 ;
  assign n564 = n563 ^ n558 ;
  assign n565 = n554 & n564 ;
  assign n566 = n565 ^ n558 ;
  assign n1533 = n1532 ^ n566 ;
  assign n518 = n517 ^ n485 ;
  assign n542 = n518 ^ n505 ;
  assign n545 = ~n473 & n542 ;
  assign n546 = n545 ^ n505 ;
  assign n547 = ~n474 & n546 ;
  assign n1534 = n1533 ^ n547 ;
  assign n1535 = n1534 ^ x1 ;
  assign n515 = n514 ^ n503 ;
  assign n1516 = n1515 ^ n515 ;
  assign n995 = n548 ^ n517 ;
  assign n996 = n995 ^ n532 ;
  assign n523 = n510 ^ n499 ;
  assign n997 = n996 ^ n523 ;
  assign n1517 = n1516 ^ n997 ;
  assign n1518 = n1517 ^ n1515 ;
  assign n1521 = ~n474 & ~n1518 ;
  assign n1522 = n1521 ^ n1515 ;
  assign n1523 = n473 & n1522 ;
  assign n1536 = n1535 ^ n1523 ;
  assign n1507 = n523 ^ n504 ;
  assign n521 = n506 ^ n500 ;
  assign n1508 = n1507 ^ n521 ;
  assign n1509 = n552 & ~n1508 ;
  assign n1537 = n1536 ^ n1509 ;
  assign n1538 = n1537 ^ x123 ;
  assign n346 = x72 ^ x8 ;
  assign n347 = x82 ^ x0 ;
  assign n348 = n346 & n347 ;
  assign n350 = x65 ^ x16 ;
  assign n351 = x120 ^ x24 ;
  assign n352 = ~n350 & ~n351 ;
  assign n353 = n352 ^ n350 ;
  assign n354 = n353 ^ n351 ;
  assign n365 = n348 & ~n354 ;
  assign n420 = n365 ^ n354 ;
  assign n349 = n348 ^ n347 ;
  assign n372 = n349 ^ n346 ;
  assign n373 = n372 ^ n347 ;
  assign n378 = ~n354 & n373 ;
  assign n355 = n349 & ~n354 ;
  assign n379 = n378 ^ n355 ;
  assign n421 = n420 ^ n379 ;
  assign n391 = n349 & ~n353 ;
  assign n422 = n421 ^ n391 ;
  assign n374 = ~n353 & n373 ;
  assign n375 = n374 ^ n355 ;
  assign n423 = n422 ^ n375 ;
  assign n424 = n423 ^ n421 ;
  assign n431 = n354 ^ n350 ;
  assign n432 = ~n372 & ~n431 ;
  assign n387 = n348 & n352 ;
  assign n388 = n387 ^ n365 ;
  assign n356 = n348 & ~n353 ;
  assign n386 = n356 ^ n348 ;
  assign n389 = n388 ^ n386 ;
  assign n433 = n432 ^ n389 ;
  assign n380 = n379 ^ n373 ;
  assign n376 = n352 & n373 ;
  assign n377 = n376 ^ n375 ;
  assign n381 = n380 ^ n377 ;
  assign n434 = n433 ^ n381 ;
  assign n1265 = n434 ^ n387 ;
  assign n358 = x96 ^ x32 ;
  assign n359 = x105 ^ x58 ;
  assign n360 = ~n358 & n359 ;
  assign n361 = n360 ^ n358 ;
  assign n1266 = n1265 ^ n361 ;
  assign n1267 = ~n424 & n1266 ;
  assign n1268 = n1267 ^ n361 ;
  assign n393 = n424 ^ n353 ;
  assign n357 = n356 ^ n355 ;
  assign n394 = n393 ^ n357 ;
  assign n446 = n394 ^ n378 ;
  assign n449 = n358 & ~n446 ;
  assign n450 = n449 ^ n378 ;
  assign n451 = ~n359 & n450 ;
  assign n1270 = n451 ^ n424 ;
  assign n362 = n361 ^ n359 ;
  assign n363 = n362 ^ n358 ;
  assign n1269 = n451 ^ n363 ;
  assign n1271 = n1270 ^ n1269 ;
  assign n1272 = ~n1268 & n1271 ;
  assign n1273 = n1272 ^ n1269 ;
  assign n385 = n359 ^ n358 ;
  assign n390 = n389 ^ n376 ;
  assign n1256 = n390 ^ n356 ;
  assign n1255 = n387 ^ n374 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1260 = n358 & n1257 ;
  assign n1261 = n1260 ^ n1255 ;
  assign n1262 = n385 & n1261 ;
  assign n1274 = n1273 ^ n1262 ;
  assign n940 = n362 & n379 ;
  assign n1275 = n1274 ^ n940 ;
  assign n435 = n434 ^ n431 ;
  assign n398 = n352 & ~n372 ;
  assign n436 = n435 ^ n398 ;
  assign n437 = n436 ^ n365 ;
  assign n440 = n358 & ~n437 ;
  assign n441 = n440 ^ n365 ;
  assign n442 = n385 & n441 ;
  assign n1276 = n1275 ^ n442 ;
  assign n382 = n349 & n352 ;
  assign n383 = n382 ^ n381 ;
  assign n941 = n436 ^ n383 ;
  assign n944 = n359 & ~n941 ;
  assign n945 = n944 ^ n383 ;
  assign n946 = ~n358 & n945 ;
  assign n444 = n363 & ~n421 ;
  assign n947 = n946 ^ n444 ;
  assign n1277 = n1276 ^ n947 ;
  assign n1249 = n433 ^ n422 ;
  assign n1252 = n359 & ~n1249 ;
  assign n1253 = n1252 ^ n433 ;
  assign n1254 = ~n358 & n1253 ;
  assign n1278 = n1277 ^ n1254 ;
  assign n467 = n360 & n376 ;
  assign n1279 = n1278 ^ n467 ;
  assign n1280 = n1279 ^ x27 ;
  assign n1281 = n1280 ^ x113 ;
  assign n1544 = n1538 ^ n1281 ;
  assign n1602 = n1489 & n1544 ;
  assign n1490 = n1468 & ~n1472 ;
  assign n1474 = n1471 ^ n1465 ;
  assign n1478 = n1474 ^ n1295 ;
  assign n1481 = ~n1470 & n1478 ;
  assign n1496 = n1490 ^ n1481 ;
  assign n1479 = n1468 & n1478 ;
  assign n1497 = n1496 ^ n1479 ;
  assign n1498 = n1497 ^ n1478 ;
  assign n1485 = n1469 & n1478 ;
  assign n1495 = n1490 ^ n1485 ;
  assign n1499 = n1498 ^ n1495 ;
  assign n1553 = n1281 & n1538 ;
  assign n1574 = n1553 ^ n1538 ;
  assign n1595 = n1574 ^ n1281 ;
  assign n1600 = n1499 & ~n1595 ;
  assign n1503 = n1468 & n1471 ;
  assign n1476 = n1474 & n1475 ;
  assign n1500 = n1499 ^ n1476 ;
  assign n1494 = n1489 ^ n1475 ;
  assign n1501 = n1500 ^ n1494 ;
  assign n1491 = n1490 ^ n1489 ;
  assign n1473 = ~n1470 & ~n1472 ;
  assign n1545 = n1491 ^ n1473 ;
  assign n1546 = n1545 ^ n1472 ;
  assign n1480 = n1479 ^ n1473 ;
  assign n1482 = n1481 ^ n1480 ;
  assign n1477 = n1476 ^ n1473 ;
  assign n1483 = n1482 ^ n1477 ;
  assign n1349 = n1348 ^ n1318 ;
  assign n1350 = n1349 ^ n1295 ;
  assign n1466 = n1465 ^ n1350 ;
  assign n1467 = n1295 & n1466 ;
  assign n1484 = n1483 ^ n1467 ;
  assign n1486 = n1485 ^ n1484 ;
  assign n1487 = n1486 ^ n1469 ;
  assign n1493 = n1546 ^ n1487 ;
  assign n1502 = n1501 ^ n1493 ;
  assign n1504 = n1503 ^ n1502 ;
  assign n1583 = n1504 ^ n1471 ;
  assign n1559 = n1502 ^ n1477 ;
  assign n1556 = n1490 ^ n1468 ;
  assign n1555 = n1503 ^ n1479 ;
  assign n1557 = n1556 ^ n1555 ;
  assign n1558 = n1557 ^ n1495 ;
  assign n1560 = n1559 ^ n1558 ;
  assign n1561 = n1560 ^ n1466 ;
  assign n1562 = n1561 ^ n1500 ;
  assign n1596 = n1583 ^ n1562 ;
  assign n1597 = ~n1595 & ~n1596 ;
  assign n1575 = n1476 & n1574 ;
  assign n1571 = n1538 & n1555 ;
  assign n1572 = n1571 ^ n1479 ;
  assign n1573 = ~n1281 & n1572 ;
  assign n1576 = n1575 ^ n1573 ;
  assign n1579 = n1501 ^ n1484 ;
  assign n1580 = n1579 ^ n1490 ;
  assign n1581 = n1580 ^ n1473 ;
  assign n1577 = n1493 ^ n1481 ;
  assign n1563 = n1562 ^ n1557 ;
  assign n1578 = n1577 ^ n1563 ;
  assign n1589 = n1581 ^ n1578 ;
  assign n1590 = n1538 & ~n1589 ;
  assign n1582 = n1497 ^ n1485 ;
  assign n1584 = n1583 ^ n1582 ;
  assign n1585 = n1538 & ~n1584 ;
  assign n1586 = n1585 ^ n1486 ;
  assign n1587 = n1586 ^ n1581 ;
  assign n1591 = n1590 ^ n1587 ;
  assign n1592 = ~n1281 & n1591 ;
  assign n1593 = n1592 ^ n1586 ;
  assign n1594 = ~n1576 & ~n1593 ;
  assign n1598 = n1597 ^ n1594 ;
  assign n1554 = n1553 ^ n1281 ;
  assign n1564 = n1554 & n1563 ;
  assign n1547 = n1546 ^ n1473 ;
  assign n1550 = n1538 & ~n1547 ;
  assign n1551 = n1550 ^ n1473 ;
  assign n1552 = n1544 & n1551 ;
  assign n1565 = n1564 ^ n1552 ;
  assign n1541 = ~n1504 & n1538 ;
  assign n1542 = n1541 ^ n1503 ;
  assign n1543 = n1281 & n1542 ;
  assign n1566 = n1565 ^ n1543 ;
  assign n1599 = n1598 ^ n1566 ;
  assign n1601 = n1600 ^ n1599 ;
  assign n1604 = n1602 ^ n1601 ;
  assign n1605 = n1546 ^ n1499 ;
  assign n1610 = ~n1538 & ~n1605 ;
  assign n1611 = n1610 ^ n1499 ;
  assign n1612 = n1281 & n1611 ;
  assign n1613 = n1604 & ~n1612 ;
  assign n1614 = n1613 ^ x2 ;
  assign n2252 = n1614 ^ x124 ;
  assign n1077 = x121 ^ x26 ;
  assign n1075 = x66 ^ x0 ;
  assign n1083 = n1077 ^ n1075 ;
  assign n1067 = x98 ^ x58 ;
  assign n1068 = x89 ^ x50 ;
  assign n1069 = n1067 & n1068 ;
  assign n1064 = x107 ^ x34 ;
  assign n1065 = x88 ^ x42 ;
  assign n1066 = n1064 & ~n1065 ;
  assign n1078 = n1066 ^ n1064 ;
  assign n1079 = n1069 & n1078 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1071 = n1066 & n1070 ;
  assign n1131 = n1079 ^ n1071 ;
  assign n1130 = n1067 ^ n1065 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1084 = n1069 ^ n1067 ;
  assign n1091 = n1078 & n1084 ;
  assign n1085 = n1078 ^ n1065 ;
  assign n1090 = n1069 & n1085 ;
  assign n1092 = n1091 ^ n1090 ;
  assign n1088 = n1066 ^ n1065 ;
  assign n1089 = n1070 & ~n1088 ;
  assign n1093 = n1092 ^ n1089 ;
  assign n1086 = n1084 & n1085 ;
  assign n1072 = n1070 ^ n1067 ;
  assign n1073 = n1066 & ~n1072 ;
  assign n1087 = n1086 ^ n1073 ;
  assign n1094 = n1093 ^ n1087 ;
  assign n1133 = n1132 ^ n1094 ;
  assign n1113 = n1070 & n1078 ;
  assign n1128 = n1113 ^ n1078 ;
  assign n1127 = n1091 ^ n1079 ;
  assign n1129 = n1128 ^ n1127 ;
  assign n1134 = n1133 ^ n1129 ;
  assign n1126 = n1073 ^ n1072 ;
  assign n1135 = n1134 ^ n1126 ;
  assign n1138 = ~n1075 & n1135 ;
  assign n1099 = n1069 & ~n1088 ;
  assign n1100 = n1099 ^ n1092 ;
  assign n1097 = n1068 ^ n1064 ;
  assign n1098 = n1067 & n1097 ;
  assign n1101 = n1100 ^ n1098 ;
  assign n1122 = n1101 ^ n1066 ;
  assign n1074 = n1073 ^ n1071 ;
  assign n1123 = n1122 ^ n1074 ;
  assign n1139 = n1138 ^ n1123 ;
  assign n1140 = n1083 & n1139 ;
  assign n1141 = n1140 ^ n1123 ;
  assign n2087 = n1141 ^ n1071 ;
  assign n1142 = n1135 ^ n1129 ;
  assign n1145 = ~n1077 & n1142 ;
  assign n1146 = n1145 ^ n1129 ;
  assign n1147 = n1075 & n1146 ;
  assign n2088 = n2087 ^ n1147 ;
  assign n1118 = n1075 & n1113 ;
  assign n1103 = n1091 ^ n1084 ;
  assign n1102 = n1101 ^ n1086 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1119 = n1118 ^ n1104 ;
  assign n1120 = n1083 & n1119 ;
  assign n1121 = n1120 ^ n1104 ;
  assign n2089 = n2088 ^ n1121 ;
  assign n1920 = n1075 & ~n1134 ;
  assign n1921 = n1920 ^ n1135 ;
  assign n1922 = n1083 & n1921 ;
  assign n1923 = n1922 ^ n1135 ;
  assign n2090 = n2089 ^ n1923 ;
  assign n1640 = n1075 & ~n1077 ;
  assign n1641 = n1640 ^ n1077 ;
  assign n1642 = n1641 ^ n1075 ;
  assign n1914 = ~n1134 & n1642 ;
  assign n1160 = n1077 & ~n1133 ;
  assign n1152 = n1086 ^ n1079 ;
  assign n1153 = n1152 ^ n1113 ;
  assign n1154 = n1077 & n1153 ;
  assign n1155 = n1154 ^ n1113 ;
  assign n1161 = n1160 ^ n1155 ;
  assign n1162 = n1075 & n1161 ;
  assign n1163 = n1162 ^ n1155 ;
  assign n1915 = n1914 ^ n1163 ;
  assign n2091 = n2090 ^ n1915 ;
  assign n2092 = n2091 ^ x23 ;
  assign n2081 = n1102 ^ n1073 ;
  assign n2084 = n2081 ^ n1071 ;
  assign n1166 = n1101 ^ n1099 ;
  assign n1904 = n1166 ^ n1091 ;
  assign n2080 = n1904 ^ n1089 ;
  assign n2082 = n2081 ^ n2080 ;
  assign n2083 = n1075 & n2082 ;
  assign n2085 = n2084 ^ n2083 ;
  assign n2086 = ~n1077 & n2085 ;
  assign n2093 = n2092 ^ n2086 ;
  assign n2079 = n1079 & ~n1083 ;
  assign n2094 = n2093 ^ n2079 ;
  assign n1096 = n1070 & n1085 ;
  assign n1167 = n1166 ^ n1096 ;
  assign n2076 = n1075 & n1167 ;
  assign n2077 = n2076 ^ n1166 ;
  assign n2078 = n1077 & n2077 ;
  assign n2095 = n2094 ^ n2078 ;
  assign n2096 = n2095 ^ x68 ;
  assign n316 = n266 ^ n257 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = n289 & ~n317 ;
  assign n312 = n311 ^ n248 ;
  assign n313 = n276 & n312 ;
  assign n302 = n258 & n276 ;
  assign n303 = n302 ^ n257 ;
  assign n304 = n226 & n303 ;
  assign n308 = n307 ^ n304 ;
  assign n309 = n308 ^ n297 ;
  assign n310 = n309 ^ x7 ;
  assign n314 = n313 ^ n310 ;
  assign n319 = n318 ^ n314 ;
  assign n290 = n289 ^ n226 ;
  assign n291 = n287 & ~n290 ;
  assign n320 = n319 ^ n291 ;
  assign n274 = n273 ^ n265 ;
  assign n270 = n269 ^ n260 ;
  assign n271 = n270 ^ n265 ;
  assign n275 = n274 ^ n271 ;
  assign n279 = ~n275 & ~n276 ;
  assign n280 = n279 ^ n271 ;
  assign n281 = n226 & ~n280 ;
  assign n321 = n320 ^ n281 ;
  assign n2097 = n321 ^ x110 ;
  assign n2098 = n2096 & ~n2097 ;
  assign n2099 = n2098 ^ n2097 ;
  assign n2100 = n2099 ^ n2096 ;
  assign n2066 = n1431 ^ n1389 ;
  assign n2067 = n1421 & ~n2066 ;
  assign n2061 = n1378 ^ n1366 ;
  assign n2052 = n1363 & ~n1448 ;
  assign n1715 = n1407 & ~n1714 ;
  assign n2051 = n1715 ^ n1425 ;
  assign n2053 = n2052 ^ n2051 ;
  assign n2062 = n2061 ^ n2053 ;
  assign n2059 = n1388 ^ n1355 ;
  assign n2060 = ~n1358 & n2059 ;
  assign n2063 = n2062 ^ n2060 ;
  assign n2064 = n1714 & n2063 ;
  assign n2054 = n2053 ^ n1422 ;
  assign n2055 = n2054 ^ n1419 ;
  assign n2056 = n2055 ^ n1404 ;
  assign n2057 = n2056 ^ x15 ;
  assign n2041 = n1406 ^ n1366 ;
  assign n2058 = n2057 ^ n2041 ;
  assign n2065 = n2064 ^ n2058 ;
  assign n2068 = n2067 ^ n2065 ;
  assign n2050 = ~n1358 & n1366 ;
  assign n2069 = n2068 ^ n2050 ;
  assign n2043 = n2041 ^ n1424 ;
  assign n2042 = n2041 ^ n1432 ;
  assign n2044 = n2043 ^ n2042 ;
  assign n2047 = ~n1358 & n2044 ;
  assign n2048 = n2047 ^ n2043 ;
  assign n2049 = ~n1391 & n2048 ;
  assign n2070 = n2069 ^ n2049 ;
  assign n2071 = n2070 ^ x117 ;
  assign n854 = n853 ^ n633 ;
  assign n855 = n854 ^ n629 ;
  assign n856 = n855 ^ n602 ;
  assign n852 = n620 ^ n597 ;
  assign n857 = n856 ^ n852 ;
  assign n862 = n861 ^ n857 ;
  assign n863 = ~n583 & ~n862 ;
  assign n864 = n863 ^ n856 ;
  assign n894 = n893 ^ n864 ;
  assign n903 = n902 ^ n894 ;
  assign n881 = ~n583 & n616 ;
  assign n882 = n881 ^ n876 ;
  assign n883 = ~n584 & n882 ;
  assign n904 = n903 ^ n883 ;
  assign n905 = n904 ^ x31 ;
  assign n650 = n618 ^ n615 ;
  assign n1676 = n650 ^ n626 ;
  assign n872 = n583 & n1676 ;
  assign n865 = n626 ^ n612 ;
  assign n866 = n865 ^ n864 ;
  assign n873 = n872 ^ n866 ;
  assign n874 = ~n584 & ~n873 ;
  assign n906 = n905 ^ n874 ;
  assign n2072 = n906 ^ x69 ;
  assign n2073 = n2071 & n2072 ;
  assign n2108 = n2073 ^ n2072 ;
  assign n2109 = n2100 & n2108 ;
  assign n2105 = n2073 & n2098 ;
  assign n2103 = n2100 ^ n2097 ;
  assign n2104 = n2073 & n2103 ;
  assign n2106 = n2105 ^ n2104 ;
  assign n2101 = n2073 & n2100 ;
  assign n2102 = n2101 ^ n2073 ;
  assign n2107 = n2106 ^ n2102 ;
  assign n2110 = n2109 ^ n2107 ;
  assign n948 = n947 ^ n940 ;
  assign n934 = n433 ^ n398 ;
  assign n931 = n382 ^ n376 ;
  assign n932 = n931 ^ n398 ;
  assign n933 = n359 & n932 ;
  assign n935 = n934 ^ n933 ;
  assign n936 = n358 & n935 ;
  assign n937 = n936 ^ n361 ;
  assign n923 = n394 ^ n365 ;
  assign n924 = n923 ^ n361 ;
  assign n925 = n435 ^ n363 ;
  assign n928 = ~n923 & n925 ;
  assign n929 = n928 ^ n435 ;
  assign n930 = n924 & n929 ;
  assign n938 = n937 ^ n930 ;
  assign n939 = n938 ^ n387 ;
  assign n949 = n948 ^ n939 ;
  assign n920 = ~n359 & n380 ;
  assign n921 = n920 ^ n381 ;
  assign n922 = ~n358 & n921 ;
  assign n950 = n949 ^ n922 ;
  assign n425 = n424 ^ n422 ;
  assign n428 = ~n358 & ~n425 ;
  assign n429 = n428 ^ n422 ;
  assign n430 = n385 & ~n429 ;
  assign n951 = n950 ^ n430 ;
  assign n952 = n951 ^ x39 ;
  assign n908 = n378 ^ n356 ;
  assign n913 = n359 & n908 ;
  assign n914 = n913 ^ n387 ;
  assign n915 = ~n358 & n914 ;
  assign n953 = n952 ^ n915 ;
  assign n2040 = n953 ^ x100 ;
  assign n337 = n182 ^ n149 ;
  assign n338 = n337 ^ n203 ;
  assign n339 = n338 ^ n207 ;
  assign n340 = ~n129 & ~n339 ;
  assign n341 = n340 ^ n203 ;
  assign n342 = ~n130 & ~n341 ;
  assign n343 = n342 ^ x57 ;
  assign n131 = n130 ^ n129 ;
  assign n324 = n323 ^ n205 ;
  assign n325 = ~n129 & n324 ;
  assign n326 = n325 ^ n205 ;
  assign n328 = n326 ^ n159 ;
  assign n327 = n326 ^ n200 ;
  assign n329 = n328 ^ n327 ;
  assign n332 = ~n129 & n329 ;
  assign n333 = n332 ^ n328 ;
  assign n334 = n131 & n333 ;
  assign n335 = n334 ^ n326 ;
  assign n336 = ~n196 & ~n335 ;
  assign n344 = n343 ^ n336 ;
  assign n2112 = n344 ^ x86 ;
  assign n2158 = n2040 & n2112 ;
  assign n2159 = n2158 ^ n2040 ;
  assign n2160 = n2159 ^ n2112 ;
  assign n2161 = n2160 ^ n2040 ;
  assign n2658 = n2110 & n2161 ;
  assign n2123 = n2112 ^ n2040 ;
  assign n2114 = ~n2099 & n2108 ;
  assign n2650 = n2114 ^ n2104 ;
  assign n2125 = n2108 ^ n2071 ;
  assign n2132 = n2100 & ~n2125 ;
  assign n2126 = n2098 & ~n2125 ;
  assign n2133 = n2132 ^ n2126 ;
  assign n2130 = ~n2099 & ~n2125 ;
  assign n2131 = n2130 ^ n2125 ;
  assign n2134 = n2133 ^ n2131 ;
  assign n2152 = n2134 ^ n2072 ;
  assign n2127 = n2125 ^ n2072 ;
  assign n2141 = n2103 & n2127 ;
  assign n2140 = n2098 & n2127 ;
  assign n2142 = n2141 ^ n2140 ;
  assign n2128 = n2100 & n2127 ;
  assign n2129 = n2128 ^ n2126 ;
  assign n2138 = n2130 ^ n2129 ;
  assign n2139 = n2138 ^ n2132 ;
  assign n2143 = n2142 ^ n2139 ;
  assign n2153 = n2152 ^ n2143 ;
  assign n2651 = n2650 ^ n2153 ;
  assign n2648 = n2141 ^ n2128 ;
  assign n2649 = n2648 ^ n2130 ;
  assign n2652 = n2651 ^ n2649 ;
  assign n2653 = n2040 & n2652 ;
  assign n2654 = n2653 ^ n2651 ;
  assign n2655 = n2123 & n2654 ;
  assign n2643 = n2105 ^ n2101 ;
  assign n2164 = n2098 & n2108 ;
  assign n2639 = n2164 ^ n2128 ;
  assign n2640 = n2639 ^ n2141 ;
  assign n2641 = n2640 ^ n2132 ;
  assign n2642 = n2112 & ~n2641 ;
  assign n2644 = n2643 ^ n2642 ;
  assign n2645 = ~n2123 & n2644 ;
  assign n2166 = n2114 ^ n2109 ;
  assign n2165 = n2164 ^ n2108 ;
  assign n2167 = n2166 ^ n2165 ;
  assign n2620 = n2107 ^ n2104 ;
  assign n2621 = n2620 ^ n2123 ;
  assign n2624 = ~n2167 & ~n2621 ;
  assign n2625 = n2624 ^ n2123 ;
  assign n2631 = n2112 & n2142 ;
  assign n2632 = n2631 ^ n2141 ;
  assign n2633 = ~n2040 & n2632 ;
  assign n2635 = n2633 ^ n2040 ;
  assign n2626 = n2167 ^ n2158 ;
  assign n2634 = n2633 ^ n2626 ;
  assign n2636 = n2635 ^ n2634 ;
  assign n2637 = n2625 & n2636 ;
  assign n2638 = n2637 ^ n2635 ;
  assign n2646 = n2645 ^ n2638 ;
  assign n2617 = n2140 ^ n2133 ;
  assign n2618 = n2617 ^ n2114 ;
  assign n2619 = ~n2160 & n2618 ;
  assign n2647 = n2646 ^ n2619 ;
  assign n2656 = n2655 ^ n2647 ;
  assign n2174 = n2159 & n2164 ;
  assign n2657 = n2656 ^ n2174 ;
  assign n2659 = n2658 ^ n2657 ;
  assign n2177 = n2167 ^ n2132 ;
  assign n2180 = ~n2112 & n2177 ;
  assign n2181 = n2180 ^ n2132 ;
  assign n2182 = ~n2040 & n2181 ;
  assign n2660 = n2659 ^ n2182 ;
  assign n2149 = n2130 ^ n2072 ;
  assign n2150 = n2149 ^ n2143 ;
  assign n2151 = n2112 & ~n2150 ;
  assign n2154 = n2153 ^ n2151 ;
  assign n2155 = n2040 & n2154 ;
  assign n2661 = n2660 ^ n2155 ;
  assign n2662 = n2661 ^ x28 ;
  assign n2663 = n2662 ^ x110 ;
  assign n2669 = ~n2252 & n2663 ;
  assign n2697 = n2669 ^ n2663 ;
  assign n664 = n611 ^ n592 ;
  assign n665 = n664 ^ n591 ;
  assign n666 = n663 & ~n665 ;
  assign n651 = n650 ^ n606 ;
  assign n655 = n654 ^ n651 ;
  assign n656 = ~n598 & n655 ;
  assign n657 = n656 ^ n651 ;
  assign n658 = n583 & n657 ;
  assign n659 = n658 ^ n651 ;
  assign n660 = ~n584 & n659 ;
  assign n661 = n660 ^ x33 ;
  assign n647 = ~n582 & ~n631 ;
  assign n648 = n647 ^ n629 ;
  assign n649 = n583 & n648 ;
  assign n662 = n661 ^ n649 ;
  assign n667 = n666 ^ n662 ;
  assign n642 = ~n583 & ~n612 ;
  assign n668 = n667 ^ n642 ;
  assign n634 = n633 ^ n620 ;
  assign n635 = n634 ^ n628 ;
  assign n636 = n635 ^ n633 ;
  assign n639 = ~n583 & n636 ;
  assign n640 = n639 ^ n633 ;
  assign n641 = ~n584 & n640 ;
  assign n669 = n668 ^ n641 ;
  assign n1943 = n669 ^ x88 ;
  assign n1905 = n1904 ^ n1071 ;
  assign n1924 = n1905 ^ n1123 ;
  assign n1175 = n1077 & n1089 ;
  assign n1168 = n1167 ^ n1113 ;
  assign n1169 = n1077 & n1168 ;
  assign n1170 = n1169 ^ n1167 ;
  assign n1176 = n1175 ^ n1170 ;
  assign n1177 = ~n1075 & n1176 ;
  assign n1178 = n1177 ^ n1170 ;
  assign n1925 = n1924 ^ n1178 ;
  assign n1926 = n1925 ^ n1923 ;
  assign n1927 = n1926 ^ n1915 ;
  assign n1928 = n1927 ^ x17 ;
  assign n1906 = n1905 ^ n1090 ;
  assign n1907 = n1906 ^ n1073 ;
  assign n1908 = n1907 ^ n1905 ;
  assign n1911 = ~n1075 & n1908 ;
  assign n1912 = n1911 ^ n1905 ;
  assign n1913 = n1083 & n1912 ;
  assign n1929 = n1928 ^ n1913 ;
  assign n1105 = n1104 ^ n1096 ;
  assign n1903 = n1105 & ~n1641 ;
  assign n1930 = n1929 ^ n1903 ;
  assign n1897 = n1131 ^ n1123 ;
  assign n1898 = n1897 ^ n1104 ;
  assign n1899 = n1898 ^ n1123 ;
  assign n1900 = n1075 & n1899 ;
  assign n1901 = n1900 ^ n1123 ;
  assign n1902 = ~n1077 & n1901 ;
  assign n1931 = n1930 ^ n1902 ;
  assign n1932 = n1931 ^ x122 ;
  assign n1933 = n1537 ^ x74 ;
  assign n1934 = ~n1932 & n1933 ;
  assign n1890 = n311 ^ n254 ;
  assign n1891 = n289 & ~n1890 ;
  assign n1887 = n270 ^ x9 ;
  assign n1880 = n253 ^ n249 ;
  assign n1881 = n1880 ^ n267 ;
  assign n1879 = n237 & n288 ;
  assign n1882 = n1881 ^ n1879 ;
  assign n1883 = ~n1296 & ~n1882 ;
  assign n1884 = n1883 ^ n249 ;
  assign n1876 = n311 ^ n269 ;
  assign n1877 = n1876 ^ n265 ;
  assign n1878 = n305 & n1877 ;
  assign n1885 = n1884 ^ n1878 ;
  assign n1886 = ~n297 & ~n1885 ;
  assign n1888 = n1887 ^ n1886 ;
  assign n1875 = n264 & ~n1296 ;
  assign n1889 = n1888 ^ n1875 ;
  assign n1892 = n1891 ^ n1889 ;
  assign n1872 = ~n226 & n316 ;
  assign n1873 = n1872 ^ n270 ;
  assign n1874 = ~n276 & ~n1873 ;
  assign n1893 = n1892 ^ n1874 ;
  assign n1894 = n1893 ^ x64 ;
  assign n717 = x108 ^ x38 ;
  assign n713 = x118 ^ x6 ;
  assign n709 = x76 ^ x22 ;
  assign n707 = x125 ^ x14 ;
  assign n708 = x77 ^ x30 ;
  assign n712 = n707 & n708 ;
  assign n758 = n709 & n712 ;
  assign n710 = ~n708 & n709 ;
  assign n757 = n710 ^ n709 ;
  assign n759 = n758 ^ n757 ;
  assign n760 = ~n713 & n759 ;
  assign n731 = ~n709 & n713 ;
  assign n732 = n708 & n731 ;
  assign n733 = n732 ^ n731 ;
  assign n743 = ~n707 & n733 ;
  assign n744 = n743 ^ n733 ;
  assign n767 = n760 ^ n744 ;
  assign n761 = n760 ^ n758 ;
  assign n711 = n707 & n710 ;
  assign n745 = n711 ^ n710 ;
  assign n746 = ~n713 & n745 ;
  assign n747 = n746 ^ n744 ;
  assign n762 = n761 ^ n747 ;
  assign n751 = n711 ^ n707 ;
  assign n752 = n751 ^ n709 ;
  assign n753 = n752 ^ n711 ;
  assign n754 = ~n713 & n753 ;
  assign n755 = n754 ^ n751 ;
  assign n714 = n713 ^ n709 ;
  assign n715 = n712 & n714 ;
  assign n756 = n755 ^ n715 ;
  assign n763 = n762 ^ n756 ;
  assign n768 = n767 ^ n763 ;
  assign n730 = n710 ^ n708 ;
  assign n734 = n733 ^ n730 ;
  assign n735 = n707 & ~n734 ;
  assign n736 = n735 ^ n734 ;
  assign n769 = n768 ^ n736 ;
  assign n770 = n717 & ~n769 ;
  assign n764 = n732 ^ n715 ;
  assign n765 = n764 ^ n763 ;
  assign n766 = n765 ^ n760 ;
  assign n771 = n770 ^ n766 ;
  assign n728 = n711 & ~n713 ;
  assign n729 = n728 ^ n711 ;
  assign n739 = n735 ^ n729 ;
  assign n723 = n715 ^ n712 ;
  assign n740 = n739 ^ n723 ;
  assign n741 = n717 & n740 ;
  assign n742 = n741 ^ n723 ;
  assign n790 = n771 ^ n742 ;
  assign n706 = x94 ^ x56 ;
  assign n725 = n717 ^ n706 ;
  assign n781 = n761 ^ n757 ;
  assign n778 = n712 ^ n708 ;
  assign n779 = n778 ^ n759 ;
  assign n780 = n779 ^ n765 ;
  assign n782 = n781 ^ n780 ;
  assign n776 = n746 ^ n745 ;
  assign n777 = n776 ^ n736 ;
  assign n783 = n782 ^ n777 ;
  assign n786 = n717 & ~n783 ;
  assign n787 = n786 ^ n777 ;
  assign n788 = n725 & ~n787 ;
  assign n791 = n790 ^ n788 ;
  assign n792 = n791 ^ x25 ;
  assign n772 = n771 ^ n759 ;
  assign n748 = n747 ^ n729 ;
  assign n749 = n748 ^ n743 ;
  assign n750 = n749 ^ n742 ;
  assign n773 = n772 ^ n750 ;
  assign n737 = n736 ^ n729 ;
  assign n738 = n717 & ~n737 ;
  assign n774 = n773 ^ n738 ;
  assign n775 = ~n725 & n774 ;
  assign n793 = n792 ^ n775 ;
  assign n724 = n706 & n717 ;
  assign n726 = n725 ^ n724 ;
  assign n727 = n723 & ~n726 ;
  assign n794 = n793 ^ n727 ;
  assign n716 = n715 ^ n711 ;
  assign n720 = n716 & ~n717 ;
  assign n721 = n720 ^ n715 ;
  assign n722 = n706 & n721 ;
  assign n795 = n794 ^ n722 ;
  assign n1895 = n795 ^ x112 ;
  assign n1896 = n1894 & ~n1895 ;
  assign n1951 = n1896 ^ n1895 ;
  assign n1952 = n1951 ^ n1894 ;
  assign n1953 = n1934 & n1952 ;
  assign n1935 = n1934 ^ n1933 ;
  assign n1939 = n1935 ^ n1932 ;
  assign n1940 = n1896 & n1939 ;
  assign n1938 = n1896 & n1934 ;
  assign n1941 = n1940 ^ n1938 ;
  assign n1970 = n1953 ^ n1941 ;
  assign n2284 = ~n1943 & n1970 ;
  assign n1936 = n1896 & n1935 ;
  assign n1937 = n1936 ^ n1896 ;
  assign n1942 = n1941 ^ n1937 ;
  assign n1944 = n1464 ^ x97 ;
  assign n1945 = ~n1943 & ~n1944 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1947 = n1946 ^ n1944 ;
  assign n1997 = n1947 ^ n1943 ;
  assign n2274 = n1942 & ~n1997 ;
  assign n1949 = n1896 ^ n1894 ;
  assign n1967 = n1935 & n1949 ;
  assign n2018 = ~n1946 & n1967 ;
  assign n2275 = n2274 ^ n2018 ;
  assign n2007 = n1944 ^ n1943 ;
  assign n1950 = n1934 & n1949 ;
  assign n1985 = n1950 ^ n1949 ;
  assign n1955 = n1934 ^ n1932 ;
  assign n1957 = n1949 & ~n1955 ;
  assign n1968 = n1967 ^ n1957 ;
  assign n1986 = n1985 ^ n1968 ;
  assign n1961 = n1935 & n1952 ;
  assign n1959 = n1955 ^ n1942 ;
  assign n1956 = ~n1951 & ~n1955 ;
  assign n1958 = n1957 ^ n1956 ;
  assign n1960 = n1959 ^ n1958 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1954 = n1953 ^ n1952 ;
  assign n1963 = n1962 ^ n1954 ;
  assign n1987 = n1986 ^ n1963 ;
  assign n2271 = n1944 & ~n1987 ;
  assign n2272 = n2271 ^ n1963 ;
  assign n2273 = ~n2007 & ~n2272 ;
  assign n2276 = n2275 ^ n2273 ;
  assign n1984 = n1940 ^ n1939 ;
  assign n1988 = n1987 ^ n1984 ;
  assign n1972 = n1933 ^ n1932 ;
  assign n1973 = n1972 ^ n1895 ;
  assign n1974 = n1973 ^ n1894 ;
  assign n1969 = n1968 ^ n1956 ;
  assign n1971 = n1970 ^ n1969 ;
  assign n1975 = n1974 ^ n1971 ;
  assign n1976 = n1975 ^ n1963 ;
  assign n1989 = n1988 ^ n1976 ;
  assign n1983 = n1956 ^ n1951 ;
  assign n1990 = n1989 ^ n1983 ;
  assign n1991 = n1990 ^ n1942 ;
  assign n2261 = n1991 ^ n1989 ;
  assign n2264 = ~n1943 & ~n2261 ;
  assign n2265 = n2264 ^ n1989 ;
  assign n2266 = ~n1944 & ~n2265 ;
  assign n2277 = n2276 ^ n2266 ;
  assign n2021 = n1988 ^ n1961 ;
  assign n2024 = ~n1943 & ~n2021 ;
  assign n2025 = n2024 ^ n1961 ;
  assign n2026 = n1944 & n2025 ;
  assign n2278 = n2277 ^ n2026 ;
  assign n2031 = n1986 ^ n1962 ;
  assign n2034 = n1944 & ~n2031 ;
  assign n2035 = n2034 ^ n1962 ;
  assign n2036 = ~n1943 & ~n2035 ;
  assign n2279 = n2278 ^ n2036 ;
  assign n2280 = n2279 ^ x52 ;
  assign n2011 = n1990 ^ n1988 ;
  assign n2258 = n2011 ^ n1969 ;
  assign n2259 = n2258 ^ n1938 ;
  assign n2260 = ~n1947 & ~n2259 ;
  assign n2281 = n2280 ^ n2260 ;
  assign n1964 = n1963 ^ n1950 ;
  assign n2255 = n1964 ^ n1936 ;
  assign n2256 = n2255 ^ n1968 ;
  assign n2257 = ~n1997 & ~n2256 ;
  assign n2282 = n2281 ^ n2257 ;
  assign n2253 = n1990 ^ n1957 ;
  assign n2254 = ~n1946 & n2253 ;
  assign n2283 = n2282 ^ n2254 ;
  assign n2285 = n2284 ^ n2283 ;
  assign n2286 = n2285 ^ x78 ;
  assign n1148 = n1075 ^ n1074 ;
  assign n1149 = n1148 ^ n1147 ;
  assign n1150 = n1149 ^ n1141 ;
  assign n1151 = n1150 ^ n1093 ;
  assign n1164 = n1163 ^ n1151 ;
  assign n1165 = n1164 ^ n1121 ;
  assign n1179 = n1178 ^ n1165 ;
  assign n1180 = n1179 ^ x5 ;
  assign n1106 = n1105 ^ n1093 ;
  assign n1107 = n1106 ^ n1094 ;
  assign n1110 = n1077 & n1107 ;
  assign n1111 = n1110 ^ n1094 ;
  assign n1112 = n1083 & n1111 ;
  assign n1181 = n1180 ^ n1112 ;
  assign n1076 = ~n1074 & n1075 ;
  assign n1182 = n1181 ^ n1076 ;
  assign n1080 = n1079 ^ n1074 ;
  assign n1081 = ~n1077 & n1080 ;
  assign n1082 = n1076 & n1081 ;
  assign n1183 = n1182 ^ n1082 ;
  assign n2353 = n1183 ^ x78 ;
  assign n1797 = n760 ^ n748 ;
  assign n1798 = ~n726 & n1797 ;
  assign n1792 = n759 ^ n711 ;
  assign n1793 = n1792 ^ n747 ;
  assign n1794 = n1793 ^ n765 ;
  assign n1795 = ~n717 & n1794 ;
  assign n1790 = n763 ^ n732 ;
  assign n1791 = n1790 ^ n728 ;
  assign n1796 = n1795 ^ n1791 ;
  assign n1799 = n1798 ^ n1796 ;
  assign n1785 = n776 ^ n723 ;
  assign n1786 = n1785 ^ n715 ;
  assign n1787 = n717 & n1786 ;
  assign n1788 = n1787 ^ n715 ;
  assign n1789 = ~n706 & n1788 ;
  assign n1800 = n1799 ^ n1789 ;
  assign n1775 = n746 ^ n735 ;
  assign n1801 = n1800 ^ n1775 ;
  assign n1783 = n780 ^ n715 ;
  assign n1784 = ~n724 & n1783 ;
  assign n1802 = n1801 ^ n1784 ;
  assign n1776 = n1775 ^ n726 ;
  assign n1777 = n733 ^ n724 ;
  assign n1780 = ~n1775 & ~n1777 ;
  assign n1781 = n1780 ^ n724 ;
  assign n1782 = ~n1776 & ~n1781 ;
  assign n1803 = n1802 ^ n1782 ;
  assign n1030 = n724 & ~n777 ;
  assign n1804 = n1803 ^ n1030 ;
  assign n1805 = n1804 ^ x29 ;
  assign n1774 = n725 & n742 ;
  assign n1806 = n1805 ^ n1774 ;
  assign n2288 = n1806 ^ x85 ;
  assign n2341 = n1378 & ~n1714 ;
  assign n2336 = n1436 ^ n1371 ;
  assign n2330 = n1377 ^ n1352 ;
  assign n2331 = n2330 ^ n1424 ;
  assign n2332 = n1358 & n2331 ;
  assign n2337 = n2336 ^ n2332 ;
  assign n2334 = n1383 ^ n1381 ;
  assign n2335 = ~n1358 & n2334 ;
  assign n2338 = n2337 ^ n2335 ;
  assign n2339 = n1391 & n2338 ;
  assign n2329 = n1455 ^ n1425 ;
  assign n2333 = n2332 ^ n2329 ;
  assign n2340 = n2339 ^ n2333 ;
  assign n2342 = n2341 ^ n2340 ;
  assign n2326 = ~n1358 & n1427 ;
  assign n2327 = n2326 ^ n1425 ;
  assign n2328 = ~n1391 & n2327 ;
  assign n2343 = n2342 ^ n2328 ;
  assign n2344 = n2343 ^ n1422 ;
  assign n2345 = n2344 ^ n1404 ;
  assign n2346 = n2345 ^ n1396 ;
  assign n2347 = n2346 ^ x13 ;
  assign n2348 = n2347 ^ x108 ;
  assign n2367 = n2288 & n2348 ;
  assign n2376 = n2367 ^ n2348 ;
  assign n2315 = n1303 ^ n269 ;
  assign n2316 = n289 & ~n2315 ;
  assign n2308 = n311 ^ n260 ;
  assign n2309 = n2308 ^ n264 ;
  assign n2300 = n267 ^ n244 ;
  assign n2301 = n2300 ^ n238 ;
  assign n2302 = n226 & ~n2301 ;
  assign n2310 = n2309 ^ n2302 ;
  assign n2311 = n2310 ^ n262 ;
  assign n2306 = n267 ^ n262 ;
  assign n2307 = ~n226 & ~n2306 ;
  assign n2312 = n2311 ^ n2307 ;
  assign n2313 = ~n1296 & ~n2312 ;
  assign n2303 = n2302 ^ n307 ;
  assign n2304 = n2303 ^ n304 ;
  assign n2305 = n2304 ^ x21 ;
  assign n2314 = n2313 ^ n2305 ;
  assign n2317 = n2316 ^ n2314 ;
  assign n2298 = n252 ^ n238 ;
  assign n2299 = ~n290 & n2298 ;
  assign n2318 = n2317 ^ n2299 ;
  assign n2292 = n311 ^ n247 ;
  assign n2295 = ~n276 & n2292 ;
  assign n2296 = n2295 ^ n247 ;
  assign n2297 = n226 & n2296 ;
  assign n2319 = n2318 ^ n2297 ;
  assign n2290 = n254 ^ n245 ;
  assign n2291 = n276 & ~n2290 ;
  assign n2320 = n2319 ^ n2291 ;
  assign n2289 = n245 & n288 ;
  assign n2321 = n2320 ^ n2289 ;
  assign n2322 = n2321 ^ x91 ;
  assign n2349 = ~n2322 & n2348 ;
  assign n2350 = n2288 & n2349 ;
  assign n2373 = n2350 ^ n2349 ;
  assign n2377 = n2376 ^ n2373 ;
  assign n2351 = ~n2288 & n2322 ;
  assign n2378 = n2377 ^ n2351 ;
  assign n2379 = ~n2353 & n2378 ;
  assign n2382 = n2379 ^ n2351 ;
  assign n2383 = n2382 ^ n2377 ;
  assign n2354 = ~n2348 & ~n2353 ;
  assign n2355 = ~n2288 & n2354 ;
  assign n2380 = n2379 ^ n2355 ;
  assign n2374 = n2373 ^ n2351 ;
  assign n2375 = n2374 ^ n2288 ;
  assign n2381 = n2380 ^ n2375 ;
  assign n2384 = n2383 ^ n2381 ;
  assign n177 = n154 ^ n136 ;
  assign n178 = n160 & ~n177 ;
  assign n180 = n179 ^ n178 ;
  assign n181 = ~n129 & n180 ;
  assign n221 = n219 ^ n181 ;
  assign n222 = n221 ^ n213 ;
  assign n223 = n222 ^ x37 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n183 ^ n129 ;
  assign n185 = n184 ^ n183 ;
  assign n150 = n149 ^ n140 ;
  assign n153 = n152 ^ n150 ;
  assign n187 = n186 ^ n153 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = n189 ^ n183 ;
  assign n191 = n190 ^ n183 ;
  assign n192 = n185 & n191 ;
  assign n193 = n192 ^ n183 ;
  assign n194 = n130 & n193 ;
  assign n224 = n223 ^ n194 ;
  assign n170 = n165 ^ n156 ;
  assign n157 = n156 ^ n153 ;
  assign n169 = n168 ^ n157 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = n170 ^ n129 ;
  assign n173 = n172 ^ n170 ;
  assign n174 = ~n171 & n173 ;
  assign n175 = n174 ^ n170 ;
  assign n176 = n131 & n175 ;
  assign n225 = n224 ^ n176 ;
  assign n2287 = n225 ^ x102 ;
  assign n993 = n512 ^ n487 ;
  assign n994 = n993 ^ n504 ;
  assign n998 = n997 ^ n994 ;
  assign n999 = n474 & ~n998 ;
  assign n1000 = n999 ^ n504 ;
  assign n1001 = ~n473 & n1000 ;
  assign n988 = n506 ^ n488 ;
  assign n989 = n988 ^ n532 ;
  assign n990 = n552 & n989 ;
  assign n976 = n514 ^ n510 ;
  assign n977 = n976 ^ n972 ;
  assign n978 = ~n550 & n977 ;
  assign n979 = n978 ^ n551 ;
  assign n984 = ~n550 & n972 ;
  assign n981 = n510 ^ n502 ;
  assign n982 = n981 ^ n548 ;
  assign n980 = n575 ^ n506 ;
  assign n983 = n982 ^ n980 ;
  assign n985 = n984 ^ n983 ;
  assign n986 = n979 & n985 ;
  assign n553 = n548 & n552 ;
  assign n567 = n566 ^ n553 ;
  assign n971 = n567 ^ x63 ;
  assign n975 = n974 ^ n971 ;
  assign n987 = n986 ^ n975 ;
  assign n991 = n990 ^ n987 ;
  assign n970 = n503 & ~n554 ;
  assign n992 = n991 ^ n970 ;
  assign n1002 = n1001 ^ n992 ;
  assign n2396 = n1002 ^ x84 ;
  assign n2417 = ~n2287 & n2396 ;
  assign n2418 = n2417 ^ n2287 ;
  assign n2419 = n2418 ^ n2396 ;
  assign n2427 = n2419 ^ n2287 ;
  assign n2450 = ~n2384 & n2427 ;
  assign n2451 = n2450 ^ x44 ;
  assign n2360 = n2353 ^ n2348 ;
  assign n2361 = n2348 ^ n2322 ;
  assign n2362 = n2360 & n2361 ;
  assign n2363 = n2362 ^ n2348 ;
  assign n2364 = n2288 & n2363 ;
  assign n2356 = n2355 ^ n2354 ;
  assign n2357 = ~n2322 & n2356 ;
  assign n2358 = n2357 ^ n2356 ;
  assign n2352 = n2351 ^ n2322 ;
  assign n2359 = n2358 ^ n2352 ;
  assign n2365 = n2364 ^ n2359 ;
  assign n2366 = n2365 ^ n2350 ;
  assign n2401 = n2366 & ~n2396 ;
  assign n2385 = n2288 & n2353 ;
  assign n2386 = n2385 ^ n2353 ;
  assign n2387 = n2386 ^ n2376 ;
  assign n2388 = n2387 ^ n2384 ;
  assign n2389 = n2388 ^ n2379 ;
  assign n2390 = n2389 ^ n2351 ;
  assign n2391 = n2390 ^ n2362 ;
  assign n2368 = n2367 ^ n2288 ;
  assign n2369 = n2368 ^ n2356 ;
  assign n2370 = ~n2322 & n2369 ;
  assign n2371 = n2370 ^ n2369 ;
  assign n2372 = n2371 ^ n2366 ;
  assign n2392 = n2391 ^ n2372 ;
  assign n2393 = n2392 ^ n2377 ;
  assign n2394 = n2393 ^ n2388 ;
  assign n2395 = n2394 ^ n2373 ;
  assign n2402 = n2401 ^ n2395 ;
  assign n2403 = n2287 & n2402 ;
  assign n2404 = n2403 ^ n2395 ;
  assign n2447 = ~n2393 & n2427 ;
  assign n2411 = n2396 ^ n2287 ;
  assign n2413 = n2385 ^ n2369 ;
  assign n2414 = n2413 ^ n2365 ;
  assign n2441 = ~n2411 & n2414 ;
  assign n2422 = n2394 ^ n2357 ;
  assign n2421 = n2387 ^ n2366 ;
  assign n2423 = n2422 ^ n2421 ;
  assign n2424 = n2396 & n2423 ;
  assign n2425 = n2424 ^ n2387 ;
  assign n2442 = n2441 ^ n2425 ;
  assign n2415 = n2414 ^ n2358 ;
  assign n2416 = n2415 ^ n2371 ;
  assign n2432 = n2416 ^ n2352 ;
  assign n2433 = n2432 ^ n2372 ;
  assign n2434 = n2433 ^ n2425 ;
  assign n2426 = n2370 ^ n2357 ;
  assign n2428 = ~n2358 & ~n2427 ;
  assign n2429 = ~n2365 & n2428 ;
  assign n2430 = ~n2426 & n2429 ;
  assign n2431 = n2430 ^ n2425 ;
  assign n2435 = n2434 ^ n2431 ;
  assign n2438 = n2396 & ~n2435 ;
  assign n2439 = n2438 ^ n2434 ;
  assign n2440 = ~n2287 & n2439 ;
  assign n2443 = n2442 ^ n2440 ;
  assign n2420 = n2416 & n2419 ;
  assign n2444 = n2443 ^ n2420 ;
  assign n2412 = n2379 & ~n2411 ;
  assign n2445 = n2444 ^ n2412 ;
  assign n2405 = n2382 ^ n2375 ;
  assign n2408 = ~n2396 & ~n2405 ;
  assign n2409 = n2408 ^ n2382 ;
  assign n2410 = ~n2287 & n2409 ;
  assign n2446 = n2445 ^ n2410 ;
  assign n2448 = n2447 ^ n2446 ;
  assign n2449 = ~n2404 & ~n2448 ;
  assign n2452 = n2451 ^ n2449 ;
  assign n2453 = n2452 ^ x93 ;
  assign n2454 = ~n2286 & ~n2453 ;
  assign n2601 = n2454 ^ n2286 ;
  assign n2604 = n2601 ^ n2453 ;
  assign n2605 = n2604 ^ n2286 ;
  assign n322 = n321 ^ x65 ;
  assign n796 = n795 ^ x72 ;
  assign n830 = n322 & n796 ;
  assign n833 = n830 ^ n796 ;
  assign n834 = n833 ^ n322 ;
  assign n345 = n344 ^ x106 ;
  assign n395 = n394 ^ n390 ;
  assign n399 = n398 ^ n383 ;
  assign n400 = n399 ^ n387 ;
  assign n396 = n390 ^ n382 ;
  assign n397 = n396 ^ n394 ;
  assign n401 = n400 ^ n397 ;
  assign n402 = n401 ^ n359 ;
  assign n403 = n402 ^ n397 ;
  assign n404 = ~n385 & n403 ;
  assign n405 = n404 ^ n385 ;
  assign n406 = n395 & ~n405 ;
  assign n407 = n406 ^ n397 ;
  assign n408 = n403 ^ n358 ;
  assign n409 = n408 ^ n404 ;
  assign n410 = ~n407 & n409 ;
  assign n411 = n410 ^ n397 ;
  assign n458 = n411 ^ n358 ;
  assign n452 = n421 ^ n374 ;
  assign n455 = n358 & ~n452 ;
  assign n456 = n455 ^ n421 ;
  assign n457 = ~n359 & ~n456 ;
  assign n459 = n458 ^ n457 ;
  assign n460 = n459 ^ n451 ;
  assign n443 = n360 & ~n394 ;
  assign n445 = n444 ^ n443 ;
  assign n461 = n460 ^ n445 ;
  assign n462 = n461 ^ n442 ;
  assign n463 = n462 ^ n430 ;
  assign n412 = n411 ^ n381 ;
  assign n413 = n412 ^ n389 ;
  assign n414 = n413 ^ n411 ;
  assign n417 = ~n359 & ~n414 ;
  assign n418 = n417 ^ n411 ;
  assign n419 = n385 & ~n418 ;
  assign n464 = n463 ^ n419 ;
  assign n384 = n360 & n383 ;
  assign n465 = n464 ^ n384 ;
  assign n364 = n363 ^ n357 ;
  assign n366 = n365 ^ n361 ;
  assign n369 = ~n357 & n366 ;
  assign n370 = n369 ^ n361 ;
  assign n371 = n364 & ~n370 ;
  assign n466 = n465 ^ n371 ;
  assign n468 = n467 ^ n466 ;
  assign n469 = n468 ^ x49 ;
  assign n470 = n469 ^ x89 ;
  assign n471 = n345 & n470 ;
  assign n472 = n471 ^ n345 ;
  assign n579 = n532 & ~n550 ;
  assign n576 = n575 ^ n504 ;
  assign n577 = ~n554 & n576 ;
  assign n526 = n525 ^ n523 ;
  assign n522 = n521 ^ n503 ;
  assign n527 = n526 ^ n522 ;
  assign n528 = ~n474 & ~n527 ;
  assign n529 = n528 ^ n526 ;
  assign n568 = n567 ^ n529 ;
  assign n569 = n568 ^ n547 ;
  assign n539 = ~n474 & n534 ;
  assign n540 = n539 ^ n506 ;
  assign n541 = n473 & n540 ;
  assign n570 = n569 ^ n541 ;
  assign n513 = n512 ^ n511 ;
  assign n516 = n515 ^ n513 ;
  assign n519 = n518 ^ n516 ;
  assign n520 = n474 & n519 ;
  assign n530 = n529 ^ n520 ;
  assign n531 = ~n473 & ~n530 ;
  assign n571 = n570 ^ n531 ;
  assign n573 = n572 ^ n571 ;
  assign n574 = n573 ^ x41 ;
  assign n578 = n577 ^ n574 ;
  assign n580 = n579 ^ n578 ;
  assign n581 = n580 ^ x115 ;
  assign n670 = n669 ^ x104 ;
  assign n671 = ~n581 & ~n670 ;
  assign n672 = n671 ^ n670 ;
  assign n673 = n672 ^ n581 ;
  assign n680 = n673 ^ n670 ;
  assign n804 = n472 & ~n680 ;
  assign n675 = n472 ^ n470 ;
  assign n676 = n675 ^ n345 ;
  assign n688 = n676 & ~n680 ;
  assign n846 = n804 ^ n688 ;
  assign n847 = ~n834 & n846 ;
  assign n677 = ~n673 & n676 ;
  assign n690 = n677 ^ n676 ;
  assign n687 = n671 & n676 ;
  assign n689 = n688 ^ n687 ;
  assign n691 = n690 ^ n689 ;
  assign n684 = n472 & ~n672 ;
  assign n683 = n471 & ~n672 ;
  assign n685 = n684 ^ n683 ;
  assign n686 = n685 ^ n672 ;
  assign n692 = n691 ^ n686 ;
  assign n843 = ~n692 & n833 ;
  assign n837 = n796 ^ n322 ;
  assign n693 = n671 & ~n675 ;
  assign n694 = n693 ^ n692 ;
  assign n681 = ~n675 & ~n680 ;
  assign n682 = n681 ^ n675 ;
  assign n695 = n694 ^ n682 ;
  assign n838 = n695 ^ n691 ;
  assign n839 = n838 ^ n688 ;
  assign n840 = ~n796 & n839 ;
  assign n841 = n840 ^ n688 ;
  assign n842 = n837 & n841 ;
  assign n844 = n843 ^ n842 ;
  assign n835 = n691 & ~n834 ;
  assign n699 = n693 ^ n687 ;
  assign n697 = n472 & n671 ;
  assign n698 = n697 ^ n671 ;
  assign n700 = n699 ^ n698 ;
  assign n674 = n472 & ~n673 ;
  assign n678 = n677 ^ n674 ;
  assign n679 = n678 ^ n673 ;
  assign n696 = n695 ^ n679 ;
  assign n701 = n700 ^ n696 ;
  assign n831 = n830 ^ n322 ;
  assign n832 = ~n701 & n831 ;
  assign n836 = n835 ^ n832 ;
  assign n845 = n844 ^ n836 ;
  assign n848 = n847 ^ n845 ;
  assign n849 = n848 ^ x60 ;
  assign n702 = n683 ^ n471 ;
  assign n703 = n702 ^ n701 ;
  assign n704 = n703 ^ n697 ;
  assign n705 = n704 ^ n688 ;
  assign n799 = ~n705 & ~n796 ;
  assign n800 = n799 ^ n688 ;
  assign n801 = n322 & n800 ;
  assign n821 = n687 ^ n678 ;
  assign n822 = n796 & n821 ;
  assign n823 = n822 ^ n687 ;
  assign n816 = n699 ^ n685 ;
  assign n817 = n796 & n816 ;
  assign n809 = n703 ^ n674 ;
  assign n810 = n796 & ~n809 ;
  assign n811 = n810 ^ n674 ;
  assign n802 = n693 ^ n681 ;
  assign n808 = n802 ^ n696 ;
  assign n812 = n811 ^ n808 ;
  assign n805 = n804 ^ n683 ;
  assign n803 = n802 ^ n700 ;
  assign n806 = n805 ^ n803 ;
  assign n807 = n796 & n806 ;
  assign n813 = n812 ^ n807 ;
  assign n814 = n813 ^ n685 ;
  assign n815 = n814 ^ n811 ;
  assign n818 = n817 ^ n815 ;
  assign n824 = n818 ^ n814 ;
  assign n825 = ~n823 & ~n824 ;
  assign n826 = n825 ^ n818 ;
  assign n827 = n322 & n826 ;
  assign n828 = n827 ^ n818 ;
  assign n829 = ~n801 & n828 ;
  assign n850 = n849 ^ n829 ;
  assign n2455 = n850 ^ x67 ;
  assign n1730 = n1410 ^ n1357 ;
  assign n1726 = n1386 ^ n1357 ;
  assign n1727 = n1726 ^ n1398 ;
  assign n1728 = n1727 ^ n1431 ;
  assign n1729 = n1358 & n1728 ;
  assign n1731 = n1730 ^ n1729 ;
  assign n1732 = ~n1391 & n1731 ;
  assign n1717 = n1371 & n1448 ;
  assign n1716 = n1376 ^ n1370 ;
  assign n1718 = n1717 ^ n1716 ;
  assign n1719 = n1718 ^ n1420 ;
  assign n1722 = n1376 & ~n1448 ;
  assign n1720 = n1450 ^ n1398 ;
  assign n1721 = n1720 ^ n1718 ;
  assign n1723 = n1722 ^ n1721 ;
  assign n1724 = n1719 & ~n1723 ;
  assign n1725 = n1724 ^ n1420 ;
  assign n1733 = n1732 ^ n1725 ;
  assign n1734 = n1733 ^ n1715 ;
  assign n1735 = n1734 ^ n1419 ;
  assign n1736 = n1735 ^ n1396 ;
  assign n1737 = n1736 ^ x61 ;
  assign n1711 = n1432 ^ n1411 ;
  assign n1712 = n1711 ^ n1362 ;
  assign n1713 = n1421 & n1712 ;
  assign n1738 = n1737 ^ n1713 ;
  assign n2456 = n1738 ^ x96 ;
  assign n2495 = n1317 ^ x114 ;
  assign n2496 = n1280 ^ x121 ;
  assign n2521 = n1511 ^ n523 ;
  assign n2522 = n551 & ~n2521 ;
  assign n2519 = n1530 ^ n541 ;
  assign n2506 = n556 ^ n479 ;
  assign n2507 = n2506 ^ n484 ;
  assign n2497 = n982 ^ n514 ;
  assign n2508 = n2507 ^ n2497 ;
  assign n2509 = n549 & ~n2508 ;
  assign n2510 = n2509 ^ n550 ;
  assign n2511 = n995 ^ n504 ;
  assign n2512 = n2511 ^ n500 ;
  assign n2513 = n2512 ^ n504 ;
  assign n2516 = ~n549 & ~n2513 ;
  assign n2517 = n2516 ^ n504 ;
  assign n2518 = ~n2510 & ~n2517 ;
  assign n2520 = n2519 ^ n2518 ;
  assign n2523 = n2522 ^ n2520 ;
  assign n2505 = ~n550 & n988 ;
  assign n2524 = n2523 ^ n2505 ;
  assign n2502 = n474 & n2497 ;
  assign n2503 = n2502 ^ n512 ;
  assign n2504 = ~n554 & n2503 ;
  assign n2525 = n2524 ^ n2504 ;
  assign n2526 = n2525 ^ n572 ;
  assign n2527 = n2526 ^ x19 ;
  assign n2528 = n2527 ^ x120 ;
  assign n2481 = n1030 ^ n780 ;
  assign n2467 = n709 ^ n708 ;
  assign n2468 = n2467 ^ n707 ;
  assign n2469 = n2468 ^ n732 ;
  assign n1021 = n743 ^ n728 ;
  assign n2457 = n1021 ^ n745 ;
  assign n2470 = n2469 ^ n2457 ;
  assign n2471 = n717 & ~n2470 ;
  assign n2472 = n2471 ^ n2457 ;
  assign n2482 = n2481 ^ n2472 ;
  assign n2483 = n2482 ^ x11 ;
  assign n2474 = n744 ^ n735 ;
  assign n2475 = n2474 ^ n2472 ;
  assign n2473 = n2472 ^ n781 ;
  assign n2476 = n2475 ^ n2473 ;
  assign n1017 = n763 ^ n712 ;
  assign n2477 = n2476 ^ n1017 ;
  assign n2478 = ~n717 & n2477 ;
  assign n2479 = n2478 ^ n2475 ;
  assign n2480 = n706 & n2479 ;
  assign n2484 = n2483 ^ n2480 ;
  assign n2466 = n724 & n761 ;
  assign n2485 = n2484 ^ n2466 ;
  assign n2465 = ~n726 & n1017 ;
  assign n2486 = n2485 ^ n2465 ;
  assign n2462 = ~n717 & n2457 ;
  assign n2463 = n2462 ^ n780 ;
  assign n2464 = n725 & n2463 ;
  assign n2487 = n2486 ^ n2464 ;
  assign n2488 = n2487 ^ x82 ;
  assign n1652 = n1100 & n1640 ;
  assign n1643 = n1091 ^ n1089 ;
  assign n1644 = n1643 ^ n1064 ;
  assign n1625 = n1135 ^ n1104 ;
  assign n1645 = n1644 ^ n1625 ;
  assign n1646 = n1642 & ~n1645 ;
  assign n1634 = n1072 ^ n1071 ;
  assign n1635 = n1634 ^ n1129 ;
  assign n1636 = ~n1077 & ~n1635 ;
  assign n1631 = n1625 ^ n1113 ;
  assign n1624 = n1129 ^ n1096 ;
  assign n1626 = n1625 ^ n1624 ;
  assign n1627 = n1624 ^ n1075 ;
  assign n1628 = n1083 & n1627 ;
  assign n1629 = n1628 ^ n1075 ;
  assign n1630 = n1626 & ~n1629 ;
  assign n1632 = n1631 ^ n1630 ;
  assign n1633 = n1632 ^ n1089 ;
  assign n1637 = n1636 ^ n1633 ;
  assign n1638 = ~n1083 & n1637 ;
  assign n1639 = n1638 ^ n1636 ;
  assign n1647 = n1646 ^ n1639 ;
  assign n1622 = n1123 ^ n1102 ;
  assign n1623 = ~n1083 & n1622 ;
  assign n1648 = n1647 ^ n1623 ;
  assign n1649 = n1648 ^ n1079 ;
  assign n1650 = n1649 ^ x3 ;
  assign n1618 = n1127 ^ n1080 ;
  assign n1619 = n1077 & n1618 ;
  assign n1620 = n1619 ^ n1127 ;
  assign n1621 = ~n1075 & n1620 ;
  assign n1651 = n1650 ^ n1621 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n2489 = n1653 ^ x73 ;
  assign n2490 = ~n2488 & n2489 ;
  assign n2491 = n2490 ^ n2488 ;
  assign n2492 = n2491 ^ n2489 ;
  assign n2569 = n2492 ^ n2488 ;
  assign n2538 = ~n2528 & n2569 ;
  assign n2539 = n2538 ^ n2491 ;
  assign n2540 = ~n2496 & ~n2539 ;
  assign n2541 = n2540 ^ n2491 ;
  assign n2542 = n2495 & ~n2541 ;
  assign n2543 = n2456 & n2542 ;
  assign n2544 = n2543 ^ n2542 ;
  assign n2493 = n2456 & n2492 ;
  assign n2494 = n2493 ^ n2492 ;
  assign n2530 = n2496 & n2528 ;
  assign n2529 = n2528 ^ n2496 ;
  assign n2531 = n2530 ^ n2529 ;
  assign n2532 = ~n2495 & ~n2531 ;
  assign n2533 = n2494 & n2532 ;
  assign n2545 = n2544 ^ n2533 ;
  assign n2570 = n2569 ^ n2491 ;
  assign n2567 = n2530 ^ n2496 ;
  assign n2549 = n2492 & ~n2496 ;
  assign n2550 = n2549 ^ n2492 ;
  assign n2568 = n2567 ^ n2550 ;
  assign n2571 = n2570 ^ n2568 ;
  assign n2585 = n2571 ^ n2456 ;
  assign n2572 = n2492 & n2530 ;
  assign n2579 = n2572 ^ n2530 ;
  assign n2573 = ~n2490 & ~n2530 ;
  assign n2574 = n2573 ^ n2529 ;
  assign n2575 = ~n2549 & ~n2574 ;
  assign n2576 = n2575 ^ n2574 ;
  assign n2577 = n2576 ^ n2572 ;
  assign n2578 = n2577 ^ n2550 ;
  assign n2580 = n2579 ^ n2578 ;
  assign n2552 = ~n2491 & ~n2496 ;
  assign n2555 = n2528 ^ n2488 ;
  assign n2556 = n2552 & ~n2555 ;
  assign n2581 = n2580 ^ n2556 ;
  assign n2582 = n2581 ^ n2571 ;
  assign n2583 = ~n2456 & n2582 ;
  assign n2584 = n2583 ^ n2581 ;
  assign n2586 = n2585 ^ n2584 ;
  assign n2587 = n2586 ^ n2581 ;
  assign n2559 = ~n2489 & n2530 ;
  assign n2553 = n2552 ^ n2531 ;
  assign n2554 = n2553 ^ n2540 ;
  assign n2557 = n2556 ^ n2554 ;
  assign n2547 = n2490 & ~n2496 ;
  assign n2546 = n2496 ^ n2488 ;
  assign n2548 = n2547 ^ n2546 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2558 = n2557 ^ n2551 ;
  assign n2560 = n2559 ^ n2558 ;
  assign n2588 = n2587 ^ n2560 ;
  assign n2562 = n2489 & n2529 ;
  assign n2563 = n2562 ^ n2551 ;
  assign n2564 = n2563 ^ n2556 ;
  assign n2561 = n2560 ^ n2550 ;
  assign n2565 = n2564 ^ n2561 ;
  assign n2566 = ~n2456 & ~n2565 ;
  assign n2589 = n2588 ^ n2566 ;
  assign n2590 = ~n2495 & ~n2589 ;
  assign n2591 = n2590 ^ n2587 ;
  assign n2592 = ~n2545 & n2591 ;
  assign n2593 = n2592 ^ x36 ;
  assign n2594 = n2593 ^ x76 ;
  assign n2595 = n2455 & n2594 ;
  assign n2607 = n2595 ^ n2455 ;
  assign n2608 = ~n2605 & n2607 ;
  assign n2606 = n2595 & ~n2605 ;
  assign n2609 = n2608 ^ n2606 ;
  assign n2743 = n2609 ^ n2605 ;
  assign n2744 = n2697 & ~n2743 ;
  assign n2670 = n2669 ^ n2252 ;
  assign n2698 = n2697 ^ n2670 ;
  assign n2672 = n2607 ^ n2594 ;
  assign n2673 = ~n2604 & ~n2672 ;
  assign n2596 = n2595 ^ n2594 ;
  assign n2602 = n2596 & ~n2601 ;
  assign n2598 = n2453 ^ n2286 ;
  assign n2599 = n2455 ^ n2286 ;
  assign n2600 = n2598 & ~n2599 ;
  assign n2603 = n2602 ^ n2600 ;
  assign n2610 = n2609 ^ n2603 ;
  assign n2597 = n2454 & n2596 ;
  assign n2611 = n2610 ^ n2597 ;
  assign n2688 = n2673 ^ n2611 ;
  assign n2686 = n2453 & ~n2455 ;
  assign n2687 = n2686 ^ n2596 ;
  assign n2689 = n2688 ^ n2687 ;
  assign n2690 = n2689 ^ n2602 ;
  assign n2691 = n2690 ^ n2597 ;
  assign n2692 = n2691 ^ n2596 ;
  assign n2683 = ~n2601 & n2607 ;
  assign n2684 = n2683 ^ n2606 ;
  assign n2677 = n2672 ^ n2602 ;
  assign n2612 = n2594 ^ n2286 ;
  assign n2613 = ~n2455 & n2612 ;
  assign n2614 = n2613 ^ n2611 ;
  assign n2678 = n2677 ^ n2614 ;
  assign n2676 = n2454 & n2595 ;
  assign n2679 = n2678 ^ n2676 ;
  assign n2675 = n2597 ^ n2454 ;
  assign n2680 = n2679 ^ n2675 ;
  assign n2681 = n2680 ^ n2609 ;
  assign n2682 = n2681 ^ n2607 ;
  assign n2685 = n2684 ^ n2682 ;
  assign n2693 = n2692 ^ n2685 ;
  assign n2674 = n2673 ^ n2604 ;
  assign n2694 = n2693 ^ n2674 ;
  assign n2738 = n2694 ^ n2681 ;
  assign n2721 = n2670 & ~n2694 ;
  assign n2725 = n2609 & ~n2721 ;
  assign n2722 = n2683 ^ n2676 ;
  assign n2723 = n2722 ^ n2721 ;
  assign n2724 = n2697 & ~n2723 ;
  assign n2726 = n2725 ^ n2724 ;
  assign n2717 = n2676 ^ n2595 ;
  assign n2716 = n2694 ^ n2606 ;
  assign n2718 = n2717 ^ n2716 ;
  assign n2727 = n2726 ^ n2718 ;
  assign n2739 = n2738 ^ n2727 ;
  assign n2699 = n2689 ^ n2678 ;
  assign n2734 = n2699 ^ n2611 ;
  assign n2735 = n2734 ^ n2681 ;
  assign n2736 = n2735 ^ n2694 ;
  assign n2737 = ~n2663 & n2736 ;
  assign n2740 = n2739 ^ n2737 ;
  assign n2741 = n2698 & ~n2740 ;
  assign n2728 = ~n2670 & ~n2680 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2671 = n2670 ^ n2663 ;
  assign n2719 = n2718 ^ n2680 ;
  assign n2720 = n2671 & ~n2719 ;
  assign n2730 = n2729 ^ n2720 ;
  assign n2711 = n2692 ^ n2252 ;
  assign n2712 = n2711 ^ n2692 ;
  assign n2713 = ~n2693 & n2712 ;
  assign n2714 = n2713 ^ n2692 ;
  assign n2715 = ~n2698 & n2714 ;
  assign n2731 = n2730 ^ n2715 ;
  assign n2701 = n2678 ^ n2605 ;
  assign n2700 = n2699 ^ n2609 ;
  assign n2702 = n2701 ^ n2700 ;
  assign n2703 = n2702 ^ n2692 ;
  assign n2704 = n2702 ^ n2663 ;
  assign n2705 = n2704 ^ n2702 ;
  assign n2706 = ~n2703 & n2705 ;
  assign n2707 = n2706 ^ n2702 ;
  assign n2708 = ~n2698 & ~n2707 ;
  assign n2732 = n2731 ^ n2708 ;
  assign n2733 = n2732 ^ n1002 ;
  assign n2742 = n2741 ^ n2733 ;
  assign n2745 = n2744 ^ n2742 ;
  assign n2695 = n2694 ^ n2685 ;
  assign n2696 = n2671 & ~n2695 ;
  assign n2746 = n2745 ^ n2696 ;
  assign n2666 = n2614 & n2663 ;
  assign n2667 = n2666 ^ n2611 ;
  assign n2668 = ~n2252 & n2667 ;
  assign n2747 = n2746 ^ n2668 ;
  assign n2748 = n2747 ^ x83 ;
  assign n1677 = n663 & n1676 ;
  assign n1667 = n623 ^ n619 ;
  assign n1668 = n1667 ^ n600 ;
  assign n1669 = n1668 ^ n860 ;
  assign n1665 = n628 ^ n616 ;
  assign n1666 = n1665 ^ n613 ;
  assign n1670 = n1669 ^ n1666 ;
  assign n1671 = n1670 ^ n860 ;
  assign n1672 = n582 & ~n1671 ;
  assign n1673 = n1672 ^ n1669 ;
  assign n1674 = n583 & ~n1673 ;
  assign n1661 = n860 ^ n620 ;
  assign n1662 = n1661 ^ n1335 ;
  assign n1663 = n1662 ^ n883 ;
  assign n1664 = n1663 ^ x45 ;
  assign n1675 = n1674 ^ n1664 ;
  assign n1678 = n1677 ^ n1675 ;
  assign n1658 = ~n583 & n618 ;
  assign n1659 = n1658 ^ n620 ;
  assign n1660 = ~n582 & n1659 ;
  assign n1679 = n1678 ^ n1660 ;
  assign n1680 = n1679 ^ x109 ;
  assign n1682 = n432 ^ n382 ;
  assign n1683 = n1682 ^ n436 ;
  assign n1686 = n1683 ^ n359 ;
  assign n1687 = ~n358 & ~n1686 ;
  assign n1688 = n1687 ^ n359 ;
  assign n1689 = n908 ^ n390 ;
  assign n1684 = n1683 ^ n908 ;
  assign n1690 = n1689 ^ n1684 ;
  assign n1691 = n1690 ^ n383 ;
  assign n1692 = n1688 & ~n1691 ;
  assign n1693 = n1692 ^ n1684 ;
  assign n1694 = n1693 ^ n391 ;
  assign n1703 = n1694 ^ n388 ;
  assign n1701 = n435 ^ n348 ;
  assign n1702 = n359 & ~n1701 ;
  assign n1704 = n1703 ^ n1702 ;
  assign n1705 = ~n358 & ~n1704 ;
  assign n1695 = n1694 ^ n445 ;
  assign n1696 = n1695 ^ n457 ;
  assign n1697 = n1696 ^ n1254 ;
  assign n1698 = n1697 ^ n922 ;
  assign n1699 = n1698 ^ n467 ;
  assign n1700 = n1699 ^ x53 ;
  assign n1706 = n1705 ^ n1700 ;
  assign n1707 = n1706 ^ x94 ;
  assign n1708 = n1680 & ~n1707 ;
  assign n1710 = n225 ^ x92 ;
  assign n1739 = n1738 ^ x83 ;
  assign n1740 = n1710 & n1739 ;
  assign n1756 = n1708 & n1740 ;
  assign n1654 = n1653 ^ x77 ;
  assign n1807 = n1806 ^ x126 ;
  assign n1813 = n1654 & ~n1807 ;
  assign n1857 = n1813 ^ n1807 ;
  assign n1858 = n1756 & ~n1857 ;
  assign n1709 = n1708 ^ n1707 ;
  assign n1758 = n1709 ^ n1680 ;
  assign n1759 = n1740 & n1758 ;
  assign n1741 = n1740 ^ n1739 ;
  assign n1748 = n1708 & n1741 ;
  assign n1743 = ~n1709 & n1740 ;
  assign n1749 = n1748 ^ n1743 ;
  assign n1750 = n1749 ^ n1741 ;
  assign n1744 = n1708 ^ n1680 ;
  assign n1745 = n1741 & n1744 ;
  assign n1746 = n1745 ^ n1743 ;
  assign n1742 = ~n1709 & n1741 ;
  assign n1747 = n1746 ^ n1742 ;
  assign n1751 = n1750 ^ n1747 ;
  assign n1822 = n1759 ^ n1751 ;
  assign n1854 = n1654 & n1822 ;
  assign n1855 = n1854 ^ n1759 ;
  assign n1856 = ~n1807 & n1855 ;
  assign n1859 = n1858 ^ n1856 ;
  assign n1767 = n1741 ^ n1710 ;
  assign n1818 = ~n1709 & ~n1767 ;
  assign n1817 = n1708 & ~n1767 ;
  assign n1819 = n1818 ^ n1817 ;
  assign n1768 = n1744 & ~n1767 ;
  assign n1816 = n1768 ^ n1767 ;
  assign n1820 = n1819 ^ n1816 ;
  assign n1821 = n1820 ^ n1758 ;
  assign n1823 = n1822 ^ n1821 ;
  assign n1752 = n1740 ^ n1710 ;
  assign n1753 = n1708 & n1752 ;
  assign n1754 = n1753 ^ n1752 ;
  assign n2753 = n1823 ^ n1754 ;
  assign n1760 = n1759 ^ n1753 ;
  assign n1761 = n1760 ^ n1745 ;
  assign n1824 = n1820 ^ n1761 ;
  assign n1834 = n1824 ^ n1818 ;
  assign n1837 = n2753 ^ n1834 ;
  assign n1838 = n1654 & n1837 ;
  assign n1860 = n1859 ^ n1838 ;
  assign n1844 = n1756 ^ n1749 ;
  assign n1847 = ~n1654 & n1844 ;
  assign n1848 = n1847 ^ n1756 ;
  assign n1849 = n1807 & n1848 ;
  assign n1861 = n1860 ^ n1849 ;
  assign n1862 = n1861 ^ x18 ;
  assign n1815 = n1807 ^ n1654 ;
  assign n1769 = n1768 ^ n1753 ;
  assign n1839 = n1817 ^ n1769 ;
  assign n1840 = n1839 ^ n1823 ;
  assign n1841 = n1840 ^ n1838 ;
  assign n1757 = n1756 ^ n1746 ;
  assign n1762 = n1761 ^ n1757 ;
  assign n1755 = n1754 ^ n1710 ;
  assign n1763 = n1762 ^ n1755 ;
  assign n1825 = n1763 ^ n1742 ;
  assign n1826 = n1825 ^ n1759 ;
  assign n1827 = n1826 ^ n1824 ;
  assign n1770 = n1769 ^ n1748 ;
  assign n1771 = n1770 ^ n1761 ;
  assign n1765 = n1739 ^ n1710 ;
  assign n1766 = n1765 ^ n1707 ;
  assign n1772 = n1771 ^ n1766 ;
  assign n1828 = n1827 ^ n1772 ;
  assign n1829 = n1828 ^ n1823 ;
  assign n1830 = n1829 ^ n1768 ;
  assign n1831 = n1830 ^ n1818 ;
  assign n1832 = n1831 ^ n1752 ;
  assign n1833 = ~n1654 & n1832 ;
  assign n1842 = n1841 ^ n1833 ;
  assign n1843 = n1815 & ~n1842 ;
  assign n1863 = n1862 ^ n1843 ;
  assign n1814 = n1747 & n1813 ;
  assign n1864 = n1863 ^ n1814 ;
  assign n1764 = n1763 ^ n1751 ;
  assign n1773 = n1772 ^ n1764 ;
  assign n1810 = n1773 & n1807 ;
  assign n1811 = n1810 ^ n1772 ;
  assign n1812 = ~n1654 & n1811 ;
  assign n1865 = n1864 ^ n1812 ;
  assign n1866 = n1865 ^ x104 ;
  assign n2037 = n2036 ^ x26 ;
  assign n1965 = ~n1946 & ~n1964 ;
  assign n1948 = n1942 & ~n1947 ;
  assign n1966 = n1965 ^ n1948 ;
  assign n2000 = n1976 ^ n1940 ;
  assign n2027 = n1945 & n2000 ;
  assign n2028 = n2027 ^ n2026 ;
  assign n2010 = n1960 ^ n1950 ;
  assign n2012 = n2011 ^ n2010 ;
  assign n2008 = n1957 ^ n1938 ;
  assign n2009 = n2008 ^ n1936 ;
  assign n2013 = n2012 ^ n2009 ;
  assign n2014 = n1943 & n2013 ;
  assign n2015 = n2014 ^ n1938 ;
  assign n2016 = ~n2007 & n2015 ;
  assign n1995 = n1945 & n1957 ;
  assign n1993 = n1967 ^ n1953 ;
  assign n1994 = n1993 ^ n1987 ;
  assign n1996 = n1995 ^ n1994 ;
  assign n1998 = n1997 ^ n1996 ;
  assign n2001 = n2000 ^ n1991 ;
  assign n2002 = n2001 ^ n1996 ;
  assign n1999 = n1945 & n1968 ;
  assign n2003 = n2002 ^ n1999 ;
  assign n2004 = n1998 & n2003 ;
  assign n2005 = n2004 ^ n1997 ;
  assign n1992 = ~n1946 & n1991 ;
  assign n2006 = n2005 ^ n1992 ;
  assign n2017 = n2016 ^ n2006 ;
  assign n2019 = n2018 ^ n2017 ;
  assign n1977 = n1976 ^ n1956 ;
  assign n1980 = n1944 & n1977 ;
  assign n1981 = n1980 ^ n1956 ;
  assign n1982 = ~n1943 & n1981 ;
  assign n2020 = n2019 ^ n1982 ;
  assign n2029 = n2028 ^ n2020 ;
  assign n2030 = ~n1966 & n2029 ;
  assign n2038 = n2037 ^ n2030 ;
  assign n2039 = n2038 ^ x105 ;
  assign n2191 = n1866 & ~n2039 ;
  assign n2202 = n2191 ^ n2039 ;
  assign n2203 = n2202 ^ n1866 ;
  assign n851 = n850 ^ x80 ;
  assign n907 = n906 ^ x75 ;
  assign n1184 = n1183 ^ x116 ;
  assign n954 = n953 ^ x70 ;
  assign n965 = n342 ^ x55 ;
  assign n959 = n180 ^ n170 ;
  assign n960 = n130 & ~n959 ;
  assign n961 = n960 ^ n170 ;
  assign n966 = n965 ^ n961 ;
  assign n962 = n961 ^ n169 ;
  assign n955 = n169 ^ n167 ;
  assign n956 = n955 ^ n189 ;
  assign n957 = n956 ^ n182 ;
  assign n958 = ~n130 & n957 ;
  assign n963 = n962 ^ n958 ;
  assign n964 = n129 & n963 ;
  assign n967 = n966 ^ n964 ;
  assign n968 = n967 ^ x93 ;
  assign n969 = ~n954 & ~n968 ;
  assign n1046 = n969 ^ n968 ;
  assign n1003 = n1002 ^ x76 ;
  assign n1012 = n755 ^ n708 ;
  assign n1013 = n1012 ^ n747 ;
  assign n1022 = n1021 ^ n1013 ;
  assign n1014 = n1013 ^ n717 ;
  assign n1015 = n725 & n1014 ;
  assign n1016 = n1015 ^ n717 ;
  assign n1018 = n1017 ^ n1013 ;
  assign n1019 = n1018 ^ n760 ;
  assign n1020 = n1016 & n1019 ;
  assign n1023 = n1022 ^ n1020 ;
  assign n1010 = n749 ^ n723 ;
  assign n1011 = ~n706 & n1010 ;
  assign n1026 = n1023 ^ n1011 ;
  assign n1027 = n725 & n1026 ;
  assign n1024 = n1023 ^ n788 ;
  assign n1028 = n1027 ^ n1024 ;
  assign n1004 = n755 ^ n739 ;
  assign n1007 = n706 & n1004 ;
  assign n1008 = n1007 ^ n739 ;
  assign n1009 = ~n717 & n1008 ;
  assign n1029 = n1028 ^ n1009 ;
  assign n1031 = n1030 ^ n1029 ;
  assign n1032 = n1031 ^ x47 ;
  assign n1033 = n1032 ^ x118 ;
  assign n1034 = ~n1003 & n1033 ;
  assign n1037 = n1034 ^ n1003 ;
  assign n1240 = n1046 ^ n1037 ;
  assign n1041 = n1037 ^ n1033 ;
  assign n1038 = n969 ^ n954 ;
  assign n1044 = n1038 ^ n968 ;
  assign n1045 = n1041 & ~n1044 ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1230 = n1045 ^ n1039 ;
  assign n1050 = n1034 ^ n1033 ;
  assign n1051 = ~n1046 & n1050 ;
  assign n1231 = n1230 ^ n1051 ;
  assign n1227 = n969 & ~n1037 ;
  assign n1047 = n1041 & ~n1046 ;
  assign n1035 = n969 & n1034 ;
  assign n1226 = n1047 ^ n1035 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1232 = n1231 ^ n1228 ;
  assign n1241 = n1240 ^ n1232 ;
  assign n1238 = n968 ^ n954 ;
  assign n1239 = n1238 ^ n1003 ;
  assign n1242 = n1241 ^ n1239 ;
  assign n1243 = ~n1184 & n1242 ;
  assign n1233 = n1184 & n1232 ;
  assign n1059 = n1034 & ~n1046 ;
  assign n1054 = n969 & n1050 ;
  assign n1053 = ~n1044 & n1050 ;
  assign n1055 = n1054 ^ n1053 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1056 = n1055 ^ n1052 ;
  assign n1048 = n1047 ^ n1045 ;
  assign n1042 = n969 & n1041 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1049 = n1048 ^ n1043 ;
  assign n1057 = n1056 ^ n1049 ;
  assign n1040 = n1039 ^ n1038 ;
  assign n1058 = n1057 ^ n1040 ;
  assign n1060 = n1059 ^ n1058 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1061 = n1060 ^ n1036 ;
  assign n1217 = n1061 ^ n1051 ;
  assign n1213 = ~n1037 & ~n1046 ;
  assign n1214 = n1213 ^ n1039 ;
  assign n1215 = n1214 ^ n1037 ;
  assign n1216 = n1215 ^ n1049 ;
  assign n1218 = n1217 ^ n1216 ;
  assign n1223 = ~n907 & n1218 ;
  assign n1224 = n1223 ^ n1053 ;
  assign n1225 = n1184 & n1224 ;
  assign n1229 = n1228 ^ n1225 ;
  assign n1234 = n1233 ^ n1229 ;
  assign n1244 = n1243 ^ n1234 ;
  assign n1245 = n1244 ^ n1225 ;
  assign n1246 = ~n907 & n1245 ;
  assign n1190 = ~n907 & n1184 ;
  assign n1210 = n1035 & n1190 ;
  assign n1207 = n1057 & n1184 ;
  assign n1208 = n1207 ^ n1056 ;
  assign n1209 = n907 & n1208 ;
  assign n1211 = n1210 ^ n1209 ;
  assign n1200 = n1049 & ~n1184 ;
  assign n1193 = n1051 ^ n1042 ;
  assign n1194 = n1184 & n1193 ;
  assign n1195 = n1194 ^ n1051 ;
  assign n1201 = n1200 ^ n1195 ;
  assign n1202 = n907 & n1201 ;
  assign n1212 = n1211 ^ n1202 ;
  assign n1235 = n1234 ^ n1212 ;
  assign n1191 = n1042 & n1190 ;
  assign n1062 = n1061 ^ n1039 ;
  assign n1063 = n1062 ^ n1060 ;
  assign n1187 = n1063 & ~n1184 ;
  assign n1188 = n1187 ^ n1060 ;
  assign n1189 = n907 & ~n1188 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n1236 = n1235 ^ n1192 ;
  assign n1237 = n1236 ^ x34 ;
  assign n1247 = n1246 ^ n1237 ;
  assign n1248 = n1247 ^ x98 ;
  assign n2172 = n2130 & n2161 ;
  assign n2168 = n2167 ^ n2101 ;
  assign n2169 = n2158 & n2168 ;
  assign n2162 = n2129 & n2161 ;
  assign n2144 = ~n2040 & n2143 ;
  assign n2145 = n2144 ^ n2142 ;
  assign n2156 = n2155 ^ n2145 ;
  assign n2135 = n2134 ^ n2129 ;
  assign n2146 = n2145 ^ n2135 ;
  assign n2124 = n2114 ^ n2102 ;
  assign n2136 = n2135 ^ n2124 ;
  assign n2137 = ~n2040 & ~n2136 ;
  assign n2147 = n2146 ^ n2137 ;
  assign n2148 = n2123 & ~n2147 ;
  assign n2157 = n2156 ^ n2148 ;
  assign n2163 = n2162 ^ n2157 ;
  assign n2170 = n2169 ^ n2163 ;
  assign n2116 = n2124 ^ n2105 ;
  assign n2117 = n2116 ^ n2102 ;
  assign n2120 = n2040 & n2117 ;
  assign n2121 = n2120 ^ n2102 ;
  assign n2122 = ~n2112 & n2121 ;
  assign n2171 = n2170 ^ n2122 ;
  assign n2173 = n2172 ^ n2171 ;
  assign n2175 = n2174 ^ n2173 ;
  assign n2111 = n2040 & n2110 ;
  assign n2176 = n2175 ^ n2111 ;
  assign n2183 = ~n2176 & ~n2182 ;
  assign n2184 = n2183 ^ x10 ;
  assign n2185 = n2184 ^ x66 ;
  assign n2244 = n1248 & ~n2185 ;
  assign n1615 = n1614 ^ x122 ;
  assign n2194 = ~n1615 & ~n2185 ;
  assign n2245 = n2244 ^ n2194 ;
  assign n2246 = ~n851 & n2245 ;
  assign n2247 = n2246 ^ n2245 ;
  assign n2248 = n2203 & n2247 ;
  assign n2195 = n2194 ^ n1615 ;
  assign n2222 = n2195 ^ n2185 ;
  assign n2205 = n2039 ^ n1866 ;
  assign n2204 = ~n1615 & ~n2203 ;
  assign n2206 = n2205 ^ n2204 ;
  assign n2198 = n1615 & n2039 ;
  assign n2200 = n2198 ^ n1615 ;
  assign n2201 = n2200 ^ n2191 ;
  assign n2207 = n2206 ^ n2201 ;
  assign n2236 = n2222 ^ n2207 ;
  assign n2219 = n2207 ^ n2205 ;
  assign n2216 = n2185 ^ n1615 ;
  assign n2217 = ~n2202 & ~n2216 ;
  assign n2213 = ~n1866 & n2194 ;
  assign n2214 = n2213 ^ n1615 ;
  assign n2215 = ~n2205 & ~n2214 ;
  assign n2218 = n2217 ^ n2215 ;
  assign n2220 = n2219 ^ n2218 ;
  assign n2192 = ~n1615 & n2191 ;
  assign n2235 = n2220 ^ n2192 ;
  assign n2237 = n2236 ^ n2235 ;
  assign n2230 = n2185 ^ n2039 ;
  assign n2229 = n2039 & ~n2195 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2232 = n1866 & ~n2231 ;
  assign n2233 = n2232 ^ n2215 ;
  assign n2234 = n2233 ^ n2220 ;
  assign n2238 = n2237 ^ n2234 ;
  assign n2239 = ~n1248 & n2238 ;
  assign n2240 = n2239 ^ n2234 ;
  assign n2223 = n2222 ^ n2198 ;
  assign n2224 = n1866 & ~n2223 ;
  assign n2208 = n2207 ^ n1615 ;
  assign n2209 = n2185 & n2208 ;
  assign n2210 = n2209 ^ n2204 ;
  assign n2221 = n2220 ^ n2210 ;
  assign n2225 = n2224 ^ n2221 ;
  assign n2197 = n2185 ^ n1866 ;
  assign n2199 = n2198 ^ n2197 ;
  assign n2226 = n2225 ^ n2199 ;
  assign n2193 = n2192 ^ n2191 ;
  assign n2196 = n2195 ^ n2193 ;
  assign n2227 = n2226 ^ n2196 ;
  assign n1867 = n1866 ^ n1615 ;
  assign n2186 = n2039 & ~n2185 ;
  assign n2187 = n2186 ^ n1866 ;
  assign n2188 = n1867 & ~n2187 ;
  assign n2189 = n2188 ^ n1866 ;
  assign n2190 = n1248 & n2189 ;
  assign n2228 = n2227 ^ n2190 ;
  assign n2241 = n2240 ^ n2228 ;
  assign n2242 = ~n851 & ~n2241 ;
  assign n2243 = n2242 ^ n2240 ;
  assign n2249 = n2248 ^ n2243 ;
  assign n2250 = n2249 ^ n225 ;
  assign n2251 = n2250 ^ x70 ;
  assign n3784 = n2748 ^ n2251 ;
  assign n3122 = n1479 & n1554 ;
  assign n3119 = n1500 & n1538 ;
  assign n3120 = n3119 ^ n1476 ;
  assign n3121 = n1544 & n3120 ;
  assign n3123 = n3122 ^ n3121 ;
  assign n3492 = n3123 ^ x4 ;
  assign n3477 = n1583 ^ n1484 ;
  assign n3478 = n3477 ^ n1546 ;
  assign n3487 = n3478 ^ n1543 ;
  assign n3481 = n1494 ^ n1350 ;
  assign n3482 = n3481 ^ n1557 ;
  assign n3483 = n3482 ^ n1605 ;
  assign n3484 = ~n1538 & ~n3483 ;
  assign n3479 = n3478 ^ n1482 ;
  assign n3124 = n1546 ^ n1496 ;
  assign n3125 = n1538 & ~n3124 ;
  assign n3126 = n3125 ^ n1496 ;
  assign n3480 = n3479 ^ n3126 ;
  assign n3485 = n3484 ^ n3480 ;
  assign n3486 = ~n1544 & n3485 ;
  assign n3488 = n3487 ^ n3486 ;
  assign n3114 = n1489 ^ n1485 ;
  assign n3476 = n1574 & n3114 ;
  assign n3489 = n3488 ^ n3476 ;
  assign n3470 = n1563 ^ n1491 ;
  assign n3473 = n1538 & n3470 ;
  assign n3474 = n3473 ^ n1491 ;
  assign n3475 = n1281 & n3474 ;
  assign n3490 = n3489 ^ n3475 ;
  assign n3491 = ~n1576 & ~n3490 ;
  assign n3493 = n3492 ^ n3491 ;
  assign n3494 = n3493 ^ x100 ;
  assign n3342 = n2167 ^ n2114 ;
  assign n3343 = n2159 & n3342 ;
  assign n3338 = n2617 ^ n2129 ;
  assign n3339 = n3338 ^ n2162 ;
  assign n3340 = ~n2159 & n3339 ;
  assign n3333 = n2109 ^ n2105 ;
  assign n3330 = n2109 ^ n2101 ;
  assign n3331 = n3330 ^ n2134 ;
  assign n3332 = ~n2040 & ~n3331 ;
  assign n3334 = n3333 ^ n3332 ;
  assign n3335 = n2112 & n3334 ;
  assign n3321 = n2651 ^ n2620 ;
  assign n3322 = n3321 ^ n2164 ;
  assign n3323 = n3322 ^ n2620 ;
  assign n3326 = ~n2112 & n3323 ;
  assign n3327 = n3326 ^ n2620 ;
  assign n3328 = ~n2040 & n3327 ;
  assign n3329 = n3328 ^ n2620 ;
  assign n3336 = n3335 ^ n3329 ;
  assign n3337 = n3336 ^ n2617 ;
  assign n3341 = n3340 ^ n3337 ;
  assign n3344 = n3343 ^ n3341 ;
  assign n3345 = n3344 ^ n2633 ;
  assign n3346 = n3345 ^ n2172 ;
  assign n3347 = n3346 ^ n2658 ;
  assign n3348 = n3347 ^ n2182 ;
  assign n3349 = n3348 ^ n2155 ;
  assign n3350 = n3349 ^ x46 ;
  assign n3351 = n3350 ^ x102 ;
  assign n2761 = n1813 ^ n1654 ;
  assign n3397 = n1751 ^ n1746 ;
  assign n3398 = n2761 & n3397 ;
  assign n3393 = n1826 ^ n1768 ;
  assign n3394 = ~n1807 & n3393 ;
  assign n2792 = n2761 ^ n1807 ;
  assign n2754 = n2753 ^ n1828 ;
  assign n2793 = n2754 ^ n1820 ;
  assign n2794 = n2792 & ~n2793 ;
  assign n3388 = n2794 ^ n1768 ;
  assign n3382 = n1819 ^ n1751 ;
  assign n3385 = ~n1654 & n3382 ;
  assign n3386 = n3385 ^ n1819 ;
  assign n3387 = ~n1815 & n3386 ;
  assign n3389 = n3388 ^ n3387 ;
  assign n3390 = n3389 ^ n1849 ;
  assign n3391 = n3390 ^ x62 ;
  assign n3375 = n1831 ^ n1826 ;
  assign n3376 = n3375 ^ n1830 ;
  assign n3379 = ~n1807 & n3376 ;
  assign n3380 = n3379 ^ n1830 ;
  assign n3381 = n1654 & n3380 ;
  assign n3392 = n3391 ^ n3381 ;
  assign n3395 = n3394 ^ n3392 ;
  assign n3374 = n1817 & n2792 ;
  assign n3396 = n3395 ^ n3374 ;
  assign n3399 = n3398 ^ n3396 ;
  assign n3373 = ~n1840 & ~n1857 ;
  assign n3400 = n3399 ^ n3373 ;
  assign n3366 = n1764 ^ n1749 ;
  assign n3365 = n1753 ^ n1742 ;
  assign n3367 = n3366 ^ n3365 ;
  assign n3370 = n1654 & n3367 ;
  assign n3371 = n3370 ^ n3365 ;
  assign n3372 = n1815 & n3371 ;
  assign n3401 = n3400 ^ n3372 ;
  assign n3402 = n3401 ^ x91 ;
  assign n3417 = ~n3351 & n3402 ;
  assign n2999 = n2493 & ~n2528 ;
  assign n3000 = ~n2495 & n2999 ;
  assign n3001 = n3000 ^ n2543 ;
  assign n3352 = n2572 ^ n2560 ;
  assign n3353 = n3352 ^ n2564 ;
  assign n3354 = n2456 & n3353 ;
  assign n3355 = n3354 ^ n2560 ;
  assign n3356 = n3355 ^ n2584 ;
  assign n3359 = n2495 & n3356 ;
  assign n3360 = n3359 ^ n3355 ;
  assign n3361 = ~n3001 & n3360 ;
  assign n3362 = n3361 ^ x54 ;
  assign n3363 = n3362 ^ x77 ;
  assign n3190 = ~n1944 & n1993 ;
  assign n3191 = n3190 ^ n1953 ;
  assign n3192 = ~n1943 & n3191 ;
  assign n3166 = n1957 ^ n1942 ;
  assign n3167 = n3166 ^ n1964 ;
  assign n3168 = n3167 ^ n1973 ;
  assign n3163 = n1976 ^ n1941 ;
  assign n3164 = n3163 ^ n1960 ;
  assign n3165 = n3164 ^ n1961 ;
  assign n3169 = n3168 ^ n3165 ;
  assign n3170 = ~n1944 & ~n3169 ;
  assign n3171 = n3170 ^ n3164 ;
  assign n3193 = n3192 ^ n3171 ;
  assign n3194 = n3193 ^ n2273 ;
  assign n3180 = n1990 ^ n1936 ;
  assign n3183 = n1943 & n3180 ;
  assign n3184 = n3183 ^ n1936 ;
  assign n3185 = n1944 & n3184 ;
  assign n3195 = n3194 ^ n3185 ;
  assign n3196 = n3195 ^ n2028 ;
  assign n3197 = n3196 ^ n2275 ;
  assign n3198 = n3197 ^ n1966 ;
  assign n3199 = n3198 ^ x38 ;
  assign n3173 = n3171 ^ n1958 ;
  assign n3172 = n3171 ^ n2012 ;
  assign n3174 = n3173 ^ n3172 ;
  assign n3177 = ~n1944 & n3174 ;
  assign n3178 = n3177 ^ n3173 ;
  assign n3179 = ~n1943 & ~n3178 ;
  assign n3200 = n3199 ^ n3179 ;
  assign n3403 = n3200 ^ x117 ;
  assign n3418 = n3363 & ~n3403 ;
  assign n3419 = n3418 ^ n3363 ;
  assign n3420 = n3419 ^ n3403 ;
  assign n3421 = n3417 & n3420 ;
  assign n3525 = n3494 ^ n3421 ;
  assign n2858 = n2370 ^ n2366 ;
  assign n2859 = n2858 ^ n2415 ;
  assign n2862 = ~n2396 & n2859 ;
  assign n2863 = n2862 ^ n2415 ;
  assign n2864 = ~n2287 & n2863 ;
  assign n2870 = n2358 & ~n2418 ;
  assign n3021 = n2432 ^ n2365 ;
  assign n3022 = n2417 & n3021 ;
  assign n3014 = n2371 ^ n2351 ;
  assign n3015 = n3014 ^ n2422 ;
  assign n3011 = n2395 ^ n2358 ;
  assign n3016 = n3015 ^ n3011 ;
  assign n3017 = ~n2396 & n3016 ;
  assign n3008 = n2390 ^ n2380 ;
  assign n3006 = n2378 ^ n2288 ;
  assign n3007 = ~n2396 & ~n3006 ;
  assign n3009 = n3008 ^ n3007 ;
  assign n3012 = n3011 ^ n3009 ;
  assign n3018 = n3017 ^ n3012 ;
  assign n3019 = n2287 & ~n3018 ;
  assign n2885 = n2375 ^ n2355 ;
  assign n2886 = n2885 ^ n2365 ;
  assign n2889 = n2396 & ~n2886 ;
  assign n2890 = n2889 ^ n2365 ;
  assign n2891 = n2287 & n2890 ;
  assign n3010 = n3009 ^ n2891 ;
  assign n3020 = n3019 ^ n3010 ;
  assign n3023 = n3022 ^ n3020 ;
  assign n3024 = ~n2441 & n3023 ;
  assign n3025 = ~n2870 & n3024 ;
  assign n3026 = ~n2864 & n3025 ;
  assign n3029 = n3026 ^ x30 ;
  assign n3005 = n2858 ^ n2432 ;
  assign n3027 = n2427 & n3026 ;
  assign n3028 = n3005 & n3027 ;
  assign n3030 = n3029 ^ n3028 ;
  assign n3320 = n3030 ^ x126 ;
  assign n3500 = n3320 & ~n3494 ;
  assign n3501 = n3500 ^ n3494 ;
  assign n3502 = n3501 ^ n3320 ;
  assign n3526 = n3525 ^ n3502 ;
  assign n3503 = n3502 ^ n3494 ;
  assign n3436 = n3417 & n3419 ;
  assign n3424 = n3417 ^ n3402 ;
  assign n3428 = n3424 ^ n3351 ;
  assign n3430 = n3428 ^ n3402 ;
  assign n3431 = n3418 & ~n3430 ;
  assign n3429 = n3418 & n3428 ;
  assign n3432 = n3431 ^ n3429 ;
  assign n3426 = n3418 & n3424 ;
  assign n3427 = n3426 ^ n3418 ;
  assign n3433 = n3432 ^ n3427 ;
  assign n3437 = n3436 ^ n3433 ;
  assign n3435 = n3421 ^ n3417 ;
  assign n3438 = n3437 ^ n3435 ;
  assign n3425 = n3420 & n3424 ;
  assign n3434 = n3433 ^ n3425 ;
  assign n3439 = n3438 ^ n3434 ;
  assign n3404 = n3402 & n3403 ;
  assign n3423 = n3417 ^ n3404 ;
  assign n3440 = n3439 ^ n3423 ;
  assign n3441 = n3440 ^ n3438 ;
  assign n3442 = n3441 ^ n3426 ;
  assign n3527 = n3494 ^ n3442 ;
  assign n3528 = n3503 & ~n3527 ;
  assign n3529 = n3528 ^ n3494 ;
  assign n3530 = n3526 & ~n3529 ;
  assign n3462 = n3420 ^ n3363 ;
  assign n3463 = n3428 & ~n3462 ;
  assign n3364 = n3363 ^ n3351 ;
  assign n3410 = n3402 ^ n3351 ;
  assign n3448 = n3410 ^ n3403 ;
  assign n3451 = n3351 & n3448 ;
  assign n3452 = n3451 ^ n3403 ;
  assign n3453 = ~n3364 & ~n3452 ;
  assign n3454 = n3453 ^ n3448 ;
  assign n3455 = n3454 ^ n3441 ;
  assign n3414 = n3403 ^ n3351 ;
  assign n3415 = n3414 ^ n3363 ;
  assign n3416 = n3415 ^ n3403 ;
  assign n3422 = n3421 ^ n3416 ;
  assign n3443 = n3442 ^ n3422 ;
  assign n3444 = n3443 ^ n3414 ;
  assign n3407 = n3403 ^ n3363 ;
  assign n3408 = n3407 ^ n3402 ;
  assign n3411 = n3363 & ~n3410 ;
  assign n3412 = ~n3408 & n3411 ;
  assign n3413 = n3412 ^ n3408 ;
  assign n3445 = n3444 ^ n3413 ;
  assign n3405 = n3404 ^ n3351 ;
  assign n3406 = ~n3364 & ~n3405 ;
  assign n3409 = n3408 ^ n3406 ;
  assign n3446 = n3445 ^ n3409 ;
  assign n3456 = n3455 ^ n3446 ;
  assign n3459 = n3456 ^ n3421 ;
  assign n3458 = n3414 ^ n3413 ;
  assign n3460 = n3459 ^ n3458 ;
  assign n3461 = n3460 ^ n3431 ;
  assign n3464 = n3463 ^ n3461 ;
  assign n3457 = n3456 ^ n3441 ;
  assign n3465 = n3464 ^ n3457 ;
  assign n3466 = n3465 ^ n3463 ;
  assign n3522 = n3466 ^ n3421 ;
  assign n3518 = n3436 ^ n3429 ;
  assign n3516 = n3433 ^ n3421 ;
  assign n3514 = n3426 ^ n3412 ;
  assign n3515 = ~n3501 & n3514 ;
  assign n3517 = n3516 ^ n3515 ;
  assign n3519 = n3518 ^ n3517 ;
  assign n3523 = n3522 ^ n3519 ;
  assign n3511 = n3461 ^ n3430 ;
  assign n3510 = n3465 ^ n3429 ;
  assign n3512 = n3511 ^ n3510 ;
  assign n3513 = ~n3501 & ~n3512 ;
  assign n3520 = n3519 ^ n3513 ;
  assign n3521 = ~n3500 & n3520 ;
  assign n3524 = n3523 ^ n3521 ;
  assign n3531 = n3530 ^ n3524 ;
  assign n3509 = n3439 & n3502 ;
  assign n3532 = n3531 ^ n3509 ;
  assign n3504 = n3503 ^ n3501 ;
  assign n3505 = n3429 ^ n3428 ;
  assign n3506 = n3505 ^ n3466 ;
  assign n3507 = n3506 ^ n3460 ;
  assign n3508 = n3504 & n3507 ;
  assign n3533 = n3532 ^ n3508 ;
  assign n3468 = n3466 ^ n3432 ;
  assign n3467 = n3466 ^ n3437 ;
  assign n3469 = n3468 ^ n3467 ;
  assign n3497 = n3469 & ~n3494 ;
  assign n3498 = n3497 ^ n3468 ;
  assign n3499 = ~n3320 & n3498 ;
  assign n3534 = n3533 ^ n3499 ;
  assign n3535 = n3426 ^ n3425 ;
  assign n3536 = n3535 ^ n3424 ;
  assign n3537 = n3536 ^ n3511 ;
  assign n3538 = n3511 ^ n3320 ;
  assign n3539 = n3538 ^ n3511 ;
  assign n3540 = ~n3537 & ~n3539 ;
  assign n3541 = n3540 ^ n3511 ;
  assign n3542 = ~n3504 & ~n3541 ;
  assign n3543 = ~n3534 & ~n3542 ;
  assign n3544 = n3543 ^ n2321 ;
  assign n3545 = n3544 ^ x126 ;
  assign n3593 = n1982 ^ n1948 ;
  assign n3576 = ~n1944 & n1986 ;
  assign n3577 = n3576 ^ n1988 ;
  assign n3578 = ~n1943 & ~n3577 ;
  assign n3579 = n3578 ^ n1971 ;
  assign n3580 = n3579 ^ n1938 ;
  assign n3581 = n3580 ^ n2010 ;
  assign n3582 = n3581 ^ n3578 ;
  assign n3583 = n1944 & ~n3582 ;
  assign n3584 = n3583 ^ n3579 ;
  assign n3594 = n3593 ^ n3584 ;
  assign n3595 = n3594 ^ n3192 ;
  assign n3596 = n3595 ^ n3185 ;
  assign n3597 = n3596 ^ n2266 ;
  assign n3598 = n3597 ^ n2036 ;
  assign n3599 = n3598 ^ x48 ;
  assign n3590 = n1944 & n3168 ;
  assign n3585 = n3584 ^ n3578 ;
  assign n3591 = n3590 ^ n3585 ;
  assign n3592 = ~n2007 & n3591 ;
  assign n3600 = n3599 ^ n3592 ;
  assign n3601 = n3600 ^ x73 ;
  assign n3621 = n1758 ^ n1756 ;
  assign n3622 = n3621 ^ n1769 ;
  assign n3623 = n3622 ^ n1822 ;
  assign n3624 = ~n1807 & n3623 ;
  assign n3625 = n3624 ^ n1769 ;
  assign n3626 = n1654 & n3625 ;
  assign n3616 = n1817 ^ n1759 ;
  assign n3617 = n3616 ^ n1828 ;
  assign n3618 = n2792 & ~n3617 ;
  assign n3609 = n2753 ^ n1769 ;
  assign n3612 = n3609 ^ n1825 ;
  assign n3608 = n1759 ^ n1747 ;
  assign n3610 = n3609 ^ n3608 ;
  assign n3611 = n1654 & ~n3610 ;
  assign n3613 = n3612 ^ n3611 ;
  assign n3614 = ~n1815 & ~n3613 ;
  assign n2778 = ~n1807 & n1819 ;
  assign n2771 = n1818 ^ n1748 ;
  assign n2772 = ~n1807 & n2771 ;
  assign n2773 = n2772 ^ n1818 ;
  assign n2779 = n2778 ^ n2773 ;
  assign n2780 = n1654 & n2779 ;
  assign n2781 = n2780 ^ n2773 ;
  assign n3603 = n2781 ^ n1825 ;
  assign n3604 = n3603 ^ n1856 ;
  assign n3605 = n3604 ^ n3387 ;
  assign n3606 = n3605 ^ n2794 ;
  assign n3607 = n3606 ^ x40 ;
  assign n3615 = n3614 ^ n3607 ;
  assign n3619 = n3618 ^ n3615 ;
  assign n3602 = n1745 & ~n1857 ;
  assign n3620 = n3619 ^ n3602 ;
  assign n3627 = n3626 ^ n3620 ;
  assign n3628 = n3627 ^ x99 ;
  assign n3629 = ~n3601 & ~n3628 ;
  assign n3630 = n3629 ^ n3628 ;
  assign n3631 = n3630 ^ n3601 ;
  assign n3002 = n3001 ^ x56 ;
  assign n2832 = n2575 ^ n2559 ;
  assign n2833 = n2832 ^ n2488 ;
  assign n2834 = n2833 ^ n2553 ;
  assign n2835 = n2834 ^ n2559 ;
  assign n2836 = n2495 & n2835 ;
  assign n2837 = n2836 ^ n2832 ;
  assign n2990 = n2837 ^ n2562 ;
  assign n2991 = n2990 ^ n2547 ;
  assign n2992 = n2991 ^ n2579 ;
  assign n2993 = n2992 ^ n2837 ;
  assign n2994 = ~n2495 & n2993 ;
  assign n2995 = n2994 ^ n2990 ;
  assign n2996 = n2456 & ~n2995 ;
  assign n2997 = n2996 ^ n2837 ;
  assign n2998 = n2576 & n2997 ;
  assign n3003 = n3002 ^ n2998 ;
  assign n3632 = n3003 ^ x90 ;
  assign n3657 = n2392 ^ n2381 ;
  assign n3658 = ~n2287 & n3657 ;
  assign n3654 = n3021 ^ n2858 ;
  assign n3655 = ~n2418 & n3654 ;
  assign n3651 = n2433 ^ n2395 ;
  assign n3652 = n2427 & n3651 ;
  assign n3648 = n2426 ^ n2390 ;
  assign n3649 = n2419 & ~n3648 ;
  assign n3641 = n2396 & n2422 ;
  assign n3642 = n3641 ^ n2395 ;
  assign n3643 = n2411 & n3642 ;
  assign n3633 = n2447 ^ n2415 ;
  assign n3634 = n3633 ^ n2380 ;
  assign n3635 = n3634 ^ n2393 ;
  assign n3636 = n3635 ^ n2447 ;
  assign n3637 = ~n2411 & ~n3636 ;
  assign n3638 = n3637 ^ n3633 ;
  assign n3644 = n3643 ^ n3638 ;
  assign n3645 = n3644 ^ n2450 ;
  assign n2851 = n2379 & n2417 ;
  assign n2852 = n2851 ^ n2447 ;
  assign n3646 = n3645 ^ n2852 ;
  assign n3647 = n3646 ^ x32 ;
  assign n3650 = n3649 ^ n3647 ;
  assign n3653 = n3652 ^ n3650 ;
  assign n3656 = n3655 ^ n3653 ;
  assign n3659 = n3658 ^ n3656 ;
  assign n3660 = n3659 ^ x88 ;
  assign n3661 = ~n3632 & n3660 ;
  assign n3662 = n3661 ^ n3632 ;
  assign n3663 = n3662 ^ n3660 ;
  assign n3679 = ~n3631 & n3663 ;
  assign n3675 = ~n3628 & n3663 ;
  assign n3678 = n3675 ^ n3663 ;
  assign n3680 = n3679 ^ n3678 ;
  assign n3550 = n2142 ^ n2105 ;
  assign n3548 = n2639 ^ n2104 ;
  assign n3546 = ~n2040 & n2073 ;
  assign n3547 = n3546 ^ n2643 ;
  assign n3549 = n3548 ^ n3547 ;
  assign n3551 = n3550 ^ n3549 ;
  assign n3552 = n2040 & n3551 ;
  assign n3553 = n3552 ^ n3549 ;
  assign n3560 = n3553 ^ n2166 ;
  assign n3559 = n2617 ^ n2134 ;
  assign n3561 = n3560 ^ n3559 ;
  assign n3555 = n2153 ^ n2134 ;
  assign n3558 = n2112 & ~n3555 ;
  assign n3562 = n3561 ^ n3558 ;
  assign n3563 = ~n2123 & ~n3562 ;
  assign n3554 = n3553 ^ n3547 ;
  assign n3556 = n3555 ^ n3554 ;
  assign n3557 = n3556 ^ n3343 ;
  assign n3564 = n3563 ^ n3557 ;
  assign n3565 = n3564 ^ n2172 ;
  assign n3566 = n3565 ^ n2174 ;
  assign n3567 = n3566 ^ n2658 ;
  assign n3568 = n3567 ^ x24 ;
  assign n3569 = n3568 ^ x121 ;
  assign n3060 = n1209 ^ n1189 ;
  assign n3041 = n1056 ^ n1051 ;
  assign n3042 = n3041 ^ n1215 ;
  assign n3035 = n1227 ^ n1059 ;
  assign n3038 = n907 & n3035 ;
  assign n3039 = n3038 ^ n1055 ;
  assign n3040 = ~n1184 & n3039 ;
  assign n3043 = n3042 ^ n3040 ;
  assign n3044 = n3043 ^ n1058 ;
  assign n3045 = n3044 ^ n1218 ;
  assign n3046 = n3045 ^ n3040 ;
  assign n3047 = ~n1184 & n3046 ;
  assign n3048 = n3047 ^ n3043 ;
  assign n3061 = n3060 ^ n3048 ;
  assign n3057 = n1048 & ~n1184 ;
  assign n3058 = n3057 ^ n1047 ;
  assign n3059 = n907 & n3058 ;
  assign n3062 = n3061 ^ n3059 ;
  assign n3063 = n3062 ^ x6 ;
  assign n3032 = n1184 ^ n907 ;
  assign n3049 = n1243 ^ n1242 ;
  assign n3050 = n3049 ^ n3040 ;
  assign n3051 = n3050 ^ n3048 ;
  assign n3052 = n3032 & ~n3051 ;
  assign n3064 = n3063 ^ n3052 ;
  assign n3570 = n3064 ^ x114 ;
  assign n3703 = ~n3569 & ~n3570 ;
  assign n3704 = n3703 ^ n3569 ;
  assign n3748 = n3680 & ~n3704 ;
  assign n3707 = ~n3631 & ~n3662 ;
  assign n3666 = n3629 ^ n3601 ;
  assign n3667 = ~n3662 & ~n3666 ;
  assign n3716 = n3707 ^ n3667 ;
  assign n3664 = n3663 ^ n3632 ;
  assign n3677 = ~n3630 & n3664 ;
  assign n3691 = n3677 ^ n3667 ;
  assign n3692 = n3691 ^ n3666 ;
  assign n3684 = ~n3630 & n3661 ;
  assign n3683 = n3629 & n3661 ;
  assign n3685 = n3684 ^ n3683 ;
  assign n3686 = n3685 ^ n3661 ;
  assign n3682 = ~n3631 & n3661 ;
  assign n3687 = n3686 ^ n3682 ;
  assign n3681 = n3680 ^ n3677 ;
  assign n3688 = n3687 ^ n3681 ;
  assign n3693 = n3692 ^ n3688 ;
  assign n3694 = n3693 ^ n3664 ;
  assign n3665 = ~n3631 & n3664 ;
  assign n3690 = n3677 ^ n3665 ;
  assign n3695 = n3694 ^ n3690 ;
  assign n3674 = ~n3630 & n3663 ;
  assign n3676 = n3675 ^ n3674 ;
  assign n3713 = n3695 ^ n3676 ;
  assign n3712 = n3683 ^ n3629 ;
  assign n3714 = n3713 ^ n3712 ;
  assign n3715 = n3714 ^ n3662 ;
  assign n3717 = n3716 ^ n3715 ;
  assign n3742 = ~n3704 & n3717 ;
  assign n3729 = n3714 ^ n3682 ;
  assign n3727 = n3707 ^ n3684 ;
  assign n3728 = n3727 ^ n3717 ;
  assign n3730 = n3729 ^ n3728 ;
  assign n3731 = n3569 & ~n3730 ;
  assign n3726 = n3707 ^ n3685 ;
  assign n3732 = n3731 ^ n3726 ;
  assign n3743 = n3742 ^ n3732 ;
  assign n3734 = n3680 ^ n3665 ;
  assign n3733 = n3732 ^ n3713 ;
  assign n3735 = n3734 ^ n3733 ;
  assign n3736 = n3735 ^ n3732 ;
  assign n3739 = n3569 & ~n3736 ;
  assign n3740 = n3739 ^ n3732 ;
  assign n3741 = ~n3570 & n3740 ;
  assign n3744 = n3743 ^ n3741 ;
  assign n3718 = n3717 ^ n3682 ;
  assign n3719 = n3718 ^ n3716 ;
  assign n3711 = n3693 ^ n3674 ;
  assign n3720 = n3719 ^ n3711 ;
  assign n3721 = n3711 ^ n3570 ;
  assign n3722 = n3721 ^ n3711 ;
  assign n3723 = ~n3720 & ~n3722 ;
  assign n3724 = n3723 ^ n3711 ;
  assign n3725 = ~n3569 & ~n3724 ;
  assign n3745 = n3744 ^ n3725 ;
  assign n3705 = n3704 ^ n3570 ;
  assign n3706 = n3705 ^ n3569 ;
  assign n3708 = n3707 ^ n3687 ;
  assign n3709 = n3708 ^ n3684 ;
  assign n3710 = ~n3706 & n3709 ;
  assign n3746 = n3745 ^ n3710 ;
  assign n3571 = n3570 ^ n3569 ;
  assign n3698 = n3693 ^ n3679 ;
  assign n3689 = n3688 ^ n3676 ;
  assign n3696 = n3695 ^ n3689 ;
  assign n3697 = n3696 ^ n3676 ;
  assign n3699 = n3698 ^ n3697 ;
  assign n3700 = ~n3569 & n3699 ;
  assign n3701 = n3700 ^ n3689 ;
  assign n3702 = ~n3571 & n3701 ;
  assign n3747 = n3746 ^ n3702 ;
  assign n3749 = n3748 ^ n3747 ;
  assign n3668 = n3667 ^ n3665 ;
  assign n3669 = n3667 ^ n3569 ;
  assign n3670 = n3669 ^ n3667 ;
  assign n3671 = n3668 & ~n3670 ;
  assign n3672 = n3671 ^ n3667 ;
  assign n3673 = n3571 & n3672 ;
  assign n3750 = n3749 ^ n3673 ;
  assign n3751 = n3750 ^ n2347 ;
  assign n3752 = n3751 ^ x76 ;
  assign n3753 = ~n3545 & ~n3752 ;
  assign n3754 = n3753 ^ n3752 ;
  assign n2795 = n2794 ^ x0 ;
  assign n2782 = n1761 ^ n1748 ;
  assign n2783 = n2782 ^ n2781 ;
  assign n2767 = n1807 ^ n1761 ;
  assign n2768 = ~n1815 & ~n2767 ;
  assign n2769 = n2768 ^ n1807 ;
  assign n2770 = n1762 & ~n2769 ;
  assign n2784 = n2783 ^ n2770 ;
  assign n2785 = n2784 ^ n2781 ;
  assign n2765 = n1831 ^ n1742 ;
  assign n2766 = ~n1807 & n2765 ;
  assign n2786 = n2785 ^ n2766 ;
  assign n2787 = ~n1815 & n2786 ;
  assign n2788 = n2787 ^ n2784 ;
  assign n2762 = n1817 ^ n1772 ;
  assign n2763 = n2762 ^ n1751 ;
  assign n2764 = n2761 & n2763 ;
  assign n2789 = n2788 ^ n2764 ;
  assign n2755 = n2754 ^ n1823 ;
  assign n2758 = n1654 & ~n2755 ;
  assign n2759 = n2758 ^ n1823 ;
  assign n2760 = n1815 & ~n2759 ;
  assign n2790 = n2789 ^ n2760 ;
  assign n2791 = ~n1859 & ~n2790 ;
  assign n2796 = n2795 ^ n2791 ;
  assign n2797 = n2796 ^ x107 ;
  assign n2752 = n2038 ^ x97 ;
  assign n2798 = n2797 ^ n2752 ;
  assign n2822 = n322 & n804 ;
  assign n2823 = n2822 ^ n701 ;
  assign n2824 = n796 & ~n2823 ;
  assign n2810 = n802 ^ n685 ;
  assign n2811 = n2810 ^ n697 ;
  assign n2814 = ~n796 & n2811 ;
  assign n2815 = n2814 ^ n697 ;
  assign n2816 = n837 & n2815 ;
  assign n2808 = n847 ^ n844 ;
  assign n2809 = n2808 ^ n823 ;
  assign n2817 = n2816 ^ n2809 ;
  assign n2825 = n2824 ^ n2817 ;
  assign n2802 = n699 ^ n683 ;
  assign n2803 = n2802 ^ n678 ;
  assign n2804 = n2803 ^ n838 ;
  assign n2805 = ~n796 & n2804 ;
  assign n2800 = n838 ^ n823 ;
  assign n2806 = n2805 ^ n2800 ;
  assign n2807 = ~n322 & n2806 ;
  assign n2826 = n2825 ^ n2807 ;
  assign n2827 = n2826 ^ n703 ;
  assign n2828 = n2827 ^ x58 ;
  assign n2799 = ~n694 & n830 ;
  assign n2829 = n2828 ^ n2799 ;
  assign n2830 = n2829 ^ x74 ;
  assign n2882 = n2394 & n2417 ;
  assign n2874 = ~n2428 & n2432 ;
  assign n2872 = n2429 ^ n2426 ;
  assign n2873 = n2872 ^ n2430 ;
  assign n2875 = n2874 ^ n2873 ;
  assign n2871 = n2870 ^ n2371 ;
  assign n2876 = n2875 ^ n2871 ;
  assign n2877 = n2876 ^ n2392 ;
  assign n2865 = n2858 ^ n2383 ;
  assign n2866 = ~n2287 & n2865 ;
  assign n2878 = n2877 ^ n2866 ;
  assign n2879 = ~n2411 & ~n2878 ;
  assign n2867 = n2866 ^ n2404 ;
  assign n2868 = n2867 ^ n2864 ;
  assign n2855 = n2364 ^ n2360 ;
  assign n2856 = n2855 ^ n2322 ;
  assign n2857 = n2419 & ~n2856 ;
  assign n2869 = n2868 ^ n2857 ;
  assign n2880 = n2879 ^ n2869 ;
  assign n2853 = n2394 ^ n2380 ;
  assign n2854 = ~n2287 & n2853 ;
  assign n2881 = n2880 ^ n2854 ;
  assign n2883 = n2882 ^ n2881 ;
  assign n2884 = ~n2852 & ~n2883 ;
  assign n2892 = n2884 & ~n2891 ;
  assign n2893 = n2892 ^ x42 ;
  assign n2894 = n2893 ^ x64 ;
  assign n2901 = ~n2830 & ~n2894 ;
  assign n2902 = n2901 ^ n2894 ;
  assign n2903 = n2902 ^ n2830 ;
  assign n2831 = n1247 ^ x112 ;
  assign n2844 = n2576 ^ n2562 ;
  assign n2845 = n2844 ^ n2837 ;
  assign n2840 = n2562 ^ n2530 ;
  assign n2841 = n2840 ^ n2547 ;
  assign n2842 = n2841 ^ n2550 ;
  assign n2843 = ~n2495 & n2842 ;
  assign n2846 = n2845 ^ n2843 ;
  assign n2847 = ~n2456 & ~n2846 ;
  assign n2838 = n2545 ^ x50 ;
  assign n2839 = n2838 ^ n2837 ;
  assign n2848 = n2847 ^ n2839 ;
  assign n2849 = n2848 ^ x65 ;
  assign n2896 = n2831 & ~n2849 ;
  assign n2905 = n2896 ^ n2831 ;
  assign n2912 = n2905 ^ n2849 ;
  assign n2913 = n2912 ^ n2831 ;
  assign n2966 = ~n2903 & ~n2913 ;
  assign n2906 = n2901 ^ n2830 ;
  assign n2920 = ~n2906 & n2912 ;
  assign n2951 = n2920 ^ n2896 ;
  assign n2850 = n2849 ^ n2831 ;
  assign n2895 = n2894 ^ n2850 ;
  assign n2897 = n2896 ^ n2895 ;
  assign n2898 = n2830 & n2897 ;
  assign n2922 = n2903 ^ n2898 ;
  assign n2921 = n2920 ^ n2912 ;
  assign n2923 = n2922 ^ n2921 ;
  assign n2909 = n2901 & n2905 ;
  assign n2927 = n2923 ^ n2909 ;
  assign n2914 = n2901 & ~n2913 ;
  assign n2907 = n2905 & ~n2906 ;
  assign n2915 = n2914 ^ n2907 ;
  assign n2928 = n2927 ^ n2915 ;
  assign n2926 = n2907 ^ n2901 ;
  assign n2929 = n2928 ^ n2926 ;
  assign n2930 = n2929 ^ n2920 ;
  assign n2911 = n2896 & ~n2906 ;
  assign n2949 = n2930 ^ n2911 ;
  assign n2904 = n2896 & ~n2903 ;
  assign n2950 = n2949 ^ n2904 ;
  assign n2952 = n2951 ^ n2950 ;
  assign n2953 = n2952 ^ n2902 ;
  assign n2941 = ~n2902 & ~n2913 ;
  assign n2940 = ~n2902 & n2905 ;
  assign n2942 = n2941 ^ n2940 ;
  assign n2954 = n2953 ^ n2942 ;
  assign n2955 = n2954 ^ n2922 ;
  assign n2976 = n2966 ^ n2955 ;
  assign n2975 = n2904 ^ n2903 ;
  assign n2977 = n2976 ^ n2975 ;
  assign n2978 = n2977 ^ n2954 ;
  assign n2931 = n2930 ^ n2927 ;
  assign n2932 = n2931 ^ n2830 ;
  assign n2916 = n2915 ^ n2911 ;
  assign n2933 = n2932 ^ n2916 ;
  assign n2979 = n2978 ^ n2933 ;
  assign n2980 = n2933 ^ n2797 ;
  assign n2981 = n2980 ^ n2933 ;
  assign n2982 = ~n2979 & ~n2981 ;
  assign n2983 = n2982 ^ n2933 ;
  assign n2984 = ~n2798 & ~n2983 ;
  assign n2965 = n2954 ^ n2952 ;
  assign n2967 = n2966 ^ n2965 ;
  assign n2968 = n2967 ^ n2966 ;
  assign n2969 = n2968 ^ n2966 ;
  assign n2970 = n2966 ^ n2752 ;
  assign n2971 = n2970 ^ n2966 ;
  assign n2972 = ~n2969 & n2971 ;
  assign n2973 = n2972 ^ n2966 ;
  assign n2974 = ~n2798 & n2973 ;
  assign n2985 = n2984 ^ n2974 ;
  assign n2956 = n2955 ^ n2930 ;
  assign n2957 = n2956 ^ n2955 ;
  assign n2958 = n2955 ^ n2752 ;
  assign n2959 = n2958 ^ n2955 ;
  assign n2960 = ~n2957 & n2959 ;
  assign n2961 = n2960 ^ n2955 ;
  assign n2962 = ~n2798 & ~n2961 ;
  assign n2963 = n2962 ^ n2955 ;
  assign n2943 = n2942 ^ n2904 ;
  assign n2917 = ~n2752 & ~n2797 ;
  assign n2918 = n2917 ^ n2752 ;
  assign n2924 = n2918 ^ n2797 ;
  assign n2925 = n2924 ^ n2752 ;
  assign n2935 = n2920 ^ n2907 ;
  assign n2934 = n2933 ^ n2923 ;
  assign n2936 = n2935 ^ n2934 ;
  assign n2937 = n2925 & ~n2936 ;
  assign n2944 = n2943 ^ n2937 ;
  assign n2919 = ~n2916 & n2918 ;
  assign n2938 = n2923 & ~n2937 ;
  assign n2939 = n2919 & n2938 ;
  assign n2945 = n2944 ^ n2939 ;
  assign n2964 = n2963 ^ n2945 ;
  assign n2986 = n2985 ^ n2964 ;
  assign n2987 = n2986 ^ n1183 ;
  assign n2908 = n2907 ^ n2904 ;
  assign n2910 = n2909 ^ n2908 ;
  assign n2946 = n2945 ^ n2910 ;
  assign n2899 = n2898 ^ n2895 ;
  assign n2900 = ~n2797 & n2899 ;
  assign n2947 = n2946 ^ n2900 ;
  assign n2948 = ~n2798 & ~n2947 ;
  assign n2988 = n2987 ^ n2948 ;
  assign n2989 = n2988 ^ x109 ;
  assign n3004 = n3003 ^ x70 ;
  assign n3201 = n3200 ^ x84 ;
  assign n3207 = ~n3004 & n3201 ;
  assign n3104 = n695 & ~n796 ;
  assign n3090 = n704 ^ n696 ;
  assign n3087 = n700 ^ n684 ;
  assign n3085 = n345 & n796 ;
  assign n3086 = n581 & n3085 ;
  assign n3088 = n3087 ^ n3086 ;
  assign n3089 = n3088 ^ n678 ;
  assign n3091 = n3090 ^ n3089 ;
  assign n3092 = n3091 ^ n3088 ;
  assign n3095 = n796 & n3092 ;
  assign n3096 = n3095 ^ n3088 ;
  assign n3097 = n837 & n3096 ;
  assign n3098 = n3097 ^ n3088 ;
  assign n3102 = n3098 ^ n687 ;
  assign n3083 = n802 ^ n691 ;
  assign n3080 = n684 ^ n672 ;
  assign n3081 = n3080 ^ n693 ;
  assign n3082 = ~n796 & ~n3081 ;
  assign n3084 = n3083 ^ n3082 ;
  assign n3099 = n3098 ^ n3084 ;
  assign n3103 = n3102 ^ n3099 ;
  assign n3105 = n3104 ^ n3103 ;
  assign n3106 = ~n322 & n3105 ;
  assign n3076 = n674 & ~n796 ;
  assign n3069 = n804 ^ n689 ;
  assign n3070 = ~n796 & n3069 ;
  assign n3071 = n3070 ^ n804 ;
  assign n3077 = n3076 ^ n3071 ;
  assign n3078 = ~n837 & n3077 ;
  assign n3079 = n3078 ^ n3071 ;
  assign n3100 = n3099 ^ n3079 ;
  assign n3101 = n3100 ^ n801 ;
  assign n3107 = n3106 ^ n3101 ;
  assign n3108 = n3107 ^ n835 ;
  assign n3109 = n3108 ^ n843 ;
  assign n3068 = ~n696 & n831 ;
  assign n3110 = n3109 ^ n3068 ;
  assign n3111 = ~n847 & ~n3110 ;
  assign n3112 = n3111 ^ x14 ;
  assign n3113 = n3112 ^ x101 ;
  assign n3031 = n3030 ^ x116 ;
  assign n3240 = n3113 ^ n3031 ;
  assign n3144 = n1495 & n1574 ;
  assign n3141 = n1563 ^ n1502 ;
  assign n3142 = ~n1595 & ~n3141 ;
  assign n3137 = n1477 & n1574 ;
  assign n3134 = n1503 ^ n1493 ;
  assign n3135 = n3134 ^ n1564 ;
  assign n3128 = n1579 ^ n1557 ;
  assign n3127 = n3126 ^ n1485 ;
  assign n3129 = n3128 ^ n3127 ;
  assign n3130 = n3129 ^ n3126 ;
  assign n3131 = n1538 & n3130 ;
  assign n3132 = n3131 ^ n3127 ;
  assign n3136 = n3135 ^ n3132 ;
  assign n3138 = n3137 ^ n3136 ;
  assign n3139 = n1544 & ~n3138 ;
  assign n3133 = n3132 ^ n1600 ;
  assign n3140 = n3139 ^ n3133 ;
  assign n3143 = n3142 ^ n3140 ;
  assign n3145 = n3144 ^ n3143 ;
  assign n3146 = ~n3123 & ~n3145 ;
  assign n3147 = ~n1612 & n3146 ;
  assign n3148 = ~n1481 & n3147 ;
  assign n3151 = n3148 ^ x22 ;
  assign n3149 = n1553 & n3148 ;
  assign n3150 = n3114 & n3149 ;
  assign n3152 = n3151 ^ n3150 ;
  assign n3153 = n3152 ^ x83 ;
  assign n3154 = ~n3113 & ~n3153 ;
  assign n3158 = n3154 ^ n3153 ;
  assign n3065 = n3064 ^ x94 ;
  assign n3066 = n3031 & ~n3065 ;
  assign n3067 = n3066 ^ n3031 ;
  assign n3220 = n3067 ^ n3065 ;
  assign n3224 = ~n3158 & n3220 ;
  assign n3155 = n3154 ^ n3113 ;
  assign n3156 = n3155 ^ n3153 ;
  assign n3214 = n3066 ^ n3065 ;
  assign n3215 = ~n3156 & ~n3214 ;
  assign n3229 = n3224 ^ n3215 ;
  assign n3223 = ~n3155 & ~n3214 ;
  assign n3225 = n3224 ^ n3223 ;
  assign n3210 = ~n3031 & n3153 ;
  assign n3226 = n3225 ^ n3210 ;
  assign n3222 = n3220 ^ n3215 ;
  assign n3227 = n3226 ^ n3222 ;
  assign n3221 = ~n3155 & n3220 ;
  assign n3228 = n3227 ^ n3221 ;
  assign n3230 = n3229 ^ n3228 ;
  assign n3241 = n3240 ^ n3230 ;
  assign n3208 = n3065 ^ n3031 ;
  assign n3209 = n3208 ^ n3153 ;
  assign n3217 = ~n3031 & n3113 ;
  assign n3218 = n3217 ^ n3158 ;
  assign n3238 = n3218 ^ n3153 ;
  assign n3239 = n3209 & n3238 ;
  assign n3242 = n3241 ^ n3239 ;
  assign n3234 = n3154 & ~n3214 ;
  assign n3235 = n3234 ^ n3228 ;
  assign n3236 = n3235 ^ n3031 ;
  assign n3237 = n3236 ^ n3155 ;
  assign n3243 = n3242 ^ n3237 ;
  assign n3244 = n3243 ^ n3067 ;
  assign n3231 = n3230 ^ n3222 ;
  assign n3159 = n3066 & ~n3158 ;
  assign n3216 = n3215 ^ n3159 ;
  assign n3219 = n3218 ^ n3216 ;
  assign n3232 = n3231 ^ n3219 ;
  assign n3157 = n3067 & ~n3156 ;
  assign n3233 = n3232 ^ n3157 ;
  assign n3245 = n3244 ^ n3233 ;
  assign n3246 = n3245 ^ n3228 ;
  assign n3211 = n3210 ^ n3209 ;
  assign n3212 = ~n3113 & ~n3211 ;
  assign n3213 = n3212 ^ n3113 ;
  assign n3247 = n3246 ^ n3213 ;
  assign n3248 = n3247 ^ n3245 ;
  assign n3249 = n3207 & ~n3248 ;
  assign n3160 = n3159 ^ n3157 ;
  assign n3204 = n3160 & ~n3201 ;
  assign n3205 = n3204 ^ n3159 ;
  assign n3206 = ~n3004 & n3205 ;
  assign n3250 = n3249 ^ n3206 ;
  assign n3274 = n3201 ^ n3004 ;
  assign n3277 = n3066 & ~n3156 ;
  assign n3278 = n3277 ^ n3248 ;
  assign n3275 = n3245 ^ n3159 ;
  assign n3276 = n3275 ^ n3066 ;
  assign n3279 = n3278 ^ n3276 ;
  assign n3280 = n3279 ^ n3243 ;
  assign n3281 = ~n3274 & n3280 ;
  assign n3258 = n3207 ^ n3004 ;
  assign n3270 = n3258 ^ n3201 ;
  assign n3271 = n3228 ^ n3160 ;
  assign n3272 = n3270 & n3271 ;
  assign n3260 = n3234 ^ n3201 ;
  assign n3261 = n3234 ^ n3215 ;
  assign n3262 = n3261 ^ n3210 ;
  assign n3263 = n3262 ^ n3261 ;
  assign n3264 = n3261 ^ n3004 ;
  assign n3265 = n3264 ^ n3261 ;
  assign n3266 = n3263 & ~n3265 ;
  assign n3267 = n3266 ^ n3261 ;
  assign n3268 = n3260 & ~n3267 ;
  assign n3269 = n3268 ^ n3201 ;
  assign n3273 = n3272 ^ n3269 ;
  assign n3282 = n3281 ^ n3273 ;
  assign n3259 = n3227 & ~n3258 ;
  assign n3283 = n3282 ^ n3259 ;
  assign n3251 = n3232 ^ n3004 ;
  assign n3252 = n3251 ^ n3232 ;
  assign n3253 = n3232 ^ n3223 ;
  assign n3254 = n3253 ^ n3232 ;
  assign n3255 = n3252 & n3254 ;
  assign n3256 = n3255 ^ n3232 ;
  assign n3257 = n3201 & ~n3256 ;
  assign n3284 = n3283 ^ n3257 ;
  assign n3285 = ~n3250 & ~n3284 ;
  assign n3286 = n3248 ^ n3229 ;
  assign n3287 = n3229 ^ n3004 ;
  assign n3288 = n3287 ^ n3229 ;
  assign n3289 = ~n3286 & n3288 ;
  assign n3290 = n3289 ^ n3229 ;
  assign n3291 = ~n3201 & n3290 ;
  assign n3292 = n3285 & ~n3291 ;
  assign n3295 = n3215 ^ n3004 ;
  assign n3296 = n3295 ^ n3215 ;
  assign n3297 = n3216 & ~n3296 ;
  assign n3298 = n3297 ^ n3215 ;
  assign n3299 = ~n3201 & n3298 ;
  assign n3300 = n3292 & ~n3299 ;
  assign n3304 = n3270 ^ n3004 ;
  assign n3305 = n3231 ^ n3223 ;
  assign n3306 = n3305 ^ n3229 ;
  assign n3307 = n3306 ^ n3236 ;
  assign n3308 = n3307 ^ n3231 ;
  assign n3309 = n3304 & ~n3308 ;
  assign n3301 = n3277 ^ n3234 ;
  assign n3302 = n3004 & n3301 ;
  assign n3303 = n3302 ^ n3234 ;
  assign n3310 = n3309 ^ n3303 ;
  assign n3311 = n3310 ^ n3309 ;
  assign n3314 = ~n3201 & n3311 ;
  assign n3315 = n3314 ^ n3309 ;
  assign n3316 = n3300 & ~n3315 ;
  assign n3317 = n3316 ^ n1806 ;
  assign n3318 = n3317 ^ x116 ;
  assign n3319 = n2989 & n3318 ;
  assign n3762 = n3319 ^ n3318 ;
  assign n3804 = ~n3754 & n3762 ;
  assign n3756 = n3319 & n3753 ;
  assign n3817 = n3804 ^ n3756 ;
  assign n3776 = n3319 ^ n2989 ;
  assign n3787 = ~n3754 & n3776 ;
  assign n3768 = n3762 ^ n2989 ;
  assign n3771 = n3753 & ~n3768 ;
  assign n3788 = n3787 ^ n3771 ;
  assign n3761 = n3754 ^ n3545 ;
  assign n3779 = n3319 & ~n3761 ;
  assign n3763 = ~n3761 & n3762 ;
  assign n3780 = n3779 ^ n3763 ;
  assign n3757 = ~n3318 & n3753 ;
  assign n3777 = n3776 ^ n3757 ;
  assign n3778 = n3777 ^ n3761 ;
  assign n3781 = n3780 ^ n3778 ;
  assign n3785 = n3781 ^ n3776 ;
  assign n3769 = ~n3761 & ~n3768 ;
  assign n3770 = n3769 ^ n3757 ;
  assign n3786 = n3785 ^ n3770 ;
  assign n3789 = n3788 ^ n3786 ;
  assign n3818 = n3817 ^ n3789 ;
  assign n3819 = ~n2748 & ~n3818 ;
  assign n2749 = n2251 & n2748 ;
  assign n3811 = n3771 ^ n3757 ;
  assign n3792 = n3545 ^ n2989 ;
  assign n3793 = n3792 ^ n3752 ;
  assign n3794 = n3793 ^ n3781 ;
  assign n3758 = n3757 ^ n3753 ;
  assign n3759 = n3758 ^ n3756 ;
  assign n3755 = n3319 & ~n3754 ;
  assign n3760 = n3759 ^ n3755 ;
  assign n3764 = n3763 ^ n3760 ;
  assign n3795 = n3794 ^ n3764 ;
  assign n3773 = n3753 ^ n3545 ;
  assign n3774 = n3762 & ~n3773 ;
  assign n3796 = n3795 ^ n3774 ;
  assign n3790 = n3789 ^ n3777 ;
  assign n3791 = n3790 ^ n3773 ;
  assign n3797 = n3796 ^ n3791 ;
  assign n3812 = n3811 ^ n3797 ;
  assign n3813 = ~n2749 & n3812 ;
  assign n3807 = n3777 ^ n3318 ;
  assign n3808 = n3807 ^ n3795 ;
  assign n3767 = n2749 ^ n2748 ;
  assign n3805 = n3804 ^ n3779 ;
  assign n3806 = n3767 & n3805 ;
  assign n3809 = n3808 ^ n3806 ;
  assign n3798 = n3797 ^ n3790 ;
  assign n3799 = n3790 ^ n2251 ;
  assign n3800 = n3799 ^ n3790 ;
  assign n3801 = ~n3798 & n3800 ;
  assign n3802 = n3801 ^ n3790 ;
  assign n3803 = ~n2748 & ~n3802 ;
  assign n3810 = n3809 ^ n3803 ;
  assign n3814 = n3813 ^ n3810 ;
  assign n3815 = n3814 ^ n3806 ;
  assign n3816 = n3815 ^ n3803 ;
  assign n3820 = n3819 ^ n3816 ;
  assign n3821 = n3784 & ~n3820 ;
  assign n3822 = n3821 ^ n3814 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3775 = n3774 ^ n3772 ;
  assign n3782 = n3781 ^ n3775 ;
  assign n3783 = n3767 & ~n3782 ;
  assign n3823 = n3822 ^ n3783 ;
  assign n2750 = n2749 ^ n2251 ;
  assign n2751 = n2750 ^ n2748 ;
  assign n3765 = n3764 ^ n3756 ;
  assign n3766 = ~n2751 & n3765 ;
  assign n3824 = n3823 ^ n3766 ;
  assign n3825 = n3763 ^ n3755 ;
  assign n3826 = n3825 ^ n3797 ;
  assign n3827 = n3797 ^ n2251 ;
  assign n3828 = n3827 ^ n3797 ;
  assign n3829 = n3826 & n3828 ;
  assign n3830 = n3829 ^ n3797 ;
  assign n3831 = n2748 & n3830 ;
  assign n3832 = n3824 & ~n3831 ;
  assign n3836 = n3832 ^ n3030 ;
  assign n3833 = n3795 ^ n3759 ;
  assign n3834 = n2251 & n3833 ;
  assign n3835 = n3832 & n3834 ;
  assign n3837 = n3836 ^ n3835 ;
  assign n5349 = n3837 ^ x94 ;
  assign n3920 = n2829 ^ x81 ;
  assign n3921 = n3659 ^ x72 ;
  assign n3922 = ~n3920 & n3921 ;
  assign n3923 = n3922 ^ n3920 ;
  assign n3924 = n3923 ^ n3921 ;
  assign n4052 = n3924 ^ n3922 ;
  assign n3925 = n2796 ^ x123 ;
  assign n3926 = n3128 ^ n1496 ;
  assign n3934 = n3926 ^ n3121 ;
  assign n3935 = n3934 ^ n1552 ;
  assign n3927 = n3926 ^ n1560 ;
  assign n3928 = n3927 ^ n3134 ;
  assign n3929 = n3928 ^ n3114 ;
  assign n3930 = n3929 ^ n3926 ;
  assign n3931 = ~n1538 & n3930 ;
  assign n3932 = n3931 ^ n3927 ;
  assign n3933 = ~n1544 & ~n3932 ;
  assign n3936 = n3935 ^ n3933 ;
  assign n3937 = ~n1573 & ~n3936 ;
  assign n3938 = ~n1597 & n3937 ;
  assign n3939 = ~n1600 & n3938 ;
  assign n3940 = ~n1612 & n3939 ;
  assign n3941 = n3940 ^ x16 ;
  assign n3942 = n3941 ^ x106 ;
  assign n3943 = ~n3925 & n3942 ;
  assign n3945 = n3568 ^ x96 ;
  assign n3976 = n1195 ^ n1047 ;
  assign n3973 = n1213 ^ n1058 ;
  assign n3972 = n3042 ^ n1048 ;
  assign n3974 = n3973 ^ n3972 ;
  assign n3975 = n1184 & n3974 ;
  assign n3977 = n3976 ^ n3975 ;
  assign n3978 = ~n907 & n3977 ;
  assign n3966 = n1211 ^ n1195 ;
  assign n3948 = n1059 ^ n1049 ;
  assign n3949 = n3948 ^ n1062 ;
  assign n3955 = n3949 ^ n1055 ;
  assign n3947 = n3035 ^ n1061 ;
  assign n3950 = n3949 ^ n3947 ;
  assign n3951 = n3947 ^ n1184 ;
  assign n3952 = n3032 & n3951 ;
  assign n3953 = n3952 ^ n1184 ;
  assign n3954 = n3950 & n3953 ;
  assign n3956 = n3955 ^ n3954 ;
  assign n3967 = n3966 ^ n3956 ;
  assign n3968 = n3967 ^ n3059 ;
  assign n3969 = n3968 ^ x8 ;
  assign n3957 = n1214 ^ n1035 ;
  assign n3958 = n3957 ^ n3956 ;
  assign n3959 = n3958 ^ n1059 ;
  assign n3960 = n3959 ^ n3956 ;
  assign n3963 = n907 & n3960 ;
  assign n3964 = n3963 ^ n3956 ;
  assign n3965 = n3032 & ~n3964 ;
  assign n3970 = n3969 ^ n3965 ;
  assign n3946 = n1042 & ~n1184 ;
  assign n3971 = n3970 ^ n3946 ;
  assign n3979 = n3978 ^ n3971 ;
  assign n3980 = n3979 ^ x113 ;
  assign n3981 = n3945 & ~n3980 ;
  assign n3998 = n3943 & n3981 ;
  assign n3982 = n3981 ^ n3945 ;
  assign n3983 = n3982 ^ n3980 ;
  assign n3944 = n3943 ^ n3925 ;
  assign n3986 = n3944 ^ n3942 ;
  assign n3990 = n3983 & n3986 ;
  assign n3988 = n3983 ^ n3945 ;
  assign n3989 = n3943 & ~n3988 ;
  assign n3991 = n3990 ^ n3989 ;
  assign n3999 = n3998 ^ n3991 ;
  assign n3994 = n3980 ^ n3925 ;
  assign n3995 = n3925 & ~n3945 ;
  assign n3996 = n3995 ^ n3942 ;
  assign n3997 = ~n3994 & n3996 ;
  assign n4000 = n3999 ^ n3997 ;
  assign n4054 = n4000 ^ n3982 ;
  assign n4001 = ~n3944 & ~n3988 ;
  assign n4002 = n4001 ^ n4000 ;
  assign n4003 = n4002 ^ n3998 ;
  assign n3987 = n3982 & n3986 ;
  assign n3992 = n3991 ^ n3987 ;
  assign n3985 = ~n3944 & n3981 ;
  assign n3993 = n3992 ^ n3985 ;
  assign n4004 = n4003 ^ n3993 ;
  assign n4005 = n4004 ^ n3994 ;
  assign n4009 = n4005 ^ n3989 ;
  assign n4008 = n3986 & ~n3988 ;
  assign n4010 = n4009 ^ n4008 ;
  assign n4006 = n4005 ^ n4001 ;
  assign n4007 = n4006 ^ n3988 ;
  assign n4011 = n4010 ^ n4007 ;
  assign n4036 = n4011 ^ n3992 ;
  assign n4029 = n3981 & n3986 ;
  assign n4030 = n4029 ^ n3998 ;
  assign n3984 = ~n3944 & n3983 ;
  assign n4035 = n4030 ^ n3984 ;
  assign n4037 = n4036 ^ n4035 ;
  assign n4033 = n3942 ^ n3925 ;
  assign n4014 = n3995 ^ n3983 ;
  assign n4034 = n4033 ^ n4014 ;
  assign n4038 = n4037 ^ n4034 ;
  assign n4039 = n4038 ^ n3987 ;
  assign n4055 = n4054 ^ n4039 ;
  assign n4031 = n4030 ^ n3981 ;
  assign n4032 = n4031 ^ n3985 ;
  assign n4065 = n4055 ^ n4032 ;
  assign n4577 = n4065 ^ n4001 ;
  assign n4578 = n4001 ^ n3920 ;
  assign n4579 = n4578 ^ n4001 ;
  assign n4580 = ~n4577 & ~n4579 ;
  assign n4581 = n4580 ^ n4001 ;
  assign n4582 = n4052 & n4581 ;
  assign n4583 = n3922 & n4001 ;
  assign n4584 = ~n4582 & n4583 ;
  assign n4585 = n4584 ^ n4582 ;
  assign n4596 = n4038 ^ n4029 ;
  assign n4597 = n3922 & n4596 ;
  assign n4623 = n4597 ^ n3922 ;
  assign n4012 = n4011 ^ n3984 ;
  assign n4617 = n4039 ^ n4012 ;
  assign n4618 = n4039 ^ n3921 ;
  assign n4619 = n4618 ^ n4039 ;
  assign n4620 = n4617 & n4619 ;
  assign n4621 = n4620 ^ n4039 ;
  assign n4622 = n3920 & ~n4621 ;
  assign n4624 = n4623 ^ n4622 ;
  assign n4598 = n4014 ^ n3990 ;
  assign n4599 = n4598 ^ n4012 ;
  assign n4600 = n3922 & ~n4599 ;
  assign n4601 = n4600 ^ n3924 ;
  assign n4625 = n4624 ^ n4601 ;
  assign n4611 = n4055 ^ n4005 ;
  assign n4612 = n4005 ^ n3920 ;
  assign n4613 = n4612 ^ n4005 ;
  assign n4614 = n4611 & ~n4613 ;
  assign n4615 = n4614 ^ n4005 ;
  assign n4616 = ~n4052 & ~n4615 ;
  assign n4626 = n4625 ^ n4616 ;
  assign n4080 = ~n3923 & ~n4006 ;
  assign n4049 = n3922 ^ n3921 ;
  assign n4079 = n3985 & n4049 ;
  assign n4081 = n4080 ^ n4079 ;
  assign n4627 = n4626 ^ n4081 ;
  assign n4605 = n4039 ^ n4030 ;
  assign n4606 = n4030 ^ n3920 ;
  assign n4607 = n4606 ^ n4030 ;
  assign n4608 = ~n4605 & n4607 ;
  assign n4609 = n4608 ^ n4030 ;
  assign n4610 = ~n4052 & n4609 ;
  assign n4628 = n4627 ^ n4610 ;
  assign n4602 = ~n4597 & n4601 ;
  assign n4603 = n3991 ^ n3922 ;
  assign n4604 = n4602 & ~n4603 ;
  assign n4629 = n4628 ^ n4604 ;
  assign n4594 = n4065 ^ n4008 ;
  assign n4595 = n3924 & ~n4594 ;
  assign n4630 = n4629 ^ n4595 ;
  assign n4587 = n4012 ^ n4000 ;
  assign n4586 = n4032 ^ n3989 ;
  assign n4588 = n4587 ^ n4586 ;
  assign n4589 = n4586 ^ n3920 ;
  assign n4590 = n4589 ^ n4586 ;
  assign n4591 = ~n4588 & ~n4590 ;
  assign n4592 = n4591 ^ n4586 ;
  assign n4593 = ~n4052 & n4592 ;
  assign n4631 = n4630 ^ n4593 ;
  assign n4632 = ~n4585 & ~n4631 ;
  assign n4633 = n4632 ^ n1280 ;
  assign n4634 = n4633 ^ x81 ;
  assign n4410 = n3441 ^ n1317 ;
  assign n4401 = ~n3320 & ~n3445 ;
  assign n4402 = n4401 ^ n3413 ;
  assign n4411 = n4410 ^ n4402 ;
  assign n4403 = n4402 ^ n3409 ;
  assign n4404 = n4403 ^ n4402 ;
  assign n4407 = n3320 & n4404 ;
  assign n4408 = n4407 ^ n4402 ;
  assign n4409 = n3494 & ~n4408 ;
  assign n4412 = n4411 ^ n4409 ;
  assign n4398 = n3454 & n3494 ;
  assign n4399 = n4398 ^ n3441 ;
  assign n4400 = ~n3320 & n4399 ;
  assign n4413 = n4412 ^ n4400 ;
  assign n4414 = n4413 ^ x96 ;
  assign n4453 = n3714 ^ n3684 ;
  assign n4454 = n4453 ^ n3687 ;
  assign n4455 = ~n3704 & ~n4454 ;
  assign n4436 = n3698 ^ n3695 ;
  assign n4445 = n4436 ^ ~n3693 ;
  assign n4446 = n4445 ^ n3690 ;
  assign n4447 = n3690 ^ n3569 ;
  assign n4448 = n4447 ^ n3690 ;
  assign n4449 = n4446 & ~n4448 ;
  assign n4450 = n4449 ^ n3690 ;
  assign n4451 = n3570 & n4450 ;
  assign n4432 = n3729 ^ n3674 ;
  assign n4430 = n3716 ^ n3684 ;
  assign n4431 = n4430 ^ n3705 ;
  assign n4433 = n4432 ^ n4431 ;
  assign n4434 = ~n3676 & ~n4433 ;
  assign n4435 = n4434 ^ n3705 ;
  assign n4441 = ~n3693 ^ n3676 ;
  assign n4440 = n3706 ^ ~n3693 ;
  assign n4442 = n4441 ^ n4440 ;
  assign n4443 = n4435 & ~n4442 ;
  assign n4444 = n4443 ^ n4441 ;
  assign n4452 = n4451 ^ n4444 ;
  assign n4456 = n4455 ^ n4452 ;
  assign n4420 = n3713 ^ n3708 ;
  assign n4419 = n3707 ^ n3677 ;
  assign n4421 = n4420 ^ n4419 ;
  assign n4417 = n3660 ^ n3632 ;
  assign n4418 = n4417 ^ n3601 ;
  assign n4422 = n4421 ^ n4418 ;
  assign n4423 = n4422 ^ n3677 ;
  assign n4415 = n3708 ^ n3683 ;
  assign n4416 = n4415 ^ n3667 ;
  assign n4424 = n4423 ^ n4416 ;
  assign n4425 = n4423 ^ n3569 ;
  assign n4426 = n4425 ^ n4423 ;
  assign n4427 = ~n4424 & n4426 ;
  assign n4428 = n4427 ^ n4423 ;
  assign n4429 = ~n3571 & ~n4428 ;
  assign n4457 = n4456 ^ n4429 ;
  assign n4458 = n4457 ^ n3748 ;
  assign n4459 = n4458 ^ n3742 ;
  assign n4460 = n4459 ^ n1464 ;
  assign n4461 = n4460 ^ x123 ;
  assign n4462 = n4414 & ~n4461 ;
  assign n4089 = n2593 ^ x86 ;
  assign n4090 = n3401 ^ x68 ;
  assign n4202 = ~n4089 & ~n4090 ;
  assign n4092 = n2662 ^ x69 ;
  assign n4114 = n3041 ^ n1047 ;
  assign n4115 = n4114 ^ n3957 ;
  assign n4116 = n1184 & n4115 ;
  assign n4106 = n1045 ^ n1035 ;
  assign n4117 = n4116 ^ n4106 ;
  assign n4118 = n3032 & n4117 ;
  assign n4093 = ~n1215 & ~n3032 ;
  assign n4105 = n4093 ^ n1061 ;
  assign n4107 = n4106 ^ n4105 ;
  assign n4108 = n4107 ^ n1202 ;
  assign n4109 = n4108 ^ n1192 ;
  assign n4110 = n4109 ^ n3059 ;
  assign n4111 = n4110 ^ x20 ;
  assign n4098 = n1053 ^ n1042 ;
  assign n4099 = n4098 ^ n3948 ;
  assign n4100 = n4099 ^ n1061 ;
  assign n4096 = n1061 ^ n1054 ;
  assign n4097 = n4096 ^ n3973 ;
  assign n4101 = n4100 ^ n4097 ;
  assign n4102 = n907 & ~n4101 ;
  assign n4103 = n4102 ^ n4100 ;
  assign n4104 = ~n1184 & ~n4103 ;
  assign n4112 = n4111 ^ n4104 ;
  assign n4094 = n907 & n1044 ;
  assign n4095 = n4093 & n4094 ;
  assign n4113 = n4112 ^ n4095 ;
  assign n4119 = n4118 ^ n4113 ;
  assign n4120 = n4119 ^ x75 ;
  assign n4121 = n4092 & n4120 ;
  assign n4122 = n4121 ^ n4092 ;
  assign n4182 = n4122 ^ n4120 ;
  assign n4123 = n3493 ^ x125 ;
  assign n4155 = n683 & n796 ;
  assign n4152 = n688 & ~n834 ;
  assign n4141 = n695 ^ n693 ;
  assign n4150 = n831 & n4141 ;
  assign n4139 = n684 ^ n677 ;
  assign n4140 = n4139 ^ n703 ;
  assign n4142 = n4141 ^ n4140 ;
  assign n4143 = n833 & ~n4142 ;
  assign n4132 = n692 ^ n681 ;
  assign n4135 = n4132 ^ n699 ;
  assign n4136 = n830 & ~n4135 ;
  assign n4137 = n4136 ^ n835 ;
  assign n4133 = n4132 ^ n677 ;
  assign n4134 = ~n834 & ~n4133 ;
  assign n4138 = n4137 ^ n4134 ;
  assign n4144 = n4143 ^ n4138 ;
  assign n4126 = n3090 ^ n805 ;
  assign n4129 = ~n796 & n4126 ;
  assign n4130 = n4129 ^ n3090 ;
  assign n4131 = n322 & n4130 ;
  assign n4145 = n4144 ^ n4131 ;
  assign n4146 = n4145 ^ n832 ;
  assign n4147 = n4146 ^ n843 ;
  assign n4148 = n4147 ^ n3079 ;
  assign n4149 = n4148 ^ x12 ;
  assign n4151 = n4150 ^ n4149 ;
  assign n4153 = n4152 ^ n4151 ;
  assign n4124 = n700 ^ n683 ;
  assign n4125 = ~n322 & n4124 ;
  assign n4154 = n4153 ^ n4125 ;
  assign n4156 = n4155 ^ n4154 ;
  assign n4157 = n4156 ^ x92 ;
  assign n4158 = n4123 & ~n4157 ;
  assign n4159 = n4158 ^ n4157 ;
  assign n4183 = n4159 ^ n4123 ;
  assign n4184 = ~n4182 & n4183 ;
  assign n4164 = n4121 ^ n4120 ;
  assign n4176 = n4158 & n4164 ;
  assign n4177 = n4176 ^ n4158 ;
  assign n4168 = n4157 ^ n4123 ;
  assign n4169 = n4120 ^ n4092 ;
  assign n4173 = n4169 ^ n4157 ;
  assign n4170 = n4169 ^ n4123 ;
  assign n4171 = n4170 ^ n4157 ;
  assign n4172 = n4092 & ~n4171 ;
  assign n4174 = n4173 ^ n4172 ;
  assign n4175 = n4168 & ~n4174 ;
  assign n4178 = n4177 ^ n4175 ;
  assign n4179 = n4178 ^ n4176 ;
  assign n4165 = n4158 ^ n4123 ;
  assign n4166 = n4164 & n4165 ;
  assign n4167 = n4166 ^ n4164 ;
  assign n4180 = n4179 ^ n4167 ;
  assign n4161 = n4121 & ~n4159 ;
  assign n4160 = n4122 & ~n4159 ;
  assign n4162 = n4161 ^ n4160 ;
  assign n4163 = n4162 ^ n4159 ;
  assign n4181 = n4180 ^ n4163 ;
  assign n4213 = n4184 ^ n4181 ;
  assign n4186 = n4158 & ~n4182 ;
  assign n4212 = n4186 ^ n4182 ;
  assign n4214 = n4213 ^ n4212 ;
  assign n4498 = n4214 ^ n4179 ;
  assign n4499 = n4202 & n4498 ;
  assign n4215 = n4214 ^ n4180 ;
  assign n4480 = n4215 ^ n4184 ;
  assign n4481 = n4480 ^ n4186 ;
  assign n4196 = n4121 & n4158 ;
  assign n4221 = n4196 ^ n4121 ;
  assign n4191 = n4121 & n4165 ;
  assign n4192 = n4191 ^ n4161 ;
  assign n4222 = n4221 ^ n4192 ;
  assign n4478 = n4222 ^ n4196 ;
  assign n4190 = n4122 & n4183 ;
  assign n4477 = n4191 ^ n4190 ;
  assign n4479 = n4478 ^ n4477 ;
  assign n4482 = n4481 ^ n4479 ;
  assign n4483 = ~n4090 & n4482 ;
  assign n4484 = n4483 ^ n4481 ;
  assign n4494 = n4484 ^ n1347 ;
  assign n4488 = n4196 ^ n4181 ;
  assign n4489 = n4196 ^ n4090 ;
  assign n4490 = n4489 ^ n4196 ;
  assign n4491 = ~n4488 & ~n4490 ;
  assign n4492 = n4491 ^ n4196 ;
  assign n4493 = ~n4089 & n4492 ;
  assign n4495 = n4494 ^ n4493 ;
  assign n4485 = n4484 ^ n4179 ;
  assign n4185 = n4184 ^ n4166 ;
  assign n4207 = n4202 ^ n4089 ;
  assign n4208 = n4207 ^ n4090 ;
  assign n4209 = ~n4185 & n4208 ;
  assign n4474 = n4186 ^ n4181 ;
  assign n4226 = n4208 ^ n4089 ;
  assign n4475 = n4474 ^ n4226 ;
  assign n4476 = ~n4209 & n4475 ;
  assign n4486 = n4485 ^ n4476 ;
  assign n4487 = n4089 & n4486 ;
  assign n4496 = n4495 ^ n4487 ;
  assign n4091 = n4090 ^ n4089 ;
  assign n4473 = n4091 & n4162 ;
  assign n4497 = n4496 ^ n4473 ;
  assign n4500 = n4499 ^ n4497 ;
  assign n4472 = n4172 & ~n4208 ;
  assign n4501 = n4500 ^ n4472 ;
  assign n4193 = n4192 ^ n4190 ;
  assign n4194 = n4193 ^ n4172 ;
  assign n4465 = n4194 ^ n4191 ;
  assign n4219 = n4160 ^ n4122 ;
  assign n4195 = n4194 ^ n4190 ;
  assign n4220 = n4219 ^ n4195 ;
  assign n4466 = n4465 ^ n4220 ;
  assign n4467 = n4220 ^ n4090 ;
  assign n4468 = n4467 ^ n4220 ;
  assign n4469 = n4466 & ~n4468 ;
  assign n4470 = n4469 ^ n4220 ;
  assign n4471 = n4091 & n4470 ;
  assign n4502 = n4501 ^ n4471 ;
  assign n4503 = n4502 ^ x113 ;
  assign n4504 = n851 & ~n2224 ;
  assign n4520 = n4504 ^ n1294 ;
  assign n4518 = n2248 ^ n1248 ;
  assign n3901 = ~n2201 & ~n2210 ;
  assign n4508 = n3901 ^ n2218 ;
  assign n4509 = ~n851 & ~n4508 ;
  assign n4510 = n4509 ^ n2218 ;
  assign n4519 = n4518 ^ n4510 ;
  assign n4521 = n4520 ^ n4519 ;
  assign n4507 = n1248 ^ n851 ;
  assign n4511 = n4510 ^ n1248 ;
  assign n4512 = n4511 ^ n4510 ;
  assign n4513 = n4510 ^ n2225 ;
  assign n4514 = n4513 ^ n4510 ;
  assign n4515 = ~n4512 & ~n4514 ;
  assign n4516 = n4515 ^ n4510 ;
  assign n4517 = ~n4507 & ~n4516 ;
  assign n4522 = n4521 ^ n4517 ;
  assign n3902 = n2235 ^ n2229 ;
  assign n4505 = n1248 & n3902 ;
  assign n4506 = n4504 & n4505 ;
  assign n4523 = n4522 ^ n4506 ;
  assign n4524 = n4523 ^ x114 ;
  assign n4525 = n4503 & ~n4524 ;
  assign n4570 = n4525 ^ n4503 ;
  assign n4642 = n4570 ^ n4524 ;
  assign n4669 = n4462 & n4642 ;
  assign n4463 = n4462 ^ n4461 ;
  assign n4526 = n4525 ^ n4524 ;
  assign n4668 = ~n4463 & ~n4526 ;
  assign n4670 = n4669 ^ n4668 ;
  assign n4464 = n4463 ^ n4414 ;
  assign n4565 = n4464 & n4525 ;
  assign n4693 = n4670 ^ n4565 ;
  assign n4562 = n2708 ^ n1537 ;
  assign n4242 = n2716 ^ n2692 ;
  assign n4243 = ~n2252 & n4242 ;
  assign n4244 = n4243 ^ n2692 ;
  assign n4246 = n4244 ^ n2684 ;
  assign n4245 = n4244 ^ n2695 ;
  assign n4247 = n4246 ^ n4245 ;
  assign n4250 = ~n2252 & ~n4247 ;
  assign n4251 = n4250 ^ n4246 ;
  assign n4252 = n2663 & n4251 ;
  assign n4253 = n4252 ^ n4244 ;
  assign n4555 = n2720 ^ n2602 ;
  assign n4537 = n2679 ^ n2608 ;
  assign n4536 = n2700 ^ n2687 ;
  assign n4538 = n4537 ^ n4536 ;
  assign n4254 = n2678 ^ n2673 ;
  assign n4255 = n4254 ^ n2602 ;
  assign n4539 = n4538 ^ n4255 ;
  assign n4540 = n2663 & ~n4539 ;
  assign n4541 = n4540 ^ n2700 ;
  assign n4556 = n4555 ^ n4541 ;
  assign n4557 = n4556 ^ n2715 ;
  assign n4549 = n2680 ^ n2673 ;
  assign n4550 = n2673 ^ n2663 ;
  assign n4551 = n4550 ^ n2673 ;
  assign n4552 = ~n4549 & n4551 ;
  assign n4553 = n4552 ^ n2673 ;
  assign n4554 = n2252 & n4553 ;
  assign n4558 = n4557 ^ n4554 ;
  assign n4535 = n2663 ^ n2252 ;
  assign n4544 = n4541 ^ n2252 ;
  assign n4545 = n4544 ^ n4541 ;
  assign n4546 = ~n2679 & n4545 ;
  assign n4547 = n4546 ^ n4541 ;
  assign n4548 = ~n4535 & ~n4547 ;
  assign n4559 = n4558 ^ n4548 ;
  assign n4528 = n2670 ^ n2602 ;
  assign n4259 = n2683 ^ n2597 ;
  assign n4260 = n4259 ^ n2673 ;
  assign n4529 = n4260 ^ n2697 ;
  assign n4530 = n2697 ^ n2602 ;
  assign n4531 = n4530 ^ n2697 ;
  assign n4532 = ~n4529 & ~n4531 ;
  assign n4533 = n4532 ^ n2697 ;
  assign n4534 = ~n4528 & ~n4533 ;
  assign n4560 = n4559 ^ n4534 ;
  assign n4561 = ~n4253 & n4560 ;
  assign n4563 = n4562 ^ n4561 ;
  assign n4564 = n4563 ^ x120 ;
  assign n4694 = n4565 ^ n4564 ;
  assign n4695 = n4694 ^ n4565 ;
  assign n4696 = n4693 & n4695 ;
  assign n4697 = n4696 ^ n4565 ;
  assign n4698 = ~n4634 & n4697 ;
  assign n4566 = n4464 ^ n4461 ;
  assign n4571 = n4566 & n4570 ;
  assign n4569 = ~n4526 & n4566 ;
  assign n4572 = n4571 ^ n4569 ;
  assign n4567 = n4525 & n4566 ;
  assign n4568 = n4567 ^ n4566 ;
  assign n4573 = n4572 ^ n4568 ;
  assign n4655 = n4564 & ~n4634 ;
  assign n4656 = n4655 ^ n4564 ;
  assign n4664 = n4656 ^ n4634 ;
  assign n4665 = n4664 ^ n4564 ;
  assign n5375 = n4573 & ~n4665 ;
  assign n4662 = n4634 ^ n4564 ;
  assign n4658 = n4567 ^ n4565 ;
  assign n4638 = n4462 & n4525 ;
  assign n4657 = n4638 ^ n4525 ;
  assign n4659 = n4658 ^ n4657 ;
  assign n4643 = n4464 & n4642 ;
  assign n4666 = n4659 ^ n4643 ;
  assign n4527 = n4464 & ~n4526 ;
  assign n4644 = n4643 ^ n4527 ;
  assign n4641 = n4565 ^ n4464 ;
  assign n4645 = n4644 ^ n4641 ;
  assign n5369 = n4666 ^ n4645 ;
  assign n5367 = n4571 ^ n4527 ;
  assign n5368 = n5367 ^ n4567 ;
  assign n5370 = n5369 ^ n5368 ;
  assign n5371 = ~n4634 & n5370 ;
  assign n4646 = n4645 ^ n4571 ;
  assign n4636 = n4462 & ~n4503 ;
  assign n4637 = n4636 ^ n4462 ;
  assign n4639 = n4638 ^ n4637 ;
  assign n4640 = n4639 ^ n4570 ;
  assign n4647 = n4646 ^ n4640 ;
  assign n4648 = n4647 ^ n4638 ;
  assign n5358 = n4670 ^ n4648 ;
  assign n5364 = n5358 ^ n4461 ;
  assign n5372 = n5371 ^ n5364 ;
  assign n5373 = n4662 & ~n5372 ;
  assign n5361 = n4569 ^ n4566 ;
  assign n5362 = n5361 ^ n4645 ;
  assign n5357 = n4641 ^ n4571 ;
  assign n5359 = n5358 ^ n5357 ;
  assign n5360 = n4664 & n5359 ;
  assign n5363 = n5362 ^ n5360 ;
  assign n5365 = n5364 ^ n5363 ;
  assign n4681 = n4645 ^ n4569 ;
  assign n5352 = n4566 ^ n4564 ;
  assign n5353 = n5352 ^ n4566 ;
  assign n5354 = n4681 & n5353 ;
  assign n5355 = n5354 ^ n4566 ;
  assign n5356 = ~n4634 & n5355 ;
  assign n5366 = n5365 ^ n5356 ;
  assign n5374 = n5373 ^ n5366 ;
  assign n5376 = n5375 ^ n5374 ;
  assign n5377 = ~n4698 & n5376 ;
  assign n5378 = n5377 ^ n3493 ;
  assign n5379 = n5378 ^ x68 ;
  assign n5768 = ~n5349 & n5379 ;
  assign n5769 = n5768 ^ n5379 ;
  assign n4197 = n4196 ^ n4195 ;
  assign n4187 = n4186 ^ n4180 ;
  assign n4188 = n4187 ^ n4185 ;
  assign n4189 = n4188 ^ n4161 ;
  assign n4198 = n4197 ^ n4189 ;
  assign n4199 = ~n4090 & n4198 ;
  assign n4200 = n4199 ^ n4188 ;
  assign n4238 = n4200 ^ n669 ;
  assign n4203 = n4181 ^ n4178 ;
  assign n4210 = n4203 & n4209 ;
  assign n4205 = n4197 ^ n4178 ;
  assign n4206 = ~n4202 & ~n4205 ;
  assign n4211 = n4210 ^ n4206 ;
  assign n4239 = n4238 ^ n4211 ;
  assign n4235 = ~n4090 & ~n4213 ;
  assign n4228 = n4220 ^ n4160 ;
  assign n4227 = n4191 ^ n4178 ;
  assign n4229 = n4228 ^ n4227 ;
  assign n4230 = n4226 & ~n4229 ;
  assign n4223 = n4207 & ~n4222 ;
  assign n4224 = ~n4192 & n4223 ;
  assign n4225 = ~n4220 & n4224 ;
  assign n4231 = n4230 ^ n4225 ;
  assign n4216 = n4215 ^ n4176 ;
  assign n4232 = n4231 ^ n4216 ;
  assign n4233 = n4232 ^ n4211 ;
  assign n4201 = n4200 ^ n4181 ;
  assign n4234 = n4233 ^ n4201 ;
  assign n4236 = n4235 ^ n4234 ;
  assign n4237 = n4091 & ~n4236 ;
  assign n4240 = n4239 ^ n4237 ;
  assign n5098 = n4240 ^ x121 ;
  assign n5099 = n4460 ^ x65 ;
  assign n5100 = ~n5098 & ~n5099 ;
  assign n5176 = n5100 ^ n5099 ;
  assign n5101 = n4563 ^ x107 ;
  assign n5131 = n3542 ^ n1893 ;
  assign n5120 = n3515 ^ n3503 ;
  assign n5121 = n3536 ^ n3517 ;
  assign n5122 = n5120 & n5121 ;
  assign n5117 = n3434 ^ n3426 ;
  assign n5118 = n5117 ^ n3436 ;
  assign n5119 = n3504 & n5118 ;
  assign n5123 = n5122 ^ n5119 ;
  assign n5110 = n3464 ^ n3421 ;
  assign n3880 = n3514 ^ n3511 ;
  assign n3881 = n3880 ^ n3506 ;
  assign n5109 = n3881 ^ n3465 ;
  assign n5111 = n5110 ^ n5109 ;
  assign n5112 = n5109 ^ n3494 ;
  assign n5113 = n5112 ^ n5109 ;
  assign n5114 = ~n5111 & ~n5113 ;
  assign n5115 = n5114 ^ n5109 ;
  assign n5116 = ~n3320 & ~n5115 ;
  assign n5124 = n5123 ^ n5116 ;
  assign n5125 = n3438 ^ n3429 ;
  assign n5128 = ~n3504 & n5125 ;
  assign n5129 = n5128 ^ n3438 ;
  assign n5130 = ~n5124 & ~n5129 ;
  assign n5132 = n5131 ^ n5130 ;
  assign n3878 = n3465 ^ n3431 ;
  assign n5104 = n3506 ^ n3494 ;
  assign n5105 = n5104 ^ n3506 ;
  assign n5106 = n3878 & ~n5105 ;
  assign n5107 = n5106 ^ n3506 ;
  assign n5108 = n3320 & n5107 ;
  assign n5133 = n5132 ^ n5108 ;
  assign n5134 = n5133 ^ x97 ;
  assign n3865 = ~n3246 & ~n3258 ;
  assign n3861 = n3279 ^ n3277 ;
  assign n3862 = n3201 & n3861 ;
  assign n3852 = n3243 ^ n3157 ;
  assign n3853 = n3852 ^ n3305 ;
  assign n3851 = n3236 ^ n3227 ;
  assign n3854 = n3853 ^ n3851 ;
  assign n3855 = n3854 ^ n3277 ;
  assign n3849 = n3277 ^ n3209 ;
  assign n3850 = n3849 ^ n3212 ;
  assign n3856 = n3855 ^ n3850 ;
  assign n3857 = ~n3201 & n3856 ;
  assign n3858 = n3857 ^ n3855 ;
  assign n3859 = n3004 & ~n3858 ;
  assign n3844 = n3207 & ~n3307 ;
  assign n3845 = n3844 ^ n3291 ;
  assign n3841 = n3207 & ~n3233 ;
  assign n3842 = n3841 ^ n3277 ;
  assign n3843 = n3842 ^ n3206 ;
  assign n3846 = n3845 ^ n3843 ;
  assign n3840 = n3247 & ~n3258 ;
  assign n3847 = n3846 ^ n3840 ;
  assign n3848 = n3847 ^ n795 ;
  assign n3860 = n3859 ^ n3848 ;
  assign n3863 = n3862 ^ n3860 ;
  assign n3839 = n3207 & n3235 ;
  assign n3864 = n3863 ^ n3839 ;
  assign n3866 = n3865 ^ n3864 ;
  assign n5135 = n3866 ^ x80 ;
  assign n5159 = n2955 ^ n2915 ;
  assign n5160 = n5159 ^ n2940 ;
  assign n5156 = n2920 ^ n2911 ;
  assign n5154 = n2914 ^ n2904 ;
  assign n5155 = n5154 ^ n2909 ;
  assign n5157 = n5156 ^ n5155 ;
  assign n5148 = n2930 ^ n2909 ;
  assign n5149 = n5148 ^ n2955 ;
  assign n5150 = ~n2797 & n5149 ;
  assign n5145 = n2977 ^ n2941 ;
  assign n5146 = n5145 ^ n2966 ;
  assign n5147 = n5146 ^ n2931 ;
  assign n5151 = n5150 ^ n5147 ;
  assign n5158 = n5157 ^ n5151 ;
  assign n5161 = n5160 ^ n5158 ;
  assign n5162 = n5161 ^ n5151 ;
  assign n5163 = n2797 & ~n5162 ;
  assign n5164 = n5163 ^ n5158 ;
  assign n5165 = ~n2798 & n5164 ;
  assign n5152 = n5151 ^ n2985 ;
  assign n5138 = n2949 ^ n2797 ;
  assign n5139 = n5138 ^ n2949 ;
  assign n5142 = ~n2950 & n5139 ;
  assign n5143 = n5142 ^ n2949 ;
  assign n5144 = n2798 & ~n5143 ;
  assign n5153 = n5152 ^ n5144 ;
  assign n5166 = n5165 ^ n5153 ;
  assign n4970 = n2911 & ~n2924 ;
  assign n5167 = n5166 ^ n4970 ;
  assign n5168 = n5167 ^ n1931 ;
  assign n5169 = n5168 ^ x90 ;
  assign n5170 = n5135 & ~n5169 ;
  assign n5171 = n5134 & n5170 ;
  assign n5231 = n5101 & n5171 ;
  assign n5254 = n5231 ^ n5171 ;
  assign n5260 = ~n5176 & n5254 ;
  assign n5261 = n5260 ^ n3200 ;
  assign n5136 = n5134 & ~n5135 ;
  assign n5137 = n5136 ^ n5134 ;
  assign n5172 = n5171 ^ n5137 ;
  assign n5173 = ~n5101 & n5172 ;
  assign n5174 = n5173 ^ n5172 ;
  assign n5175 = n5100 & n5174 ;
  assign n5177 = n5176 ^ n5098 ;
  assign n5178 = n5177 ^ n5099 ;
  assign n5255 = n5254 ^ n5174 ;
  assign n5256 = ~n5178 & n5255 ;
  assign n5189 = ~n5101 & n5136 ;
  assign n5197 = n5189 ^ n5136 ;
  assign n5182 = ~n5101 & ~n5134 ;
  assign n5183 = ~n5135 & n5182 ;
  assign n5193 = ~n5169 & n5183 ;
  assign n5194 = n5193 ^ n5183 ;
  assign n5190 = n5169 & n5189 ;
  assign n5191 = n5190 ^ n5189 ;
  assign n5185 = n5136 ^ n5135 ;
  assign n5186 = n5185 ^ n5183 ;
  assign n5187 = ~n5169 & ~n5186 ;
  assign n5188 = n5187 ^ n5186 ;
  assign n5192 = n5191 ^ n5188 ;
  assign n5195 = n5194 ^ n5192 ;
  assign n5180 = n5169 ^ n5101 ;
  assign n5181 = ~n5135 & ~n5180 ;
  assign n5184 = n5183 ^ n5181 ;
  assign n5196 = n5195 ^ n5184 ;
  assign n5198 = n5197 ^ n5196 ;
  assign n5250 = n5198 ^ n5194 ;
  assign n5251 = ~n5178 & ~n5250 ;
  assign n5244 = n5189 ^ n5186 ;
  assign n5245 = ~n5177 & n5244 ;
  assign n5235 = n5191 ^ n5187 ;
  assign n5234 = n5192 ^ n5181 ;
  assign n5238 = n5234 ^ n5099 ;
  assign n5239 = n5238 ^ n5234 ;
  assign n5240 = ~n5235 & ~n5239 ;
  assign n5241 = n5240 ^ n5234 ;
  assign n5242 = ~n5098 & n5241 ;
  assign n5243 = n5242 ^ n5099 ;
  assign n5246 = n5245 ^ n5243 ;
  assign n5179 = n5178 ^ n5176 ;
  assign n5199 = n5170 ^ n5135 ;
  assign n5201 = n5182 & n5199 ;
  assign n5232 = n5231 ^ n5201 ;
  assign n5233 = ~n5179 & n5232 ;
  assign n5247 = n5246 ^ n5233 ;
  assign n5211 = n5201 ^ n5182 ;
  assign n5212 = n5211 ^ n5183 ;
  assign n5200 = n5199 ^ n5172 ;
  assign n5202 = n5201 ^ n5200 ;
  assign n5223 = n5212 ^ n5202 ;
  assign n5221 = n5190 ^ n5188 ;
  assign n5222 = n5221 ^ n5173 ;
  assign n5224 = n5223 ^ n5222 ;
  assign n5225 = n5224 ^ n5173 ;
  assign n5226 = n5173 ^ n5099 ;
  assign n5227 = n5226 ^ n5173 ;
  assign n5228 = ~n5225 & ~n5227 ;
  assign n5229 = n5228 ^ n5173 ;
  assign n5230 = n5098 & n5229 ;
  assign n5248 = n5247 ^ n5230 ;
  assign n5210 = n5171 ^ n5170 ;
  assign n5213 = n5212 ^ n5210 ;
  assign n5249 = n5248 ^ n5213 ;
  assign n5252 = n5251 ^ n5249 ;
  assign n5214 = n5213 ^ n5099 ;
  assign n5215 = n5214 ^ n5213 ;
  assign n5216 = n5213 ^ n5194 ;
  assign n5217 = n5216 ^ n5213 ;
  assign n5218 = ~n5215 & n5217 ;
  assign n5219 = n5218 ^ n5213 ;
  assign n5220 = ~n5098 & n5219 ;
  assign n5253 = n5252 ^ n5220 ;
  assign n5257 = n5256 ^ n5253 ;
  assign n5203 = n5202 ^ n5173 ;
  assign n5204 = n5203 ^ n5198 ;
  assign n5205 = n5203 ^ n5098 ;
  assign n5206 = n5205 ^ n5203 ;
  assign n5207 = ~n5204 & n5206 ;
  assign n5208 = n5207 ^ n5203 ;
  assign n5209 = n5179 & n5208 ;
  assign n5258 = n5257 ^ n5209 ;
  assign n5259 = ~n5175 & ~n5258 ;
  assign n5262 = n5261 ^ n5259 ;
  assign n5554 = n5262 ^ x85 ;
  assign n4759 = n4000 ^ n3985 ;
  assign n4760 = n4759 ^ n3922 ;
  assign n4013 = n4012 ^ n4008 ;
  assign n4761 = n4013 ^ n3924 ;
  assign n4764 = ~n4759 & n4761 ;
  assign n4765 = n4764 ^ n3924 ;
  assign n4766 = n4760 & n4765 ;
  assign n4752 = n4029 ^ n3991 ;
  assign n4753 = n4752 ^ n4039 ;
  assign n4757 = ~n3923 & n4753 ;
  assign n4754 = n4616 ^ n3920 ;
  assign n4758 = n4757 ^ n4754 ;
  assign n4767 = n4766 ^ n4758 ;
  assign n4747 = n4035 ^ n3921 ;
  assign n4748 = n4747 ^ n4035 ;
  assign n4749 = ~n4037 & ~n4748 ;
  assign n4750 = n4749 ^ n4035 ;
  assign n4751 = n3920 & n4750 ;
  assign n4768 = n4767 ^ n4751 ;
  assign n4769 = n4768 ^ n4080 ;
  assign n4066 = n4065 ^ n4038 ;
  assign n4015 = n4014 ^ n4013 ;
  assign n4067 = n4066 ^ n4015 ;
  assign n4068 = n4015 ^ n3920 ;
  assign n4069 = n4068 ^ n4015 ;
  assign n4070 = ~n4067 & n4069 ;
  assign n4071 = n4070 ^ n4015 ;
  assign n4072 = n3921 & ~n4071 ;
  assign n4770 = n4769 ^ n4072 ;
  assign n4771 = n4770 ^ n4582 ;
  assign n4016 = n3924 & ~n4015 ;
  assign n4772 = n4771 ^ n4016 ;
  assign n4050 = n4008 & n4049 ;
  assign n4773 = n4772 ^ n4050 ;
  assign n4774 = n4773 ^ n953 ;
  assign n5556 = n4774 ^ x68 ;
  assign n3914 = n2203 & n2246 ;
  assign n3903 = n3902 ^ n3901 ;
  assign n3904 = n851 & n3903 ;
  assign n3905 = n3904 ^ n3902 ;
  assign n3915 = n3914 ^ n3905 ;
  assign n3907 = n3905 ^ n2218 ;
  assign n3906 = n3905 ^ n2221 ;
  assign n3908 = n3907 ^ n3906 ;
  assign n3911 = n851 & n3908 ;
  assign n3912 = n3911 ^ n3907 ;
  assign n3913 = ~n1248 & n3912 ;
  assign n3916 = n3915 ^ n3913 ;
  assign n3917 = ~n2224 & ~n3916 ;
  assign n3918 = n3917 ^ n344 ;
  assign n5557 = n3918 ^ x117 ;
  assign n5558 = n5556 & ~n5557 ;
  assign n5559 = n5558 ^ n5556 ;
  assign n5560 = n5559 ^ n5557 ;
  assign n5581 = n4970 ^ n2095 ;
  assign n5575 = n5146 ^ n2923 ;
  assign n5576 = n2917 & ~n5575 ;
  assign n5571 = n5155 ^ n2954 ;
  assign n5572 = ~n2925 & n5571 ;
  assign n5569 = n2934 ^ n2917 ;
  assign n5570 = ~n2919 & n5569 ;
  assign n5573 = n5572 ^ n5570 ;
  assign n5574 = n5573 ^ n2929 ;
  assign n5577 = n5576 ^ n5574 ;
  assign n5561 = n2977 ^ n2967 ;
  assign n5562 = n5561 ^ n2914 ;
  assign n5563 = n5562 ^ n2967 ;
  assign n5564 = n2967 ^ n2752 ;
  assign n5565 = n5564 ^ n2967 ;
  assign n5566 = n5563 & n5565 ;
  assign n5567 = n5566 ^ n2967 ;
  assign n5568 = n2797 & ~n5567 ;
  assign n5578 = n5577 ^ n5568 ;
  assign n5579 = n2963 & n5578 ;
  assign n5580 = ~n5144 & n5579 ;
  assign n5582 = n5581 ^ n5580 ;
  assign n5583 = n5582 ^ x67 ;
  assign n4728 = n4166 ^ n4160 ;
  assign n4729 = n4728 ^ n4478 ;
  assign n4727 = n4194 ^ n4187 ;
  assign n4730 = n4729 ^ n4727 ;
  assign n4731 = ~n4090 & n4730 ;
  assign n4732 = n4731 ^ n4727 ;
  assign n4733 = ~n4089 & n4732 ;
  assign n4723 = n4215 ^ n4181 ;
  assign n4724 = ~n4226 & ~n4723 ;
  assign n4707 = ~n4195 & n4223 ;
  assign n4709 = ~n4193 & n4208 ;
  assign n4710 = ~n4707 & n4709 ;
  assign n4708 = n4707 ^ n4220 ;
  assign n4711 = n4710 ^ n4708 ;
  assign n4720 = n4711 ^ n906 ;
  assign n4713 = n4711 ^ n4182 ;
  assign n4712 = n4711 ^ n4172 ;
  assign n4714 = n4713 ^ n4712 ;
  assign n4715 = n4713 ^ n4089 ;
  assign n4716 = n4715 ^ n4713 ;
  assign n4717 = ~n4714 & n4716 ;
  assign n4718 = n4717 ^ n4713 ;
  assign n4719 = ~n4090 & n4718 ;
  assign n4721 = n4720 ^ n4719 ;
  assign n4704 = n4123 ^ n4120 ;
  assign n4705 = ~n4092 & ~n4208 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4722 = n4721 ^ n4706 ;
  assign n4725 = n4724 ^ n4722 ;
  assign n4703 = n4091 & n4178 ;
  assign n4726 = n4725 ^ n4703 ;
  assign n4734 = n4733 ^ n4726 ;
  assign n5584 = n4734 ^ x100 ;
  assign n5585 = ~n5583 & n5584 ;
  assign n5586 = n5585 ^ n5583 ;
  assign n3892 = n3441 ^ n3436 ;
  assign n3877 = n3536 ^ n3440 ;
  assign n3883 = n3463 ^ n3430 ;
  assign n3884 = n3883 ^ n3514 ;
  assign n3885 = n3884 ^ n3878 ;
  assign n3886 = ~n3494 & ~n3885 ;
  assign n3879 = n3878 ^ n3877 ;
  assign n3882 = n3881 ^ n3879 ;
  assign n3887 = n3886 ^ n3882 ;
  assign n3888 = ~n3877 & n3887 ;
  assign n3889 = n3320 & n3888 ;
  assign n3893 = ~n3494 & n3889 ;
  assign n3894 = n3892 & n3893 ;
  assign n3890 = n3889 ^ n3320 ;
  assign n3876 = n3535 ^ n321 ;
  assign n3891 = n3890 ^ n3876 ;
  assign n3895 = n3894 ^ n3891 ;
  assign n3896 = n3895 ^ n3421 ;
  assign n3875 = ~n3320 & n3459 ;
  assign n3897 = n3896 ^ n3875 ;
  assign n3868 = n3535 ^ n3421 ;
  assign n3869 = n3868 ^ n3456 ;
  assign n3870 = n3869 ^ n3535 ;
  assign n3871 = n3870 ^ n3454 ;
  assign n3872 = ~n3320 & n3871 ;
  assign n3873 = n3872 ^ n3868 ;
  assign n3874 = ~n3494 & n3873 ;
  assign n3898 = n3897 ^ n3874 ;
  assign n5587 = n3898 ^ x78 ;
  assign n5607 = n3742 ^ n3691 ;
  assign n5608 = n5607 ^ n3673 ;
  assign n5609 = n5608 ^ n2070 ;
  assign n5602 = n4420 ^ n3681 ;
  assign n5603 = n5602 ^ n3729 ;
  assign n5604 = ~n3569 & n5603 ;
  assign n5605 = n5604 ^ n3691 ;
  assign n5606 = ~n3570 & ~n5605 ;
  assign n5610 = n5609 ^ n5606 ;
  assign n5595 = n4436 ^ n3683 ;
  assign n5596 = n5595 ^ n3676 ;
  assign n5597 = n5596 ^ n4436 ;
  assign n5598 = n5597 ^ n3718 ;
  assign n5599 = n3569 & ~n5598 ;
  assign n5600 = n5599 ^ n5595 ;
  assign n5601 = n3571 & ~n5600 ;
  assign n5611 = n5610 ^ n5601 ;
  assign n5588 = n4453 ^ n3674 ;
  assign n5589 = n5588 ^ n3706 ;
  assign n5590 = n5589 ^ n3734 ;
  assign n5591 = ~n3687 & ~n5590 ;
  assign n5592 = n5591 ^ n3706 ;
  assign n5593 = n3705 ^ n3687 ;
  assign n5594 = ~n5592 & ~n5593 ;
  assign n5612 = n5611 ^ n5594 ;
  assign n5613 = n5612 ^ x85 ;
  assign n5614 = ~n5587 & ~n5613 ;
  assign n5615 = n5614 ^ n5587 ;
  assign n5616 = n5615 ^ n5613 ;
  assign n5617 = ~n5586 & ~n5616 ;
  assign n5618 = n5560 & n5617 ;
  assign n5637 = n5585 & n5614 ;
  assign n5619 = n5614 ^ n5613 ;
  assign n5627 = n5584 & ~n5619 ;
  assign n5628 = n5583 & n5627 ;
  assign n5677 = n5637 ^ n5628 ;
  assign n5620 = n5587 ^ n5583 ;
  assign n5621 = n5587 ^ n5584 ;
  assign n5622 = n5620 & n5621 ;
  assign n5630 = n5622 ^ n5587 ;
  assign n5631 = n5620 ^ n5613 ;
  assign n5632 = ~n5630 & ~n5631 ;
  assign n5638 = n5637 ^ n5632 ;
  assign n5635 = ~n5586 & n5614 ;
  assign n5636 = n5635 ^ n5617 ;
  assign n5639 = n5638 ^ n5636 ;
  assign n5624 = n5586 ^ n5584 ;
  assign n5634 = n5614 & n5624 ;
  assign n5640 = n5639 ^ n5634 ;
  assign n5641 = n5640 ^ n5617 ;
  assign n5633 = n5632 ^ n5614 ;
  assign n5642 = n5641 ^ n5633 ;
  assign n5629 = n5628 ^ n5627 ;
  assign n5643 = n5642 ^ n5629 ;
  assign n5625 = n5624 ^ n5583 ;
  assign n5626 = ~n5615 & n5625 ;
  assign n5644 = n5643 ^ n5626 ;
  assign n5645 = n5644 ^ n5628 ;
  assign n5646 = n5645 ^ n5617 ;
  assign n5623 = n5622 ^ n5619 ;
  assign n5647 = n5646 ^ n5623 ;
  assign n5648 = n5647 ^ n5619 ;
  assign n5649 = n5648 ^ n5627 ;
  assign n5650 = n5649 ^ n5641 ;
  assign n5651 = n5650 ^ n5620 ;
  assign n5652 = n5651 ^ n5644 ;
  assign n5696 = n5677 ^ n5652 ;
  assign n5683 = n5627 ^ n5625 ;
  assign n5695 = n5683 ^ n5584 ;
  assign n5697 = n5696 ^ n5695 ;
  assign n5698 = n5697 ^ n5629 ;
  assign n5699 = n5560 & n5698 ;
  assign n5684 = n5683 ^ n5644 ;
  assign n5685 = n5684 ^ n5635 ;
  assign n5686 = n5685 ^ n5649 ;
  assign n5687 = n5686 ^ n5642 ;
  assign n5688 = n5687 ^ n5634 ;
  assign n5666 = n5647 ^ n5624 ;
  assign n5667 = n5666 ^ n5640 ;
  assign n5682 = n5667 ^ n5626 ;
  assign n5689 = n5688 ^ n5682 ;
  assign n5668 = n5649 ^ n5586 ;
  assign n5669 = n5668 ^ n5636 ;
  assign n5678 = n5677 ^ n5669 ;
  assign n5679 = n5678 ^ n5647 ;
  assign n5690 = n5689 ^ n5679 ;
  assign n5691 = ~n5557 & ~n5690 ;
  assign n5670 = n5649 ^ n5647 ;
  assign n5671 = n5670 ^ n5669 ;
  assign n5672 = n5671 ^ n5667 ;
  assign n5664 = n5613 ^ n5584 ;
  assign n5663 = n5650 ^ n5630 ;
  assign n5665 = n5664 ^ n5663 ;
  assign n5673 = n5672 ^ n5665 ;
  assign n5674 = n5557 & n5673 ;
  assign n5675 = n5674 ^ n5672 ;
  assign n5680 = n5679 ^ n5675 ;
  assign n5692 = n5691 ^ n5680 ;
  assign n5693 = ~n5556 & ~n5692 ;
  assign n5661 = n5558 & n5644 ;
  assign n5653 = n5652 ^ n5556 ;
  assign n5654 = n5653 ^ n5652 ;
  assign n5657 = n5639 & ~n5654 ;
  assign n5658 = n5657 ^ n5652 ;
  assign n5659 = n5557 & n5658 ;
  assign n5660 = n5659 ^ n5652 ;
  assign n5662 = n5661 ^ n5660 ;
  assign n5676 = n5675 ^ n5662 ;
  assign n5694 = n5693 ^ n5676 ;
  assign n5700 = n5699 ^ n5694 ;
  assign n5701 = ~n5618 & n5700 ;
  assign n5702 = n5701 ^ n3350 ;
  assign n5703 = n5702 ^ x70 ;
  assign n5704 = n5554 & ~n5703 ;
  assign n5705 = n5704 ^ n5703 ;
  assign n5706 = n5705 ^ n5554 ;
  assign n5055 = n3570 & ~n4420 ;
  assign n5051 = n4432 ^ n3665 ;
  assign n5052 = ~n3705 & ~n5051 ;
  assign n5044 = n4453 ^ n3677 ;
  assign n5041 = n3693 ^ n3675 ;
  assign n5042 = n5041 ^ n4453 ;
  assign n5043 = ~n3569 & n5042 ;
  assign n5045 = n5044 ^ n5043 ;
  assign n5047 = n3703 ^ n3570 ;
  assign n5046 = n3703 ^ n3677 ;
  assign n5048 = n5047 ^ n5046 ;
  assign n5049 = n5045 & ~n5048 ;
  assign n5050 = n5049 ^ n5047 ;
  assign n5053 = n5052 ^ n5050 ;
  assign n5039 = n4436 ^ n3680 ;
  assign n5040 = ~n3706 & n5039 ;
  assign n5054 = n5053 ^ n5040 ;
  assign n5056 = n5055 ^ n5054 ;
  assign n5033 = n3703 ^ n3667 ;
  assign n5034 = n4415 ^ n3569 ;
  assign n5036 = ~n3667 & n5034 ;
  assign n5037 = n5036 ^ n3569 ;
  assign n5038 = n5033 & ~n5037 ;
  assign n5057 = n5056 ^ n5038 ;
  assign n5058 = ~n3748 & n5057 ;
  assign n5059 = ~n3742 & n5058 ;
  assign n5060 = ~n3673 & n5059 ;
  assign n5061 = n5060 ^ n1738 ;
  assign n5062 = n5061 ^ x64 ;
  assign n5006 = n4413 ^ x82 ;
  assign n4901 = n4633 ^ x89 ;
  assign n4966 = n2728 ^ n2527 ;
  assign n4967 = n4966 ^ n2708 ;
  assign n4963 = n2684 & n2697 ;
  assign n4932 = n2722 ^ n2609 ;
  assign n4933 = n2669 & n4932 ;
  assign n4934 = n2698 & ~n4933 ;
  assign n4939 = n4255 & n4537 ;
  assign n4940 = n4939 ^ n2685 ;
  assign n4941 = n4934 & n4940 ;
  assign n4942 = n4941 ^ n4933 ;
  assign n4257 = n2718 ^ n2685 ;
  assign n4931 = ~n2670 & ~n4257 ;
  assign n4943 = n4942 ^ n4931 ;
  assign n4944 = n2702 ^ n2611 ;
  assign n4945 = n4944 ^ n2252 ;
  assign n4946 = n4535 & n4945 ;
  assign n4947 = n4946 ^ n2252 ;
  assign n4950 = n4944 ^ n2691 ;
  assign n4951 = n4947 & ~n4950 ;
  assign n4948 = n2694 ^ n2691 ;
  assign n4952 = n4951 ^ n4948 ;
  assign n4953 = n4952 ^ n2690 ;
  assign n4954 = n4953 ^ n2610 ;
  assign n4955 = n4954 ^ n4952 ;
  assign n4958 = n2252 & n4955 ;
  assign n4959 = n4958 ^ n4952 ;
  assign n4960 = n4535 & n4959 ;
  assign n4961 = n4960 ^ n4952 ;
  assign n4962 = ~n4943 & ~n4961 ;
  assign n4964 = n4963 ^ n4962 ;
  assign n4965 = ~n4554 & n4964 ;
  assign n4968 = n4967 ^ n4965 ;
  assign n4969 = n4968 ^ x88 ;
  assign n4994 = n2923 ^ n2901 ;
  assign n4995 = n4994 ^ n2904 ;
  assign n4996 = ~n2797 & ~n4995 ;
  assign n4992 = n2976 ^ n2928 ;
  assign n4984 = n2977 ^ n2942 ;
  assign n4985 = n4984 ^ n2952 ;
  assign n4986 = n4985 ^ n2949 ;
  assign n4987 = n4986 ^ n2933 ;
  assign n4988 = ~n2797 & ~n4987 ;
  assign n4989 = n4988 ^ n4985 ;
  assign n4993 = n4992 ^ n4989 ;
  assign n4997 = n4996 ^ n4993 ;
  assign n4998 = n2798 & ~n4997 ;
  assign n4971 = n2920 ^ n2909 ;
  assign n4972 = n4971 ^ n2952 ;
  assign n4973 = n4972 ^ n2941 ;
  assign n4974 = ~n2752 & ~n4973 ;
  assign n4975 = n4974 ^ n4971 ;
  assign n4990 = n4989 ^ n4975 ;
  assign n4991 = n4990 ^ n2984 ;
  assign n4999 = n4998 ^ n4991 ;
  assign n4976 = n4975 ^ n2942 ;
  assign n4979 = n4976 ^ n2902 ;
  assign n4980 = n4979 ^ n4976 ;
  assign n4981 = n2752 & ~n4980 ;
  assign n4982 = n4981 ^ n4976 ;
  assign n4983 = ~n2797 & n4982 ;
  assign n5000 = n4999 ^ n4983 ;
  assign n5001 = n5000 ^ n4970 ;
  assign n5002 = n5001 ^ n1653 ;
  assign n5003 = n5002 ^ x106 ;
  assign n5004 = ~n4969 & n5003 ;
  assign n5074 = n5004 ^ n4969 ;
  assign n5075 = n4901 & ~n5074 ;
  assign n4927 = n3243 & ~n3258 ;
  assign n4925 = n3270 & n3306 ;
  assign n4917 = n3234 ^ n3227 ;
  assign n4905 = n3004 & n3853 ;
  assign n4906 = n4905 ^ n3305 ;
  assign n4918 = n4917 ^ n4906 ;
  assign n4919 = n4918 ^ n3275 ;
  assign n4920 = n4919 ^ n3861 ;
  assign n4912 = n3222 ^ n3210 ;
  assign n4913 = n4912 ^ n3221 ;
  assign n4914 = n4913 ^ n3234 ;
  assign n4915 = n4914 ^ n3279 ;
  assign n4916 = ~n3004 & n4915 ;
  assign n4921 = n4920 ^ n4916 ;
  assign n4922 = n3201 & ~n4921 ;
  assign n4904 = n3845 ^ n3309 ;
  assign n4907 = n4906 ^ n4904 ;
  assign n4908 = n4907 ^ n3275 ;
  assign n4909 = n4908 ^ n3841 ;
  assign n4910 = n4909 ^ n2487 ;
  assign n4911 = n4910 ^ n3247 ;
  assign n4923 = n4922 ^ n4911 ;
  assign n4902 = n3275 ^ n3247 ;
  assign n4903 = n3004 & ~n4902 ;
  assign n4924 = n4923 ^ n4903 ;
  assign n4926 = n4925 ^ n4924 ;
  assign n4928 = n4927 ^ n4926 ;
  assign n4929 = n4928 ^ x115 ;
  assign n4930 = n4929 ^ n4901 ;
  assign n5005 = ~n4930 & n5004 ;
  assign n5081 = n5075 ^ n5005 ;
  assign n5007 = n5003 ^ n4901 ;
  assign n5008 = n5007 ^ n5003 ;
  assign n5009 = n5003 ^ n4929 ;
  assign n5010 = n5009 ^ n5003 ;
  assign n5011 = ~n5008 & ~n5010 ;
  assign n5012 = n5011 ^ n5003 ;
  assign n5013 = n4969 & n5012 ;
  assign n5084 = n5081 ^ n5013 ;
  assign n5027 = n4969 ^ n4930 ;
  assign n5019 = n4969 ^ n4901 ;
  assign n5020 = n5019 ^ n5003 ;
  assign n5021 = n5020 ^ n4969 ;
  assign n5024 = n5003 & n5009 ;
  assign n5022 = n5004 ^ n5003 ;
  assign n5023 = n5022 ^ n4929 ;
  assign n5025 = n5024 ^ n5023 ;
  assign n5026 = ~n5021 & ~n5025 ;
  assign n5028 = n5027 ^ n5026 ;
  assign n5085 = n5084 ^ n5028 ;
  assign n5386 = n5006 & n5085 ;
  assign n5387 = n5386 ^ n5028 ;
  assign n5014 = ~n4901 & ~n4969 ;
  assign n5015 = n5014 ^ n5003 ;
  assign n5016 = n4969 ^ n4929 ;
  assign n5017 = n5015 & n5016 ;
  assign n5018 = n5017 ^ n4930 ;
  assign n5382 = n5018 ^ n5009 ;
  assign n5380 = n5024 ^ n4969 ;
  assign n5381 = n4901 & n5380 ;
  assign n5383 = n5382 ^ n5381 ;
  assign n5384 = n5006 & n5383 ;
  assign n5385 = n5384 ^ n5018 ;
  assign n5388 = n5387 ^ n5385 ;
  assign n5389 = n5062 & ~n5388 ;
  assign n5390 = n5389 ^ n5385 ;
  assign n5391 = n5390 ^ n3362 ;
  assign n5392 = n5391 ^ x108 ;
  assign n5394 = n5061 ^ x118 ;
  assign n5447 = ~n3920 & n4004 ;
  assign n5441 = n4011 ^ n4003 ;
  assign n4073 = n4008 ^ n3984 ;
  assign n4074 = n4008 ^ n3920 ;
  assign n4075 = n4074 ^ n4008 ;
  assign n4076 = n4073 & ~n4075 ;
  assign n4077 = n4076 ^ n4008 ;
  assign n4078 = ~n3921 & n4077 ;
  assign n5442 = n5441 ^ n4078 ;
  assign n5443 = n5442 ^ n4622 ;
  assign n5444 = n5443 ^ n4610 ;
  assign n5445 = n5444 ^ n4585 ;
  assign n4042 = n3921 ^ n3920 ;
  assign n5434 = n3997 ^ n3942 ;
  assign n5435 = n5434 ^ n4011 ;
  assign n5436 = n4011 ^ n3921 ;
  assign n5437 = n5436 ^ n4011 ;
  assign n5438 = ~n5435 & ~n5437 ;
  assign n5439 = n5438 ^ n4011 ;
  assign n5440 = ~n4042 & ~n5439 ;
  assign n5446 = n5445 ^ n5440 ;
  assign n5448 = n5447 ^ n5446 ;
  assign n5427 = n4030 ^ n4003 ;
  assign n5425 = n4004 ^ n4003 ;
  assign n5428 = n5427 ^ n5425 ;
  assign n5429 = n5425 ^ n3920 ;
  assign n5430 = n5429 ^ n5425 ;
  assign n5431 = n5428 & n5430 ;
  assign n5432 = n5431 ^ n5425 ;
  assign n5433 = ~n3921 & n5432 ;
  assign n5449 = n5448 ^ n5433 ;
  assign n5450 = n5449 ^ n4016 ;
  assign n5451 = ~n4050 & n5450 ;
  assign n5452 = n5451 ^ n1706 ;
  assign n5453 = n5452 ^ x125 ;
  assign n5422 = n4091 & n4477 ;
  assign n5414 = n4175 ^ n4169 ;
  assign n5415 = n5414 ^ n4196 ;
  assign n5416 = n5415 ^ n4191 ;
  assign n5417 = n4090 & ~n5416 ;
  assign n5418 = n5417 ^ n4166 ;
  assign n5419 = n4089 & n5418 ;
  assign n5410 = n4493 ^ n4166 ;
  assign n5396 = n4187 ^ n4179 ;
  assign n5397 = n5396 ^ n4187 ;
  assign n5398 = n5397 ^ n4181 ;
  assign n5399 = n5398 ^ n4214 ;
  assign n5400 = n4090 & ~n5399 ;
  assign n5401 = n5400 ^ n5396 ;
  assign n5411 = n5410 ^ n5401 ;
  assign n5412 = n5411 ^ n1679 ;
  assign n5402 = n5401 ^ n4170 ;
  assign n5403 = n5402 ^ n4175 ;
  assign n5404 = n5403 ^ n5401 ;
  assign n5405 = n5401 ^ n4089 ;
  assign n5406 = n5405 ^ n5401 ;
  assign n5407 = n5404 & ~n5406 ;
  assign n5408 = n5407 ^ n5401 ;
  assign n5409 = ~n4091 & n5408 ;
  assign n5413 = n5412 ^ n5409 ;
  assign n5420 = n5419 ^ n5413 ;
  assign n5395 = ~n4226 & n4228 ;
  assign n5421 = n5420 ^ n5395 ;
  assign n5423 = n5422 ^ n5421 ;
  assign n5424 = n5423 ^ x77 ;
  assign n5474 = n5453 ^ n5424 ;
  assign n5475 = n5394 & ~n5474 ;
  assign n5476 = n5475 ^ n5474 ;
  assign n5457 = n2250 ^ x91 ;
  assign n5458 = ~n5394 & n5457 ;
  assign n5459 = n5458 ^ n5394 ;
  assign n5454 = ~n5424 & n5453 ;
  assign n5460 = n5454 ^ n5453 ;
  assign n5462 = n5460 ^ n5424 ;
  assign n5463 = n5462 ^ n5453 ;
  assign n5466 = ~n5459 & ~n5463 ;
  assign n5464 = n5458 & ~n5463 ;
  assign n5461 = ~n5459 & n5460 ;
  assign n5465 = n5464 ^ n5461 ;
  assign n5467 = n5466 ^ n5465 ;
  assign n5477 = n5476 ^ n5467 ;
  assign n5393 = n3317 ^ x94 ;
  assign n5481 = n5002 ^ x108 ;
  assign n5482 = ~n5393 & n5481 ;
  assign n5541 = n5482 ^ n5393 ;
  assign n5540 = n5453 ^ n5394 ;
  assign n5542 = n5541 ^ n5540 ;
  assign n5493 = n5457 ^ n5453 ;
  assign n5494 = n5493 ^ n5424 ;
  assign n5495 = n5424 ^ n5394 ;
  assign n5497 = n5453 & ~n5495 ;
  assign n5498 = n5497 ^ n5424 ;
  assign n5499 = n5494 & n5498 ;
  assign n5543 = n5542 ^ n5499 ;
  assign n5544 = n5477 & n5543 ;
  assign n5545 = n5544 ^ n5541 ;
  assign n5507 = n5482 ^ n5481 ;
  assign n5546 = n5507 ^ n5477 ;
  assign n5547 = ~n5545 & ~n5546 ;
  assign n5548 = n5547 ^ n3401 ;
  assign n5470 = n5454 & ~n5459 ;
  assign n5500 = n5499 ^ n5470 ;
  assign n5469 = n5466 ^ n5464 ;
  assign n5471 = n5470 ^ n5469 ;
  assign n5472 = n5471 ^ n5459 ;
  assign n5473 = n5472 ^ n5465 ;
  assign n5478 = n5477 ^ n5473 ;
  assign n5501 = n5500 ^ n5478 ;
  assign n5484 = n5458 ^ n5457 ;
  assign n5487 = ~n5463 & n5484 ;
  assign n5491 = n5487 ^ n5463 ;
  assign n5492 = n5491 ^ n5469 ;
  assign n5502 = n5501 ^ n5492 ;
  assign n5485 = n5454 & n5484 ;
  assign n5503 = n5502 ^ n5485 ;
  assign n5489 = n5459 ^ n5457 ;
  assign n5455 = ~n5394 & n5454 ;
  assign n5483 = n5455 ^ n5454 ;
  assign n5490 = n5489 ^ n5483 ;
  assign n5504 = n5503 ^ n5490 ;
  assign n5505 = n5504 ^ n5485 ;
  assign n5513 = n5505 ^ n5487 ;
  assign n5514 = n5513 ^ n5501 ;
  assign n5515 = n5514 ^ n5475 ;
  assign n5516 = n5515 ^ n5503 ;
  assign n5527 = n5516 ^ n5487 ;
  assign n5526 = n5485 ^ n5484 ;
  assign n5528 = n5527 ^ n5526 ;
  assign n5517 = n5516 ^ n5492 ;
  assign n5520 = n5492 ^ n5393 ;
  assign n5521 = n5520 ^ n5492 ;
  assign n5522 = ~n5517 & n5521 ;
  assign n5523 = n5522 ^ n5492 ;
  assign n5524 = ~n5481 & ~n5523 ;
  assign n5525 = n5524 ^ n5505 ;
  assign n5529 = n5528 ^ n5525 ;
  assign n5537 = n5529 ^ n5471 ;
  assign n5534 = n5503 & ~n5516 ;
  assign n5535 = n5534 ^ n5529 ;
  assign n5536 = n5393 & n5535 ;
  assign n5538 = n5537 ^ n5536 ;
  assign n5539 = ~n5481 & n5538 ;
  assign n5549 = n5548 ^ n5539 ;
  assign n5456 = n5455 ^ n5394 ;
  assign n5468 = n5467 ^ n5456 ;
  assign n5479 = n5478 ^ n5468 ;
  assign n5508 = n5479 & ~n5507 ;
  assign n5509 = n5508 ^ n5478 ;
  assign n5510 = ~n5470 & n5509 ;
  assign n5486 = n5485 ^ n5483 ;
  assign n5488 = n5487 ^ n5486 ;
  assign n5506 = n5505 ^ n5488 ;
  assign n5511 = n5510 ^ n5506 ;
  assign n5512 = n5482 & ~n5511 ;
  assign n5550 = n5549 ^ n5512 ;
  assign n5480 = n5393 & ~n5479 ;
  assign n5551 = n5550 ^ n5480 ;
  assign n5552 = n5551 ^ x126 ;
  assign n5712 = n5392 & n5552 ;
  assign n5738 = n5706 & n5712 ;
  assign n5739 = n5738 ^ n5712 ;
  assign n5736 = ~n5705 & n5712 ;
  assign n5707 = n5706 ^ n5703 ;
  assign n5722 = n5707 & n5712 ;
  assign n5737 = n5736 ^ n5722 ;
  assign n5740 = n5739 ^ n5737 ;
  assign n5713 = n5712 ^ n5392 ;
  assign n5714 = n5713 ^ n5552 ;
  assign n5724 = n5714 ^ n5392 ;
  assign n5725 = n5706 & n5724 ;
  assign n5774 = n5740 ^ n5725 ;
  assign n5775 = n5769 & n5774 ;
  assign n5770 = n5738 & n5769 ;
  assign n5729 = n5554 ^ n5552 ;
  assign n5730 = ~n5703 & ~n5729 ;
  assign n5731 = n5730 ^ n5552 ;
  assign n5732 = n5703 ^ n5392 ;
  assign n5733 = ~n5731 & n5732 ;
  assign n5553 = n5552 ^ n5392 ;
  assign n5555 = n5554 ^ n5553 ;
  assign n5754 = n5733 ^ n5555 ;
  assign n5726 = n5704 & n5713 ;
  assign n5718 = ~n5705 & ~n5714 ;
  assign n5750 = n5726 ^ n5718 ;
  assign n5743 = n5707 & n5713 ;
  assign n5719 = n5718 ^ n5714 ;
  assign n5716 = n5706 & ~n5714 ;
  assign n5715 = n5704 & ~n5714 ;
  assign n5717 = n5716 ^ n5715 ;
  assign n5720 = n5719 ^ n5717 ;
  assign n5748 = n5743 ^ n5720 ;
  assign n5747 = n5722 ^ n5707 ;
  assign n5749 = n5748 ^ n5747 ;
  assign n5751 = n5750 ^ n5749 ;
  assign n5752 = n5751 ^ n5743 ;
  assign n5741 = n5740 ^ n5730 ;
  assign n5728 = n5719 ^ n5704 ;
  assign n5734 = n5733 ^ n5728 ;
  assign n5735 = n5734 ^ n5718 ;
  assign n5742 = n5741 ^ n5735 ;
  assign n5744 = n5743 ^ n5742 ;
  assign n5727 = n5726 ^ n5713 ;
  assign n5745 = n5744 ^ n5727 ;
  assign n5746 = n5745 ^ n5725 ;
  assign n5753 = n5752 ^ n5746 ;
  assign n5755 = n5754 ^ n5753 ;
  assign n5756 = n5379 & n5755 ;
  assign n5757 = n5756 ^ n5754 ;
  assign n5771 = n5770 ^ n5757 ;
  assign n5761 = n5745 ^ n5720 ;
  assign n5762 = n5761 ^ n5744 ;
  assign n5763 = n5744 ^ n5379 ;
  assign n5764 = n5763 ^ n5744 ;
  assign n5765 = ~n5762 & ~n5764 ;
  assign n5766 = n5765 ^ n5744 ;
  assign n5767 = n5349 & ~n5766 ;
  assign n5772 = n5771 ^ n5767 ;
  assign n5721 = n5720 ^ n5718 ;
  assign n5723 = n5722 ^ n5721 ;
  assign n5758 = n5757 ^ n5723 ;
  assign n5708 = n5707 ^ n5552 ;
  assign n5709 = n5555 & n5708 ;
  assign n5710 = n5709 ^ n5552 ;
  assign n5711 = ~n5379 & n5710 ;
  assign n5759 = n5758 ^ n5711 ;
  assign n5760 = n5349 & ~n5759 ;
  assign n5773 = n5772 ^ n5760 ;
  assign n5776 = n5775 ^ n5773 ;
  assign n5777 = n5379 ^ n5349 ;
  assign n5778 = n5737 ^ n5726 ;
  assign n5779 = n5737 ^ n5349 ;
  assign n5780 = n5779 ^ n5737 ;
  assign n5781 = n5778 & n5780 ;
  assign n5782 = n5781 ^ n5737 ;
  assign n5783 = n5777 & n5782 ;
  assign n5784 = ~n5776 & ~n5783 ;
  assign n5785 = n5784 ^ n3898 ;
  assign n5786 = n5785 ^ x66 ;
  assign n5066 = ~n4929 & ~n5019 ;
  assign n5067 = n5066 ^ n4901 ;
  assign n5068 = n5009 & ~n5067 ;
  assign n5082 = n5081 ^ n5068 ;
  assign n5083 = n5082 ^ n4930 ;
  assign n5086 = n5085 ^ n5083 ;
  assign n5069 = n5022 ^ n4969 ;
  assign n5070 = n5069 ^ n5015 ;
  assign n5071 = n5070 ^ n5003 ;
  assign n5072 = ~n4929 & n5071 ;
  assign n5073 = n5072 ^ n5020 ;
  assign n5076 = n5075 ^ n5073 ;
  assign n5077 = n5076 ^ n5068 ;
  assign n5078 = n5062 & ~n5077 ;
  assign n5079 = n5078 ^ n5073 ;
  assign n5087 = n5086 ^ n5079 ;
  assign n5029 = n5028 ^ n5018 ;
  assign n5030 = n5029 ^ n5024 ;
  assign n5031 = n5030 ^ n5013 ;
  assign n5032 = n5031 ^ n5027 ;
  assign n5080 = n5079 ^ n5032 ;
  assign n5088 = n5087 ^ n5080 ;
  assign n5089 = n5087 ^ n5062 ;
  assign n5090 = n5089 ^ n5087 ;
  assign n5091 = n5088 & ~n5090 ;
  assign n5092 = n5091 ^ n5087 ;
  assign n5093 = n5006 & ~n5092 ;
  assign n5094 = n5093 ^ n5079 ;
  assign n5095 = ~n5005 & n5094 ;
  assign n5096 = n5095 ^ n3003 ;
  assign n5097 = n5096 ^ x101 ;
  assign n5263 = n5262 ^ x83 ;
  assign n5264 = ~n5097 & n5263 ;
  assign n5265 = n5264 ^ n5263 ;
  assign n5266 = n5265 ^ n5097 ;
  assign n3838 = n3837 ^ x84 ;
  assign n3867 = n3866 ^ x105 ;
  assign n3899 = n3898 ^ x98 ;
  assign n3900 = n3867 & n3899 ;
  assign n3919 = n3918 ^ x74 ;
  assign n4082 = n4081 ^ n4078 ;
  assign n4083 = n4082 ^ n4072 ;
  assign n4017 = n3920 & ~n4010 ;
  assign n4018 = n4017 ^ n4008 ;
  assign n4019 = n4018 ^ n4011 ;
  assign n4020 = n4019 ^ n4002 ;
  assign n4021 = n4020 ^ n4018 ;
  assign n4022 = n4018 ^ n3920 ;
  assign n4023 = n4022 ^ n4018 ;
  assign n4024 = ~n4021 & ~n4023 ;
  assign n4025 = n4024 ^ n4018 ;
  assign n4026 = n3921 & n4025 ;
  assign n4027 = n4026 ^ n4018 ;
  assign n4060 = n3924 & n3985 ;
  assign n4058 = n3922 & n4029 ;
  assign n4053 = n3998 ^ n3987 ;
  assign n4056 = n4055 ^ n4053 ;
  assign n4040 = n4039 ^ n4032 ;
  assign n4047 = n4040 ^ n4000 ;
  assign n4028 = n4015 ^ n4011 ;
  assign n4041 = n4040 ^ n4028 ;
  assign n4043 = n4028 ^ n3921 ;
  assign n4044 = n4042 & ~n4043 ;
  assign n4045 = n4044 ^ n3921 ;
  assign n4046 = ~n4041 & n4045 ;
  assign n4048 = n4047 ^ n4046 ;
  assign n4057 = n4056 ^ n4048 ;
  assign n4059 = n4058 ^ n4057 ;
  assign n4061 = n4060 ^ n4059 ;
  assign n4062 = n4052 & n4061 ;
  assign n4051 = n4050 ^ n4048 ;
  assign n4063 = n4062 ^ n4051 ;
  assign n4064 = ~n4027 & n4063 ;
  assign n4084 = n4083 ^ n4064 ;
  assign n4085 = ~n4016 & n4084 ;
  assign n4086 = n4085 ^ n469 ;
  assign n4087 = n4086 ^ x122 ;
  assign n4088 = ~n3919 & n4087 ;
  assign n4241 = n4240 ^ x72 ;
  assign n4290 = n2728 ^ n580 ;
  assign n4265 = n2718 ^ n2606 ;
  assign n4266 = n2700 ^ n2605 ;
  assign n4267 = n4266 ^ n2690 ;
  assign n4268 = n2669 & ~n4267 ;
  assign n4269 = ~n4265 & n4268 ;
  assign n4270 = n4269 ^ n2669 ;
  assign n4276 = n4270 ^ n2608 ;
  assign n4271 = n2699 & n2721 ;
  assign n4272 = ~n2610 & n4271 ;
  assign n4273 = n4272 ^ n2698 ;
  assign n4274 = ~n2698 & ~n4273 ;
  assign n4275 = ~n4270 & n4274 ;
  assign n4277 = n4276 ^ n4275 ;
  assign n4278 = n4277 ^ n4270 ;
  assign n4279 = n4278 ^ n4275 ;
  assign n4280 = n4279 ^ n4278 ;
  assign n4281 = n4278 ^ n2687 ;
  assign n4282 = n4281 ^ n4278 ;
  assign n4283 = n4280 & n4282 ;
  assign n4284 = n4283 ^ n4278 ;
  assign n4285 = ~n2697 & n4284 ;
  assign n4286 = n4285 ^ n4277 ;
  assign n4287 = n4286 ^ n2676 ;
  assign n4256 = n4255 ^ n2608 ;
  assign n4258 = n4257 ^ n4256 ;
  assign n4261 = n4260 ^ n4258 ;
  assign n4262 = n2252 & n4261 ;
  assign n4263 = n4262 ^ n2676 ;
  assign n4264 = n2698 & n4263 ;
  assign n4288 = n4287 ^ n4264 ;
  assign n4289 = ~n4253 & ~n4288 ;
  assign n4291 = n4290 ^ n4289 ;
  assign n4292 = n4291 ^ x112 ;
  assign n4293 = n4241 & ~n4292 ;
  assign n4294 = n4293 ^ n4292 ;
  assign n4295 = n4294 ^ n4241 ;
  assign n4296 = n4295 ^ n4292 ;
  assign n4297 = n4088 & n4296 ;
  assign n4298 = n3900 & n4297 ;
  assign n4299 = n4088 ^ n3919 ;
  assign n4300 = ~n4294 & ~n4299 ;
  assign n4377 = n3900 ^ n3899 ;
  assign n4378 = n4300 & n4377 ;
  assign n4328 = n4294 ^ n4088 ;
  assign n4304 = n4299 ^ n4087 ;
  assign n4305 = n4304 ^ n3919 ;
  assign n4311 = n4293 & n4305 ;
  assign n4309 = n4088 & n4295 ;
  assign n4310 = n4309 ^ n4297 ;
  assign n4312 = n4311 ^ n4310 ;
  assign n4307 = n4292 ^ n3919 ;
  assign n4308 = n4087 & n4307 ;
  assign n4313 = n4312 ^ n4308 ;
  assign n4327 = n4313 ^ n4309 ;
  assign n4329 = n4328 ^ n4327 ;
  assign n4302 = n4088 & ~n4294 ;
  assign n4320 = n4302 ^ n4088 ;
  assign n4321 = n4320 ^ n4310 ;
  assign n4325 = n4321 ^ n4300 ;
  assign n4326 = n4325 ^ n4297 ;
  assign n4330 = n4329 ^ n4326 ;
  assign n4323 = n4296 & n4304 ;
  assign n4353 = n4330 ^ n4323 ;
  assign n4335 = n4295 & n4304 ;
  assign n4352 = n4335 ^ n4304 ;
  assign n4354 = n4353 ^ n4352 ;
  assign n4317 = n4296 & ~n4299 ;
  assign n4340 = n4317 ^ n4295 ;
  assign n4306 = n4295 & n4305 ;
  assign n4314 = n4313 ^ n4306 ;
  assign n4338 = n4314 ^ n4300 ;
  assign n4333 = n4317 ^ n4300 ;
  assign n4336 = n4335 ^ n4333 ;
  assign n4337 = n4336 ^ n4327 ;
  assign n4339 = n4338 ^ n4337 ;
  assign n4341 = n4340 ^ n4339 ;
  assign n4334 = n4333 ^ n4299 ;
  assign n4342 = n4341 ^ n4334 ;
  assign n4343 = n4342 ^ n4302 ;
  assign n4324 = n4323 ^ n4306 ;
  assign n4331 = n4330 ^ n4324 ;
  assign n4322 = n4321 ^ n4309 ;
  assign n4332 = n4331 ^ n4322 ;
  assign n4344 = n4343 ^ n4332 ;
  assign n4345 = n3867 & n4344 ;
  assign n4346 = n4345 ^ n4321 ;
  assign n4373 = n4354 ^ n4346 ;
  assign n4369 = n3899 ^ n3867 ;
  assign n4370 = n4309 & n4369 ;
  assign n4363 = n4323 ^ n4297 ;
  assign n4364 = n4297 ^ n3899 ;
  assign n4365 = n4364 ^ n4297 ;
  assign n4366 = n4363 & n4365 ;
  assign n4367 = n4366 ^ n4297 ;
  assign n4368 = ~n3867 & n4367 ;
  assign n4371 = n4370 ^ n4368 ;
  assign n4360 = n3900 ^ n3867 ;
  assign n4361 = n4360 ^ n3899 ;
  assign n4362 = ~n4354 & ~n4361 ;
  assign n4372 = n4371 ^ n4362 ;
  assign n4374 = n4373 ^ n4372 ;
  assign n4349 = n4311 ^ n4305 ;
  assign n4350 = n4349 ^ n4314 ;
  assign n4348 = n4335 ^ n4311 ;
  assign n4351 = n4350 ^ n4348 ;
  assign n4359 = ~n3867 & n4351 ;
  assign n4375 = n4374 ^ n4359 ;
  assign n4355 = n4354 ^ n4351 ;
  assign n4318 = n4317 ^ n4302 ;
  assign n4319 = n4318 ^ n4314 ;
  assign n4347 = n4346 ^ n4319 ;
  assign n4356 = n4355 ^ n4347 ;
  assign n4301 = n4300 ^ n4297 ;
  assign n4303 = n4302 ^ n4301 ;
  assign n4315 = n4314 ^ n4303 ;
  assign n4316 = n3867 & n4315 ;
  assign n4357 = n4356 ^ n4316 ;
  assign n4358 = ~n3899 & ~n4357 ;
  assign n4376 = n4375 ^ n4358 ;
  assign n4379 = n4378 ^ n4376 ;
  assign n4380 = ~n4298 & n4379 ;
  assign n4381 = n4341 ^ n4311 ;
  assign n4382 = n4381 ^ n4313 ;
  assign n4383 = n4313 ^ n3867 ;
  assign n4384 = n4383 ^ n4313 ;
  assign n4385 = n4382 & ~n4384 ;
  assign n4386 = n4385 ^ n4313 ;
  assign n4387 = ~n3899 & n4386 ;
  assign n4388 = n4380 & ~n4387 ;
  assign n4389 = n4388 ^ n3112 ;
  assign n4390 = n4389 ^ x69 ;
  assign n4391 = ~n3838 & n4390 ;
  assign n4574 = n4573 ^ n4565 ;
  assign n4575 = ~n4564 & n4574 ;
  assign n4576 = n4575 ^ n4573 ;
  assign n4651 = n4576 ^ n4572 ;
  assign n4635 = n4565 ^ n4527 ;
  assign n4649 = n4648 ^ n4635 ;
  assign n4650 = n4564 & n4649 ;
  assign n4652 = n4651 ^ n4650 ;
  assign n4653 = ~n4634 & n4652 ;
  assign n4654 = n4653 ^ n4576 ;
  assign n4676 = n4669 ^ n4636 ;
  assign n4677 = n4676 ^ n4647 ;
  assign n4678 = n4677 ^ n4573 ;
  assign n4679 = n4678 ^ n4638 ;
  assign n4663 = n4659 ^ n4524 ;
  assign n4671 = n4670 ^ n4637 ;
  assign n4667 = ~n4665 & n4666 ;
  assign n4672 = n4671 ^ n4667 ;
  assign n4673 = ~n4656 & n4672 ;
  assign n4674 = ~n4663 & n4673 ;
  assign n4675 = n4674 ^ n4672 ;
  assign n4680 = n4679 ^ n4675 ;
  assign n4682 = n4681 ^ n4680 ;
  assign n4683 = n4682 ^ n4675 ;
  assign n4684 = n4675 ^ n4634 ;
  assign n4685 = n4684 ^ n4675 ;
  assign n4686 = n4683 & n4685 ;
  assign n4687 = n4686 ^ n4675 ;
  assign n4688 = n4662 & n4687 ;
  assign n4689 = n4688 ^ n4675 ;
  assign n4660 = n4659 ^ n4567 ;
  assign n4661 = n4656 & n4660 ;
  assign n4690 = n4689 ^ n4661 ;
  assign n4691 = ~n4654 & ~n4690 ;
  assign n4692 = ~n4527 & n4691 ;
  assign n4699 = n4692 & ~n4698 ;
  assign n4700 = n4699 ^ n3152 ;
  assign n4701 = n4700 ^ x118 ;
  assign n4735 = n4734 ^ x110 ;
  assign n4702 = n2988 ^ x84 ;
  assign n4739 = n2240 ^ n851 ;
  assign n4740 = n4739 ^ n2243 ;
  assign n4741 = n4740 ^ n2228 ;
  assign n4742 = n4741 ^ n3914 ;
  assign n4743 = n4742 ^ n967 ;
  assign n4744 = n4743 ^ x124 ;
  assign n4775 = n4774 ^ x101 ;
  assign n4776 = n4744 & ~n4775 ;
  assign n4808 = n4776 ^ n4744 ;
  assign n4809 = n4808 ^ n4775 ;
  assign n4777 = n2747 ^ x75 ;
  assign n4796 = n3303 ^ n3157 ;
  assign n4797 = n4796 ^ n3243 ;
  assign n4798 = n4797 ^ n3278 ;
  assign n4799 = n4798 ^ n3303 ;
  assign n4800 = n3004 & ~n4799 ;
  assign n4801 = n4800 ^ n4796 ;
  assign n4802 = n3201 & n4801 ;
  assign n4788 = n3299 ^ n3225 ;
  assign n4789 = n4788 ^ n3303 ;
  assign n4790 = n4789 ^ n3250 ;
  assign n4791 = n4790 ^ n3840 ;
  assign n4792 = n4791 ^ n3309 ;
  assign n4793 = n4792 ^ n1032 ;
  assign n4780 = n3230 ^ n3225 ;
  assign n4781 = n4780 ^ n3004 ;
  assign n4782 = n4781 ^ n4780 ;
  assign n4783 = n4780 ^ n3242 ;
  assign n4784 = n4783 ^ n4780 ;
  assign n4785 = n4782 & n4784 ;
  assign n4786 = n4785 ^ n4780 ;
  assign n4787 = n3274 & n4786 ;
  assign n4794 = n4793 ^ n4787 ;
  assign n4778 = n3232 ^ n3221 ;
  assign n4779 = ~n3258 & ~n4778 ;
  assign n4795 = n4794 ^ n4779 ;
  assign n4803 = n4802 ^ n4795 ;
  assign n4804 = n4803 ^ x86 ;
  assign n4805 = ~n4777 & n4804 ;
  assign n4806 = n4805 ^ n4804 ;
  assign n4824 = n4806 ^ n4777 ;
  assign n4825 = n4809 & n4824 ;
  assign n4810 = n4806 & n4809 ;
  assign n4826 = n4825 ^ n4810 ;
  assign n4818 = n4805 ^ n4777 ;
  assign n4819 = n4809 & ~n4818 ;
  assign n4823 = n4819 ^ n4809 ;
  assign n4827 = n4826 ^ n4823 ;
  assign n4816 = n4776 & n4805 ;
  assign n4815 = n4805 & n4808 ;
  assign n4817 = n4816 ^ n4815 ;
  assign n4830 = n4827 ^ n4817 ;
  assign n4831 = n4830 ^ n4805 ;
  assign n4829 = n4808 & ~n4818 ;
  assign n4832 = n4831 ^ n4829 ;
  assign n4813 = n4775 ^ n4744 ;
  assign n4833 = n4832 ^ n4813 ;
  assign n4822 = n4776 & ~n4818 ;
  assign n4828 = n4827 ^ n4822 ;
  assign n4834 = n4833 ^ n4828 ;
  assign n4820 = n4819 ^ n4817 ;
  assign n4814 = n4813 ^ n4777 ;
  assign n4821 = n4820 ^ n4814 ;
  assign n4835 = n4834 ^ n4821 ;
  assign n4891 = n4835 ^ n4832 ;
  assign n4892 = n4702 & ~n4891 ;
  assign n4893 = n4892 ^ n4832 ;
  assign n4894 = n4735 & n4893 ;
  assign n4836 = n4835 ^ n4815 ;
  assign n4852 = n4836 ^ n4808 ;
  assign n4850 = n4835 ^ n4829 ;
  assign n4849 = n4806 & n4808 ;
  assign n4851 = n4850 ^ n4849 ;
  assign n4853 = n4852 ^ n4851 ;
  assign n4807 = n4776 & n4806 ;
  assign n4854 = n4853 ^ n4807 ;
  assign n4880 = n4854 ^ n4825 ;
  assign n4844 = n4804 ^ n4775 ;
  assign n4845 = n4777 & n4844 ;
  assign n4881 = n4880 ^ n4845 ;
  assign n4884 = n4881 ^ n4825 ;
  assign n4867 = n4853 ^ n4831 ;
  assign n4843 = n4777 ^ n4744 ;
  assign n4846 = n4845 ^ n4775 ;
  assign n4847 = ~n4843 & ~n4846 ;
  assign n4866 = n4847 ^ n4835 ;
  assign n4868 = n4867 ^ n4866 ;
  assign n4879 = n4868 ^ n4824 ;
  assign n4882 = n4881 ^ n4879 ;
  assign n4883 = ~n4702 & ~n4882 ;
  assign n4885 = n4884 ^ n4883 ;
  assign n4886 = n4735 & n4885 ;
  assign n4736 = n4702 & ~n4735 ;
  assign n4737 = n4736 ^ n4735 ;
  assign n4738 = n4737 ^ n4702 ;
  assign n4877 = n4738 ^ n4735 ;
  assign n4878 = n4828 & n4877 ;
  assign n4887 = n4886 ^ n4878 ;
  assign n4855 = n4854 ^ n4819 ;
  assign n4811 = n4810 ^ n4807 ;
  assign n4812 = n4811 ^ n4738 ;
  assign n4837 = n4836 ^ n4736 ;
  assign n4838 = n4836 ^ n4738 ;
  assign n4839 = n4838 ^ n4836 ;
  assign n4840 = n4837 & ~n4839 ;
  assign n4841 = n4840 ^ n4836 ;
  assign n4842 = n4812 & n4841 ;
  assign n4856 = n4855 ^ n4842 ;
  assign n4848 = n4847 ^ n4804 ;
  assign n4857 = n4856 ^ n4848 ;
  assign n4858 = n4857 ^ n4842 ;
  assign n4859 = ~n4735 & ~n4858 ;
  assign n4860 = n4859 ^ n4856 ;
  assign n4888 = n4887 ^ n4860 ;
  assign n4889 = n4888 ^ n3064 ;
  assign n4865 = n4853 ^ n4811 ;
  assign n4869 = n4868 ^ n4865 ;
  assign n4864 = n4827 ^ n4807 ;
  assign n4870 = n4869 ^ n4864 ;
  assign n4871 = n4870 ^ n4814 ;
  assign n4874 = ~n4735 & n4871 ;
  assign n4861 = n4860 ^ n4842 ;
  assign n4875 = n4874 ^ n4861 ;
  assign n4876 = ~n4702 & ~n4875 ;
  assign n4890 = n4889 ^ n4876 ;
  assign n4895 = n4894 ^ n4890 ;
  assign n4896 = n4895 ^ x125 ;
  assign n4897 = ~n4701 & n4896 ;
  assign n5296 = n4391 & n4897 ;
  assign n4392 = n4391 ^ n4390 ;
  assign n4393 = n4392 ^ n3838 ;
  assign n5291 = n4393 & n4701 ;
  assign n5293 = n5291 ^ n4393 ;
  assign n4394 = n4393 ^ n4390 ;
  assign n5268 = n4897 ^ n4701 ;
  assign n5273 = ~n4394 & ~n5268 ;
  assign n5269 = n4391 & ~n5268 ;
  assign n5274 = n5273 ^ n5269 ;
  assign n5271 = n4392 & ~n5268 ;
  assign n5272 = n5271 ^ n5268 ;
  assign n5275 = n5274 ^ n5272 ;
  assign n5294 = n5293 ^ n5275 ;
  assign n5320 = n5296 ^ n5294 ;
  assign n4898 = n4897 ^ n4896 ;
  assign n5282 = n4391 & n4898 ;
  assign n5286 = n5282 ^ n4394 ;
  assign n5283 = n5282 ^ n5273 ;
  assign n4899 = n4898 ^ n4701 ;
  assign n4900 = ~n4394 & n4899 ;
  assign n5284 = n5283 ^ n4900 ;
  assign n5281 = ~n4394 & n4898 ;
  assign n5285 = n5284 ^ n5281 ;
  assign n5287 = n5286 ^ n5285 ;
  assign n5319 = n5287 ^ n4897 ;
  assign n5321 = n5320 ^ n5319 ;
  assign n5322 = n5321 ^ n5271 ;
  assign n5277 = n4392 & n4898 ;
  assign n5318 = n5277 ^ n4392 ;
  assign n5323 = n5322 ^ n5318 ;
  assign n5290 = n4393 & n4898 ;
  assign n5324 = n5323 ^ n5290 ;
  assign n5345 = n5266 & n5324 ;
  assign n5346 = n5345 ^ n3866 ;
  assign n5267 = n4900 & n5266 ;
  assign n5327 = n5277 ^ n5271 ;
  assign n5328 = n5327 ^ n5287 ;
  assign n5329 = n5328 ^ n5291 ;
  assign n5330 = n5263 & ~n5329 ;
  assign n5331 = n5330 ^ n5274 ;
  assign n5340 = n5331 ^ n5263 ;
  assign n5341 = n5097 & n5340 ;
  assign n5334 = n5282 ^ n5275 ;
  assign n5333 = n5323 ^ n5291 ;
  assign n5335 = n5334 ^ n5333 ;
  assign n5336 = n5097 & ~n5335 ;
  assign n5292 = n5291 ^ n5290 ;
  assign n5325 = n5321 ^ n5292 ;
  assign n5326 = n5325 ^ n5324 ;
  assign n5332 = n5331 ^ n5326 ;
  assign n5337 = n5336 ^ n5332 ;
  assign n5338 = ~n5263 & ~n5337 ;
  assign n5307 = n5263 ^ n5097 ;
  assign n5309 = n5296 ^ n5281 ;
  assign n5297 = n5296 ^ n5269 ;
  assign n5298 = n5297 ^ n3838 ;
  assign n5299 = n5298 ^ n5286 ;
  assign n5308 = n5299 ^ n5281 ;
  assign n5310 = n5309 ^ n5308 ;
  assign n5311 = n5309 ^ n5263 ;
  assign n5312 = n5311 ^ n5309 ;
  assign n5313 = n5310 & ~n5312 ;
  assign n5314 = n5313 ^ n5309 ;
  assign n5315 = n5307 & n5314 ;
  assign n5316 = n5315 ^ n5281 ;
  assign n5295 = n5294 ^ n5292 ;
  assign n5300 = n5299 ^ n5295 ;
  assign n5301 = n5300 ^ n5299 ;
  assign n5302 = n5299 ^ n5263 ;
  assign n5303 = n5302 ^ n5299 ;
  assign n5304 = ~n5301 & n5303 ;
  assign n5305 = n5304 ^ n5299 ;
  assign n5306 = ~n5097 & n5305 ;
  assign n5317 = n5316 ^ n5306 ;
  assign n5339 = n5338 ^ n5317 ;
  assign n5342 = n5341 ^ n5339 ;
  assign n5270 = n5269 ^ n5266 ;
  assign n5276 = n5275 ^ n5270 ;
  assign n5278 = n5277 ^ n5276 ;
  assign n5279 = n5264 & n5278 ;
  assign n5280 = n5279 ^ n5266 ;
  assign n5288 = n5287 ^ n5264 ;
  assign n5289 = n5280 & ~n5288 ;
  assign n5343 = n5342 ^ n5289 ;
  assign n5344 = ~n5267 & n5343 ;
  assign n5347 = n5346 ^ n5344 ;
  assign n5348 = n5347 ^ x73 ;
  assign n6841 = n5786 ^ n5348 ;
  assign n5951 = n5213 ^ n5201 ;
  assign n5952 = ~n5176 & n5951 ;
  assign n5953 = n5952 ^ n5251 ;
  assign n5950 = ~n5176 & n5255 ;
  assign n5954 = n5953 ^ n5950 ;
  assign n5955 = n5954 ^ n5209 ;
  assign n5956 = n5955 ^ n2038 ;
  assign n5920 = n5100 & n5172 ;
  assign n5941 = n5194 ^ n5188 ;
  assign n5939 = n5100 & n5193 ;
  assign n5937 = n5254 ^ n5196 ;
  assign n5938 = n5937 ^ n5213 ;
  assign n5940 = n5939 ^ n5938 ;
  assign n5942 = n5941 ^ n5940 ;
  assign n5936 = ~n5177 & n5191 ;
  assign n5943 = n5942 ^ n5936 ;
  assign n5944 = n5099 ^ n5098 ;
  assign n5945 = ~n5943 & ~n5944 ;
  assign n5946 = n5945 ^ n5098 ;
  assign n5930 = n5203 ^ n5193 ;
  assign n5931 = n5203 ^ n5099 ;
  assign n5932 = n5931 ^ n5203 ;
  assign n5933 = ~n5930 & ~n5932 ;
  assign n5934 = n5933 ^ n5203 ;
  assign n5935 = n5098 & ~n5934 ;
  assign n5947 = n5946 ^ n5935 ;
  assign n5921 = n5190 ^ n5187 ;
  assign n5922 = n5921 ^ n5178 ;
  assign n5923 = n5231 ^ n5212 ;
  assign n5924 = n5923 ^ n5176 ;
  assign n5927 = ~n5921 & n5924 ;
  assign n5928 = n5927 ^ n5176 ;
  assign n5929 = ~n5922 & ~n5928 ;
  assign n5948 = n5947 ^ n5929 ;
  assign n5949 = ~n5920 & n5948 ;
  assign n5957 = n5956 ^ n5949 ;
  assign n5958 = n5957 ^ x73 ;
  assign n5916 = n5375 ^ n1614 ;
  assign n5897 = n4643 ^ n4571 ;
  assign n5887 = ~n4463 & n4642 ;
  assign n5888 = n5887 ^ n4677 ;
  assign n5898 = n5897 ^ n5888 ;
  assign n5899 = n5888 ^ n4634 ;
  assign n5900 = n5899 ^ n5888 ;
  assign n5901 = n5898 & ~n5900 ;
  assign n5902 = n5901 ^ n5888 ;
  assign n5903 = n4662 & n5902 ;
  assign n5891 = n4669 ^ n4658 ;
  assign n5892 = n4669 ^ n4634 ;
  assign n5893 = n5892 ^ n4669 ;
  assign n5894 = n5891 & ~n5893 ;
  assign n5895 = n5894 ^ n4669 ;
  assign n5896 = n4662 & n5895 ;
  assign n5904 = n5903 ^ n5896 ;
  assign n5889 = n5888 ^ n4668 ;
  assign n5890 = n4655 & n5889 ;
  assign n5905 = n5904 ^ n5890 ;
  assign n5880 = n4671 ^ n4636 ;
  assign n5881 = n5880 ^ n4671 ;
  assign n5882 = n4671 ^ n4634 ;
  assign n5883 = n5882 ^ n4671 ;
  assign n5884 = n5881 & n5883 ;
  assign n5885 = n5884 ^ n4671 ;
  assign n5886 = ~n4662 & n5885 ;
  assign n5906 = n5905 ^ n5886 ;
  assign n5878 = n4659 ^ n4527 ;
  assign n5879 = ~n4665 & n5878 ;
  assign n5907 = n5906 ^ n5879 ;
  assign n5870 = n4645 ^ n4643 ;
  assign n5871 = n5870 ^ n4569 ;
  assign n5872 = n5871 ^ n4645 ;
  assign n5873 = n4645 ^ n4634 ;
  assign n5874 = n5873 ^ n4645 ;
  assign n5875 = n5872 & n5874 ;
  assign n5876 = n5875 ^ n4645 ;
  assign n5877 = ~n4662 & n5876 ;
  assign n5908 = n5907 ^ n5877 ;
  assign n5917 = n5916 ^ n5908 ;
  assign n5911 = ~n4564 & ~n5908 ;
  assign n5912 = n5368 & n5911 ;
  assign n5913 = n5912 ^ n5368 ;
  assign n5866 = n5368 ^ n4576 ;
  assign n5914 = n5913 ^ n5866 ;
  assign n5915 = n4634 & n5914 ;
  assign n5918 = n5917 ^ n5915 ;
  assign n5919 = n5918 ^ x90 ;
  assign n5968 = n5958 ^ n5919 ;
  assign n5790 = n5669 ^ n5667 ;
  assign n5791 = n5790 ^ n5684 ;
  assign n5792 = n5684 ^ n5556 ;
  assign n5793 = n5792 ^ n5684 ;
  assign n5794 = n5791 & ~n5793 ;
  assign n5795 = n5794 ^ n5684 ;
  assign n5796 = ~n5557 & n5795 ;
  assign n5819 = n5584 ^ n5583 ;
  assign n5820 = n5613 & n5819 ;
  assign n5818 = n5646 ^ n5642 ;
  assign n5821 = n5820 ^ n5818 ;
  assign n5822 = n5556 & n5821 ;
  assign n5816 = n5646 ^ n5635 ;
  assign n5811 = n5664 ^ n5632 ;
  assign n5808 = n5637 ^ n5626 ;
  assign n5809 = n5808 ^ n5647 ;
  assign n5810 = n5809 ^ n5698 ;
  assign n5812 = n5811 ^ n5810 ;
  assign n5813 = ~n5556 & ~n5812 ;
  assign n5814 = n5813 ^ n5810 ;
  assign n5817 = n5816 ^ n5814 ;
  assign n5823 = n5822 ^ n5817 ;
  assign n5824 = ~n5557 & ~n5823 ;
  assign n5797 = ~n5557 & n5650 ;
  assign n5798 = n5797 ^ n5641 ;
  assign n5801 = n5798 ^ n5652 ;
  assign n5802 = n5801 ^ n5798 ;
  assign n5803 = n5557 & n5802 ;
  assign n5804 = n5803 ^ n5798 ;
  assign n5805 = ~n5556 & n5804 ;
  assign n5806 = n5805 ^ n5798 ;
  assign n5807 = n5806 ^ n5618 ;
  assign n5815 = n5814 ^ n5807 ;
  assign n5825 = n5824 ^ n5815 ;
  assign n5826 = ~n5796 & n5825 ;
  assign n5827 = n5826 ^ n2184 ;
  assign n5828 = n5827 ^ x99 ;
  assign n5963 = n5919 ^ n5828 ;
  assign n5829 = n5479 ^ n5470 ;
  assign n5830 = n5541 ^ n5507 ;
  assign n5832 = n5524 ^ n5507 ;
  assign n5844 = n5492 & n5529 ;
  assign n5845 = n5832 & n5844 ;
  assign n5835 = n5486 ^ n5473 ;
  assign n5833 = n5470 ^ n5455 ;
  assign n5834 = n5833 ^ n5466 ;
  assign n5836 = n5835 ^ n5834 ;
  assign n5837 = n5836 ^ n5482 ;
  assign n5838 = n5504 ^ n5501 ;
  assign n5839 = n5838 ^ n5836 ;
  assign n5840 = ~n5837 & ~n5839 ;
  assign n5841 = n5840 ^ n5482 ;
  assign n5843 = n5841 ^ n5832 ;
  assign n5846 = n5845 ^ n5843 ;
  assign n5831 = ~n5393 & n5527 ;
  assign n5847 = n5846 ^ n5831 ;
  assign n5849 = n5836 ^ n5501 ;
  assign n5848 = n5485 ^ n5478 ;
  assign n5850 = n5849 ^ n5848 ;
  assign n5851 = n5848 ^ n5393 ;
  assign n5852 = n5851 ^ n5848 ;
  assign n5853 = ~n5850 & n5852 ;
  assign n5854 = n5853 ^ n5848 ;
  assign n5855 = ~n5481 & n5854 ;
  assign n5856 = ~n5847 & ~n5855 ;
  assign n5857 = ~n5830 & n5856 ;
  assign n5858 = ~n5829 & n5857 ;
  assign n5859 = n5858 ^ n5856 ;
  assign n5862 = n5859 ^ n1865 ;
  assign n5860 = n5393 & n5465 ;
  assign n5861 = n5859 & n5860 ;
  assign n5863 = n5862 ^ n5861 ;
  assign n5864 = n5863 ^ x72 ;
  assign n5975 = n5963 ^ n5864 ;
  assign n5976 = n5958 & ~n5975 ;
  assign n5977 = n5976 ^ n5864 ;
  assign n5978 = ~n5968 & n5977 ;
  assign n5979 = n5978 ^ n5977 ;
  assign n5865 = n5864 ^ n5828 ;
  assign n5965 = ~n5864 & n5919 ;
  assign n5971 = n5965 ^ n5864 ;
  assign n5969 = ~n5864 & ~n5968 ;
  assign n5970 = n5969 ^ n5919 ;
  assign n5972 = n5971 ^ n5970 ;
  assign n5973 = ~n5865 & ~n5972 ;
  assign n5974 = ~n5963 & n5973 ;
  assign n5980 = n5979 ^ n5974 ;
  assign n5966 = n5965 ^ n5919 ;
  assign n5959 = n5958 ^ n5864 ;
  assign n5960 = n5919 & n5959 ;
  assign n5967 = n5966 ^ n5960 ;
  assign n5981 = n5980 ^ n5967 ;
  assign n5982 = n5981 ^ n5864 ;
  assign n5993 = n5982 ^ n5828 ;
  assign n5994 = n5993 ^ n5974 ;
  assign n5987 = n5958 ^ n5828 ;
  assign n5990 = n5987 ^ n5973 ;
  assign n5961 = n5960 ^ n5958 ;
  assign n5962 = n5865 & ~n5961 ;
  assign n5989 = n5978 ^ n5962 ;
  assign n5991 = n5990 ^ n5989 ;
  assign n5983 = n5959 ^ n5919 ;
  assign n5992 = n5991 ^ n5983 ;
  assign n5995 = n5994 ^ n5992 ;
  assign n5984 = ~n5982 & ~n5983 ;
  assign n5985 = n5984 ^ n5919 ;
  assign n5964 = n5963 ^ n5962 ;
  assign n5986 = n5985 ^ n5964 ;
  assign n5988 = n5987 ^ n5986 ;
  assign n5996 = n5995 ^ n5988 ;
  assign n6013 = ~n4868 & n4877 ;
  assign n6007 = n4871 ^ n4834 ;
  assign n6008 = n4702 & ~n6007 ;
  assign n6009 = n6008 ^ n4834 ;
  assign n6014 = n6013 ^ n6009 ;
  assign n6015 = n6014 ^ n4886 ;
  assign n6016 = n6015 ^ n1247 ;
  assign n6003 = n4827 ^ n4816 ;
  assign n6004 = n6003 ^ n4819 ;
  assign n6005 = n6004 ^ n4881 ;
  assign n6006 = n6005 ^ n4893 ;
  assign n6010 = n6009 ^ n6006 ;
  assign n5997 = n4804 ^ n4777 ;
  assign n5998 = n4777 ^ n4775 ;
  assign n5999 = n5998 ^ n4777 ;
  assign n6000 = ~n5997 & ~n5999 ;
  assign n6001 = n6000 ^ n4777 ;
  assign n6002 = n4702 & ~n6001 ;
  assign n6011 = n6010 ^ n6002 ;
  assign n6012 = n4735 & n6011 ;
  assign n6017 = n6016 ^ n6012 ;
  assign n6018 = n6017 ^ x66 ;
  assign n6046 = n4297 & n4377 ;
  assign n6047 = n6046 ^ n4378 ;
  assign n6033 = n4314 ^ n4311 ;
  assign n6034 = n6033 ^ n4341 ;
  assign n6026 = n4353 ^ n3867 ;
  assign n6027 = n6026 ^ n4383 ;
  assign n6028 = n6027 ^ n3867 ;
  assign n6029 = n4369 ^ n3867 ;
  assign n6030 = n6028 & ~n6029 ;
  assign n6031 = n6030 ^ n3867 ;
  assign n6032 = ~n4331 & n6031 ;
  assign n6035 = n6034 ^ n6032 ;
  assign n6048 = n6047 ^ n6035 ;
  assign n6040 = n4350 ^ n4318 ;
  assign n6041 = n4350 ^ n3867 ;
  assign n6042 = n6041 ^ n4350 ;
  assign n6043 = n6040 & n6042 ;
  assign n6044 = n6043 ^ n4350 ;
  assign n6045 = ~n4369 & n6044 ;
  assign n6049 = n6048 ^ n6045 ;
  assign n6036 = n6035 ^ n4355 ;
  assign n6023 = n4343 ^ n4306 ;
  assign n6037 = n6036 ^ n6023 ;
  assign n6020 = n4341 ^ n4327 ;
  assign n6021 = n6020 ^ n4321 ;
  assign n6019 = n4355 ^ n4330 ;
  assign n6022 = n6021 ^ n6019 ;
  assign n6024 = n6023 ^ n6022 ;
  assign n6025 = ~n3867 & ~n6024 ;
  assign n6038 = n6037 ^ n6025 ;
  assign n6039 = ~n3899 & n6038 ;
  assign n6050 = n6049 ^ n6039 ;
  assign n6051 = ~n4371 & ~n6050 ;
  assign n6052 = n6051 ^ n4362 ;
  assign n6053 = ~n4298 & n6052 ;
  assign n6054 = n6053 ^ n850 ;
  assign n6055 = n6054 ^ x113 ;
  assign n6056 = n5828 & ~n5970 ;
  assign n6057 = n6056 ^ n5983 ;
  assign n6058 = n6057 ^ n5964 ;
  assign n6059 = n6055 & ~n6058 ;
  assign n6060 = n6059 ^ n5964 ;
  assign n6063 = n6060 ^ n5985 ;
  assign n6061 = n5978 ^ n5975 ;
  assign n6062 = n6061 ^ n6060 ;
  assign n6064 = n6063 ^ n6062 ;
  assign n6067 = n6055 & ~n6064 ;
  assign n6068 = n6067 ^ n6063 ;
  assign n6069 = n6018 & n6068 ;
  assign n6070 = n6069 ^ n6060 ;
  assign n6071 = n5996 & n6070 ;
  assign n6072 = n6071 ^ n3918 ;
  assign n6073 = n6072 ^ x107 ;
  assign n6074 = n5387 ^ n5062 ;
  assign n6075 = n6074 ^ n5389 ;
  assign n6076 = n6075 ^ n2593 ;
  assign n6077 = n6076 ^ x117 ;
  assign n6078 = n5551 ^ x67 ;
  assign n6079 = ~n6077 & n6078 ;
  assign n6083 = n5378 ^ x93 ;
  assign n6109 = n3899 & n4321 ;
  assign n6091 = n4334 ^ n4310 ;
  assign n6092 = n6091 ^ n4331 ;
  assign n6093 = n6092 ^ n4334 ;
  assign n6094 = n6093 ^ n4350 ;
  assign n6095 = ~n3867 & ~n6094 ;
  assign n6096 = n6095 ^ n6091 ;
  assign n6103 = n4311 ^ n3900 ;
  assign n6104 = n6103 ^ n4324 ;
  assign n6105 = n4360 & n6104 ;
  assign n6097 = n3900 & ~n4354 ;
  assign n6098 = n6097 ^ n4298 ;
  assign n6099 = n6098 ^ n4369 ;
  assign n6100 = n6099 ^ n6045 ;
  assign n6101 = n6100 ^ n6098 ;
  assign n6102 = n6101 ^ n6045 ;
  assign n6106 = n6105 ^ n6102 ;
  assign n6107 = n6096 & n6106 ;
  assign n6108 = n6107 ^ n6100 ;
  assign n6110 = n6109 ^ n6108 ;
  assign n6084 = n4338 ^ n3899 ;
  assign n6085 = n6084 ^ n4338 ;
  assign n6088 = n4339 & ~n6085 ;
  assign n6089 = n6088 ^ n4338 ;
  assign n6090 = ~n4369 & n6089 ;
  assign n6111 = n6110 ^ n6090 ;
  assign n6112 = ~n4378 & ~n6111 ;
  assign n6113 = ~n4387 & n6112 ;
  assign n6114 = n6113 ^ n4156 ;
  assign n6115 = n6114 ^ x91 ;
  assign n6116 = n6083 & n6115 ;
  assign n6117 = n6116 ^ n6115 ;
  assign n6121 = n4735 ^ n4702 ;
  assign n6122 = ~n4737 & n4849 ;
  assign n6131 = n4868 ^ n4702 ;
  assign n6133 = n4868 ^ n4830 ;
  assign n6132 = n4884 ^ n4868 ;
  assign n6134 = n6133 ^ n6132 ;
  assign n6135 = n6133 ^ n4735 ;
  assign n6136 = n6135 ^ n6133 ;
  assign n6137 = n6134 & ~n6136 ;
  assign n6138 = n6137 ^ n6133 ;
  assign n6139 = n6131 & n6138 ;
  assign n6140 = n6139 ^ n4702 ;
  assign n6130 = n4832 & n4877 ;
  assign n6141 = n6140 ^ n6130 ;
  assign n6123 = n6004 ^ n4831 ;
  assign n6124 = n6123 ^ n4826 ;
  assign n6125 = n4826 ^ n4735 ;
  assign n6126 = n6125 ^ n4826 ;
  assign n6127 = n6124 & ~n6126 ;
  assign n6128 = n6127 ^ n4826 ;
  assign n6129 = n6121 & n6128 ;
  assign n6142 = n6141 ^ n6129 ;
  assign n6143 = ~n6122 & n6142 ;
  assign n6144 = ~n4878 & n6143 ;
  assign n6145 = ~n6121 & n6144 ;
  assign n6146 = n4825 ^ n4824 ;
  assign n6119 = n4868 ^ n4853 ;
  assign n6147 = n6146 ^ n6119 ;
  assign n6148 = n6147 ^ n4817 ;
  assign n6149 = n4817 ^ n4735 ;
  assign n6150 = n6149 ^ n4817 ;
  assign n6151 = ~n6148 & n6150 ;
  assign n6152 = n6151 ^ n4817 ;
  assign n6153 = n6145 & n6152 ;
  assign n6154 = n6153 ^ n6144 ;
  assign n6155 = n4850 ^ n4735 ;
  assign n6156 = n6155 ^ n4850 ;
  assign n6159 = ~n4851 & n6156 ;
  assign n6160 = n6159 ^ n4850 ;
  assign n6161 = ~n6121 & ~n6160 ;
  assign n6162 = n6154 & ~n6161 ;
  assign n6163 = ~n4886 & n6162 ;
  assign n6166 = n6163 ^ n4119 ;
  assign n6120 = n6119 ^ n4811 ;
  assign n6164 = n4736 & n6163 ;
  assign n6165 = ~n6120 & n6164 ;
  assign n6167 = n6166 ^ n6165 ;
  assign n6168 = n6167 ^ x110 ;
  assign n6189 = n5558 & n5636 ;
  assign n6179 = n5626 ^ n5556 ;
  assign n6180 = n5696 ^ n5626 ;
  assign n6181 = n6180 ^ n5557 ;
  assign n6182 = n6181 ^ n6180 ;
  assign n6183 = n5671 ^ n5626 ;
  assign n6184 = n6183 ^ n6180 ;
  assign n6185 = n6182 & n6184 ;
  assign n6186 = n6185 ^ n6180 ;
  assign n6187 = ~n6179 & ~n6186 ;
  assign n6188 = n6187 ^ n5556 ;
  assign n6190 = n6189 ^ n6188 ;
  assign n6177 = n5685 ^ n5678 ;
  assign n6178 = n5559 & ~n6177 ;
  assign n6191 = n6190 ^ n6178 ;
  assign n6176 = n5560 & n5642 ;
  assign n6192 = n6191 ^ n6176 ;
  assign n6171 = n5634 ^ n5556 ;
  assign n6172 = n6171 ^ n5634 ;
  assign n6173 = ~n5647 & ~n6172 ;
  assign n6174 = n6173 ^ n5634 ;
  assign n6175 = ~n5557 & n6174 ;
  assign n6193 = n6192 ^ n6175 ;
  assign n6194 = ~n5806 & n6193 ;
  assign n6195 = ~n5661 & n6194 ;
  assign n6196 = ~n5699 & n6195 ;
  assign n6197 = ~n5796 & n6196 ;
  assign n6198 = n6197 ^ n2662 ;
  assign n6199 = n6198 ^ x100 ;
  assign n6200 = ~n6168 & n6199 ;
  assign n6201 = n6200 ^ n6168 ;
  assign n6207 = n6117 & ~n6201 ;
  assign n6208 = n6079 & n6207 ;
  assign n6080 = n6079 ^ n6077 ;
  assign n6081 = n6080 ^ n6078 ;
  assign n6082 = n6081 ^ n6077 ;
  assign n6202 = n6201 ^ n6199 ;
  assign n6204 = n6116 & n6202 ;
  assign n6118 = n6117 ^ n6083 ;
  assign n6203 = ~n6118 & n6202 ;
  assign n6205 = n6204 ^ n6203 ;
  assign n6206 = n6082 & n6205 ;
  assign n6209 = n6208 ^ n6206 ;
  assign n6229 = n6116 ^ n6083 ;
  assign n6251 = n6200 & n6229 ;
  assign n6216 = n6200 ^ n6199 ;
  assign n6239 = n6216 & n6229 ;
  assign n6252 = n6251 ^ n6239 ;
  assign n6253 = n6079 & n6252 ;
  assign n6213 = n6082 ^ n6080 ;
  assign n6230 = ~n6201 & n6229 ;
  assign n6228 = ~n6118 & ~n6201 ;
  assign n6231 = n6230 ^ n6228 ;
  assign n6223 = n6117 & n6200 ;
  assign n6222 = ~n6118 & n6200 ;
  assign n6224 = n6223 ^ n6222 ;
  assign n6217 = ~n6118 & n6216 ;
  assign n6220 = n6217 ^ n6207 ;
  assign n6219 = n6116 & n6216 ;
  assign n6221 = n6220 ^ n6219 ;
  assign n6225 = n6224 ^ n6221 ;
  assign n6226 = ~n6078 & n6225 ;
  assign n6214 = n6116 & n6200 ;
  assign n6215 = n6214 ^ n6207 ;
  assign n6218 = n6217 ^ n6215 ;
  assign n6227 = n6226 ^ n6218 ;
  assign n6232 = n6231 ^ n6227 ;
  assign n6233 = ~n6213 & n6232 ;
  assign n6210 = n6117 & n6202 ;
  assign n6211 = n6210 ^ n6204 ;
  assign n6212 = ~n6080 & n6211 ;
  assign n6234 = n6233 ^ n6212 ;
  assign n6243 = n6116 & ~n6201 ;
  assign n6244 = n6243 ^ n6228 ;
  assign n6240 = n6239 ^ n6210 ;
  assign n6241 = n6078 & n6240 ;
  assign n6242 = n6241 ^ n6239 ;
  assign n6245 = n6244 ^ n6242 ;
  assign n6235 = n6228 ^ n6117 ;
  assign n6236 = n6235 ^ n6203 ;
  assign n6237 = n6236 ^ n6224 ;
  assign n6238 = ~n6078 & n6237 ;
  assign n6246 = n6245 ^ n6238 ;
  assign n6247 = n6213 & ~n6242 ;
  assign n6248 = ~n6246 & n6247 ;
  assign n6249 = n6248 ^ n6213 ;
  assign n6250 = ~n6234 & ~n6249 ;
  assign n6254 = n6253 ^ n6250 ;
  assign n6255 = n6230 ^ n6229 ;
  assign n6256 = n6255 ^ n6252 ;
  assign n6257 = n6256 ^ n6251 ;
  assign n6260 = n6251 ^ n6078 ;
  assign n6261 = n6260 ^ n6251 ;
  assign n6262 = n6257 & n6261 ;
  assign n6263 = n6262 ^ n6251 ;
  assign n6264 = n6213 & n6263 ;
  assign n6265 = n6254 & ~n6264 ;
  assign n6266 = ~n6209 & n6265 ;
  assign n6268 = n6210 ^ n6207 ;
  assign n6267 = n6223 ^ n6117 ;
  assign n6269 = n6268 ^ n6267 ;
  assign n6270 = n6269 ^ n6219 ;
  assign n6271 = n6269 ^ n6077 ;
  assign n6272 = n6271 ^ n6269 ;
  assign n6273 = n6270 & n6272 ;
  assign n6274 = n6273 ^ n6269 ;
  assign n6275 = n6078 & n6274 ;
  assign n6276 = n6266 & ~n6275 ;
  assign n6277 = n6276 ^ n4240 ;
  assign n6278 = n6277 ^ x105 ;
  assign n6279 = ~n6073 & ~n6278 ;
  assign n6365 = n6198 ^ x78 ;
  assign n6364 = n5918 ^ x92 ;
  assign n6412 = n6365 ^ n6364 ;
  assign n6309 = n6076 ^ x75 ;
  assign n6340 = n3774 ^ n3756 ;
  assign n6341 = n6340 ^ n3769 ;
  assign n6335 = n3795 ^ n3780 ;
  assign n6336 = n6335 ^ n3804 ;
  assign n6317 = n3812 ^ n3769 ;
  assign n6327 = n6317 ^ n3787 ;
  assign n6337 = n6336 ^ n6327 ;
  assign n6338 = ~n2748 & n6337 ;
  assign n6339 = n6338 ^ n6327 ;
  assign n6342 = n6341 ^ n6339 ;
  assign n6343 = n6342 ^ n3790 ;
  assign n6344 = n6343 ^ n6339 ;
  assign n6347 = n2748 & ~n6344 ;
  assign n6348 = n6347 ^ n6339 ;
  assign n6349 = ~n3784 & n6348 ;
  assign n6350 = n6349 ^ n6339 ;
  assign n6328 = n6327 ^ n3779 ;
  assign n6318 = n6317 ^ n3807 ;
  assign n6326 = n6318 ^ n3757 ;
  assign n6329 = n6328 ^ n6326 ;
  assign n6330 = n6326 ^ n2251 ;
  assign n6331 = n6330 ^ n6326 ;
  assign n6332 = ~n6329 & ~n6331 ;
  assign n6333 = n6332 ^ n6326 ;
  assign n6334 = ~n2748 & ~n6333 ;
  assign n6351 = n6350 ^ n6334 ;
  assign n6352 = n6351 ^ n3760 ;
  assign n6319 = n6318 ^ n3786 ;
  assign n6320 = n6319 ^ n3760 ;
  assign n6321 = n3760 ^ n2251 ;
  assign n6322 = n6321 ^ n3760 ;
  assign n6323 = n6320 & n6322 ;
  assign n6324 = n6323 ^ n3760 ;
  assign n6325 = n2748 & n6324 ;
  assign n6353 = n6352 ^ n6325 ;
  assign n6354 = n6353 ^ n3803 ;
  assign n6355 = n6354 ^ n2452 ;
  assign n6312 = n3760 ^ n2748 ;
  assign n6313 = n6312 ^ n3760 ;
  assign n6314 = n3796 & n6313 ;
  assign n6315 = n6314 ^ n3760 ;
  assign n6316 = n3784 & n6315 ;
  assign n6356 = n6355 ^ n6316 ;
  assign n6357 = n6356 ^ x124 ;
  assign n6358 = n6309 & n6357 ;
  assign n6359 = n6358 ^ n6309 ;
  assign n6360 = n6359 ^ n6357 ;
  assign n6377 = n6360 ^ n6309 ;
  assign n6302 = ~n5177 & n5951 ;
  assign n6299 = n5254 ^ n5223 ;
  assign n6300 = ~n5098 & n6299 ;
  assign n6282 = n5098 & n5181 ;
  assign n6281 = n5195 ^ n5187 ;
  assign n6283 = n6282 ^ n6281 ;
  assign n6296 = n6283 ^ n5950 ;
  assign n6290 = n5213 ^ n5172 ;
  assign n6291 = n5172 ^ n5098 ;
  assign n6292 = n6291 ^ n5172 ;
  assign n6293 = n6290 & ~n6292 ;
  assign n6294 = n6293 ^ n5172 ;
  assign n6295 = n5099 & n6294 ;
  assign n6297 = n6296 ^ n6295 ;
  assign n6285 = n5923 ^ n5197 ;
  assign n6286 = n6285 ^ n6281 ;
  assign n6287 = n5098 & ~n6286 ;
  assign n6284 = n6283 ^ n5136 ;
  assign n6288 = n6287 ^ n6284 ;
  assign n6289 = n5179 & ~n6288 ;
  assign n6298 = n6297 ^ n6289 ;
  assign n6301 = n6300 ^ n6298 ;
  assign n6303 = n6302 ^ n6301 ;
  assign n6304 = ~n5175 & n6303 ;
  assign n6305 = n6304 ^ n2285 ;
  assign n6306 = n6305 ^ x109 ;
  assign n6307 = n6054 ^ x102 ;
  assign n6308 = ~n6306 & n6307 ;
  assign n6384 = n6308 ^ n6307 ;
  assign n6385 = n6384 ^ n6306 ;
  assign n6386 = n6377 & n6385 ;
  assign n6378 = n6308 & n6377 ;
  assign n6379 = n6378 ^ n6308 ;
  assign n6362 = n6308 & n6358 ;
  assign n6361 = n6308 & ~n6360 ;
  assign n6363 = n6362 ^ n6361 ;
  assign n6380 = n6379 ^ n6363 ;
  assign n6376 = n6307 & ~n6357 ;
  assign n6381 = n6380 ^ n6376 ;
  assign n6371 = n6309 ^ n6306 ;
  assign n6372 = n6371 ^ n6357 ;
  assign n6373 = n6309 & n6372 ;
  assign n6374 = n6373 ^ n6357 ;
  assign n6375 = n6307 & ~n6374 ;
  assign n6382 = n6381 ^ n6375 ;
  assign n6455 = n6386 ^ n6382 ;
  assign n6388 = n6359 & n6385 ;
  assign n6387 = ~n6360 & n6385 ;
  assign n6389 = n6388 ^ n6387 ;
  assign n6390 = n6389 ^ n6385 ;
  assign n6391 = n6390 ^ n6386 ;
  assign n6399 = n6391 ^ n6380 ;
  assign n6398 = n6382 ^ n6373 ;
  assign n6400 = n6399 ^ n6398 ;
  assign n6456 = n6455 ^ n6400 ;
  assign n6457 = ~n6365 & n6456 ;
  assign n6458 = n6457 ^ n6382 ;
  assign n6459 = n6458 ^ n6391 ;
  assign n6460 = n6459 ^ n6458 ;
  assign n6463 = ~n6365 & n6460 ;
  assign n6464 = n6463 ^ n6458 ;
  assign n6465 = ~n6412 & n6464 ;
  assign n6466 = n6465 ^ n6458 ;
  assign n6445 = n6308 ^ n6306 ;
  assign n6446 = n6377 & ~n6445 ;
  assign n6401 = n6400 ^ n6382 ;
  assign n6397 = n6380 ^ n6378 ;
  assign n6402 = n6401 ^ n6397 ;
  assign n6396 = n6389 ^ n6378 ;
  assign n6403 = n6402 ^ n6396 ;
  assign n6404 = n6403 ^ n6357 ;
  assign n6405 = n6404 ^ n6375 ;
  assign n6392 = n6391 ^ n6358 ;
  assign n6383 = n6382 ^ n6362 ;
  assign n6393 = n6392 ^ n6383 ;
  assign n6395 = n6393 ^ n6387 ;
  assign n6406 = n6405 ^ n6395 ;
  assign n6407 = n6406 ^ n6361 ;
  assign n6394 = n6393 ^ n6360 ;
  assign n6408 = n6407 ^ n6394 ;
  assign n6409 = n6408 ^ n6400 ;
  assign n6444 = n6409 ^ n6389 ;
  assign n6447 = n6446 ^ n6444 ;
  assign n6448 = n6365 & n6447 ;
  assign n6420 = ~n6372 & n6376 ;
  assign n6421 = n6420 ^ n6361 ;
  assign n6449 = n6448 ^ n6421 ;
  assign n6450 = ~n6364 & n6449 ;
  assign n6451 = n6450 ^ n6421 ;
  assign n6437 = n6407 ^ n6380 ;
  assign n6438 = n6437 ^ n6383 ;
  assign n6439 = n6383 ^ n6364 ;
  assign n6440 = n6439 ^ n6383 ;
  assign n6441 = ~n6438 & ~n6440 ;
  assign n6442 = n6441 ^ n6383 ;
  assign n6443 = ~n6365 & n6442 ;
  assign n6452 = n6451 ^ n6443 ;
  assign n6453 = n6452 ^ n6378 ;
  assign n6423 = n6384 ^ n6382 ;
  assign n6422 = n6421 ^ n6408 ;
  assign n6424 = n6423 ^ n6422 ;
  assign n6431 = n6424 ^ n6405 ;
  assign n6432 = n6405 ^ n6365 ;
  assign n6433 = n6432 ^ n6405 ;
  assign n6434 = ~n6431 & n6433 ;
  assign n6435 = n6434 ^ n6405 ;
  assign n6436 = n6364 & ~n6435 ;
  assign n6454 = n6453 ^ n6436 ;
  assign n6467 = n6466 ^ n6454 ;
  assign n6425 = n6424 ^ n6408 ;
  assign n6426 = n6408 ^ n6365 ;
  assign n6427 = n6426 ^ n6408 ;
  assign n6428 = n6425 & n6427 ;
  assign n6429 = n6428 ^ n6408 ;
  assign n6430 = ~n6364 & n6429 ;
  assign n6468 = n6467 ^ n6430 ;
  assign n6413 = n6378 ^ n6365 ;
  assign n6414 = n6413 ^ n6378 ;
  assign n6417 = n6395 & n6414 ;
  assign n6418 = n6417 ^ n6378 ;
  assign n6419 = ~n6412 & n6418 ;
  assign n6469 = n6468 ^ n6419 ;
  assign n6470 = n6446 ^ n6424 ;
  assign n6471 = n6424 ^ n6364 ;
  assign n6472 = n6471 ^ n6424 ;
  assign n6473 = n6470 & n6472 ;
  assign n6474 = n6473 ^ n6424 ;
  assign n6475 = ~n6365 & n6474 ;
  assign n6476 = ~n6469 & ~n6475 ;
  assign n6366 = ~n6364 & ~n6365 ;
  assign n6367 = n6366 ^ n6364 ;
  assign n6368 = n6367 ^ n6365 ;
  assign n6410 = ~n6368 & n6409 ;
  assign n6369 = n6363 & ~n6368 ;
  assign n6370 = n6369 ^ n4291 ;
  assign n6411 = n6410 ^ n6370 ;
  assign n6477 = n6476 ^ n6411 ;
  assign n6478 = n6477 ^ x80 ;
  assign n6781 = n6279 & ~n6478 ;
  assign n6794 = n6781 ^ n6279 ;
  assign n6615 = n6318 ^ n3833 ;
  assign n6616 = n6615 ^ n3779 ;
  assign n6613 = n3797 ^ n3788 ;
  assign n6614 = n3767 & n6613 ;
  assign n6617 = n6616 ^ n6614 ;
  assign n6620 = n2751 & ~n6617 ;
  assign n6621 = n6620 ^ n3770 ;
  assign n6622 = ~n2749 & n6621 ;
  assign n6623 = n6622 ^ n3770 ;
  assign n6612 = ~n2751 & n6317 ;
  assign n6624 = n6623 ^ n6612 ;
  assign n6641 = n3786 ^ n2749 ;
  assign n6633 = n2749 & ~n3817 ;
  assign n6634 = n6633 ^ n3784 ;
  assign n6635 = n6318 ^ n3763 ;
  assign n6636 = n6635 ^ n6340 ;
  assign n6637 = ~n6634 & n6636 ;
  assign n6638 = n6637 ^ n3825 ;
  assign n6639 = n6634 ^ n2749 ;
  assign n6640 = ~n6638 & ~n6639 ;
  assign n6642 = n6641 ^ n6640 ;
  assign n6632 = n2750 & ~n3781 ;
  assign n6643 = n6642 ^ n6632 ;
  assign n6625 = n3786 ^ n2748 ;
  assign n6626 = n6625 ^ n3786 ;
  assign n6629 = n3780 & n6626 ;
  assign n6630 = n6629 ^ n3786 ;
  assign n6631 = n3784 & ~n6630 ;
  assign n6644 = n6643 ^ n6631 ;
  assign n6645 = ~n6624 & n6644 ;
  assign n6646 = n6645 ^ n3659 ;
  assign n6647 = n6646 ^ x105 ;
  assign n6661 = n6098 ^ n6047 ;
  assign n6650 = n6023 ^ n4348 ;
  assign n6649 = n6021 ^ n4323 ;
  assign n6651 = n6650 ^ n6649 ;
  assign n6652 = ~n3867 & ~n6651 ;
  assign n6653 = n6652 ^ n6649 ;
  assign n6662 = n6661 ^ n6653 ;
  assign n6663 = n6662 ^ n4362 ;
  assign n6664 = n6663 ^ n4387 ;
  assign n6655 = n4329 ^ n3919 ;
  assign n6656 = n6655 ^ n6653 ;
  assign n6648 = n4325 ^ n4324 ;
  assign n6654 = n6653 ^ n6648 ;
  assign n6657 = n6656 ^ n6654 ;
  assign n6658 = ~n3867 & n6657 ;
  assign n6659 = n6658 ^ n6656 ;
  assign n6660 = ~n3899 & n6659 ;
  assign n6665 = n6664 ^ n6660 ;
  assign n6666 = ~n4350 & ~n6665 ;
  assign n6667 = n6666 ^ n2829 ;
  assign n6668 = n6667 ^ x114 ;
  assign n6669 = n6647 & n6668 ;
  assign n6670 = n6669 ^ n6668 ;
  assign n6671 = n6670 ^ n6647 ;
  assign n6562 = n5697 ^ n5643 ;
  assign n6554 = n5670 ^ n5640 ;
  assign n6555 = n6554 ^ n5808 ;
  assign n6556 = n6555 ^ n5670 ;
  assign n6557 = n5670 ^ n5556 ;
  assign n6558 = n6557 ^ n5670 ;
  assign n6559 = n6556 & n6558 ;
  assign n6560 = n6559 ^ n5670 ;
  assign n6561 = ~n5557 & ~n6560 ;
  assign n6563 = n6562 ^ n6561 ;
  assign n6564 = n6563 ^ n5820 ;
  assign n6565 = n6564 ^ n5679 ;
  assign n6566 = n6565 ^ n6561 ;
  assign n6567 = n5556 & n6566 ;
  assign n6568 = n6567 ^ n6563 ;
  assign n6577 = n6568 ^ n5660 ;
  assign n6553 = n5557 ^ n5556 ;
  assign n6569 = n6568 ^ n6561 ;
  assign n6570 = n6569 ^ n5687 ;
  assign n6571 = n6570 ^ n6569 ;
  assign n6572 = n6569 ^ n5557 ;
  assign n6573 = n6572 ^ n6569 ;
  assign n6574 = n6571 & n6573 ;
  assign n6575 = n6574 ^ n6569 ;
  assign n6576 = n6553 & n6575 ;
  assign n6578 = n6577 ^ n6576 ;
  assign n6579 = n6578 ^ n5699 ;
  assign n6580 = n6579 ^ n5618 ;
  assign n6581 = n6580 ^ n5796 ;
  assign n6582 = n6581 ^ n3568 ;
  assign n6583 = n6582 ^ x64 ;
  assign n6604 = n5375 ^ n3941 ;
  assign n6598 = n4677 ^ n4637 ;
  assign n6599 = ~n4665 & n6598 ;
  assign n6587 = n4648 ^ n4569 ;
  assign n6588 = n6587 ^ n4565 ;
  assign n6594 = n6588 ^ n4527 ;
  assign n6590 = n5887 ^ n4681 ;
  assign n6591 = n6590 ^ n4639 ;
  assign n6589 = n6588 ^ n4571 ;
  assign n6592 = n6591 ^ n6589 ;
  assign n6593 = ~n4634 & n6592 ;
  assign n6595 = n6594 ^ n6593 ;
  assign n6596 = n4662 & n6595 ;
  assign n6586 = n5896 ^ n5367 ;
  assign n6597 = n6596 ^ n6586 ;
  assign n6600 = n6599 ^ n6597 ;
  assign n6585 = n4634 & n4666 ;
  assign n6601 = n6600 ^ n6585 ;
  assign n6584 = n4656 & n4679 ;
  assign n6602 = n6601 ^ n6584 ;
  assign n6603 = ~n4698 & ~n6602 ;
  assign n6605 = n6604 ^ n6603 ;
  assign n6606 = n6605 ^ x74 ;
  assign n6607 = ~n6583 & n6606 ;
  assign n6608 = n6607 ^ n6606 ;
  assign n6609 = n6608 ^ n6583 ;
  assign n6610 = n6609 ^ n6606 ;
  assign n6502 = n6003 ^ n4850 ;
  assign n6503 = n4877 & ~n6502 ;
  assign n6498 = n4880 ^ n4831 ;
  assign n6499 = n4738 & n6498 ;
  assign n6495 = n4868 ^ n4827 ;
  assign n6496 = ~n4737 & ~n6495 ;
  assign n6488 = n6013 ^ n4884 ;
  assign n6489 = n6488 ^ n4867 ;
  assign n6490 = n6119 ^ n4881 ;
  assign n6491 = n4877 & ~n6490 ;
  assign n6492 = n6491 ^ n4736 ;
  assign n6493 = n6489 & n6492 ;
  assign n6494 = n6493 ^ n6161 ;
  assign n6497 = n6496 ^ n6494 ;
  assign n6500 = n6499 ^ n6497 ;
  assign n6479 = n4822 ^ n4820 ;
  assign n6501 = n6500 ^ n6479 ;
  assign n6504 = n6503 ^ n6501 ;
  assign n6480 = n6479 ^ n6147 ;
  assign n6481 = n6480 ^ n4811 ;
  assign n6482 = n6481 ^ n6479 ;
  assign n6483 = n6479 ^ n4702 ;
  assign n6484 = n6483 ^ n6479 ;
  assign n6485 = ~n6482 & ~n6484 ;
  assign n6486 = n6485 ^ n6479 ;
  assign n6487 = ~n6121 & n6486 ;
  assign n6505 = n6504 ^ n6487 ;
  assign n6506 = n6505 ^ n6122 ;
  assign n6507 = n6506 ^ n3979 ;
  assign n6508 = n6507 ^ x81 ;
  assign n6540 = n5835 ^ n5513 ;
  assign n6541 = n5513 ^ n5481 ;
  assign n6542 = n6541 ^ n5513 ;
  assign n6543 = ~n6540 & n6542 ;
  assign n6544 = n6543 ^ n5513 ;
  assign n6545 = n5393 & n6544 ;
  assign n6525 = n5510 ^ n5470 ;
  assign n6526 = n6525 ^ n5509 ;
  assign n6523 = n5508 ^ n5485 ;
  assign n6524 = ~n5541 & ~n6523 ;
  assign n6527 = n6526 ^ n6524 ;
  assign n6528 = n6527 ^ n5465 ;
  assign n6522 = ~n5508 & n5833 ;
  assign n6529 = n6528 ^ n6522 ;
  assign n6519 = n5473 ^ n5466 ;
  assign n6509 = n5528 ^ n5516 ;
  assign n6520 = n6519 ^ n6509 ;
  assign n6521 = n6520 ^ n5494 ;
  assign n6530 = n6529 ^ n6521 ;
  assign n6517 = n5834 ^ n5479 ;
  assign n6518 = n6517 ^ n5473 ;
  assign n6531 = n6530 ^ n6518 ;
  assign n6532 = n6531 ^ n6529 ;
  assign n6533 = ~n5481 & ~n6532 ;
  assign n6534 = n6533 ^ n6530 ;
  assign n6536 = n6529 ^ n5393 ;
  assign n6535 = n6529 ^ n5481 ;
  assign n6537 = n6536 ^ n6535 ;
  assign n6538 = n6534 & n6537 ;
  assign n6539 = n6538 ^ n6536 ;
  assign n6546 = n6545 ^ n6539 ;
  assign n6510 = n6509 ^ n5541 ;
  assign n6511 = n5507 ^ n5501 ;
  assign n6514 = ~n6509 & ~n6511 ;
  assign n6515 = n6514 ^ n5507 ;
  assign n6516 = ~n6510 & n6515 ;
  assign n6547 = n6546 ^ n6516 ;
  assign n6548 = ~n5524 & n6547 ;
  assign n6549 = n6548 ^ n2796 ;
  assign n6550 = n6549 ^ x120 ;
  assign n6551 = ~n6508 & ~n6550 ;
  assign n6678 = n6551 ^ n6508 ;
  assign n6700 = ~n6610 & ~n6678 ;
  assign n6552 = n6551 ^ n6550 ;
  assign n6611 = ~n6552 & ~n6610 ;
  assign n6701 = n6700 ^ n6611 ;
  assign n6673 = n6551 & ~n6610 ;
  assign n6699 = n6673 ^ n6610 ;
  assign n6702 = n6701 ^ n6699 ;
  assign n6771 = ~n6671 & ~n6702 ;
  assign n6772 = n6771 ^ n4086 ;
  assign n6687 = n6551 & n6609 ;
  assign n6682 = ~n6552 & n6583 ;
  assign n6683 = n6682 ^ n6552 ;
  assign n6684 = n6683 ^ n6611 ;
  assign n6685 = n6684 ^ n6673 ;
  assign n6679 = n6607 & ~n6678 ;
  assign n6675 = n6552 ^ n6508 ;
  assign n6676 = n6607 & ~n6675 ;
  assign n6677 = n6676 ^ n6673 ;
  assign n6680 = n6679 ^ n6677 ;
  assign n6681 = n6680 ^ n6607 ;
  assign n6686 = n6685 ^ n6681 ;
  assign n6688 = n6687 ^ n6686 ;
  assign n6674 = n6673 ^ n6551 ;
  assign n6689 = n6688 ^ n6674 ;
  assign n6690 = n6670 & ~n6689 ;
  assign n6672 = n6611 & ~n6671 ;
  assign n6691 = n6690 ^ n6672 ;
  assign n6692 = n6689 ^ n6679 ;
  assign n6693 = n6679 ^ n6647 ;
  assign n6694 = n6693 ^ n6679 ;
  assign n6695 = ~n6692 & n6694 ;
  assign n6696 = n6695 ^ n6679 ;
  assign n6697 = n6668 & n6696 ;
  assign n6698 = n6668 ^ n6647 ;
  assign n6720 = n6687 ^ n6682 ;
  assign n6716 = ~n6552 & n6609 ;
  assign n6717 = n6716 ^ n6682 ;
  assign n6704 = n6609 & ~n6675 ;
  assign n6718 = n6717 ^ n6704 ;
  assign n6719 = n6718 ^ n6609 ;
  assign n6721 = n6720 ^ n6719 ;
  assign n6722 = n6721 ^ n6716 ;
  assign n6723 = n6722 ^ n6704 ;
  assign n6714 = n6608 & ~n6678 ;
  assign n6705 = n6704 ^ n6611 ;
  assign n6713 = n6705 ^ n6687 ;
  assign n6715 = n6714 ^ n6713 ;
  assign n6724 = n6723 ^ n6715 ;
  assign n6727 = n6723 ^ n6647 ;
  assign n6728 = ~n6698 & n6727 ;
  assign n6729 = n6728 ^ n6647 ;
  assign n6730 = n6724 & n6729 ;
  assign n6731 = n6730 ^ n6723 ;
  assign n6732 = n6731 ^ n6676 ;
  assign n6733 = n6732 ^ n6700 ;
  assign n6707 = n6608 & ~n6675 ;
  assign n6708 = n6707 ^ n6685 ;
  assign n6709 = n6708 ^ n6689 ;
  assign n6703 = n6702 ^ n6680 ;
  assign n6706 = n6705 ^ n6703 ;
  assign n6710 = n6709 ^ n6706 ;
  assign n6711 = n6647 & ~n6710 ;
  assign n6712 = n6711 ^ n6709 ;
  assign n6734 = n6733 ^ n6712 ;
  assign n6741 = n6734 ^ n6684 ;
  assign n6742 = n6741 ^ n6734 ;
  assign n6745 = n6734 ^ n6668 ;
  assign n6746 = n6745 ^ n6734 ;
  assign n6747 = ~n6733 & ~n6746 ;
  assign n6748 = ~n6742 & n6747 ;
  assign n6749 = n6748 ^ n6742 ;
  assign n6750 = n6749 ^ n6741 ;
  assign n6751 = n6698 & n6750 ;
  assign n6752 = n6751 ^ n6712 ;
  assign n6753 = ~n6697 & ~n6752 ;
  assign n6754 = n6687 ^ n6668 ;
  assign n6755 = n6754 ^ n6687 ;
  assign n6758 = ~n6688 & ~n6755 ;
  assign n6759 = n6758 ^ n6687 ;
  assign n6760 = n6647 & n6759 ;
  assign n6761 = n6753 & ~n6760 ;
  assign n6762 = ~n6691 & n6761 ;
  assign n6763 = n6716 ^ n6714 ;
  assign n6764 = n6763 ^ n6684 ;
  assign n6765 = n6684 ^ n6668 ;
  assign n6766 = n6765 ^ n6684 ;
  assign n6767 = ~n6764 & ~n6766 ;
  assign n6768 = n6767 ^ n6684 ;
  assign n6769 = ~n6647 & ~n6768 ;
  assign n6770 = n6762 & ~n6769 ;
  assign n6773 = n6772 ^ n6770 ;
  assign n6774 = n6773 ^ x90 ;
  assign n6775 = n6478 & n6774 ;
  assign n6792 = n6279 & n6775 ;
  assign n6795 = n6794 ^ n6792 ;
  assign n6778 = n6775 ^ n6774 ;
  assign n6779 = n6778 ^ n6478 ;
  assign n6780 = n6279 & ~n6779 ;
  assign n6782 = n6781 ^ n6780 ;
  assign n6796 = n6795 ^ n6782 ;
  assign n6280 = n6279 ^ n6073 ;
  assign n6790 = ~n6280 & ~n6779 ;
  assign n10080 = n6796 ^ n6790 ;
  assign n6786 = ~n6280 & n6775 ;
  assign n6797 = n6796 ^ n6786 ;
  assign n6791 = n6790 ^ n6780 ;
  assign n6793 = n6792 ^ n6791 ;
  assign n6798 = n6797 ^ n6793 ;
  assign n6776 = n6775 ^ n6478 ;
  assign n6777 = ~n6280 & n6776 ;
  assign n6789 = n6777 ^ n6073 ;
  assign n6799 = n6798 ^ n6789 ;
  assign n10081 = n10080 ^ n6799 ;
  assign n10082 = ~n5786 & ~n10081 ;
  assign n6807 = n6279 ^ n6278 ;
  assign n6808 = n6807 ^ n6073 ;
  assign n6809 = n6776 & ~n6808 ;
  assign n10083 = n10082 ^ n6809 ;
  assign n10084 = n6841 & n10083 ;
  assign n5787 = ~n5348 & n5786 ;
  assign n5788 = n5787 ^ n5348 ;
  assign n5789 = n5788 ^ n5786 ;
  assign n6785 = n5789 ^ n5348 ;
  assign n6833 = n6775 & ~n6807 ;
  assign n6800 = n6799 ^ n6782 ;
  assign n6819 = n6800 ^ n6778 ;
  assign n6811 = n6778 & ~n6808 ;
  assign n6820 = n6819 ^ n6811 ;
  assign n6834 = n6833 ^ n6820 ;
  assign n6835 = n6834 ^ n6809 ;
  assign n6836 = n6835 ^ n6073 ;
  assign n6813 = ~n6779 & ~n6807 ;
  assign n6814 = n6813 ^ n6779 ;
  assign n6815 = n6814 ^ n6791 ;
  assign n6816 = n6815 ^ n6809 ;
  assign n6812 = n6811 ^ n6808 ;
  assign n6817 = n6816 ^ n6812 ;
  assign n6831 = n6817 ^ n6815 ;
  assign n6830 = n6813 ^ n6811 ;
  assign n6832 = n6831 ^ n6830 ;
  assign n6837 = n6836 ^ n6832 ;
  assign n8744 = n6837 ^ n6815 ;
  assign n9307 = n8744 ^ n6820 ;
  assign n10078 = n6785 & n9307 ;
  assign n9297 = n6833 ^ n6830 ;
  assign n10073 = n5789 & n9297 ;
  assign n9301 = ~n6785 & ~n6791 ;
  assign n10067 = n9301 ^ n6792 ;
  assign n10068 = ~n6841 & n10067 ;
  assign n6783 = n6782 ^ n6777 ;
  assign n10066 = n6783 & ~n9301 ;
  assign n10069 = n10068 ^ n10066 ;
  assign n8754 = n6817 ^ n6799 ;
  assign n8755 = n6799 ^ n5786 ;
  assign n8756 = n8755 ^ n6799 ;
  assign n8757 = ~n8754 & ~n8756 ;
  assign n8758 = n8757 ^ n6799 ;
  assign n8759 = n5348 & ~n8758 ;
  assign n10070 = n10069 ^ n8759 ;
  assign n10065 = ~n5788 & n6799 ;
  assign n10071 = n10070 ^ n10065 ;
  assign n10062 = n6808 ^ n6797 ;
  assign n10063 = n10062 ^ n6813 ;
  assign n10064 = n5787 & ~n10063 ;
  assign n10072 = n10071 ^ n10064 ;
  assign n10074 = n10073 ^ n10072 ;
  assign n10060 = n6834 ^ n6817 ;
  assign n10061 = ~n5788 & ~n10060 ;
  assign n10075 = n10074 ^ n10061 ;
  assign n10076 = n10075 ^ n6809 ;
  assign n10077 = n10076 ^ n4389 ;
  assign n10079 = n10078 ^ n10077 ;
  assign n10085 = n10084 ^ n10079 ;
  assign n10086 = n10085 ^ x100 ;
  assign n7787 = n6219 ^ n6205 ;
  assign n7788 = n7787 ^ n6257 ;
  assign n7789 = ~n6078 & n7788 ;
  assign n7786 = n6219 ^ n6210 ;
  assign n7790 = n7789 ^ n7786 ;
  assign n7791 = n6213 & n7790 ;
  assign n7473 = n6078 ^ n6077 ;
  assign n7772 = n6239 ^ n6223 ;
  assign n7773 = n6239 ^ n6078 ;
  assign n7774 = n7773 ^ n6239 ;
  assign n7775 = n7772 & ~n7774 ;
  assign n7776 = n7775 ^ n6239 ;
  assign n7777 = n7473 & n7776 ;
  assign n7778 = n7777 ^ n6275 ;
  assign n7754 = n6207 ^ n6205 ;
  assign n7751 = n6243 ^ n6204 ;
  assign n7750 = n6230 ^ n6207 ;
  assign n7752 = n7751 ^ n7750 ;
  assign n7753 = n6078 & n7752 ;
  assign n7755 = n7754 ^ n7753 ;
  assign n7779 = n7778 ^ n7755 ;
  assign n7764 = n6222 ^ n6080 ;
  assign n7765 = n6239 ^ n6082 ;
  assign n7768 = ~n6222 & ~n7765 ;
  assign n7769 = n7768 ^ n6082 ;
  assign n7770 = ~n7764 & n7769 ;
  assign n7771 = n7770 ^ n6080 ;
  assign n7780 = n7779 ^ n7771 ;
  assign n7454 = n6228 ^ n6077 ;
  assign n7455 = n7454 ^ n6228 ;
  assign n7456 = n6244 & n7455 ;
  assign n7457 = n7456 ^ n6228 ;
  assign n7458 = ~n6078 & n7457 ;
  assign n7781 = n7780 ^ n7458 ;
  assign n7459 = n6269 ^ n6214 ;
  assign n7475 = n7459 ^ n6223 ;
  assign n7474 = n7459 ^ n6217 ;
  assign n7476 = n7475 ^ n7474 ;
  assign n7477 = n7475 ^ n6078 ;
  assign n7478 = n7477 ^ n7475 ;
  assign n7479 = n7476 & ~n7478 ;
  assign n7480 = n7479 ^ n7475 ;
  assign n7481 = n7473 & n7480 ;
  assign n7482 = n7481 ^ n7459 ;
  assign n7782 = n7781 ^ n7482 ;
  assign n7435 = n6256 ^ n6228 ;
  assign n7485 = n6082 & n7435 ;
  assign n7783 = n7782 ^ n7485 ;
  assign n7784 = n7783 ^ n4734 ;
  assign n7756 = n7755 ^ n6207 ;
  assign n7757 = n7756 ^ n6239 ;
  assign n7758 = n7757 ^ n7755 ;
  assign n7759 = n7755 ^ n6078 ;
  assign n7760 = n7759 ^ n7755 ;
  assign n7761 = n7758 & n7760 ;
  assign n7762 = n7761 ^ n7755 ;
  assign n7763 = n6077 & n7762 ;
  assign n7785 = n7784 ^ n7763 ;
  assign n7792 = n7791 ^ n7785 ;
  assign n7793 = n7792 ^ x78 ;
  assign n6883 = n3780 ^ n3757 ;
  assign n6884 = n6883 ^ n6341 ;
  assign n6885 = ~n2751 & n6884 ;
  assign n6881 = n2750 & n3794 ;
  assign n6875 = n6325 ^ n3806 ;
  assign n6876 = n6875 ^ n3831 ;
  assign n6877 = n6876 ^ n3803 ;
  assign n6878 = n6877 ^ n2893 ;
  assign n6868 = n3796 ^ n3788 ;
  assign n6869 = n6868 ^ n3811 ;
  assign n6870 = n3811 ^ n2251 ;
  assign n6871 = n6870 ^ n3811 ;
  assign n6872 = n6869 & n6871 ;
  assign n6873 = n6872 ^ n3811 ;
  assign n6874 = n2748 & n6873 ;
  assign n6879 = n6878 ^ n6874 ;
  assign n6861 = n6319 ^ n2748 ;
  assign n6862 = n6861 ^ n6319 ;
  assign n6863 = n6319 ^ n3790 ;
  assign n6864 = n6863 ^ n6319 ;
  assign n6865 = ~n6862 & ~n6864 ;
  assign n6866 = n6865 ^ n6319 ;
  assign n6867 = n3784 & n6866 ;
  assign n6880 = n6879 ^ n6867 ;
  assign n6882 = n6881 ^ n6880 ;
  assign n6886 = n6885 ^ n6882 ;
  assign n6887 = n6886 ^ x97 ;
  assign n6889 = n5073 ^ n5032 ;
  assign n6890 = n5006 & ~n6889 ;
  assign n6891 = n6890 ^ n5073 ;
  assign n6893 = n6891 ^ n5082 ;
  assign n6894 = n6893 ^ n5005 ;
  assign n6895 = n6894 ^ n5086 ;
  assign n6896 = n6895 ^ n6891 ;
  assign n6897 = n5006 & n6896 ;
  assign n6898 = n6897 ^ n6893 ;
  assign n6899 = ~n5062 & n6898 ;
  assign n6892 = n6891 ^ n2848 ;
  assign n6900 = n6899 ^ n6892 ;
  assign n6901 = n6900 ^ x98 ;
  assign n6906 = ~n6887 & n6901 ;
  assign n6888 = n6667 ^ x107 ;
  assign n6909 = n6017 ^ x80 ;
  assign n6910 = ~n6888 & n6909 ;
  assign n6911 = n6906 & n6910 ;
  assign n6923 = n6549 ^ x104 ;
  assign n6860 = n5957 ^ x65 ;
  assign n6963 = n6923 ^ n6860 ;
  assign n7001 = n6911 & ~n6963 ;
  assign n7002 = n7001 ^ n2988 ;
  assign n6917 = n6901 & n6910 ;
  assign n6968 = n6917 ^ n6911 ;
  assign n6918 = n6917 ^ n6910 ;
  assign n6903 = ~n6888 & ~n6901 ;
  assign n6934 = n6918 ^ n6903 ;
  assign n6914 = n6887 & ~n6909 ;
  assign n6931 = n6901 & n6914 ;
  assign n6932 = n6931 ^ n6914 ;
  assign n6902 = n6901 ^ n6888 ;
  assign n6904 = n6903 ^ n6902 ;
  assign n6913 = n6904 ^ n6888 ;
  assign n6915 = ~n6913 & n6914 ;
  assign n6933 = n6932 ^ n6915 ;
  assign n6935 = n6934 ^ n6933 ;
  assign n6969 = n6968 ^ n6935 ;
  assign n6905 = n6887 & ~n6904 ;
  assign n6946 = n6905 & n6909 ;
  assign n6945 = n6931 ^ n6905 ;
  assign n6947 = n6946 ^ n6945 ;
  assign n6966 = n6947 ^ n6931 ;
  assign n6964 = n6887 & ~n6913 ;
  assign n6965 = n6964 ^ n6915 ;
  assign n6967 = n6966 ^ n6965 ;
  assign n6970 = n6969 ^ n6967 ;
  assign n6971 = ~n6860 & n6970 ;
  assign n6972 = n6971 ^ n6969 ;
  assign n6982 = n6968 & ~n6972 ;
  assign n6975 = n6964 ^ n6913 ;
  assign n6976 = n6909 & ~n6975 ;
  assign n6977 = n6976 ^ n6975 ;
  assign n6907 = n6906 ^ n6904 ;
  assign n6908 = n6907 ^ n6905 ;
  assign n6912 = n6911 ^ n6908 ;
  assign n6936 = n6935 ^ n6912 ;
  assign n6930 = n6914 ^ n6909 ;
  assign n6937 = n6936 ^ n6930 ;
  assign n6929 = n6908 ^ n6906 ;
  assign n6938 = n6937 ^ n6929 ;
  assign n6978 = n6977 ^ n6938 ;
  assign n6979 = n6978 ^ n6929 ;
  assign n6980 = n6979 ^ n6976 ;
  assign n6973 = n6972 ^ n6947 ;
  assign n6974 = n6973 ^ n6915 ;
  assign n6981 = n6980 ^ n6974 ;
  assign n6983 = n6982 ^ n6981 ;
  assign n6984 = ~n6963 & ~n6983 ;
  assign n6985 = n6984 ^ n6973 ;
  assign n6956 = n6947 ^ n6938 ;
  assign n6955 = n6947 ^ n6946 ;
  assign n6957 = n6956 ^ n6955 ;
  assign n6958 = n6956 ^ n6923 ;
  assign n6959 = n6958 ^ n6956 ;
  assign n6960 = ~n6957 & ~n6959 ;
  assign n6961 = n6960 ^ n6956 ;
  assign n6962 = ~n6860 & ~n6961 ;
  assign n6986 = n6985 ^ n6962 ;
  assign n6919 = ~n6887 & n6918 ;
  assign n6948 = n6947 ^ n6919 ;
  assign n6949 = n6948 ^ n6936 ;
  assign n6950 = n6936 ^ n6860 ;
  assign n6951 = n6950 ^ n6936 ;
  assign n6952 = ~n6949 & n6951 ;
  assign n6953 = n6952 ^ n6936 ;
  assign n6954 = n6923 & ~n6953 ;
  assign n6987 = n6986 ^ n6954 ;
  assign n6920 = n6919 ^ n6918 ;
  assign n6988 = n6987 ^ n6920 ;
  assign n6939 = n6938 ^ n6933 ;
  assign n6940 = n6933 ^ n6923 ;
  assign n6941 = n6940 ^ n6933 ;
  assign n6942 = ~n6939 & ~n6941 ;
  assign n6943 = n6942 ^ n6933 ;
  assign n6944 = n6860 & n6943 ;
  assign n6989 = n6988 ^ n6944 ;
  assign n6916 = n6915 ^ n6912 ;
  assign n6921 = n6920 ^ n6916 ;
  assign n6922 = n6921 ^ n6920 ;
  assign n6926 = ~n6922 & ~n6923 ;
  assign n6927 = n6926 ^ n6920 ;
  assign n6928 = n6860 & n6927 ;
  assign n6990 = n6989 ^ n6928 ;
  assign n6991 = ~n6860 & n6923 ;
  assign n6992 = n6991 ^ n6860 ;
  assign n6993 = n6992 ^ n6923 ;
  assign n6994 = n6920 & n6993 ;
  assign n6996 = n6991 ^ n6923 ;
  assign n6997 = n6946 & n6996 ;
  assign n6995 = n6911 & n6991 ;
  assign n6998 = n6997 ^ n6995 ;
  assign n6999 = ~n6994 & ~n6998 ;
  assign n7000 = ~n6990 & n6999 ;
  assign n7003 = n7002 ^ n7000 ;
  assign n7749 = n7003 ^ x83 ;
  assign n7794 = n7793 ^ n7749 ;
  assign n7073 = n5321 ^ n5275 ;
  assign n7849 = n7073 ^ n5296 ;
  assign n7850 = n7849 ^ n5295 ;
  assign n7848 = n5321 ^ n5274 ;
  assign n7851 = n7850 ^ n7848 ;
  assign n7852 = n7850 ^ n5263 ;
  assign n7853 = n7852 ^ n7850 ;
  assign n7854 = n7851 & n7853 ;
  assign n7855 = n7854 ^ n7850 ;
  assign n7856 = ~n5097 & n7855 ;
  assign n7840 = n5322 ^ n5283 ;
  assign n7841 = n7840 ^ n5324 ;
  assign n7842 = n7841 ^ n5283 ;
  assign n7843 = n5283 ^ n5263 ;
  assign n7844 = n7843 ^ n5283 ;
  assign n7845 = n7842 & n7844 ;
  assign n7846 = n7845 ^ n5283 ;
  assign n7847 = ~n5307 & n7846 ;
  assign n7857 = n7856 ^ n7847 ;
  assign n7858 = n7857 ^ n5281 ;
  assign n7859 = n7858 ^ n5306 ;
  assign n7064 = n5266 ^ n5264 ;
  assign n7089 = n5323 ^ n5269 ;
  assign n7090 = n5269 ^ n5263 ;
  assign n7091 = n7090 ^ n5269 ;
  assign n7092 = n7089 & n7091 ;
  assign n7093 = n7092 ^ n5269 ;
  assign n7094 = n7064 & n7093 ;
  assign n7860 = n7859 ^ n7094 ;
  assign n7832 = n5328 ^ n5307 ;
  assign n7833 = n5328 ^ n5281 ;
  assign n7834 = n7833 ^ n5281 ;
  assign n7835 = n5281 ^ n5263 ;
  assign n7836 = n7835 ^ n5281 ;
  assign n7837 = ~n7834 & ~n7836 ;
  assign n7838 = n7837 ^ n5281 ;
  assign n7839 = n7832 & n7838 ;
  assign n7861 = n7860 ^ n7839 ;
  assign n7862 = n7861 ^ n5267 ;
  assign n7081 = n5287 ^ n4900 ;
  assign n7082 = n5265 & ~n7081 ;
  assign n7863 = n7862 ^ n7082 ;
  assign n7864 = n7863 ^ n5345 ;
  assign n7865 = n7864 ^ n4803 ;
  assign n7866 = n7865 ^ x117 ;
  assign n7566 = n6721 ^ n6717 ;
  assign n7818 = n7566 ^ n6684 ;
  assign n7557 = n6700 ^ n6686 ;
  assign n7816 = n7557 ^ n6677 ;
  assign n7817 = n7816 ^ n6716 ;
  assign n7819 = n7818 ^ n7817 ;
  assign n7820 = n6647 & ~n7819 ;
  assign n7821 = n7820 ^ n7818 ;
  assign n7822 = ~n6698 & n7821 ;
  assign n7796 = n6671 ^ n6668 ;
  assign n7813 = ~n6689 & n7796 ;
  assign n7814 = n7813 ^ n6769 ;
  assign n7804 = n6686 ^ n6676 ;
  assign n7805 = n7804 ^ n7566 ;
  assign n7806 = n7566 ^ n6668 ;
  assign n7807 = n7806 ^ n7566 ;
  assign n7808 = ~n7805 & ~n7807 ;
  assign n7809 = n7808 ^ n7566 ;
  assign n7810 = ~n6647 & n7809 ;
  assign n7811 = n7810 ^ n6668 ;
  assign n7812 = n7811 ^ n6697 ;
  assign n7815 = n7814 ^ n7812 ;
  assign n7823 = n7822 ^ n7815 ;
  assign n7797 = n7796 ^ n6713 ;
  assign n7798 = n6707 ^ n6670 ;
  assign n7801 = ~n6713 & ~n7798 ;
  assign n7802 = n7801 ^ n6670 ;
  assign n7803 = n7797 & n7802 ;
  assign n7824 = n7823 ^ n7803 ;
  assign n7825 = n7824 ^ n6771 ;
  assign n7586 = n6714 ^ n6702 ;
  assign n7587 = n6714 ^ n6647 ;
  assign n7588 = n7587 ^ n6714 ;
  assign n7589 = ~n7586 & n7588 ;
  assign n7590 = n7589 ^ n6714 ;
  assign n7591 = n6668 & n7590 ;
  assign n7826 = n7825 ^ n7591 ;
  assign n7827 = n7826 ^ n4774 ;
  assign n7547 = n6707 ^ n6680 ;
  assign n7548 = ~n6668 & n7547 ;
  assign n7549 = n7548 ^ n6707 ;
  assign n7795 = n6647 & n7549 ;
  assign n7828 = n7827 ^ n7795 ;
  assign n7829 = n7828 ^ x69 ;
  assign n7888 = n7866 ^ n7829 ;
  assign n7112 = ~n5995 & ~n6018 ;
  assign n7113 = n7112 ^ n5992 ;
  assign n7867 = n7113 ^ n6055 ;
  assign n7105 = n5919 ^ n5864 ;
  assign n7106 = n5828 & n5958 ;
  assign n7107 = n7106 ^ n5919 ;
  assign n7108 = ~n7105 & ~n7107 ;
  assign n7109 = n7108 ^ n5919 ;
  assign n7110 = n6018 & n7109 ;
  assign n7111 = n7110 ^ n5990 ;
  assign n7114 = n7113 ^ n7111 ;
  assign n7115 = ~n6055 & ~n7114 ;
  assign n7116 = n7115 ^ n7113 ;
  assign n7868 = n7867 ^ n7116 ;
  assign n7869 = n7868 ^ n7111 ;
  assign n7870 = n7869 ^ n4743 ;
  assign n7871 = n7870 ^ x92 ;
  assign n7872 = n7866 & n7871 ;
  assign n7873 = n7872 ^ n7866 ;
  assign n7874 = n7873 ^ n7871 ;
  assign n7147 = n6412 & n6424 ;
  assign n7141 = n6405 ^ n6388 ;
  assign n7139 = n6399 ^ n6393 ;
  assign n7136 = n6422 ^ n6397 ;
  assign n7140 = n7139 ^ n7136 ;
  assign n7142 = n7141 ^ n7140 ;
  assign n7143 = n6365 & ~n7142 ;
  assign n7137 = n7136 ^ n6393 ;
  assign n7131 = ~n6365 & n6403 ;
  assign n7132 = n7131 ^ n6396 ;
  assign n7138 = n7137 ^ n7132 ;
  assign n7144 = n7143 ^ n7138 ;
  assign n7145 = ~n6364 & n7144 ;
  assign n7125 = n6386 ^ n6365 ;
  assign n7126 = n7125 ^ n6386 ;
  assign n7127 = n6455 ^ n6386 ;
  assign n7128 = n7126 & n7127 ;
  assign n7129 = n7128 ^ n6386 ;
  assign n7130 = ~n6412 & n7129 ;
  assign n7133 = n7132 ^ n7130 ;
  assign n7134 = n7133 ^ n6436 ;
  assign n7119 = n6422 ^ n6395 ;
  assign n7120 = n6395 ^ n6365 ;
  assign n7121 = n7120 ^ n6395 ;
  assign n7122 = n7119 & n7121 ;
  assign n7123 = n7122 ^ n6395 ;
  assign n7124 = n6412 & n7123 ;
  assign n7135 = n7134 ^ n7124 ;
  assign n7146 = n7145 ^ n7135 ;
  assign n7148 = n7147 ^ n7146 ;
  assign n7149 = ~n6369 & ~n7148 ;
  assign n7150 = n7141 ^ n6446 ;
  assign n7151 = n6446 ^ n6365 ;
  assign n7152 = n7151 ^ n6446 ;
  assign n7153 = ~n7150 & ~n7152 ;
  assign n7154 = n7153 ^ n6446 ;
  assign n7155 = ~n6364 & n7154 ;
  assign n7156 = n7149 & ~n7155 ;
  assign n7157 = n7156 ^ n2747 ;
  assign n7830 = n7157 ^ x110 ;
  assign n7895 = n7874 ^ n7830 ;
  assign n7896 = ~n7888 & ~n7895 ;
  assign n7831 = n7829 & ~n7830 ;
  assign n7882 = n7872 ^ n7871 ;
  assign n7883 = n7831 & n7882 ;
  assign n7880 = n7831 & n7872 ;
  assign n7876 = n7831 ^ n7829 ;
  assign n7877 = n7876 ^ n7830 ;
  assign n7878 = n7877 ^ n7829 ;
  assign n7879 = n7873 & ~n7878 ;
  assign n7881 = n7880 ^ n7879 ;
  assign n7884 = n7883 ^ n7881 ;
  assign n7875 = n7831 & ~n7874 ;
  assign n7885 = n7884 ^ n7875 ;
  assign n7926 = n7896 ^ n7885 ;
  assign n7925 = n7873 & n7876 ;
  assign n7927 = n7926 ^ n7925 ;
  assign n7908 = ~n7878 & n7882 ;
  assign n7921 = n7908 ^ n7880 ;
  assign n7889 = ~n7830 & ~n7888 ;
  assign n7886 = n7885 ^ n7831 ;
  assign n7887 = n7886 ^ n7879 ;
  assign n7890 = n7889 ^ n7887 ;
  assign n7922 = n7921 ^ n7890 ;
  assign n7923 = n7922 ^ n7884 ;
  assign n7919 = n7872 & n7876 ;
  assign n7920 = n7919 ^ n7875 ;
  assign n7924 = n7923 ^ n7920 ;
  assign n7928 = n7927 ^ n7924 ;
  assign n7918 = ~n7874 & n7876 ;
  assign n7929 = n7928 ^ n7918 ;
  assign n9574 = n7794 & n7929 ;
  assign n7904 = ~n7749 & ~n7793 ;
  assign n7931 = n7904 ^ n7749 ;
  assign n7932 = n7931 ^ n7793 ;
  assign n8793 = n7928 & ~n7932 ;
  assign n7905 = n7873 & n7877 ;
  assign n8786 = n7919 ^ n7905 ;
  assign n7941 = ~n7874 & n7877 ;
  assign n7942 = n7941 ^ n7925 ;
  assign n8787 = n8786 ^ n7942 ;
  assign n8788 = n7942 ^ n7749 ;
  assign n8789 = n8788 ^ n7942 ;
  assign n8790 = n8787 & ~n8789 ;
  assign n8791 = n8790 ^ n7942 ;
  assign n8792 = n7793 & n8791 ;
  assign n8794 = n8793 ^ n8792 ;
  assign n7933 = n7879 & ~n7932 ;
  assign n9572 = n8794 ^ n7933 ;
  assign n7955 = n7904 ^ n7793 ;
  assign n9568 = n7925 ^ n7905 ;
  assign n9569 = n9568 ^ n7880 ;
  assign n9570 = ~n7955 & n9569 ;
  assign n7891 = n7890 ^ n7878 ;
  assign n7892 = n7891 ^ n7881 ;
  assign n7893 = n7892 ^ n7887 ;
  assign n9571 = n9570 ^ n7893 ;
  assign n9573 = n9572 ^ n9571 ;
  assign n9575 = n9574 ^ n9573 ;
  assign n9563 = n7920 ^ n7749 ;
  assign n9564 = n9563 ^ n7920 ;
  assign n9565 = n7924 & ~n9564 ;
  assign n9566 = n9565 ^ n7920 ;
  assign n9567 = n7793 & n9566 ;
  assign n9576 = n9575 ^ n9567 ;
  assign n9556 = n7893 ^ n7793 ;
  assign n9557 = n9556 ^ n7893 ;
  assign n9558 = ~n7926 & ~n9557 ;
  assign n9559 = n9558 ^ n7893 ;
  assign n9560 = ~n7749 & ~n9559 ;
  assign n9577 = n9576 ^ n9560 ;
  assign n7956 = n7922 & ~n7955 ;
  assign n9578 = n9577 ^ n7956 ;
  assign n9579 = n9578 ^ n4895 ;
  assign n10087 = n9579 ^ x93 ;
  assign n10088 = n10086 & ~n10087 ;
  assign n7117 = n7116 ^ n2250 ;
  assign n7118 = n7117 ^ x101 ;
  assign n7049 = n5750 & n5768 ;
  assign n7043 = n5736 & n5769 ;
  assign n7044 = n7043 ^ n5767 ;
  assign n7032 = ~n5349 & ~n5748 ;
  assign n7033 = n7032 ^ n5743 ;
  assign n7034 = n7033 ^ n5749 ;
  assign n7035 = n7034 ^ n5738 ;
  assign n7036 = n7035 ^ n7033 ;
  assign n7037 = n7033 ^ n5379 ;
  assign n7038 = n7037 ^ n7033 ;
  assign n7039 = ~n7036 & ~n7038 ;
  assign n7040 = n7039 ^ n7033 ;
  assign n7041 = ~n5777 & n7040 ;
  assign n7042 = n7041 ^ n7033 ;
  assign n7045 = n7044 ^ n7042 ;
  assign n7013 = n5720 ^ n5709 ;
  assign n7014 = n7013 ^ n5774 ;
  assign n7015 = n7014 ^ n5740 ;
  assign n7016 = n7015 ^ n5716 ;
  assign n7031 = n7016 ^ n5734 ;
  assign n7046 = n7045 ^ n7031 ;
  assign n7025 = n7014 ^ n5749 ;
  assign n7026 = n7014 ^ n5349 ;
  assign n7027 = n7026 ^ n7014 ;
  assign n7028 = n7025 & n7027 ;
  assign n7029 = n7028 ^ n7014 ;
  assign n7030 = ~n5777 & ~n7029 ;
  assign n7047 = n7046 ^ n7030 ;
  assign n7017 = n7016 ^ n5717 ;
  assign n7018 = n7017 ^ n5744 ;
  assign n7019 = n7018 ^ n7016 ;
  assign n7020 = n7016 ^ n5379 ;
  assign n7021 = n7020 ^ n7016 ;
  assign n7022 = ~n7019 & ~n7021 ;
  assign n7023 = n7022 ^ n7016 ;
  assign n7024 = ~n5777 & ~n7023 ;
  assign n7048 = n7047 ^ n7024 ;
  assign n7050 = n7049 ^ n7048 ;
  assign n7005 = n5745 ^ n5715 ;
  assign n7008 = n5734 ^ n5349 ;
  assign n7009 = n7008 ^ n5734 ;
  assign n7010 = ~n7005 & n7009 ;
  assign n7011 = n7010 ^ n5734 ;
  assign n7012 = n5379 & ~n7011 ;
  assign n7051 = n7050 ^ n7012 ;
  assign n7052 = n7051 ^ n5775 ;
  assign n7053 = ~n5783 & ~n7052 ;
  assign n7054 = n7053 ^ n3544 ;
  assign n7055 = n7054 ^ x94 ;
  assign n7161 = n4895 ^ x82 ;
  assign n7162 = n6582 ^ x89 ;
  assign n7163 = ~n7161 & n7162 ;
  assign n7164 = n5221 ^ n5201 ;
  assign n7165 = n5099 & ~n7164 ;
  assign n7166 = n7165 ^ n5201 ;
  assign n7185 = n7166 ^ n5202 ;
  assign n7182 = n5203 ^ n5191 ;
  assign n7183 = n7182 ^ n5186 ;
  assign n7184 = ~n5099 & ~n7183 ;
  assign n7186 = n7185 ^ n7184 ;
  assign n7187 = n5098 & n7186 ;
  assign n7172 = n5235 ^ n5231 ;
  assign n7173 = ~n5100 & ~n7172 ;
  assign n7168 = n5231 ^ n5194 ;
  assign n7169 = n7168 ^ n5212 ;
  assign n7174 = n7173 ^ n7169 ;
  assign n7175 = n7174 ^ n5923 ;
  assign n7176 = n5197 ^ n5181 ;
  assign n7177 = n5177 & ~n7176 ;
  assign n7178 = ~n7175 & n7177 ;
  assign n7179 = n7178 ^ n7174 ;
  assign n7180 = ~n5179 & ~n7179 ;
  assign n7167 = n7166 ^ n5231 ;
  assign n7181 = n7180 ^ n7167 ;
  assign n7188 = n7187 ^ n7181 ;
  assign n7189 = n7188 ^ n5256 ;
  assign n7190 = ~n5920 & ~n7189 ;
  assign n7191 = ~n6295 & n7190 ;
  assign n7192 = n7191 ^ n5953 ;
  assign n7193 = ~n5260 & n7192 ;
  assign n7194 = n7193 ^ n3600 ;
  assign n7195 = n7194 ^ x106 ;
  assign n7196 = n5833 ^ n5478 ;
  assign n7197 = n7196 ^ n5483 ;
  assign n7198 = n7197 ^ n5833 ;
  assign n7199 = n7198 ^ n6509 ;
  assign n7200 = n5481 & n7199 ;
  assign n7201 = n7200 ^ n7196 ;
  assign n7202 = n5830 & n7201 ;
  assign n7203 = n7202 ^ n5833 ;
  assign n7205 = n5501 ^ n5483 ;
  assign n7206 = n7205 ^ n5479 ;
  assign n7207 = n5393 & ~n7206 ;
  assign n7208 = n7207 ^ n5514 ;
  assign n7209 = ~n5830 & ~n7208 ;
  assign n7204 = n5479 ^ n5464 ;
  assign n7210 = n7209 ^ n7204 ;
  assign n7218 = n7210 ^ n5456 ;
  assign n7211 = n5470 ^ n5393 ;
  assign n7212 = n7211 ^ n5470 ;
  assign n7213 = n5517 ^ n5488 ;
  assign n7214 = n7213 ^ n5470 ;
  assign n7215 = n7212 & ~n7214 ;
  assign n7216 = n7215 ^ n5470 ;
  assign n7217 = n7210 & ~n7216 ;
  assign n7219 = n7218 ^ n7217 ;
  assign n7220 = n7219 ^ n7204 ;
  assign n7221 = n7220 ^ n5456 ;
  assign n7222 = n7221 ^ n7219 ;
  assign n7223 = n7219 ^ n5393 ;
  assign n7224 = n7223 ^ n7219 ;
  assign n7225 = n7222 & n7224 ;
  assign n7226 = n7225 ^ n7219 ;
  assign n7227 = n5481 & ~n7226 ;
  assign n7228 = n7227 ^ n7217 ;
  assign n7229 = ~n7203 & n7228 ;
  assign n7231 = n5467 & n5507 ;
  assign n7232 = n7229 & n7231 ;
  assign n7230 = n7229 ^ n3627 ;
  assign n7233 = n7232 ^ n7230 ;
  assign n7234 = n7233 ^ x96 ;
  assign n7235 = n6646 ^ x121 ;
  assign n7236 = n5096 ^ x123 ;
  assign n7237 = n7235 & ~n7236 ;
  assign n7238 = n7234 & n7237 ;
  assign n7239 = ~n7195 & n7238 ;
  assign n7281 = n7239 ^ n7238 ;
  assign n7317 = n7163 & n7281 ;
  assign n7245 = ~n7234 & n7236 ;
  assign n7260 = n7245 ^ n7236 ;
  assign n7246 = n7235 & n7245 ;
  assign n7247 = n7246 ^ n7235 ;
  assign n7248 = n7247 ^ n7237 ;
  assign n7288 = n7260 ^ n7248 ;
  assign n7240 = n7195 & ~n7235 ;
  assign n7266 = n7240 ^ n7235 ;
  assign n7267 = n7234 & ~n7266 ;
  assign n7268 = n7267 ^ n7266 ;
  assign n7289 = n7288 ^ n7268 ;
  assign n7290 = n7289 ^ n7235 ;
  assign n7261 = n7240 & n7260 ;
  assign n7262 = n7261 ^ n7240 ;
  assign n7291 = n7290 ^ n7262 ;
  assign n7292 = n7291 ^ n7267 ;
  assign n7249 = ~n7195 & n7248 ;
  assign n7307 = n7292 ^ n7249 ;
  assign n7308 = n7307 ^ n7268 ;
  assign n7258 = n7195 & n7246 ;
  assign n7309 = n7308 ^ n7258 ;
  assign n7310 = n7309 ^ n7292 ;
  assign n7311 = ~n7162 & ~n7310 ;
  assign n7312 = n7311 ^ n7307 ;
  assign n7313 = n7161 & n7312 ;
  assign n7293 = n7292 ^ n7239 ;
  assign n7269 = n7246 ^ n7245 ;
  assign n7241 = ~n7236 & n7240 ;
  assign n7263 = n7262 ^ n7241 ;
  assign n7270 = n7269 ^ n7263 ;
  assign n7255 = n7236 ^ n7235 ;
  assign n7256 = n7255 ^ n7195 ;
  assign n7257 = ~n7234 & ~n7256 ;
  assign n7287 = n7270 ^ n7257 ;
  assign n7294 = n7293 ^ n7287 ;
  assign n7295 = ~n7161 & n7294 ;
  assign n7296 = n7295 ^ n7257 ;
  assign n7314 = n7313 ^ n7296 ;
  assign n7277 = n7162 ^ n7161 ;
  assign n7303 = n7277 ^ n7162 ;
  assign n7304 = n7234 & ~n7303 ;
  assign n7305 = n7304 ^ n7162 ;
  assign n7306 = n7241 & n7305 ;
  assign n7315 = n7314 ^ n7306 ;
  assign n7259 = n7258 ^ n7246 ;
  assign n7297 = n7296 ^ n7259 ;
  assign n7283 = n7270 ^ n7258 ;
  assign n7284 = n7283 ^ n7261 ;
  assign n7298 = n7297 ^ n7284 ;
  assign n7242 = n7234 & n7241 ;
  assign n7278 = n7242 ^ n7241 ;
  assign n7271 = n7270 ^ n7268 ;
  assign n7264 = n7263 ^ n7259 ;
  assign n7265 = n7264 ^ n7257 ;
  assign n7272 = n7271 ^ n7265 ;
  assign n7254 = n7238 ^ n7237 ;
  assign n7273 = n7272 ^ n7254 ;
  assign n7279 = n7278 ^ n7273 ;
  assign n7280 = n7279 ^ n7259 ;
  assign n7282 = n7281 ^ n7280 ;
  assign n7285 = n7284 ^ n7282 ;
  assign n7286 = ~n7162 & ~n7285 ;
  assign n7299 = n7298 ^ n7286 ;
  assign n7300 = n7277 & n7299 ;
  assign n7316 = n7315 ^ n7300 ;
  assign n7318 = n7317 ^ n7316 ;
  assign n7319 = n7272 ^ n7267 ;
  assign n7320 = n7319 ^ n7249 ;
  assign n7323 = n7249 ^ n7161 ;
  assign n7324 = n7323 ^ n7249 ;
  assign n7325 = ~n7320 & ~n7324 ;
  assign n7326 = n7325 ^ n7249 ;
  assign n7327 = ~n7162 & n7326 ;
  assign n7328 = ~n7318 & ~n7327 ;
  assign n7251 = n7163 ^ n7161 ;
  assign n7274 = ~n7251 & ~n7273 ;
  assign n7250 = n7249 ^ n7248 ;
  assign n7252 = n7250 & ~n7251 ;
  assign n7243 = n7242 ^ n7239 ;
  assign n7244 = n7163 & n7243 ;
  assign n7253 = n7252 ^ n7244 ;
  assign n7275 = n7274 ^ n7253 ;
  assign n7276 = n7275 ^ n3751 ;
  assign n7329 = n7328 ^ n7276 ;
  assign n7330 = n7329 ^ x75 ;
  assign n7335 = n7055 & n7330 ;
  assign n7336 = n7335 ^ n7330 ;
  assign n7337 = n7336 ^ n7055 ;
  assign n7004 = n7003 ^ x77 ;
  assign n7074 = n7073 ^ n5281 ;
  assign n7075 = n5263 & ~n7074 ;
  assign n7076 = n7075 ^ n5281 ;
  assign n7077 = n7076 ^ n5294 ;
  assign n7095 = n7077 ^ n5316 ;
  assign n7096 = n7095 ^ n7094 ;
  assign n7083 = n5325 ^ n5299 ;
  assign n7084 = n5325 ^ n5263 ;
  assign n7085 = n7084 ^ n5325 ;
  assign n7086 = n7083 & n7085 ;
  assign n7087 = n7086 ^ n5325 ;
  assign n7088 = n7064 & n7087 ;
  assign n7097 = n7096 ^ n7088 ;
  assign n7098 = n7097 ^ n7082 ;
  assign n7078 = n7077 ^ n5296 ;
  assign n7065 = n5295 ^ n5263 ;
  assign n7066 = n5307 & ~n7065 ;
  assign n7067 = n7066 ^ n5263 ;
  assign n7070 = n5334 ^ n5295 ;
  assign n7071 = ~n7067 & n7070 ;
  assign n7068 = n5334 ^ n5327 ;
  assign n7072 = n7071 ^ n7068 ;
  assign n7079 = n7078 ^ n7072 ;
  assign n7080 = ~n7064 & n7079 ;
  assign n7099 = n7098 ^ n7080 ;
  assign n7057 = n5274 ^ n5263 ;
  assign n7058 = n7057 ^ n5274 ;
  assign n7059 = n5282 ^ n4900 ;
  assign n7060 = n7059 ^ n5274 ;
  assign n7061 = n7058 & n7060 ;
  assign n7062 = n7061 ^ n5274 ;
  assign n7063 = ~n5097 & n7062 ;
  assign n7100 = n7099 ^ n7063 ;
  assign n7101 = n7100 ^ n5345 ;
  assign n7102 = n7101 ^ n3317 ;
  assign n7103 = n7102 ^ x84 ;
  assign n7338 = ~n7004 & n7103 ;
  assign n7374 = ~n7337 & n7338 ;
  assign n7339 = n7338 ^ n7103 ;
  assign n7373 = n7336 & n7339 ;
  assign n7375 = n7374 ^ n7373 ;
  assign n7369 = n7337 ^ n7330 ;
  assign n7370 = n7338 & n7369 ;
  assign n7351 = n7103 & ~n7330 ;
  assign n7371 = n7370 ^ n7351 ;
  assign n7372 = n7371 ^ n7339 ;
  assign n7376 = n7375 ^ n7372 ;
  assign n8863 = n7118 & n7376 ;
  assign n7158 = n7157 ^ x118 ;
  assign n7159 = ~n7118 & ~n7158 ;
  assign n7362 = n7159 ^ n7158 ;
  assign n7160 = n7159 ^ n7118 ;
  assign n7389 = n7362 ^ n7160 ;
  assign n7392 = n7370 ^ n7369 ;
  assign n7352 = n7351 ^ n7330 ;
  assign n7353 = n7352 ^ n7103 ;
  assign n7344 = n7338 ^ n7004 ;
  assign n7345 = n7336 & ~n7344 ;
  assign n7340 = n7339 ^ n7004 ;
  assign n7343 = n7335 & n7340 ;
  assign n7346 = n7345 ^ n7343 ;
  assign n7342 = n7336 & n7340 ;
  assign n7347 = n7346 ^ n7342 ;
  assign n7354 = n7353 ^ n7347 ;
  assign n7349 = ~n7337 & ~n7344 ;
  assign n7350 = n7349 ^ n7342 ;
  assign n7355 = n7354 ^ n7350 ;
  assign n7356 = n7355 ^ n7343 ;
  assign n7348 = n7347 ^ n7344 ;
  assign n7357 = n7356 ^ n7348 ;
  assign n7341 = ~n7337 & n7340 ;
  assign n7358 = n7357 ^ n7341 ;
  assign n7359 = n7358 ^ n7349 ;
  assign n7390 = n7359 ^ n7352 ;
  assign n7391 = n7390 ^ n7357 ;
  assign n7393 = n7392 ^ n7391 ;
  assign n7394 = n7393 ^ n7374 ;
  assign n7395 = n7394 ^ n7371 ;
  assign n7377 = n7336 & n7338 ;
  assign n7396 = n7395 ^ n7377 ;
  assign n7397 = n7396 ^ n7393 ;
  assign n7398 = n7393 ^ n7158 ;
  assign n7399 = n7398 ^ n7393 ;
  assign n7400 = n7397 & n7399 ;
  assign n7401 = n7400 ^ n7393 ;
  assign n7402 = ~n7389 & ~n7401 ;
  assign n8864 = n8863 ^ n7402 ;
  assign n9714 = n8864 ^ n7158 ;
  assign n9697 = ~n7362 & ~n7394 ;
  assign n9695 = n7370 ^ n7354 ;
  assign n9686 = n7158 ^ n7118 ;
  assign n7407 = n7395 ^ n7370 ;
  assign n9687 = n7407 ^ n7349 ;
  assign n7378 = n7377 ^ n7376 ;
  assign n9688 = n9687 ^ n7378 ;
  assign n9689 = n9688 ^ n7349 ;
  assign n9690 = n7349 ^ n7158 ;
  assign n9691 = n9690 ^ n7349 ;
  assign n9692 = ~n9689 & ~n9691 ;
  assign n9693 = n9692 ^ n7349 ;
  assign n9694 = ~n9686 & n9693 ;
  assign n9696 = n9695 ^ n9694 ;
  assign n9698 = n9697 ^ n9696 ;
  assign n9715 = n9714 ^ n9698 ;
  assign n8884 = ~n7160 & n7375 ;
  assign n7421 = n7390 ^ n7354 ;
  assign n8883 = ~n7160 & n7421 ;
  assign n8885 = n8884 ^ n8883 ;
  assign n7403 = n7362 ^ n7118 ;
  assign n7404 = n7390 ^ n7345 ;
  assign n7405 = ~n7403 & n7404 ;
  assign n9713 = n8885 ^ n7405 ;
  assign n9716 = n9715 ^ n9713 ;
  assign n8869 = n7353 ^ n7330 ;
  assign n7379 = n7378 ^ n7373 ;
  assign n8870 = n8869 ^ n7379 ;
  assign n9707 = n8870 ^ n7346 ;
  assign n9708 = n7346 ^ n7158 ;
  assign n9709 = n9708 ^ n7346 ;
  assign n9710 = n9707 & n9709 ;
  assign n9711 = n9710 ^ n7346 ;
  assign n9712 = ~n7118 & n9711 ;
  assign n9717 = n9716 ^ n9712 ;
  assign n9718 = n9717 ^ n3837 ;
  assign n9699 = n9698 ^ n9694 ;
  assign n9700 = n9699 ^ n7343 ;
  assign n9701 = n9700 ^ n9699 ;
  assign n9702 = n9699 ^ n7158 ;
  assign n9703 = n9702 ^ n9699 ;
  assign n9704 = ~n9701 & n9703 ;
  assign n9705 = n9704 ^ n9699 ;
  assign n9706 = ~n7118 & ~n9705 ;
  assign n9719 = n9718 ^ n9706 ;
  assign n9679 = n7362 ^ n7358 ;
  assign n9680 = n7342 ^ n7160 ;
  assign n9683 = n7362 & n9680 ;
  assign n9684 = n9683 ^ n7342 ;
  assign n9685 = n9679 & ~n9684 ;
  assign n9720 = n9719 ^ n9685 ;
  assign n10089 = n9720 ^ x83 ;
  assign n7999 = n5996 ^ n4523 ;
  assign n7990 = n5986 & ~n6018 ;
  assign n7991 = n7990 ^ n5985 ;
  assign n8000 = n7999 ^ n7991 ;
  assign n7992 = n7991 ^ n6018 ;
  assign n7993 = n7992 ^ n7991 ;
  assign n7994 = n7991 ^ n6061 ;
  assign n7995 = n7994 ^ n7991 ;
  assign n7996 = n7993 & ~n7995 ;
  assign n7997 = n7996 ^ n7991 ;
  assign n7998 = ~n6055 & ~n7997 ;
  assign n8001 = n8000 ^ n7998 ;
  assign n7987 = ~n6018 & ~n6057 ;
  assign n7988 = n7987 ^ n5996 ;
  assign n7989 = ~n6055 & ~n7988 ;
  assign n8002 = n8001 ^ n7989 ;
  assign n8003 = n8002 ^ x82 ;
  assign n8020 = n6078 & n6217 ;
  assign n8016 = n6230 ^ n6214 ;
  assign n8017 = n8016 ^ n6217 ;
  assign n8018 = ~n6077 & n8017 ;
  assign n8004 = n6268 ^ n6243 ;
  assign n8005 = n8004 ^ n6203 ;
  assign n8006 = ~n6078 & n8005 ;
  assign n8007 = n8006 ^ n6203 ;
  assign n8019 = n8018 ^ n8007 ;
  assign n8021 = n8020 ^ n8019 ;
  assign n8009 = n8007 ^ n6211 ;
  assign n8008 = n8007 ^ n7750 ;
  assign n8010 = n8009 ^ n8008 ;
  assign n8013 = ~n6078 & n8010 ;
  assign n8014 = n8013 ^ n8009 ;
  assign n8015 = n6077 & n8014 ;
  assign n8022 = n8021 ^ n8015 ;
  assign n8023 = n8022 ^ n6208 ;
  assign n8024 = n8023 ^ n6264 ;
  assign n8025 = n8024 ^ n7778 ;
  assign n8026 = n8025 ^ n7771 ;
  assign n7460 = n7459 ^ n6251 ;
  assign n7461 = n7460 ^ n6205 ;
  assign n7462 = ~n6078 & n7461 ;
  assign n7463 = n7462 ^ n6251 ;
  assign n7464 = n7463 ^ n6222 ;
  assign n7465 = n7464 ^ n7463 ;
  assign n7468 = n6078 & n7465 ;
  assign n7469 = n7468 ^ n7463 ;
  assign n7470 = ~n6077 & n7469 ;
  assign n7471 = n7470 ^ n7463 ;
  assign n8027 = n8026 ^ n7471 ;
  assign n8028 = ~n7485 & n8027 ;
  assign n8029 = n8028 ^ n4502 ;
  assign n8030 = n8029 ^ x81 ;
  assign n8031 = n8003 & n8030 ;
  assign n8032 = n8031 ^ n8003 ;
  assign n8033 = n8032 ^ n8030 ;
  assign n8034 = n8033 ^ n8003 ;
  assign n7522 = n7271 ^ n7250 ;
  assign n7523 = n7271 ^ n7162 ;
  assign n7524 = n7523 ^ n7271 ;
  assign n7525 = ~n7522 & n7524 ;
  assign n7526 = n7525 ^ n7271 ;
  assign n7527 = n7161 & ~n7526 ;
  assign n7490 = n7292 ^ n7258 ;
  assign n7491 = ~n7251 & n7490 ;
  assign n8064 = n7491 ^ n7252 ;
  assign n8037 = n7319 ^ n7238 ;
  assign n8036 = n7278 ^ n7239 ;
  assign n8038 = n8037 ^ n8036 ;
  assign n8039 = n8036 ^ n7162 ;
  assign n8040 = n8039 ^ n8036 ;
  assign n8041 = ~n8038 & ~n8040 ;
  assign n8042 = n8041 ^ n8036 ;
  assign n8043 = n7277 & n8042 ;
  assign n8044 = n8043 ^ n8036 ;
  assign n8045 = n7249 ^ n7242 ;
  assign n8046 = n8045 ^ n7162 ;
  assign n8051 = n7283 ^ n7162 ;
  assign n8047 = n7263 ^ n7258 ;
  assign n8048 = n8047 ^ n7273 ;
  assign n7502 = n7291 ^ n7281 ;
  assign n8049 = n8048 ^ n7502 ;
  assign n8050 = ~n7161 & ~n8049 ;
  assign n8052 = n8051 ^ n8050 ;
  assign n8053 = n8046 & n8052 ;
  assign n8054 = n8053 ^ n7162 ;
  assign n8055 = ~n8044 & ~n8054 ;
  assign n7528 = n7251 ^ n7162 ;
  assign n8035 = n7261 & n7528 ;
  assign n8056 = n8055 ^ n8035 ;
  assign n8057 = n7292 ^ n7271 ;
  assign n8058 = n7271 ^ n7161 ;
  assign n8059 = n8058 ^ n7271 ;
  assign n8060 = ~n8057 & n8059 ;
  assign n8061 = n8060 ^ n7271 ;
  assign n8062 = ~n7162 & ~n8061 ;
  assign n8063 = n8056 & ~n8062 ;
  assign n8065 = n8064 ^ n8063 ;
  assign n8066 = ~n7274 & n8065 ;
  assign n8067 = ~n7259 & n8066 ;
  assign n8068 = ~n7527 & n8067 ;
  assign n8069 = n8068 ^ n4460 ;
  assign n8070 = n8069 ^ x120 ;
  assign n8086 = n5768 ^ n5349 ;
  assign n8087 = n5716 & ~n8086 ;
  assign n8088 = n8087 ^ n5770 ;
  assign n8089 = n8088 ^ n7044 ;
  assign n8072 = n7015 ^ n5749 ;
  assign n8073 = n8072 ^ n5742 ;
  assign n8074 = n8073 ^ n5752 ;
  assign n8075 = n8073 ^ n5349 ;
  assign n8076 = n8075 ^ n8073 ;
  assign n8077 = n8074 & ~n8076 ;
  assign n8078 = n8077 ^ n8073 ;
  assign n8079 = ~n5737 & n8078 ;
  assign n8090 = n8089 ^ n8079 ;
  assign n8091 = n8090 ^ n7030 ;
  assign n8092 = n8091 ^ n4413 ;
  assign n8080 = n8079 ^ n5754 ;
  assign n8071 = n5735 ^ n5716 ;
  assign n8081 = n8080 ^ n8071 ;
  assign n8082 = n8081 ^ n8079 ;
  assign n8083 = n5349 & ~n8082 ;
  assign n8084 = n8083 ^ n8080 ;
  assign n8085 = n5379 & ~n8084 ;
  assign n8093 = n8092 ^ n8085 ;
  assign n8094 = n8093 ^ x64 ;
  assign n8095 = n8070 & n8094 ;
  assign n8096 = n8095 ^ n8094 ;
  assign n8100 = n8096 ^ n8070 ;
  assign n8108 = n8100 ^ n8094 ;
  assign n8113 = n8034 & n8108 ;
  assign n7973 = n6708 ^ n6679 ;
  assign n7974 = n7973 ^ n6722 ;
  assign n7975 = n6647 & ~n7974 ;
  assign n7967 = n6702 ^ n6677 ;
  assign n7976 = n7975 ^ n7967 ;
  assign n7977 = ~n6698 & ~n7976 ;
  assign n7968 = n7967 ^ n6760 ;
  assign n7969 = n7968 ^ n7810 ;
  assign n7579 = n6714 ^ n6707 ;
  assign n7580 = n6707 ^ n6647 ;
  assign n7581 = n7580 ^ n6707 ;
  assign n7582 = n7579 & n7581 ;
  assign n7583 = n7582 ^ n6707 ;
  assign n7584 = ~n6668 & n7583 ;
  assign n7970 = n7969 ^ n7584 ;
  assign n7971 = n7970 ^ n7814 ;
  assign n7972 = n7971 ^ n6691 ;
  assign n7978 = n7977 ^ n7972 ;
  assign n7960 = n6700 ^ n6687 ;
  assign n7961 = n7960 ^ n6718 ;
  assign n7962 = n6718 ^ n6647 ;
  assign n7963 = n7962 ^ n6718 ;
  assign n7964 = n7961 & ~n7963 ;
  assign n7965 = n7964 ^ n6718 ;
  assign n7966 = ~n6668 & n7965 ;
  assign n7979 = n7978 ^ n7966 ;
  assign n7980 = ~n7591 & n7979 ;
  assign n7981 = n7980 ^ n4633 ;
  assign n7982 = n7981 ^ x114 ;
  assign n8188 = n8034 & n8095 ;
  assign n8111 = n8032 & n8108 ;
  assign n8104 = n8034 & ~n8100 ;
  assign n8105 = n8104 ^ n8100 ;
  assign n8102 = n8032 & ~n8100 ;
  assign n8101 = n8031 & ~n8100 ;
  assign n8103 = n8102 ^ n8101 ;
  assign n8106 = n8105 ^ n8103 ;
  assign n8112 = n8111 ^ n8106 ;
  assign n8114 = n8113 ^ n8112 ;
  assign n8115 = n8114 ^ n8108 ;
  assign n8109 = n8031 & n8108 ;
  assign n8110 = n8109 ^ n8106 ;
  assign n8116 = n8115 ^ n8110 ;
  assign n10112 = n8188 ^ n8116 ;
  assign n8173 = n8032 & n8095 ;
  assign n8174 = n8173 ^ n8113 ;
  assign n10113 = n10112 ^ n8174 ;
  assign n10114 = ~n7982 & n10113 ;
  assign n8117 = ~n8033 & n8095 ;
  assign n8118 = n8117 ^ n8116 ;
  assign n8107 = n8106 ^ n8033 ;
  assign n8119 = n8118 ^ n8107 ;
  assign n8176 = n8119 ^ n8102 ;
  assign n8098 = n8031 & n8096 ;
  assign n10099 = n8176 ^ n8098 ;
  assign n8097 = n8034 & n8096 ;
  assign n10100 = n10099 ^ n8097 ;
  assign n10101 = n10100 ^ n10099 ;
  assign n8145 = n6430 ^ n6410 ;
  assign n8129 = n6446 ^ n6387 ;
  assign n8130 = n8129 ^ n7136 ;
  assign n8125 = n6387 ^ n6360 ;
  assign n8126 = n8125 ^ n6397 ;
  assign n8127 = n8126 ^ n6393 ;
  assign n8128 = n6365 & ~n8127 ;
  assign n8131 = n8130 ^ n8128 ;
  assign n8132 = n6412 & n8131 ;
  assign n8133 = n8132 ^ n6446 ;
  assign n8123 = n6424 ^ n6362 ;
  assign n8124 = n6366 & n8123 ;
  assign n8134 = n8133 ^ n8124 ;
  assign n8137 = n6380 ^ n6365 ;
  assign n8138 = n8137 ^ n6380 ;
  assign n8139 = n6399 & ~n8138 ;
  assign n8140 = n8139 ^ n6380 ;
  assign n8141 = n6364 & n8140 ;
  assign n8142 = ~n8134 & ~n8141 ;
  assign n8143 = n8142 ^ n7130 ;
  assign n8144 = ~n6466 & n8143 ;
  assign n8146 = n8145 ^ n8144 ;
  assign n8147 = ~n6369 & n8146 ;
  assign n8148 = ~n7155 & n8147 ;
  assign n8149 = n8148 ^ n4563 ;
  assign n8150 = n8149 ^ x88 ;
  assign n10102 = n10099 ^ n8150 ;
  assign n10103 = n10102 ^ n10099 ;
  assign n10104 = ~n10101 & n10103 ;
  assign n10105 = n10104 ^ n10099 ;
  assign n10107 = n8098 ^ n7982 ;
  assign n8158 = n8031 & n8095 ;
  assign n8178 = ~n7982 & n8150 ;
  assign n8184 = n8178 ^ n8150 ;
  assign n9211 = n8158 & n8184 ;
  assign n8159 = n8104 ^ n8098 ;
  assign n8160 = n8159 ^ n8158 ;
  assign n8161 = n8159 ^ n7982 ;
  assign n8162 = n8161 ^ n8159 ;
  assign n8163 = n8160 & n8162 ;
  assign n8164 = n8163 ^ n8159 ;
  assign n8165 = ~n8150 & n8164 ;
  assign n9212 = n9211 ^ n8165 ;
  assign n10108 = n10107 ^ n9212 ;
  assign n8168 = n8150 ^ n8098 ;
  assign n10106 = n9212 ^ n8168 ;
  assign n10109 = n10108 ^ n10106 ;
  assign n10110 = n10105 & ~n10109 ;
  assign n10111 = n10110 ^ n10108 ;
  assign n10115 = n10114 ^ n10111 ;
  assign n10091 = n8106 ^ n7982 ;
  assign n10092 = n10091 ^ n8117 ;
  assign n9206 = n8184 ^ n7982 ;
  assign n8702 = n8119 ^ n8104 ;
  assign n8189 = n8188 ^ n8111 ;
  assign n10093 = n8702 ^ n8189 ;
  assign n10096 = n9206 & ~n10093 ;
  assign n10097 = n10096 ^ n8189 ;
  assign n10098 = ~n10092 & n10097 ;
  assign n10116 = n10115 ^ n10098 ;
  assign n8185 = n8116 & n8184 ;
  assign n10117 = n10116 ^ n8185 ;
  assign n8120 = n8119 ^ n8096 ;
  assign n8099 = n8098 ^ n8097 ;
  assign n8121 = n8120 ^ n8099 ;
  assign n8166 = n8150 ^ n7982 ;
  assign n8693 = n8121 & n8166 ;
  assign n10118 = n10117 ^ n8693 ;
  assign n10090 = ~n8110 & n8178 ;
  assign n10119 = n10118 ^ n10090 ;
  assign n10120 = ~n8113 & ~n10119 ;
  assign n10121 = n10120 ^ n4700 ;
  assign n10122 = n10121 ^ x86 ;
  assign n10123 = n10089 & ~n10122 ;
  assign n10171 = n10088 & n10123 ;
  assign n10128 = n10088 ^ n10086 ;
  assign n10139 = n10123 ^ n10089 ;
  assign n10164 = n10128 & n10139 ;
  assign n10173 = n10171 ^ n10164 ;
  assign n10129 = n10128 ^ n10087 ;
  assign n10162 = n10129 & n10139 ;
  assign n10180 = n10173 ^ n10162 ;
  assign n10160 = n10088 & n10139 ;
  assign n10165 = n10164 ^ n10160 ;
  assign n10166 = n10165 ^ n10162 ;
  assign n10167 = n10166 ^ n10139 ;
  assign n10181 = n10180 ^ n10167 ;
  assign n7636 = n6978 & n6991 ;
  assign n7637 = n7636 ^ n6997 ;
  assign n7638 = ~n6994 & ~n7637 ;
  assign n7688 = n6933 & n6993 ;
  assign n7687 = n6946 & ~n6992 ;
  assign n7689 = n7688 ^ n7687 ;
  assign n7682 = ~n6909 & n6991 ;
  assign n7683 = n7682 ^ n6860 ;
  assign n7684 = ~n6975 & ~n7683 ;
  assign n7672 = n6965 ^ n6938 ;
  assign n7673 = n7672 ^ n6965 ;
  assign n7674 = n6965 ^ n6923 ;
  assign n7675 = n7674 ^ n6965 ;
  assign n7676 = ~n7673 & n7675 ;
  assign n7677 = n7676 ^ n6965 ;
  assign n7678 = ~n6963 & n7677 ;
  assign n7685 = n7684 ^ n7678 ;
  assign n7639 = n6979 ^ n6966 ;
  assign n7660 = n7639 ^ n6975 ;
  assign n7657 = n6969 ^ n6920 ;
  assign n7643 = n6947 ^ n6915 ;
  assign n7644 = n7643 ^ n6919 ;
  assign n7645 = n7644 ^ n6912 ;
  assign n7646 = n7645 ^ n6947 ;
  assign n7647 = ~n6860 & ~n7646 ;
  assign n7648 = n7647 ^ n7643 ;
  assign n7658 = n7657 ^ n7648 ;
  assign n7661 = n7660 ^ n7658 ;
  assign n7662 = n7661 ^ n7648 ;
  assign n7663 = n6860 & n7662 ;
  assign n7659 = n7658 ^ n6911 ;
  assign n7664 = n7663 ^ n7659 ;
  assign n7665 = n6963 & n7664 ;
  assign n7650 = n6933 ^ n6860 ;
  assign n7651 = n7650 ^ n6933 ;
  assign n7653 = n6934 & n7651 ;
  assign n7654 = n7653 ^ n6933 ;
  assign n7655 = n6923 & n7654 ;
  assign n7649 = n7648 ^ n6911 ;
  assign n7656 = n7655 ^ n7649 ;
  assign n7666 = n7665 ^ n7656 ;
  assign n7686 = n7685 ^ n7666 ;
  assign n7690 = n7689 ^ n7686 ;
  assign n7640 = n7639 ^ n6923 ;
  assign n7641 = n7640 ^ n7639 ;
  assign n7642 = n6968 ^ n6912 ;
  assign n7667 = ~n7642 & ~n7666 ;
  assign n7668 = n7667 ^ n7639 ;
  assign n7669 = ~n7641 & ~n7668 ;
  assign n7670 = n7669 ^ n7639 ;
  assign n7671 = n6963 & ~n7670 ;
  assign n7691 = n7690 ^ n7671 ;
  assign n7692 = n7638 & ~n7691 ;
  assign n7693 = n7692 ^ n5002 ;
  assign n8897 = n7693 ^ x74 ;
  assign n8920 = n7155 ^ n4968 ;
  assign n8907 = n6375 ^ n6372 ;
  assign n8905 = n6421 ^ n6401 ;
  assign n8904 = n6391 ^ n6361 ;
  assign n8906 = n8905 ^ n8904 ;
  assign n8908 = n8907 ^ n8906 ;
  assign n8909 = n8906 ^ n6365 ;
  assign n8910 = n8909 ^ n8906 ;
  assign n8911 = n8908 & ~n8910 ;
  assign n8912 = n8911 ^ n8906 ;
  assign n8913 = ~n6412 & n8912 ;
  assign n8914 = n8913 ^ n8906 ;
  assign n8901 = n6420 ^ n6372 ;
  assign n8902 = n8901 ^ n6408 ;
  assign n8903 = ~n6368 & ~n8902 ;
  assign n8915 = n8914 ^ n8903 ;
  assign n8900 = n6362 & ~n6367 ;
  assign n8916 = n8915 ^ n8900 ;
  assign n8917 = ~n8141 & ~n8916 ;
  assign n8918 = n8917 ^ n6475 ;
  assign n8919 = ~n7124 & n8918 ;
  assign n8921 = n8920 ^ n8919 ;
  assign n8922 = n8921 ^ x121 ;
  assign n8898 = n7981 ^ x122 ;
  assign n8969 = n8922 ^ n8898 ;
  assign n8951 = n5323 ^ n5294 ;
  assign n8952 = ~n7064 & ~n8951 ;
  assign n8946 = n5273 ^ n4394 ;
  assign n8947 = n5263 & ~n8946 ;
  assign n8939 = n5297 ^ n5271 ;
  assign n8940 = n8939 ^ n5323 ;
  assign n8941 = ~n5263 & n8940 ;
  assign n8942 = n8941 ^ n5297 ;
  assign n8945 = n8942 ^ n5285 ;
  assign n8948 = n8947 ^ n8945 ;
  assign n8949 = ~n5097 & n8948 ;
  assign n8943 = n8942 ^ n7082 ;
  assign n8944 = n8943 ^ n7088 ;
  assign n8950 = n8949 ^ n8944 ;
  assign n8953 = n8952 ^ n8950 ;
  assign n8931 = n4393 & n5263 ;
  assign n8936 = n4899 & n5097 ;
  assign n8937 = n8936 ^ n4701 ;
  assign n8938 = n8931 & n8937 ;
  assign n8954 = n8953 ^ n8938 ;
  assign n8930 = n5265 & n5277 ;
  assign n8955 = n8954 ^ n8930 ;
  assign n8925 = n5283 ^ n5097 ;
  assign n8926 = n8925 ^ n5283 ;
  assign n8927 = n7840 & ~n8926 ;
  assign n8928 = n8927 ^ n5283 ;
  assign n8929 = ~n5263 & n8928 ;
  assign n8956 = n8955 ^ n8929 ;
  assign n8957 = n8956 ^ n5267 ;
  assign n8958 = n8957 ^ n4928 ;
  assign n8924 = n7064 & n7076 ;
  assign n8959 = n8958 ^ n8924 ;
  assign n8960 = n8959 ^ x112 ;
  assign n8978 = n8969 ^ n8960 ;
  assign n8999 = n8960 ^ n8898 ;
  assign n9000 = ~n8978 & n8999 ;
  assign n9001 = n9000 ^ n8922 ;
  assign n9002 = ~n8897 & n9001 ;
  assign n8894 = n8093 ^ x115 ;
  assign n7529 = n7264 & n7528 ;
  assign n7530 = n7529 ^ n7274 ;
  assign n7531 = n7530 ^ n5061 ;
  assign n7532 = n7531 ^ n7527 ;
  assign n7511 = n7261 ^ n7242 ;
  assign n7512 = n7511 ^ n7261 ;
  assign n7513 = n7261 ^ n7162 ;
  assign n7514 = n7513 ^ n7261 ;
  assign n7515 = n7512 & n7514 ;
  assign n7516 = n7515 ^ n7261 ;
  assign n7517 = n7277 & n7516 ;
  assign n7518 = n7517 ^ n7327 ;
  assign n7498 = n7293 ^ n7259 ;
  assign n7497 = n7279 ^ n7271 ;
  assign n7499 = n7498 ^ n7497 ;
  assign n7493 = n7263 ^ n7245 ;
  assign n7494 = n7493 ^ n7249 ;
  assign n7495 = n7494 ^ n7239 ;
  assign n7496 = ~n7161 & n7495 ;
  assign n7500 = n7499 ^ n7496 ;
  assign n7510 = n7500 ^ n7261 ;
  assign n7519 = n7518 ^ n7510 ;
  assign n7503 = n7502 ^ n7270 ;
  assign n7504 = n7503 ^ n7250 ;
  assign n7505 = n7504 ^ n7500 ;
  assign n7492 = n7278 ^ n7249 ;
  assign n7501 = n7500 ^ n7492 ;
  assign n7506 = n7505 ^ n7501 ;
  assign n7507 = ~n7161 & n7506 ;
  assign n7508 = n7507 ^ n7505 ;
  assign n7509 = ~n7162 & n7508 ;
  assign n7520 = n7519 ^ n7509 ;
  assign n7521 = ~n7491 & ~n7520 ;
  assign n7533 = n7532 ^ n7521 ;
  assign n8895 = n7533 ^ x97 ;
  assign n8980 = n8960 & n8969 ;
  assign n8968 = n8922 ^ n8897 ;
  assign n8970 = n8968 & ~n8969 ;
  assign n8979 = n8978 ^ n8970 ;
  assign n8981 = n8980 ^ n8979 ;
  assign n8961 = n8960 ^ n8897 ;
  assign n8982 = n8981 ^ n8961 ;
  assign n8991 = n8960 ^ n8922 ;
  assign n9008 = n8982 & n8991 ;
  assign n9009 = n9008 ^ n8961 ;
  assign n8899 = n8898 ^ n8897 ;
  assign n8976 = ~n8899 & n8960 ;
  assign n8973 = n8897 & ~n8898 ;
  assign n8974 = ~n8960 & n8973 ;
  assign n8971 = n8968 ^ n8960 ;
  assign n8972 = ~n8970 & ~n8971 ;
  assign n8975 = n8974 ^ n8972 ;
  assign n8977 = n8976 ^ n8975 ;
  assign n8983 = n8982 ^ n8977 ;
  assign n9514 = n9009 ^ n8983 ;
  assign n9515 = n8895 & ~n9514 ;
  assign n9516 = n9515 ^ n8983 ;
  assign n8923 = n8922 ^ n8899 ;
  assign n8964 = n8899 & n8961 ;
  assign n8965 = n8964 ^ n8897 ;
  assign n8966 = n8923 & n8965 ;
  assign n8967 = n8966 ^ n8897 ;
  assign n9517 = n9516 ^ n8967 ;
  assign n8995 = n8976 ^ n8974 ;
  assign n8992 = n8980 ^ n8897 ;
  assign n8993 = ~n8991 & n8992 ;
  assign n8994 = n8993 ^ n8969 ;
  assign n8996 = n8995 ^ n8994 ;
  assign n8990 = n8898 & n8922 ;
  assign n8997 = n8996 ^ n8990 ;
  assign n8998 = n8997 ^ n8975 ;
  assign n9136 = n9002 ^ n8998 ;
  assign n9137 = n9136 ^ n8967 ;
  assign n9518 = n9517 ^ n9137 ;
  assign n9519 = n9518 ^ n9517 ;
  assign n9522 = ~n8895 & ~n9519 ;
  assign n9523 = n9522 ^ n9517 ;
  assign n9524 = n8894 & n9523 ;
  assign n9525 = n9524 ^ n9516 ;
  assign n9526 = ~n9002 & ~n9525 ;
  assign n9527 = n9526 ^ n5096 ;
  assign n10131 = n9527 ^ x69 ;
  assign n10142 = n10088 ^ n10087 ;
  assign n10175 = n10123 & ~n10142 ;
  assign n10159 = n10123 & n10128 ;
  assign n10161 = n10160 ^ n10159 ;
  assign n10163 = n10162 ^ n10161 ;
  assign n10168 = n10167 ^ n10163 ;
  assign n10176 = n10175 ^ n10168 ;
  assign n10174 = n10173 ^ n10089 ;
  assign n10177 = n10176 ^ n10174 ;
  assign n10172 = n10171 ^ n10162 ;
  assign n10178 = n10177 ^ n10172 ;
  assign n10179 = ~n10131 & n10178 ;
  assign n10182 = n10181 ^ n10179 ;
  assign n8465 = n8069 ^ x98 ;
  assign n8466 = n6277 ^ x89 ;
  assign n8467 = n8465 & n8466 ;
  assign n8468 = n8467 ^ n8465 ;
  assign n8469 = n8468 ^ n8466 ;
  assign n8481 = n5724 ^ n5707 ;
  assign n8482 = n8481 ^ n5748 ;
  assign n8478 = n7005 ^ n5740 ;
  assign n8479 = n8478 ^ n5750 ;
  assign n8480 = ~n8086 & ~n8479 ;
  assign n8483 = n8482 ^ n8480 ;
  assign n8473 = n5744 ^ n5736 ;
  assign n8492 = n8483 ^ n8473 ;
  assign n8487 = n8073 ^ n5719 ;
  assign n8488 = n5349 & n8487 ;
  assign n8489 = n8488 ^ n8482 ;
  assign n8484 = n8483 ^ n5736 ;
  assign n8485 = n8484 ^ n8483 ;
  assign n8490 = n8489 ^ n8485 ;
  assign n8491 = n8490 ^ n8484 ;
  assign n8493 = n8492 ^ n8491 ;
  assign n8471 = n5744 ^ n5721 ;
  assign n8477 = ~n5379 & n8471 ;
  assign n8494 = n8493 ^ n8477 ;
  assign n8495 = n5777 & n8494 ;
  assign n8496 = n8495 ^ n8491 ;
  assign n8497 = ~n8088 & ~n8496 ;
  assign n8470 = n7042 ^ n5133 ;
  assign n8498 = n8497 ^ n8470 ;
  assign n8499 = n8498 ^ x65 ;
  assign n8500 = n8149 ^ x104 ;
  assign n8501 = n8499 & ~n8500 ;
  assign n8502 = n8501 ^ n8499 ;
  assign n8503 = n5347 ^ x113 ;
  assign n8525 = n7001 ^ n5168 ;
  assign n8210 = n6915 & ~n6992 ;
  assign n8211 = n8210 ^ n7655 ;
  assign n8522 = n8211 ^ n7637 ;
  assign n8212 = n6968 & n6996 ;
  assign n8213 = n8212 ^ n6944 ;
  assign n8504 = ~n7688 & ~n8213 ;
  assign n8519 = n6935 & ~n6992 ;
  assign n8517 = ~n6963 & n6976 ;
  assign n8515 = n6967 & n6996 ;
  assign n8512 = n6919 ^ n6915 ;
  assign n8513 = n6991 & n8512 ;
  assign n8508 = n7642 ^ n6967 ;
  assign n8505 = n6979 ^ n6946 ;
  assign n8506 = n8505 ^ n6948 ;
  assign n8507 = ~n6923 & ~n8506 ;
  assign n8509 = n8508 ^ n8507 ;
  assign n8510 = ~n6860 & ~n8509 ;
  assign n8511 = n8510 ^ n8507 ;
  assign n8514 = n8513 ^ n8511 ;
  assign n8516 = n8515 ^ n8514 ;
  assign n8518 = n8517 ^ n8516 ;
  assign n8520 = n8519 ^ n8518 ;
  assign n8521 = n8504 & ~n8520 ;
  assign n8523 = n8522 ^ n8521 ;
  assign n8524 = ~n6994 & n8523 ;
  assign n8526 = n8525 ^ n8524 ;
  assign n8527 = n8526 ^ x123 ;
  assign n8528 = n8503 & ~n8527 ;
  assign n8555 = n8502 & n8528 ;
  assign n8556 = n8555 ^ n8528 ;
  assign n8532 = n8501 ^ n8500 ;
  assign n8551 = n8532 ^ n8499 ;
  assign n8552 = n8528 & n8551 ;
  assign n8533 = n8528 & ~n8532 ;
  assign n8554 = n8552 ^ n8533 ;
  assign n8557 = n8556 ^ n8554 ;
  assign n8547 = n8528 ^ n8503 ;
  assign n8548 = n8502 & n8547 ;
  assign n8558 = n8557 ^ n8548 ;
  assign n8596 = n8558 ^ n8551 ;
  assign n8529 = n8528 ^ n8527 ;
  assign n8562 = n8502 & ~n8529 ;
  assign n8543 = n8501 & ~n8529 ;
  assign n8563 = n8562 ^ n8543 ;
  assign n8537 = ~n8529 & ~n8532 ;
  assign n8564 = n8563 ^ n8537 ;
  assign n8550 = n8501 & n8547 ;
  assign n8553 = n8552 ^ n8550 ;
  assign n8559 = n8558 ^ n8553 ;
  assign n8541 = n8527 ^ n8500 ;
  assign n8542 = n8503 & n8541 ;
  assign n8544 = n8543 ^ n8542 ;
  assign n8539 = n8527 ^ n8503 ;
  assign n8540 = n8539 ^ n8500 ;
  assign n8545 = n8544 ^ n8540 ;
  assign n8530 = n8529 ^ n8503 ;
  assign n8531 = n8502 & n8530 ;
  assign n8538 = n8537 ^ n8531 ;
  assign n8546 = n8545 ^ n8538 ;
  assign n8549 = n8548 ^ n8546 ;
  assign n8560 = n8559 ^ n8549 ;
  assign n8561 = n8560 ^ n8539 ;
  assign n8565 = n8564 ^ n8561 ;
  assign n8597 = n8596 ^ n8565 ;
  assign n9753 = n8597 ^ n8562 ;
  assign n9752 = n8555 ^ n8533 ;
  assign n9754 = n9753 ^ n9752 ;
  assign n9755 = ~n8469 & n9754 ;
  assign n8536 = n8466 ^ n8465 ;
  assign n8578 = n8547 & n8551 ;
  assign n9465 = n8578 ^ n8543 ;
  assign n9466 = n8543 ^ n8466 ;
  assign n9467 = n9466 ^ n8543 ;
  assign n9468 = n9465 & ~n9467 ;
  assign n9469 = n9468 ^ n8543 ;
  assign n9470 = n8536 & n9469 ;
  assign n8588 = n8564 ^ n8529 ;
  assign n8610 = n8469 ^ n8465 ;
  assign n8611 = ~n8588 & n8610 ;
  assign n9750 = n9470 ^ n8611 ;
  assign n9751 = n9750 ^ n8538 ;
  assign n9756 = n9755 ^ n9751 ;
  assign n9742 = n8578 ^ n8538 ;
  assign n8585 = n8501 & n8530 ;
  assign n8586 = n8585 ^ n8546 ;
  assign n8584 = n8531 ^ n8530 ;
  assign n8587 = n8586 ^ n8584 ;
  assign n9743 = n9742 ^ n8587 ;
  assign n9744 = n9743 ^ n8538 ;
  assign n9745 = n8538 ^ n8465 ;
  assign n9746 = n9745 ^ n8538 ;
  assign n9747 = ~n9744 & ~n9746 ;
  assign n9748 = n9747 ^ n8538 ;
  assign n9749 = n8466 & n9748 ;
  assign n9757 = n9756 ^ n9749 ;
  assign n9735 = n8588 ^ n8544 ;
  assign n9736 = n9735 ^ n8556 ;
  assign n9737 = n8556 ^ n8466 ;
  assign n9738 = n9737 ^ n8556 ;
  assign n9739 = ~n9736 & n9738 ;
  assign n9740 = n9739 ^ n8556 ;
  assign n9741 = n8465 & n9740 ;
  assign n9758 = n9757 ^ n9741 ;
  assign n9759 = n9758 ^ n8585 ;
  assign n8572 = n8562 ^ n8546 ;
  assign n8573 = n8562 ^ n8466 ;
  assign n8574 = n8573 ^ n8562 ;
  assign n8575 = ~n8572 & n8574 ;
  assign n8576 = n8575 ^ n8562 ;
  assign n8577 = n8465 & n8576 ;
  assign n9760 = n9759 ^ n8577 ;
  assign n9761 = n9760 ^ n5262 ;
  assign n9734 = n8559 & n8610 ;
  assign n9762 = n9761 ^ n9734 ;
  assign n9733 = n8468 & ~n8587 ;
  assign n9763 = n9762 ^ n9733 ;
  assign n9726 = n8585 ^ n8469 ;
  assign n9727 = n8546 ^ n8467 ;
  assign n9730 = ~n8585 & n9727 ;
  assign n9731 = n9730 ^ n8467 ;
  assign n9732 = ~n9726 & ~n9731 ;
  assign n9764 = n9763 ^ n9732 ;
  assign n10126 = n9764 ^ x118 ;
  assign n10190 = n10182 ^ n10126 ;
  assign n10186 = n10126 & n10131 ;
  assign n10140 = n10139 ^ n10122 ;
  assign n10145 = n10088 & n10140 ;
  assign n10143 = n10140 & ~n10142 ;
  assign n10141 = n10128 & n10140 ;
  assign n10144 = n10143 ^ n10141 ;
  assign n10146 = n10145 ^ n10144 ;
  assign n10124 = n10123 ^ n10122 ;
  assign n10130 = ~n10124 & n10129 ;
  assign n10187 = n10146 ^ n10130 ;
  assign n10188 = n10187 ^ n10163 ;
  assign n10189 = n10186 & n10188 ;
  assign n10191 = n10190 ^ n10189 ;
  assign n10138 = n10131 ^ n10126 ;
  assign n10185 = ~n10138 & ~n10175 ;
  assign n10192 = n10191 ^ n10185 ;
  assign n10169 = n10131 & n10168 ;
  assign n10170 = n10169 ^ n10168 ;
  assign n10183 = n10182 ^ n10170 ;
  assign n10184 = n10126 & n10183 ;
  assign n10193 = n10192 ^ n10184 ;
  assign n10149 = ~n10124 & n10128 ;
  assign n10125 = n10088 & ~n10124 ;
  assign n10150 = n10149 ^ n10125 ;
  assign n10148 = n10130 ^ n10124 ;
  assign n10151 = n10150 ^ n10148 ;
  assign n10147 = n10146 ^ n10140 ;
  assign n10152 = n10151 ^ n10147 ;
  assign n10153 = n10152 ^ n10145 ;
  assign n10154 = n10145 ^ n10131 ;
  assign n10155 = n10154 ^ n10145 ;
  assign n10156 = ~n10153 & n10155 ;
  assign n10157 = n10156 ^ n10145 ;
  assign n10158 = n10138 & ~n10157 ;
  assign n10194 = n10193 ^ n10158 ;
  assign n10127 = n10126 ^ n10125 ;
  assign n10132 = n10131 ^ n10130 ;
  assign n10133 = n10131 ^ n10125 ;
  assign n10134 = n10133 ^ n10131 ;
  assign n10135 = n10132 & ~n10134 ;
  assign n10136 = n10135 ^ n10131 ;
  assign n10137 = ~n10127 & ~n10136 ;
  assign n10195 = n10194 ^ n10137 ;
  assign n10196 = n10149 ^ n10145 ;
  assign n10197 = n10196 ^ n10152 ;
  assign n10198 = n10196 ^ n10126 ;
  assign n10199 = n10198 ^ n10196 ;
  assign n10200 = ~n10197 & n10199 ;
  assign n10201 = n10200 ^ n10196 ;
  assign n10202 = ~n10131 & n10201 ;
  assign n10203 = ~n10195 & ~n10202 ;
  assign n10204 = n10203 ^ n5347 ;
  assign n10205 = n10204 ^ x81 ;
  assign n9135 = n8995 ^ n8973 ;
  assign n9138 = n9137 ^ n9135 ;
  assign n9139 = n9138 ^ n8972 ;
  assign n9140 = n9139 ^ n9138 ;
  assign n9141 = n9138 ^ n9000 ;
  assign n9142 = n9141 ^ n9138 ;
  assign n9143 = ~n9140 & ~n9142 ;
  assign n9144 = n9143 ^ n9138 ;
  assign n9145 = ~n8894 & n9144 ;
  assign n9146 = n9145 ^ n9138 ;
  assign n9133 = n8894 & n8997 ;
  assign n9134 = n9133 ^ n8994 ;
  assign n9147 = n9146 ^ n9134 ;
  assign n9148 = ~n8895 & ~n9147 ;
  assign n9149 = n9148 ^ n9146 ;
  assign n9150 = n9149 ^ n8895 ;
  assign n9151 = n9150 ^ n9146 ;
  assign n9152 = n9151 ^ n9134 ;
  assign n9153 = n9152 ^ n6076 ;
  assign n10206 = n9153 ^ x110 ;
  assign n8589 = n8588 ^ n8587 ;
  assign n8590 = n8589 ^ n8578 ;
  assign n8591 = n8578 ^ n8466 ;
  assign n8592 = n8591 ^ n8578 ;
  assign n8593 = n8590 & ~n8592 ;
  assign n8594 = n8593 ^ n8578 ;
  assign n8595 = n8536 & n8594 ;
  assign n10221 = ~n8469 & n8533 ;
  assign n8579 = ~n8468 & ~n8578 ;
  assign n10218 = n8550 ^ n8469 ;
  assign n10219 = ~n8579 & ~n10218 ;
  assign n10210 = n9752 ^ n8553 ;
  assign n10209 = n8585 ^ n8563 ;
  assign n10211 = n10210 ^ n10209 ;
  assign n10212 = n10210 ^ n8466 ;
  assign n10213 = n10212 ^ n10210 ;
  assign n10214 = n10211 & ~n10213 ;
  assign n10215 = n10214 ^ n10210 ;
  assign n10216 = ~n8536 & n10215 ;
  assign n10217 = n10216 ^ n8558 ;
  assign n10220 = n10219 ^ n10217 ;
  assign n10222 = n10221 ^ n10220 ;
  assign n10231 = n10222 ^ n9750 ;
  assign n10223 = n10222 ^ n10216 ;
  assign n9481 = n8585 ^ n8562 ;
  assign n10226 = n10223 ^ n9481 ;
  assign n10227 = n10226 ^ n10223 ;
  assign n10228 = ~n8465 & n10227 ;
  assign n10229 = n10228 ^ n10223 ;
  assign n10230 = n8466 & n10229 ;
  assign n10232 = n10231 ^ n10230 ;
  assign n10207 = n9481 ^ n8538 ;
  assign n10208 = n8467 & n10207 ;
  assign n10233 = n10232 ^ n10208 ;
  assign n9483 = n8548 ^ n8533 ;
  assign n10234 = n9483 ^ n8597 ;
  assign n10235 = n10234 ^ n8537 ;
  assign n10236 = n8537 ^ n8466 ;
  assign n10237 = n10236 ^ n8537 ;
  assign n10238 = n10235 & n10237 ;
  assign n10239 = n10238 ^ n8537 ;
  assign n10240 = n8536 & n10239 ;
  assign n10241 = ~n10233 & ~n10240 ;
  assign n10242 = ~n8595 & n10241 ;
  assign n10244 = ~n8466 & ~n8546 ;
  assign n10245 = n10242 & n10244 ;
  assign n10243 = n10242 ^ n6305 ;
  assign n10246 = n10245 ^ n10243 ;
  assign n10247 = n10246 ^ x77 ;
  assign n10248 = n10206 & ~n10247 ;
  assign n10303 = n10248 ^ n10247 ;
  assign n10304 = n10303 ^ n10206 ;
  assign n7422 = n7421 ^ n7370 ;
  assign n7423 = n7370 ^ n7158 ;
  assign n7424 = n7423 ^ n7370 ;
  assign n7425 = n7422 & ~n7424 ;
  assign n7426 = n7425 ^ n7370 ;
  assign n7427 = ~n7118 & n7426 ;
  assign n10249 = ~n7427 & ~n9712 ;
  assign n10267 = n7345 ^ n7341 ;
  assign n10266 = n7378 ^ n7375 ;
  assign n10268 = n10267 ^ n10266 ;
  assign n10269 = ~n7158 & n10268 ;
  assign n10270 = n10269 ^ n10267 ;
  assign n10274 = n10270 ^ n8883 ;
  assign n10252 = n7395 ^ n7376 ;
  assign n10251 = n7391 ^ n7354 ;
  assign n10253 = n10252 ^ n10251 ;
  assign n10254 = n10251 ^ n7158 ;
  assign n10255 = n10254 ^ n10251 ;
  assign n10256 = n10253 & n10255 ;
  assign n10257 = n10256 ^ n10251 ;
  assign n10258 = n7389 & ~n10257 ;
  assign n10275 = n10274 ^ n10258 ;
  assign n10264 = n8870 ^ n7393 ;
  assign n10265 = n10264 ^ n7407 ;
  assign n10271 = n10270 ^ n10265 ;
  assign n10260 = n7393 ^ n7341 ;
  assign n10261 = n10260 ^ n7373 ;
  assign n10262 = n10261 ^ n8870 ;
  assign n10263 = ~n7158 & ~n10262 ;
  assign n10272 = n10271 ^ n10263 ;
  assign n10273 = ~n7389 & n10272 ;
  assign n10276 = n10275 ^ n10273 ;
  assign n10259 = n7347 & ~n7403 ;
  assign n10277 = n10276 ^ n10259 ;
  assign n10250 = n7118 & n7349 ;
  assign n10282 = n10277 ^ n10250 ;
  assign n10283 = n10249 & ~n10282 ;
  assign n10284 = n10283 ^ n6356 ;
  assign n10285 = n10284 ^ x92 ;
  assign n8745 = n8744 ^ n6817 ;
  assign n8746 = n8745 ^ n6833 ;
  assign n6787 = n6786 ^ n6780 ;
  assign n8741 = n6811 ^ n6787 ;
  assign n8739 = n6809 ^ n6800 ;
  assign n6838 = n6837 ^ n6833 ;
  assign n8740 = n8739 ^ n6838 ;
  assign n8742 = n8741 ^ n8740 ;
  assign n8743 = ~n5348 & ~n8742 ;
  assign n8747 = n8746 ^ n8743 ;
  assign n8735 = n6834 ^ n6799 ;
  assign n8736 = n8735 ^ n6780 ;
  assign n8733 = n6833 ^ n6796 ;
  assign n8734 = n8733 ^ n6837 ;
  assign n8737 = n8736 ^ n8734 ;
  assign n8738 = ~n5348 & n8737 ;
  assign n8748 = n8747 ^ n8738 ;
  assign n8749 = n5786 & ~n8748 ;
  assign n8750 = n8749 ^ n8743 ;
  assign n6821 = n6820 ^ n6792 ;
  assign n8730 = n6821 ^ n6809 ;
  assign n8731 = n8730 ^ n6830 ;
  assign n8732 = n5789 & ~n8731 ;
  assign n8751 = n8750 ^ n8732 ;
  assign n6784 = n5789 & n6783 ;
  assign n8752 = n8751 ^ n6784 ;
  assign n8729 = n6785 & n6793 ;
  assign n8753 = n8752 ^ n8729 ;
  assign n8760 = ~n8753 & ~n8759 ;
  assign n8761 = n8760 ^ n6054 ;
  assign n10286 = n8761 ^ x70 ;
  assign n10287 = ~n10285 & n10286 ;
  assign n10289 = n10287 ^ n10286 ;
  assign n10290 = n10248 & n10289 ;
  assign n10291 = n10290 ^ n10289 ;
  assign n10308 = n10291 ^ n10286 ;
  assign n10309 = ~n10304 & n10308 ;
  assign n10310 = n10309 ^ n10308 ;
  assign n10298 = n10289 ^ n10285 ;
  assign n10305 = n10298 & n10304 ;
  assign n10301 = n10248 ^ n10206 ;
  assign n10302 = n10298 & n10301 ;
  assign n10306 = n10305 ^ n10302 ;
  assign n10299 = n10248 & n10298 ;
  assign n10300 = n10299 ^ n10298 ;
  assign n10307 = n10306 ^ n10300 ;
  assign n10311 = n10310 ^ n10307 ;
  assign n8205 = n6072 ^ x85 ;
  assign n8204 = n7828 ^ x67 ;
  assign n8638 = n8205 ^ n8204 ;
  assign n8261 = n7320 ^ n7279 ;
  assign n8262 = n7162 & ~n7277 ;
  assign n8263 = n8261 & n8262 ;
  assign n8264 = n8263 ^ n7277 ;
  assign n8266 = n7284 & ~n8264 ;
  assign n8269 = n7251 & ~n7270 ;
  assign n8270 = n8266 & n8269 ;
  assign n8267 = n8266 ^ n7244 ;
  assign n8268 = n8267 ^ n8263 ;
  assign n8271 = n8270 ^ n8268 ;
  assign n8259 = n8045 ^ n7254 ;
  assign n8260 = n7528 & n8259 ;
  assign n8272 = n8271 ^ n8260 ;
  assign n8252 = n7289 ^ n7236 ;
  assign n8253 = n8252 ^ n7502 ;
  assign n8254 = n7502 ^ n7162 ;
  assign n8255 = n8254 ^ n7502 ;
  assign n8256 = ~n8253 & n8255 ;
  assign n8257 = n8256 ^ n7502 ;
  assign n8258 = ~n7161 & n8257 ;
  assign n8273 = n8272 ^ n8258 ;
  assign n8274 = ~n8062 & ~n8273 ;
  assign n8275 = ~n7530 & n8274 ;
  assign n8276 = ~n7252 & n8275 ;
  assign n8277 = ~n7527 & n8276 ;
  assign n8278 = n8277 ^ n5612 ;
  assign n8279 = n8278 ^ x116 ;
  assign n8280 = n7792 ^ x68 ;
  assign n8281 = n8279 & ~n8280 ;
  assign n8231 = n7689 ^ n6998 ;
  assign n8218 = n7672 ^ n6978 ;
  assign n8219 = n8218 ^ n6916 ;
  assign n8220 = n6860 & n8219 ;
  assign n8221 = n8220 ^ n7672 ;
  assign n8232 = n8231 ^ n8221 ;
  assign n8217 = n6972 ^ n6919 ;
  assign n8222 = n8221 ^ n8217 ;
  assign n8223 = n8222 ^ n6919 ;
  assign n8224 = n8223 ^ n6976 ;
  assign n8225 = n8224 ^ n8222 ;
  assign n8226 = n8222 ^ n6923 ;
  assign n8227 = n8226 ^ n8222 ;
  assign n8228 = n8225 & n8227 ;
  assign n8229 = n8228 ^ n8222 ;
  assign n8230 = n6963 & ~n8229 ;
  assign n8233 = n8232 ^ n8230 ;
  assign n8215 = n6920 ^ n6911 ;
  assign n8216 = ~n6992 & n8215 ;
  assign n8234 = n8233 ^ n8216 ;
  assign n8214 = n6967 & n6993 ;
  assign n8235 = n8234 ^ n8214 ;
  assign n8236 = n6991 ^ n6919 ;
  assign n8237 = n8236 ^ n8235 ;
  assign n8238 = n6947 ^ n6923 ;
  assign n8239 = ~n6991 & ~n8238 ;
  assign n8240 = n8239 ^ n6947 ;
  assign n8241 = ~n8237 & ~n8240 ;
  assign n8242 = n8241 ^ n6991 ;
  assign n8243 = n8235 & ~n8242 ;
  assign n8244 = ~n8213 & n8243 ;
  assign n8245 = ~n8211 & n8244 ;
  assign n8246 = ~n6935 & n8245 ;
  assign n8247 = n8246 ^ n5582 ;
  assign n8248 = n8247 ^ x102 ;
  assign n8249 = n5785 ^ x109 ;
  assign n8250 = n8248 & n8249 ;
  assign n8251 = n8250 ^ n8248 ;
  assign n8284 = n8251 ^ n8249 ;
  assign n8289 = n8281 & ~n8284 ;
  assign n8282 = n8281 ^ n8280 ;
  assign n8285 = n8284 ^ n8248 ;
  assign n8286 = ~n8282 & n8285 ;
  assign n8307 = n8289 ^ n8286 ;
  assign n8291 = n8282 ^ n8279 ;
  assign n8293 = n8291 ^ n8280 ;
  assign n8302 = n8250 & n8293 ;
  assign n8294 = ~n8284 & n8293 ;
  assign n8303 = n8302 ^ n8294 ;
  assign n8297 = n8285 & n8293 ;
  assign n8296 = ~n8284 & n8291 ;
  assign n8298 = n8297 ^ n8296 ;
  assign n8304 = n8303 ^ n8298 ;
  assign n8301 = n8296 ^ n8293 ;
  assign n8305 = n8304 ^ n8301 ;
  assign n8306 = n8305 ^ n8297 ;
  assign n8308 = n8307 ^ n8306 ;
  assign n8292 = n8251 & n8291 ;
  assign n8295 = n8294 ^ n8292 ;
  assign n8299 = n8298 ^ n8295 ;
  assign n8300 = n8299 ^ n8249 ;
  assign n8309 = n8308 ^ n8300 ;
  assign n9270 = n8309 ^ n8303 ;
  assign n8313 = n8281 & n8285 ;
  assign n8311 = n8250 & ~n8282 ;
  assign n8310 = n8309 ^ n8282 ;
  assign n8312 = n8311 ^ n8310 ;
  assign n8314 = n8313 ^ n8312 ;
  assign n8290 = n8289 ^ n8281 ;
  assign n8315 = n8314 ^ n8290 ;
  assign n8349 = n8315 ^ n8312 ;
  assign n9265 = n8349 ^ n8309 ;
  assign n9266 = n8349 ^ n8205 ;
  assign n9267 = n8638 & n9266 ;
  assign n9268 = n9267 ^ n8205 ;
  assign n9269 = ~n9265 & ~n9268 ;
  assign n9271 = n9270 ^ n9269 ;
  assign n9272 = n9271 ^ n8314 ;
  assign n9273 = n9272 ^ n8308 ;
  assign n9274 = n9273 ^ n9271 ;
  assign n9275 = n9271 ^ n8205 ;
  assign n9276 = n9275 ^ n9271 ;
  assign n9277 = n9274 & ~n9276 ;
  assign n9278 = n9277 ^ n9271 ;
  assign n9279 = n8638 & ~n9278 ;
  assign n9280 = n9279 ^ n9271 ;
  assign n9256 = n8315 ^ n8311 ;
  assign n8283 = n8251 & ~n8282 ;
  assign n8287 = n8286 ^ n8283 ;
  assign n8288 = n8287 ^ n8282 ;
  assign n9257 = n9256 ^ n8288 ;
  assign n8318 = n8250 & n8291 ;
  assign n8324 = n8318 ^ n8295 ;
  assign n8323 = n8303 ^ n8296 ;
  assign n8325 = n8324 ^ n8323 ;
  assign n8326 = n8325 ^ n8291 ;
  assign n8327 = n8326 ^ n8302 ;
  assign n9258 = n9257 ^ n8327 ;
  assign n9259 = n8205 & ~n9258 ;
  assign n9260 = n9259 ^ n8327 ;
  assign n9261 = ~n8204 & n9260 ;
  assign n9255 = ~n8205 & n8292 ;
  assign n9262 = n9261 ^ n9255 ;
  assign n9263 = n9262 ^ n6198 ;
  assign n8328 = n8327 ^ n8306 ;
  assign n8648 = n8328 ^ n8288 ;
  assign n8649 = n8288 ^ n8205 ;
  assign n8650 = n8649 ^ n8288 ;
  assign n8651 = ~n8648 & n8650 ;
  assign n8652 = n8651 ^ n8288 ;
  assign n8653 = ~n8204 & ~n8652 ;
  assign n9264 = n9263 ^ n8653 ;
  assign n9281 = n9280 ^ n9264 ;
  assign n8616 = n8292 ^ n8289 ;
  assign n8344 = n8313 ^ n8296 ;
  assign n9251 = n8616 ^ n8344 ;
  assign n9252 = ~n8204 & n9251 ;
  assign n9253 = n9252 ^ n8289 ;
  assign n9254 = n8205 & n9253 ;
  assign n9284 = n9281 ^ n9254 ;
  assign n9285 = n9284 ^ n9264 ;
  assign n9286 = n8204 & n8318 ;
  assign n9287 = n9285 & n9286 ;
  assign n9288 = n9287 ^ n9284 ;
  assign n10293 = n9288 ^ x109 ;
  assign n8715 = n8174 ^ n8117 ;
  assign n8716 = n8150 & n8715 ;
  assign n8706 = n8150 ^ n8097 ;
  assign n8707 = n8706 ^ n8097 ;
  assign n8709 = n8098 & n8707 ;
  assign n8710 = n8709 ^ n8097 ;
  assign n8711 = ~n7982 & n8710 ;
  assign n8167 = n8118 ^ n8098 ;
  assign n8170 = ~n8150 & n8167 ;
  assign n8171 = n8170 ^ n8098 ;
  assign n8172 = ~n8166 & n8171 ;
  assign n8712 = n8711 ^ n8172 ;
  assign n8697 = n8070 ^ n8003 ;
  assign n8698 = n8095 ^ n8030 ;
  assign n8699 = ~n8150 & n8698 ;
  assign n8700 = ~n8697 & n8699 ;
  assign n8705 = n8700 ^ n8097 ;
  assign n8713 = n8712 ^ n8705 ;
  assign n8714 = n8713 ^ n8103 ;
  assign n8717 = n8716 ^ n8714 ;
  assign n8722 = n8717 ^ n8185 ;
  assign n8694 = n8189 ^ n8109 ;
  assign n8703 = n8702 ^ n8694 ;
  assign n8701 = n8700 ^ n8158 ;
  assign n8704 = n8703 ^ n8701 ;
  assign n8718 = n8717 ^ n8704 ;
  assign n8719 = n8718 ^ n8713 ;
  assign n8695 = n8694 ^ n8114 ;
  assign n8696 = n8150 & ~n8695 ;
  assign n8720 = n8719 ^ n8696 ;
  assign n8721 = n8166 & n8720 ;
  assign n8723 = n8722 ^ n8721 ;
  assign n8724 = ~n8693 & ~n8723 ;
  assign n8725 = n8724 ^ n5918 ;
  assign n10294 = n8725 ^ x91 ;
  assign n10295 = n10293 & n10294 ;
  assign n10296 = n10295 ^ n10293 ;
  assign n10313 = n10298 ^ n10286 ;
  assign n10314 = n10248 & ~n10313 ;
  assign n10321 = n10295 & n10314 ;
  assign n10297 = n10296 ^ n10294 ;
  assign n10312 = n10297 ^ n10293 ;
  assign n10317 = n10301 & ~n10313 ;
  assign n10316 = ~n10303 & ~n10313 ;
  assign n10318 = n10317 ^ n10316 ;
  assign n10315 = n10314 ^ n10313 ;
  assign n10319 = n10318 ^ n10315 ;
  assign n10320 = n10312 & ~n10319 ;
  assign n10322 = n10321 ^ n10320 ;
  assign n10323 = n10317 ^ n10312 ;
  assign n10324 = n10305 ^ n10296 ;
  assign n10327 = n10312 & ~n10324 ;
  assign n10328 = n10327 ^ n10296 ;
  assign n10329 = n10323 & ~n10328 ;
  assign n10330 = n10329 ^ n10317 ;
  assign n10339 = n10287 & n10301 ;
  assign n10340 = n10294 & ~n10339 ;
  assign n10334 = n10319 ^ n10305 ;
  assign n10335 = n10334 ^ n10304 ;
  assign n10336 = n10335 ^ n10310 ;
  assign n10350 = n10336 ^ n10290 ;
  assign n10351 = n10350 ^ n10310 ;
  assign n10288 = n10248 & n10287 ;
  assign n10347 = n10310 ^ n10288 ;
  assign n10346 = n10339 ^ n10287 ;
  assign n10348 = n10347 ^ n10346 ;
  assign n10342 = n10316 ^ n10302 ;
  assign n10343 = n10342 ^ n10339 ;
  assign n10341 = n10318 ^ n10301 ;
  assign n10344 = n10343 ^ n10341 ;
  assign n10345 = n10344 ^ n10299 ;
  assign n10349 = n10348 ^ n10345 ;
  assign n10352 = n10351 ^ n10349 ;
  assign n10353 = ~n10293 & ~n10352 ;
  assign n10354 = n10353 ^ n10351 ;
  assign n10355 = n10340 & n10354 ;
  assign n10356 = n10355 ^ n10294 ;
  assign n10337 = n10336 ^ n10289 ;
  assign n10338 = n10296 & ~n10337 ;
  assign n10357 = n10356 ^ n10338 ;
  assign n10331 = n10319 ^ n10307 ;
  assign n10332 = n10331 ^ n10302 ;
  assign n10333 = ~n10297 & ~n10332 ;
  assign n10358 = n10357 ^ n10333 ;
  assign n10359 = n10348 ^ n10317 ;
  assign n10360 = n10317 ^ n10293 ;
  assign n10361 = n10360 ^ n10317 ;
  assign n10362 = n10359 & n10361 ;
  assign n10363 = n10362 ^ n10317 ;
  assign n10364 = ~n10294 & n10363 ;
  assign n10365 = ~n10358 & ~n10364 ;
  assign n10366 = n10294 ^ n10293 ;
  assign n10369 = n10342 ^ n10299 ;
  assign n10370 = n10294 & n10369 ;
  assign n10371 = n10370 ^ n10314 ;
  assign n10372 = ~n10366 & n10371 ;
  assign n10373 = n10372 ^ n10314 ;
  assign n10374 = n10365 & n10373 ;
  assign n10375 = n10374 ^ n10365 ;
  assign n10376 = ~n10330 & n10375 ;
  assign n10377 = ~n10322 & n10376 ;
  assign n10378 = n10296 & n10377 ;
  assign n10379 = n10311 & n10378 ;
  assign n10380 = n10379 ^ n10377 ;
  assign n10383 = n10380 ^ n8149 ;
  assign n10292 = n10291 ^ n10288 ;
  assign n10381 = ~n10297 & n10380 ;
  assign n10382 = n10292 & n10381 ;
  assign n10384 = n10383 ^ n10382 ;
  assign n10385 = n10384 ^ x72 ;
  assign n10386 = n10205 & n10385 ;
  assign n10392 = n10386 ^ n10205 ;
  assign n10395 = n10392 ^ n10385 ;
  assign n7534 = n7533 ^ x86 ;
  assign n7472 = n7471 ^ n7458 ;
  assign n7483 = n7482 ^ n7472 ;
  assign n7484 = n7483 ^ n6209 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7487 = n7486 ^ n5423 ;
  assign n7436 = n7435 ^ n6239 ;
  assign n7437 = n7436 ^ n6269 ;
  assign n7434 = n6199 ^ n6168 ;
  assign n7438 = n7437 ^ n7434 ;
  assign n7439 = ~n6078 & ~n7438 ;
  assign n7440 = n7439 ^ n6243 ;
  assign n7433 = n6242 ^ n6228 ;
  assign n7441 = n7440 ^ n7433 ;
  assign n7442 = n7441 ^ n6205 ;
  assign n7443 = n7442 ^ n6228 ;
  assign n7444 = n7443 ^ n7441 ;
  assign n7447 = n6078 & n7444 ;
  assign n7448 = n7447 ^ n7441 ;
  assign n7449 = n6213 & n7448 ;
  assign n7450 = n7449 ^ n7440 ;
  assign n7451 = ~n6253 & ~n7450 ;
  assign n7488 = n7487 ^ n7451 ;
  assign n7489 = n7488 ^ x108 ;
  assign n7610 = n7534 ^ n7489 ;
  assign n7538 = n7117 ^ x126 ;
  assign n7558 = n7557 ^ n6673 ;
  assign n7559 = n7558 ^ n7549 ;
  assign n7555 = n6701 ^ n6610 ;
  assign n7556 = n6668 & ~n7555 ;
  assign n7560 = n7559 ^ n7556 ;
  assign n7561 = ~n6647 & ~n7560 ;
  assign n7550 = n7549 ^ n6684 ;
  assign n7544 = n6689 ^ n6687 ;
  assign n7545 = n7544 ^ n6714 ;
  assign n7546 = n6647 & ~n7545 ;
  assign n7551 = n7550 ^ n7546 ;
  assign n7552 = n7551 ^ n7549 ;
  assign n7553 = ~n6698 & ~n7552 ;
  assign n7554 = n7553 ^ n7550 ;
  assign n7562 = n7561 ^ n7554 ;
  assign n7563 = n7562 ^ n6771 ;
  assign n7564 = n6704 ^ n6647 ;
  assign n7565 = n7564 ^ n6704 ;
  assign n7567 = ~n6668 & n7566 ;
  assign n7568 = n7567 ^ n6704 ;
  assign n7569 = n7565 & n7568 ;
  assign n7570 = n7569 ^ n6704 ;
  assign n7571 = n7563 & n7570 ;
  assign n7572 = n7571 ^ n7563 ;
  assign n7575 = n7572 ^ n6687 ;
  assign n7543 = n6701 ^ n6684 ;
  assign n7573 = n6669 & n7572 ;
  assign n7574 = ~n7543 & n7573 ;
  assign n7576 = n7575 ^ n7574 ;
  assign n7539 = n6720 ^ n6687 ;
  assign n7540 = ~n6755 & n7539 ;
  assign n7541 = n7540 ^ n6687 ;
  assign n7542 = ~n6698 & n7541 ;
  assign n7577 = n7576 ^ n7542 ;
  assign n7578 = n7577 ^ n6690 ;
  assign n7585 = n7578 & ~n7584 ;
  assign n7592 = n7585 & ~n7591 ;
  assign n7593 = n7592 ^ n5452 ;
  assign n7594 = n7593 ^ x93 ;
  assign n7611 = n7594 ^ n7489 ;
  assign n7612 = n7538 & n7611 ;
  assign n7613 = n7612 ^ n7489 ;
  assign n7614 = ~n7610 & n7613 ;
  assign n7615 = n7614 ^ n7534 ;
  assign n7535 = n7489 & ~n7534 ;
  assign n7536 = n7535 ^ n7489 ;
  assign n7595 = n7538 & n7594 ;
  assign n7601 = n7595 ^ n7538 ;
  assign n7602 = n7536 & n7601 ;
  assign n7537 = n7536 ^ n7534 ;
  assign n7609 = n7602 ^ n7537 ;
  assign n7616 = n7615 ^ n7609 ;
  assign n7604 = n7535 ^ n7534 ;
  assign n7596 = n7595 ^ n7594 ;
  assign n7607 = n7596 ^ n7538 ;
  assign n7608 = ~n7604 & ~n7607 ;
  assign n7617 = n7616 ^ n7608 ;
  assign n7605 = n7596 & ~n7604 ;
  assign n7606 = n7605 ^ n7604 ;
  assign n7618 = n7617 ^ n7606 ;
  assign n7432 = n7102 ^ x125 ;
  assign n7694 = n7693 ^ x76 ;
  assign n7730 = n7432 & ~n7694 ;
  assign n8689 = ~n7618 & n7730 ;
  assign n9183 = n8689 ^ n5551 ;
  assign n7700 = n7694 ^ n7432 ;
  assign n7701 = n7594 ^ n7538 ;
  assign n7702 = n7534 & ~n7701 ;
  assign n7703 = n7702 ^ n7534 ;
  assign n7621 = n7535 & n7601 ;
  assign n7627 = n7621 ^ n7618 ;
  assign n7628 = n7627 ^ n7605 ;
  assign n7598 = n7536 & n7595 ;
  assign n7629 = n7628 ^ n7598 ;
  assign n7623 = n7535 & n7595 ;
  assign n7624 = n7623 ^ n7535 ;
  assign n7620 = n7535 & ~n7607 ;
  assign n7622 = n7621 ^ n7620 ;
  assign n7625 = n7624 ^ n7622 ;
  assign n7626 = n7625 ^ n7621 ;
  assign n7630 = n7629 ^ n7626 ;
  assign n7619 = n7618 ^ n7596 ;
  assign n7631 = n7630 ^ n7619 ;
  assign n7597 = n7537 & n7596 ;
  assign n7599 = n7598 ^ n7597 ;
  assign n7632 = n7631 ^ n7599 ;
  assign n7603 = n7602 ^ n7597 ;
  assign n7633 = n7632 ^ n7603 ;
  assign n7704 = n7703 ^ n7633 ;
  assign n7705 = n7700 & n7704 ;
  assign n7600 = n7599 ^ n7536 ;
  assign n7634 = n7633 ^ n7600 ;
  assign n7635 = n7634 ^ n7632 ;
  assign n7697 = n7635 & n7694 ;
  assign n7698 = n7697 ^ n7632 ;
  assign n7699 = ~n7432 & n7698 ;
  assign n7706 = n7705 ^ n7699 ;
  assign n9169 = n7617 ^ n7599 ;
  assign n7711 = n7624 ^ n7616 ;
  assign n9170 = n9169 ^ n7711 ;
  assign n9171 = n9170 ^ n7617 ;
  assign n9172 = n7617 ^ n7432 ;
  assign n9173 = n9172 ^ n7617 ;
  assign n9174 = n9171 & ~n9173 ;
  assign n9175 = n9174 ^ n7617 ;
  assign n9176 = n7694 & ~n9175 ;
  assign n9177 = n9176 ^ n7617 ;
  assign n7714 = n7634 ^ n7602 ;
  assign n9163 = n7714 ^ n7702 ;
  assign n9164 = n7702 ^ n7694 ;
  assign n9165 = n9164 ^ n7702 ;
  assign n9166 = ~n9163 & ~n9165 ;
  assign n9167 = n9166 ^ n7702 ;
  assign n9168 = n7432 & n9167 ;
  assign n9178 = n9177 ^ n9168 ;
  assign n8682 = n7625 ^ n7618 ;
  assign n7734 = n7730 ^ n7694 ;
  assign n9155 = n8682 ^ n7734 ;
  assign n9156 = n7602 ^ n7599 ;
  assign n7735 = n7734 ^ n7432 ;
  assign n8658 = n7735 ^ n7694 ;
  assign n9157 = n9156 ^ n8658 ;
  assign n9158 = n9156 ^ n8682 ;
  assign n9159 = n9158 ^ n9156 ;
  assign n9160 = ~n9157 & ~n9159 ;
  assign n9161 = n9160 ^ n9156 ;
  assign n9162 = n9155 & ~n9161 ;
  assign n9179 = n9178 ^ n9162 ;
  assign n8659 = n7622 & n8658 ;
  assign n9180 = n9179 ^ n8659 ;
  assign n7739 = n7623 ^ n7605 ;
  assign n7740 = n7730 & n7739 ;
  assign n9181 = n9180 ^ n7740 ;
  assign n9182 = ~n7706 & n9181 ;
  assign n9184 = n9183 ^ n9182 ;
  assign n9724 = n9184 ^ x94 ;
  assign n9722 = n9149 ^ n5391 ;
  assign n9723 = n9722 ^ x76 ;
  assign n9765 = n9764 ^ x116 ;
  assign n8206 = ~n8204 & n8205 ;
  assign n8208 = n8206 ^ n8205 ;
  assign n8207 = n8206 ^ n8204 ;
  assign n8209 = n8208 ^ n8207 ;
  assign n9775 = n8311 ^ n8289 ;
  assign n9771 = n8207 & ~n8287 ;
  assign n9774 = n8314 & ~n9771 ;
  assign n9776 = n9775 ^ n9774 ;
  assign n9777 = n9776 ^ n8304 ;
  assign n9778 = n9777 ^ n8313 ;
  assign n9779 = n9778 ^ n9776 ;
  assign n8316 = n8315 ^ n8288 ;
  assign n9780 = n9779 ^ n8316 ;
  assign n9781 = n8204 & ~n9780 ;
  assign n9782 = n9781 ^ n9777 ;
  assign n9783 = n8209 & n9782 ;
  assign n9784 = n9783 ^ n9776 ;
  assign n9770 = n8302 ^ n8298 ;
  assign n9772 = n9771 ^ n9770 ;
  assign n9773 = n8208 & ~n9772 ;
  assign n9785 = n9784 ^ n9773 ;
  assign n9769 = ~n8209 & n8305 ;
  assign n9786 = n9785 ^ n9769 ;
  assign n9787 = n8318 ^ n8287 ;
  assign n9788 = ~n8205 & n9787 ;
  assign n9789 = n9788 ^ n8287 ;
  assign n9790 = n9789 ^ n8204 ;
  assign n9791 = n9790 ^ n9789 ;
  assign n9792 = ~n8205 & n8328 ;
  assign n9793 = n9792 ^ n9789 ;
  assign n9794 = n9791 & n9793 ;
  assign n9795 = n9794 ^ n9789 ;
  assign n9796 = ~n9786 & n9795 ;
  assign n9797 = n9796 ^ n9786 ;
  assign n9798 = ~n9262 & ~n9797 ;
  assign n9799 = n9798 ^ n5702 ;
  assign n9800 = n9799 ^ x101 ;
  assign n9804 = n9765 & n9800 ;
  assign n9805 = n9723 & n9804 ;
  assign n9842 = ~n9724 & n9805 ;
  assign n9207 = n8173 & n9206 ;
  assign n9195 = n8106 ^ n8101 ;
  assign n9196 = n9195 ^ n8097 ;
  assign n9203 = n9196 ^ n8693 ;
  assign n9200 = n8176 ^ n8113 ;
  assign n9201 = n9200 ^ n8159 ;
  assign n9202 = n8184 & n9201 ;
  assign n9204 = n9203 ^ n9202 ;
  assign n9197 = n9196 ^ n8109 ;
  assign n9193 = n8715 ^ n8112 ;
  assign n9194 = ~n8150 & ~n9193 ;
  assign n9198 = n9197 ^ n9194 ;
  assign n9199 = ~n8166 & ~n9198 ;
  assign n9205 = n9204 ^ n9199 ;
  assign n9208 = n9207 ^ n9205 ;
  assign n9192 = n8178 & n8188 ;
  assign n9209 = n9208 ^ n9192 ;
  assign n9190 = n8111 & n8166 ;
  assign n9189 = n7982 & n8117 ;
  assign n9191 = n9190 ^ n9189 ;
  assign n9210 = n9209 ^ n9191 ;
  assign n8179 = n8158 ^ n8116 ;
  assign n8180 = n8178 & n8179 ;
  assign n9213 = ~n8180 & ~n9212 ;
  assign n9214 = n9210 & n9213 ;
  assign n9215 = n9214 ^ n5378 ;
  assign n9819 = n9215 ^ x67 ;
  assign n9721 = n9720 ^ x125 ;
  assign n9992 = n9819 ^ n9721 ;
  assign n10017 = n9842 & ~n9992 ;
  assign n9725 = n9723 & n9724 ;
  assign n9827 = n9725 & ~n9800 ;
  assign n9809 = n9765 ^ n9723 ;
  assign n9767 = n9723 & ~n9765 ;
  assign n9810 = n9809 ^ n9767 ;
  assign n9812 = n9810 ^ n9723 ;
  assign n9814 = n9724 & ~n9812 ;
  assign n9826 = ~n9800 & n9814 ;
  assign n9828 = n9827 ^ n9826 ;
  assign n9801 = ~n9724 & ~n9800 ;
  assign n9825 = n9801 ^ n9800 ;
  assign n9829 = n9828 ^ n9825 ;
  assign n9830 = n9721 & n9819 ;
  assign n9831 = n9830 ^ n9721 ;
  assign n9832 = ~n9829 & n9831 ;
  assign n10018 = n10017 ^ n9832 ;
  assign n9802 = n9767 & n9801 ;
  assign n9766 = n9725 & ~n9765 ;
  assign n9768 = n9767 ^ n9766 ;
  assign n9803 = n9802 ^ n9768 ;
  assign n10005 = n9829 ^ n9803 ;
  assign n9815 = n9814 ^ n9812 ;
  assign n9813 = n9801 & ~n9812 ;
  assign n9816 = n9815 ^ n9813 ;
  assign n9811 = n9801 & n9810 ;
  assign n9817 = n9816 ^ n9811 ;
  assign n10006 = n10005 ^ n9817 ;
  assign n10007 = ~n9831 & ~n10006 ;
  assign n9843 = n9842 ^ n9805 ;
  assign n9841 = n9826 ^ n9814 ;
  assign n9844 = n9843 ^ n9841 ;
  assign n10000 = n9844 ^ n9827 ;
  assign n10011 = n10007 ^ n10000 ;
  assign n9835 = n9811 ^ n9802 ;
  assign n9834 = n9813 ^ n9801 ;
  assign n9836 = n9835 ^ n9834 ;
  assign n9837 = n9836 ^ n9803 ;
  assign n9848 = n9830 ^ n9819 ;
  assign n10008 = n9816 & ~n9848 ;
  assign n10009 = ~n9837 & n10008 ;
  assign n10010 = ~n10007 & n10009 ;
  assign n10012 = n10011 ^ n10010 ;
  assign n10019 = n10018 ^ n10012 ;
  assign n10001 = n10000 ^ n9725 ;
  assign n10002 = n10001 ^ n9814 ;
  assign n9806 = n9805 ^ n9804 ;
  assign n9807 = ~n9724 & n9806 ;
  assign n9839 = n9807 ^ n9806 ;
  assign n10003 = n10002 ^ n9839 ;
  assign n9993 = n9843 ^ n9725 ;
  assign n9994 = n9993 ^ n9766 ;
  assign n10004 = n10003 ^ n9994 ;
  assign n10013 = n10012 ^ n10004 ;
  assign n9998 = n9811 ^ n9768 ;
  assign n9999 = n9830 & n9998 ;
  assign n10014 = n10013 ^ n9999 ;
  assign n9995 = n9994 ^ n9807 ;
  assign n9846 = n9836 ^ n9813 ;
  assign n9996 = n9995 ^ n9846 ;
  assign n9997 = ~n9721 & n9996 ;
  assign n10015 = n10014 ^ n9997 ;
  assign n10016 = ~n9992 & ~n10015 ;
  assign n10020 = n10019 ^ n10016 ;
  assign n10021 = n10002 ^ n9802 ;
  assign n10022 = n10002 ^ n9721 ;
  assign n10023 = n10022 ^ n10002 ;
  assign n10024 = n10021 & ~n10023 ;
  assign n10025 = n10024 ^ n10002 ;
  assign n10026 = ~n9992 & n10025 ;
  assign n10027 = n10020 & ~n10026 ;
  assign n10028 = n10027 ^ n8498 ;
  assign n10029 = n10028 ^ x98 ;
  assign n8604 = n8558 ^ n8552 ;
  assign n8605 = n8604 ^ n8585 ;
  assign n8606 = ~n8466 & n8605 ;
  assign n8580 = n8467 & n8557 ;
  assign n8581 = n8580 ^ n8579 ;
  assign n8582 = n8581 ^ n8553 ;
  assign n8607 = n8606 ^ n8582 ;
  assign n8608 = n8536 & ~n8607 ;
  assign n8598 = n8468 & n8597 ;
  assign n8599 = n8598 ^ n8595 ;
  assign n8583 = n8582 ^ n8564 ;
  assign n8600 = n8599 ^ n8583 ;
  assign n8601 = n8600 ^ n8577 ;
  assign n8566 = n8565 ^ n8564 ;
  assign n8567 = n8564 ^ n8466 ;
  assign n8568 = n8567 ^ n8564 ;
  assign n8569 = ~n8566 & n8568 ;
  assign n8570 = n8569 ^ n8564 ;
  assign n8571 = n8536 & n8570 ;
  assign n8602 = n8601 ^ n8571 ;
  assign n8534 = n8533 ^ n8531 ;
  assign n8535 = ~n8469 & n8534 ;
  assign n8603 = n8602 ^ n8535 ;
  assign n8609 = n8608 ^ n8603 ;
  assign n8612 = n8611 ^ n8609 ;
  assign n8613 = n8612 ^ n5957 ;
  assign n9067 = n8613 ^ x98 ;
  assign n7738 = n7704 & ~n7734 ;
  assign n7741 = n7740 ^ n7738 ;
  assign n7716 = n7537 & n7595 ;
  assign n7715 = n7714 ^ n7598 ;
  assign n7717 = n7716 ^ n7715 ;
  assign n7713 = n7702 ^ n7537 ;
  assign n7718 = n7717 ^ n7713 ;
  assign n7719 = n7718 ^ n7609 ;
  assign n7712 = n7711 ^ n7602 ;
  assign n7720 = n7719 ^ n7712 ;
  assign n7707 = n7594 ^ n7534 ;
  assign n7708 = n7707 ^ n7613 ;
  assign n7709 = n7708 ^ n7702 ;
  assign n7710 = n7432 & ~n7709 ;
  assign n7721 = n7720 ^ n7710 ;
  assign n7742 = n7741 ^ n7721 ;
  assign n7736 = n7719 ^ n7716 ;
  assign n7737 = n7735 & n7736 ;
  assign n7743 = n7742 ^ n7737 ;
  assign n7731 = n7716 ^ n7632 ;
  assign n7732 = n7731 ^ n7608 ;
  assign n7733 = n7730 & n7732 ;
  assign n7744 = n7743 ^ n7733 ;
  assign n7722 = n7721 ^ n7626 ;
  assign n7723 = n7722 ^ n7630 ;
  assign n7724 = n7723 ^ n7722 ;
  assign n7725 = n7722 ^ n7694 ;
  assign n7726 = n7725 ^ n7722 ;
  assign n7727 = ~n7724 & n7726 ;
  assign n7728 = n7727 ^ n7722 ;
  assign n7729 = n7700 & n7728 ;
  assign n7745 = n7744 ^ n7729 ;
  assign n7746 = ~n7706 & ~n7745 ;
  assign n7747 = n7746 ^ n6549 ;
  assign n9066 = n7747 ^ x72 ;
  assign n9109 = n9067 ^ n9066 ;
  assign n8888 = n7377 ^ n7118 ;
  assign n8889 = ~n7158 & ~n8888 ;
  assign n8872 = n7356 ^ n7158 ;
  assign n8873 = n8872 ^ n7356 ;
  assign n8874 = ~n7342 & n7359 ;
  assign n8875 = n8874 ^ n7356 ;
  assign n8876 = n8873 & ~n8875 ;
  assign n8877 = n8876 ^ n7356 ;
  assign n8878 = n7118 & ~n8877 ;
  assign n8879 = n8878 ^ n7118 ;
  assign n8871 = ~n7389 & n8870 ;
  assign n8880 = n8879 ^ n8871 ;
  assign n8866 = n7391 ^ n7346 ;
  assign n8867 = n8866 ^ n7373 ;
  assign n8868 = n7159 & ~n8867 ;
  assign n8881 = n8880 ^ n8868 ;
  assign n8865 = n8864 ^ n7118 ;
  assign n8882 = n8881 ^ n8865 ;
  assign n8886 = n8885 ^ n8882 ;
  assign n8887 = n8886 ^ n6886 ;
  assign n8890 = n8889 ^ n8887 ;
  assign n8856 = n7407 ^ n7160 ;
  assign n8857 = n7362 ^ n7350 ;
  assign n8858 = n7350 ^ n7160 ;
  assign n8859 = n8858 ^ n7350 ;
  assign n8860 = n8857 & n8859 ;
  assign n8861 = n8860 ^ n7350 ;
  assign n8862 = n8856 & ~n8861 ;
  assign n8891 = n8890 ^ n8862 ;
  assign n8892 = n8891 ^ x65 ;
  assign n9003 = n9002 ^ n8895 ;
  assign n9004 = n9003 ^ n8894 ;
  assign n9005 = n9004 ^ n9003 ;
  assign n9006 = n8998 & n9005 ;
  assign n9007 = n9006 ^ n8895 ;
  assign n9012 = n9005 & ~n9009 ;
  assign n9010 = n9009 ^ n9003 ;
  assign n9013 = n9012 ^ n9010 ;
  assign n9014 = n8895 & ~n9013 ;
  assign n9015 = n9007 & n9014 ;
  assign n9016 = n9015 ^ n9012 ;
  assign n9017 = n9016 ^ n9010 ;
  assign n9018 = n9017 ^ n6900 ;
  assign n8896 = n8895 ^ n8894 ;
  assign n8984 = n8983 ^ n8967 ;
  assign n8985 = n8983 ^ n8894 ;
  assign n8986 = n8985 ^ n8983 ;
  assign n8987 = ~n8984 & n8986 ;
  assign n8988 = n8987 ^ n8983 ;
  assign n8989 = n8896 & ~n8988 ;
  assign n9019 = n9018 ^ n8989 ;
  assign n9020 = n9019 ^ x66 ;
  assign n9023 = ~n8892 & n9020 ;
  assign n6850 = n6795 ^ n6777 ;
  assign n6851 = n5787 & n6850 ;
  assign n6852 = n6851 ^ n6811 ;
  assign n6843 = n6831 ^ n6820 ;
  assign n6842 = n6833 ^ n6816 ;
  assign n6844 = n6843 ^ n6842 ;
  assign n6845 = n6842 ^ n5786 ;
  assign n6846 = n6845 ^ n6842 ;
  assign n6847 = ~n6844 & ~n6846 ;
  assign n6848 = n6847 ^ n6842 ;
  assign n6849 = ~n6841 & ~n6848 ;
  assign n6853 = n6852 ^ n6849 ;
  assign n6839 = n6838 ^ n6793 ;
  assign n6840 = n5789 & ~n6839 ;
  assign n6854 = n6853 ^ n6840 ;
  assign n6822 = n6821 ^ n6799 ;
  assign n6818 = n6817 ^ n6813 ;
  assign n6823 = n6822 ^ n6818 ;
  assign n6810 = n6809 ^ n6795 ;
  assign n6824 = n6823 ^ n6810 ;
  assign n6825 = n6823 ^ n5786 ;
  assign n6826 = n6825 ^ n6823 ;
  assign n6827 = n6824 & ~n6826 ;
  assign n6828 = n6827 ^ n6823 ;
  assign n6829 = ~n5348 & ~n6828 ;
  assign n6855 = n6854 ^ n6829 ;
  assign n6788 = n6787 ^ n6785 ;
  assign n6801 = n6800 ^ n5788 ;
  assign n6802 = n6785 ^ n5788 ;
  assign n6803 = n6802 ^ n5788 ;
  assign n6804 = ~n6801 & n6803 ;
  assign n6805 = n6804 ^ n5788 ;
  assign n6806 = n6788 & ~n6805 ;
  assign n6856 = n6855 ^ n6806 ;
  assign n6857 = ~n6784 & n6856 ;
  assign n6858 = n6857 ^ n6667 ;
  assign n8893 = n6858 ^ x104 ;
  assign n7936 = n7872 & n7877 ;
  assign n8763 = n7936 ^ n7883 ;
  assign n8800 = n8763 ^ n7941 ;
  assign n8801 = ~n7931 & n8800 ;
  assign n7930 = n7904 & n7929 ;
  assign n7934 = n7933 ^ n7930 ;
  assign n8795 = n8794 ^ n7934 ;
  assign n8796 = n8795 ^ n8763 ;
  assign n8779 = n7908 ^ n7890 ;
  assign n8780 = n8779 ^ n7936 ;
  assign n8781 = n7936 ^ n7749 ;
  assign n8782 = n8781 ^ n7936 ;
  assign n8783 = n8780 & n8782 ;
  assign n8784 = n8783 ^ n7936 ;
  assign n8785 = ~n7794 & n8784 ;
  assign n8797 = n8796 ^ n8785 ;
  assign n8798 = n8797 ^ n6017 ;
  assign n8772 = n7889 ^ n7875 ;
  assign n8773 = n8772 ^ n7889 ;
  assign n8774 = n7889 ^ n7793 ;
  assign n8775 = n8774 ^ n7889 ;
  assign n8776 = n8773 & n8775 ;
  assign n8777 = n8776 ^ n7889 ;
  assign n8778 = ~n7749 & n8777 ;
  assign n8799 = n8798 ^ n8778 ;
  assign n8802 = n8801 ^ n8799 ;
  assign n8764 = n8763 ^ n7926 ;
  assign n8765 = n8764 ^ n7927 ;
  assign n8766 = n8765 ^ n8764 ;
  assign n8767 = n8764 ^ n7749 ;
  assign n8768 = n8767 ^ n8764 ;
  assign n8769 = ~n8766 & ~n8768 ;
  assign n8770 = n8769 ^ n8764 ;
  assign n8771 = ~n7793 & ~n8770 ;
  assign n8803 = n8802 ^ n8771 ;
  assign n9025 = n8803 ^ x113 ;
  assign n9026 = n8893 & n9025 ;
  assign n9034 = n9023 & n9026 ;
  assign n9095 = n9034 ^ n9023 ;
  assign n9027 = n9026 ^ n8893 ;
  assign n9028 = n9027 ^ n9025 ;
  assign n9039 = n9023 & ~n9028 ;
  assign n9031 = n9026 ^ n9025 ;
  assign n9032 = n9023 & n9031 ;
  assign n9040 = n9039 ^ n9032 ;
  assign n9096 = n9095 ^ n9040 ;
  assign n9029 = n9023 ^ n9020 ;
  assign n9057 = n9029 ^ n8892 ;
  assign n9058 = n9026 & n9057 ;
  assign n9059 = n9058 ^ n9057 ;
  assign n9045 = n9025 ^ n9020 ;
  assign n9046 = n9045 ^ n8892 ;
  assign n9047 = n8893 & ~n9046 ;
  assign n9048 = n9047 ^ n9046 ;
  assign n9041 = n9040 ^ n9028 ;
  assign n9035 = n9025 ^ n8892 ;
  assign n9021 = n9020 ^ n8893 ;
  assign n9022 = ~n8892 & ~n9021 ;
  assign n9036 = n9022 ^ n8893 ;
  assign n9037 = n9035 & ~n9036 ;
  assign n9038 = n9037 ^ n9034 ;
  assign n9042 = n9041 ^ n9038 ;
  assign n9030 = ~n9028 & n9029 ;
  assign n9033 = n9032 ^ n9030 ;
  assign n9043 = n9042 ^ n9033 ;
  assign n9049 = n9048 ^ n9043 ;
  assign n9044 = n9043 ^ n9041 ;
  assign n9050 = n9049 ^ n9044 ;
  assign n9060 = n9059 ^ n9050 ;
  assign n9056 = n9026 & n9029 ;
  assign n9061 = n9060 ^ n9056 ;
  assign n9062 = n9061 ^ n9047 ;
  assign n9063 = n9062 ^ n8892 ;
  assign n9051 = n9050 ^ n9030 ;
  assign n9052 = n9051 ^ n8893 ;
  assign n9024 = n9023 ^ n9022 ;
  assign n9053 = n9052 ^ n9024 ;
  assign n9054 = n9053 ^ n9034 ;
  assign n9055 = n9054 ^ n9051 ;
  assign n9064 = n9063 ^ n9055 ;
  assign n9097 = n9096 ^ n9064 ;
  assign n9112 = n9096 ^ n9066 ;
  assign n9113 = n9112 ^ n9096 ;
  assign n9114 = ~n9097 & ~n9113 ;
  assign n9115 = n9114 ^ n9096 ;
  assign n9116 = n9109 & n9115 ;
  assign n9068 = n9066 & n9067 ;
  assign n9069 = n9068 ^ n9067 ;
  assign n9070 = n9069 ^ n9066 ;
  assign n9085 = n9047 ^ n8893 ;
  assign n9118 = n9085 ^ n9061 ;
  assign n9119 = ~n9070 & n9118 ;
  assign n9117 = n9033 & n9068 ;
  assign n9120 = n9119 ^ n9117 ;
  assign n10045 = n9060 & ~n9070 ;
  assign n9072 = n9053 ^ n9042 ;
  assign n10038 = n9072 ^ n9041 ;
  assign n10039 = n9066 & ~n10038 ;
  assign n10040 = n10039 ^ n9048 ;
  assign n10041 = n10040 ^ n9034 ;
  assign n10046 = n10045 ^ n10041 ;
  assign n9073 = n9072 ^ n9032 ;
  assign n10034 = n9073 ^ n9044 ;
  assign n10035 = n10034 ^ n9096 ;
  assign n10042 = n10041 ^ n10035 ;
  assign n9126 = n9049 ^ n9034 ;
  assign n10031 = n9126 ^ n9063 ;
  assign n9098 = n9060 ^ n9027 ;
  assign n9099 = n9098 ^ n9097 ;
  assign n9100 = n9099 ^ n9044 ;
  assign n9094 = n9072 ^ n9033 ;
  assign n9101 = n9100 ^ n9094 ;
  assign n10032 = n10031 ^ n9101 ;
  assign n10030 = n8893 ^ n8892 ;
  assign n10033 = n10032 ^ n10030 ;
  assign n10036 = n10035 ^ n10033 ;
  assign n10037 = n9066 & n10036 ;
  assign n10043 = n10042 ^ n10037 ;
  assign n10044 = n9067 & ~n10043 ;
  assign n10047 = n10046 ^ n10044 ;
  assign n10048 = ~n9120 & n10047 ;
  assign n10049 = ~n9116 & n10048 ;
  assign n10055 = n10049 ^ n8526 ;
  assign n10050 = n9096 ^ n9061 ;
  assign n10051 = n10050 ^ n9085 ;
  assign n10052 = n10051 ^ n9099 ;
  assign n10053 = n9109 & ~n10052 ;
  assign n10054 = n10049 & n10053 ;
  assign n10056 = n10055 ^ n10054 ;
  assign n10057 = n10056 ^ x120 ;
  assign n10058 = n10029 & n10057 ;
  assign n10397 = n10058 ^ n10057 ;
  assign n10402 = ~n10395 & n10397 ;
  assign n9485 = n8587 ^ n8543 ;
  assign n9486 = n9485 ^ n8531 ;
  assign n9487 = n9486 ^ n9483 ;
  assign n9482 = n9481 ^ n8597 ;
  assign n9484 = n9483 ^ n9482 ;
  assign n9488 = n9487 ^ n9484 ;
  assign n9489 = n9484 ^ n9483 ;
  assign n9490 = n9489 ^ n8466 ;
  assign n9491 = n8536 & ~n9490 ;
  assign n9492 = n9491 ^ n8466 ;
  assign n9493 = ~n9488 & n9492 ;
  assign n9494 = n9493 ^ n9487 ;
  assign n9495 = ~n8552 & n9494 ;
  assign n9496 = n8546 & n9495 ;
  assign n9478 = n8563 ^ n8533 ;
  assign n9479 = n9478 ^ n8550 ;
  assign n9480 = ~n8466 & n9479 ;
  assign n9497 = n9496 ^ n9480 ;
  assign n9498 = n8536 & ~n9497 ;
  assign n9499 = n9498 ^ n9496 ;
  assign n9471 = n8586 ^ n8542 ;
  assign n9472 = n9471 ^ n8555 ;
  assign n9473 = n8555 ^ n8466 ;
  assign n9474 = n9473 ^ n8555 ;
  assign n9475 = ~n9472 & n9474 ;
  assign n9476 = n9475 ^ n8555 ;
  assign n9477 = ~n8465 & n9476 ;
  assign n9500 = n9499 ^ n9477 ;
  assign n9501 = n9500 ^ n8580 ;
  assign n9502 = n9501 ^ n8599 ;
  assign n9503 = n9502 ^ n9470 ;
  assign n9504 = n9503 ^ n7194 ;
  assign n9505 = n9504 ^ x74 ;
  assign n7419 = ~n7394 & ~n7403 ;
  assign n7411 = n7346 ^ n7341 ;
  assign n7408 = n7407 ^ n7338 ;
  assign n7056 = ~n7004 & ~n7055 ;
  assign n7409 = n7408 ^ n7056 ;
  assign n7412 = n7411 ^ n7409 ;
  assign n7413 = n7118 & ~n7412 ;
  assign n7410 = n7409 ^ n7342 ;
  assign n7414 = n7413 ^ n7410 ;
  assign n7415 = ~n7158 & n7414 ;
  assign n7406 = n7405 ^ n7402 ;
  assign n7416 = n7415 ^ n7406 ;
  assign n7386 = n7357 ^ n7342 ;
  assign n7387 = n7386 ^ n7158 ;
  assign n7388 = n7118 & ~n7387 ;
  assign n7417 = n7416 ^ n7388 ;
  assign n7104 = n7103 ^ n7056 ;
  assign n7331 = n7330 ^ n7004 ;
  assign n7332 = n7160 & ~n7331 ;
  assign n7333 = n7104 & n7332 ;
  assign n7334 = n7333 ^ n7160 ;
  assign n7363 = n7362 ^ n7354 ;
  assign n7364 = n7363 ^ n7354 ;
  assign n7365 = n7359 & n7364 ;
  assign n7366 = n7365 ^ n7354 ;
  assign n7367 = ~n7334 & ~n7366 ;
  assign n7368 = n7367 ^ n7160 ;
  assign n7380 = n7379 ^ n7362 ;
  assign n7383 = ~n7367 & n7380 ;
  assign n7384 = n7383 ^ n7362 ;
  assign n7385 = ~n7368 & ~n7384 ;
  assign n7418 = n7417 ^ n7385 ;
  assign n7420 = n7419 ^ n7418 ;
  assign n7428 = n7420 & ~n7427 ;
  assign n7429 = n7428 ^ n6646 ;
  assign n9507 = n7429 ^ x89 ;
  assign n9510 = n9505 & ~n9507 ;
  assign n9511 = n9510 ^ n9505 ;
  assign n9513 = n9511 ^ n9507 ;
  assign n9429 = n7700 ^ n7621 ;
  assign n9430 = n7621 ^ n7535 ;
  assign n9431 = n9430 ^ n7618 ;
  assign n9432 = ~n7432 & ~n9431 ;
  assign n9433 = n9432 ^ n7622 ;
  assign n9434 = n9429 & n9433 ;
  assign n9435 = n9434 ^ n7621 ;
  assign n9448 = n7714 ^ n7627 ;
  assign n9449 = n9448 ^ n7734 ;
  assign n9450 = n9449 ^ n7731 ;
  assign n9451 = ~n7617 & ~n9450 ;
  assign n9452 = n9451 ^ n7734 ;
  assign n9453 = n8658 ^ n7617 ;
  assign n9454 = ~n9452 & n9453 ;
  assign n9436 = n7719 ^ n7633 ;
  assign n9437 = n9436 ^ n9156 ;
  assign n9438 = ~n7432 & n9437 ;
  assign n9439 = n9438 ^ n7633 ;
  assign n9455 = n9454 ^ n9439 ;
  assign n9440 = n9439 ^ n7605 ;
  assign n9441 = n9440 ^ n7620 ;
  assign n9442 = n9441 ^ n9439 ;
  assign n9443 = n9439 ^ n7694 ;
  assign n9444 = n9443 ^ n9439 ;
  assign n9445 = ~n9442 & ~n9444 ;
  assign n9446 = n9445 ^ n9439 ;
  assign n9447 = ~n7700 & ~n9446 ;
  assign n9456 = n9455 ^ n9447 ;
  assign n9457 = ~n8689 & ~n9456 ;
  assign n9458 = ~n7741 & n9457 ;
  assign n9459 = ~n9435 & n9458 ;
  assign n9462 = n9459 ^ n7233 ;
  assign n9428 = n7731 ^ n7598 ;
  assign n9460 = ~n7734 & n9459 ;
  assign n9461 = n9428 & n9460 ;
  assign n9463 = n9462 ^ n9461 ;
  assign n9464 = n9463 ^ x64 ;
  assign n9528 = n9527 ^ x120 ;
  assign n9529 = ~n9464 & ~n9528 ;
  assign n9530 = n9529 ^ n9528 ;
  assign n9531 = n9530 ^ n9464 ;
  assign n9597 = n9513 & ~n9531 ;
  assign n9535 = n9511 & ~n9531 ;
  assign n8331 = n8327 ^ n8204 ;
  assign n8332 = n8327 ^ n8324 ;
  assign n8335 = n8332 ^ n8205 ;
  assign n8336 = n8335 ^ n8332 ;
  assign n8337 = n8325 & n8336 ;
  assign n8338 = n8337 ^ n8332 ;
  assign n8339 = n8331 & ~n8338 ;
  assign n8340 = n8339 ^ n8204 ;
  assign n8329 = n8328 ^ n8296 ;
  assign n8330 = ~n8207 & n8329 ;
  assign n8341 = n8340 ^ n8330 ;
  assign n8320 = n8313 ^ n8283 ;
  assign n8319 = n8318 ^ n8308 ;
  assign n8321 = n8320 ^ n8319 ;
  assign n8322 = n8206 & n8321 ;
  assign n8342 = n8341 ^ n8322 ;
  assign n8317 = ~n8209 & ~n8316 ;
  assign n8343 = n8342 ^ n8317 ;
  assign n8345 = n8205 & n8344 ;
  assign n8346 = n8345 ^ n8313 ;
  assign n8347 = n8346 ^ n8204 ;
  assign n8348 = n8347 ^ n8346 ;
  assign n8350 = ~n8205 & n8349 ;
  assign n8351 = n8350 ^ n8346 ;
  assign n8352 = n8348 & n8351 ;
  assign n8353 = n8352 ^ n8346 ;
  assign n8354 = ~n8343 & n8353 ;
  assign n8355 = n8354 ^ n8343 ;
  assign n8356 = n8283 ^ n8205 ;
  assign n8357 = n8356 ^ n8283 ;
  assign n8359 = n8313 & ~n8357 ;
  assign n8360 = n8359 ^ n8283 ;
  assign n8361 = n8204 & n8360 ;
  assign n8362 = ~n8355 & ~n8361 ;
  assign n8363 = n8362 ^ n6582 ;
  assign n9581 = n8363 ^ x122 ;
  assign n9580 = n9579 ^ x115 ;
  assign n9618 = n9581 ^ n9580 ;
  assign n9987 = n9535 & ~n9618 ;
  assign n9582 = ~n9580 & n9581 ;
  assign n9608 = n9582 ^ n9581 ;
  assign n9506 = n9505 ^ n9464 ;
  assign n9590 = n9506 & ~n9507 ;
  assign n9552 = n9513 & n9529 ;
  assign n9542 = n9528 ^ n9464 ;
  assign n9543 = n9542 ^ n9507 ;
  assign n9544 = n9505 & n9543 ;
  assign n9545 = n9544 ^ n9535 ;
  assign n9540 = n9510 & ~n9530 ;
  assign n9539 = n9511 & n9529 ;
  assign n9541 = n9540 ^ n9539 ;
  assign n9546 = n9545 ^ n9541 ;
  assign n9532 = n9531 ^ n9528 ;
  assign n9547 = n9546 ^ n9532 ;
  assign n9508 = n9507 ^ n9505 ;
  assign n9509 = ~n9506 & ~n9508 ;
  assign n9536 = n9535 ^ n9509 ;
  assign n9534 = n9509 & ~n9528 ;
  assign n9537 = n9536 ^ n9534 ;
  assign n9533 = n9513 & ~n9532 ;
  assign n9538 = n9537 ^ n9533 ;
  assign n9548 = n9547 ^ n9538 ;
  assign n9549 = n9548 ^ n9537 ;
  assign n9512 = n9511 ^ n9509 ;
  assign n9550 = n9549 ^ n9512 ;
  assign n9551 = n9550 ^ n9529 ;
  assign n9553 = n9552 ^ n9551 ;
  assign n9591 = n9590 ^ n9553 ;
  assign n9587 = n9513 ^ n9505 ;
  assign n9588 = ~n9530 & ~n9587 ;
  assign n9589 = n9588 ^ n9546 ;
  assign n9592 = n9591 ^ n9589 ;
  assign n9593 = n9592 ^ n9533 ;
  assign n9983 = n9593 ^ n9553 ;
  assign n9984 = n9983 ^ n9548 ;
  assign n9985 = n9608 & ~n9984 ;
  assign n9610 = n9553 ^ n9534 ;
  assign n9611 = n9610 ^ n9552 ;
  assign n9594 = n9593 ^ n9537 ;
  assign n9595 = n9594 ^ n9535 ;
  assign n9612 = n9611 ^ n9595 ;
  assign n9613 = n9612 ^ n9545 ;
  assign n9598 = n9597 ^ n9538 ;
  assign n9596 = n9595 ^ n9531 ;
  assign n9599 = n9598 ^ n9596 ;
  assign n9600 = n9599 ^ n9588 ;
  assign n9601 = n9600 ^ n9548 ;
  assign n9609 = n9601 ^ n9597 ;
  assign n9614 = n9613 ^ n9609 ;
  assign n9981 = ~n9580 & n9614 ;
  assign n9977 = n9593 ^ n9550 ;
  assign n9978 = n9977 ^ n9599 ;
  assign n9979 = n9582 & n9978 ;
  assign n9639 = n9552 ^ n9540 ;
  assign n9640 = n9639 ^ n9534 ;
  assign n9641 = n9640 ^ n9589 ;
  assign n9642 = n9641 ^ n9639 ;
  assign n9643 = n9639 ^ n9581 ;
  assign n9644 = n9643 ^ n9639 ;
  assign n9645 = n9642 & ~n9644 ;
  assign n9646 = n9645 ^ n9639 ;
  assign n9647 = n9618 & n9646 ;
  assign n9973 = n9647 ^ n9639 ;
  assign n9670 = n9588 ^ n9537 ;
  assign n9673 = ~n9580 & n9670 ;
  assign n9674 = n9673 ^ n9537 ;
  assign n9675 = ~n9581 & n9674 ;
  assign n9974 = n9973 ^ n9675 ;
  assign n9967 = n9549 ^ n9541 ;
  assign n9970 = ~n9580 & ~n9967 ;
  assign n9971 = n9970 ^ n9541 ;
  assign n9972 = ~n9581 & n9971 ;
  assign n9975 = n9974 ^ n9972 ;
  assign n9583 = ~n9553 & n9582 ;
  assign n9976 = n9975 ^ n9583 ;
  assign n9980 = n9979 ^ n9976 ;
  assign n9982 = n9981 ^ n9980 ;
  assign n9986 = n9985 ^ n9982 ;
  assign n9988 = n9987 ^ n9986 ;
  assign n9989 = ~n9597 & ~n9988 ;
  assign n9990 = n9989 ^ n8069 ;
  assign n9991 = n9990 ^ x66 ;
  assign n9154 = n9153 ^ x85 ;
  assign n9185 = n9184 ^ x102 ;
  assign n9186 = ~n9154 & n9185 ;
  assign n9187 = n9186 ^ n9185 ;
  assign n9289 = n9288 ^ x68 ;
  assign n9319 = n6784 ^ n6114 ;
  assign n9320 = n9319 ^ n8759 ;
  assign n9302 = n6793 ^ n6786 ;
  assign n9303 = ~n9301 & n9302 ;
  assign n9304 = n9303 ^ n6796 ;
  assign n9300 = n5788 & n6781 ;
  assign n9305 = n9304 ^ n9300 ;
  assign n9306 = n9305 ^ n8741 ;
  assign n9308 = n9307 ^ n9306 ;
  assign n9309 = n9308 ^ n9305 ;
  assign n9310 = n9305 ^ n5786 ;
  assign n9311 = n9310 ^ n9305 ;
  assign n9312 = n9309 & n9311 ;
  assign n9313 = n9312 ^ n9305 ;
  assign n9314 = n6841 & n9313 ;
  assign n9315 = n9314 ^ n9305 ;
  assign n9298 = n9297 ^ n6817 ;
  assign n9299 = ~n5788 & n9298 ;
  assign n9316 = n9315 ^ n9299 ;
  assign n9290 = n8736 ^ n6815 ;
  assign n9291 = n9290 ^ n6835 ;
  assign n9292 = n6835 ^ n5786 ;
  assign n9293 = n9292 ^ n6835 ;
  assign n9294 = n9291 & ~n9293 ;
  assign n9295 = n9294 ^ n6835 ;
  assign n9296 = n5348 & ~n9295 ;
  assign n9317 = n9316 ^ n9296 ;
  assign n9318 = ~n6851 & ~n9317 ;
  assign n9321 = n9320 ^ n9318 ;
  assign n9322 = n9321 ^ x126 ;
  assign n9323 = n9289 & n9322 ;
  assign n9325 = n9323 ^ n9289 ;
  assign n9333 = n9325 ^ n9322 ;
  assign n9334 = n9333 ^ n9289 ;
  assign n9216 = n9215 ^ x124 ;
  assign n7910 = n7908 ^ n7875 ;
  assign n7907 = n7876 & n7882 ;
  assign n7909 = n7908 ^ n7907 ;
  assign n7911 = n7910 ^ n7909 ;
  assign n7912 = n7910 ^ n7749 ;
  assign n7913 = n7912 ^ n7910 ;
  assign n7914 = n7911 & ~n7913 ;
  assign n7915 = n7914 ^ n7910 ;
  assign n7916 = ~n7794 & n7915 ;
  assign n7917 = n7916 ^ n7908 ;
  assign n9242 = n7794 & n7875 ;
  assign n9237 = n7925 ^ n7887 ;
  assign n9234 = n7905 ^ n7893 ;
  assign n9235 = n9234 ^ n7907 ;
  assign n9236 = n7793 & ~n9235 ;
  assign n9238 = n9237 ^ n9236 ;
  assign n9239 = n7749 & n9238 ;
  assign n9219 = n7929 ^ n7919 ;
  assign n9220 = n9219 ^ n7936 ;
  assign n9218 = n7908 ^ n7884 ;
  assign n9221 = n9220 ^ n9218 ;
  assign n9222 = ~n7749 & n9221 ;
  assign n9223 = n9222 ^ n9220 ;
  assign n9232 = n9223 ^ n7925 ;
  assign n9224 = n9223 ^ n7918 ;
  assign n9225 = n9224 ^ n8763 ;
  assign n9226 = n9225 ^ n9223 ;
  assign n9229 = ~n7749 & n9226 ;
  assign n9230 = n9229 ^ n9223 ;
  assign n9231 = n7793 & n9230 ;
  assign n9233 = n9232 ^ n9231 ;
  assign n9240 = n9239 ^ n9233 ;
  assign n9217 = n7904 & n7941 ;
  assign n9241 = n9240 ^ n9217 ;
  assign n9243 = n9242 ^ n9241 ;
  assign n9244 = ~n8792 & ~n9243 ;
  assign n9245 = ~n7917 & n9244 ;
  assign n9246 = ~n7956 & n9245 ;
  assign n9247 = ~n8785 & n9246 ;
  assign n9248 = n9247 ^ n6167 ;
  assign n9249 = n9248 ^ x78 ;
  assign n9250 = n9216 & n9249 ;
  assign n9326 = n9250 ^ n9249 ;
  assign n9338 = n9326 ^ n9216 ;
  assign n9349 = n9334 & ~n9338 ;
  assign n9339 = n9338 ^ n9249 ;
  assign n9340 = n9325 & n9339 ;
  assign n9327 = n9325 & n9326 ;
  assign n9324 = n9250 & n9323 ;
  assign n9328 = n9327 ^ n9324 ;
  assign n9341 = n9340 ^ n9328 ;
  assign n9342 = n9341 ^ n9289 ;
  assign n9343 = n9250 & n9342 ;
  assign n9337 = n9250 & n9334 ;
  assign n9344 = n9343 ^ n9337 ;
  assign n9330 = n9322 ^ n9289 ;
  assign n9331 = n9289 ^ n9249 ;
  assign n9332 = n9330 & ~n9331 ;
  assign n9335 = n9334 ^ n9332 ;
  assign n9336 = n9335 ^ n9327 ;
  assign n9345 = n9344 ^ n9336 ;
  assign n9362 = n9349 ^ n9345 ;
  assign n9363 = n9362 ^ n9337 ;
  assign n10436 = ~n9187 & ~n9363 ;
  assign n9359 = n9344 ^ n9324 ;
  assign n9360 = n9359 ^ n9250 ;
  assign n9369 = n9360 ^ n9333 ;
  assign n9367 = n9326 & ~n9333 ;
  assign n9351 = ~n9333 & n9339 ;
  assign n9368 = n9367 ^ n9351 ;
  assign n9370 = n9369 ^ n9368 ;
  assign n10437 = n10436 ^ n9370 ;
  assign n9374 = n9323 & n9326 ;
  assign n9371 = n9363 ^ n9334 ;
  assign n9372 = n9371 ^ n9370 ;
  assign n9373 = n9372 ^ n9345 ;
  assign n9375 = n9374 ^ n9373 ;
  assign n9365 = n9343 ^ n9327 ;
  assign n9366 = n9365 ^ n9340 ;
  assign n9376 = n9375 ^ n9366 ;
  assign n9377 = n9376 ^ n9368 ;
  assign n9355 = n9289 ^ n9216 ;
  assign n9356 = n9355 ^ n9322 ;
  assign n9357 = n9333 ^ n9332 ;
  assign n9358 = n9356 & n9357 ;
  assign n9361 = n9360 ^ n9358 ;
  assign n9364 = n9363 ^ n9361 ;
  assign n9378 = n9377 ^ n9364 ;
  assign n10439 = n9378 ^ n9340 ;
  assign n10438 = n9345 ^ n9343 ;
  assign n10440 = n10439 ^ n10438 ;
  assign n10441 = n9187 & n10440 ;
  assign n9348 = n9186 ^ n9154 ;
  assign n10442 = n10441 ^ n9348 ;
  assign n10443 = n10437 & ~n10442 ;
  assign n10446 = n9368 ^ n9337 ;
  assign n10447 = n9187 & n10446 ;
  assign n10448 = ~n10443 & n10447 ;
  assign n9354 = n9185 ^ n9154 ;
  assign n9400 = n9374 ^ n9349 ;
  assign n9399 = n9323 & n9339 ;
  assign n9401 = n9400 ^ n9399 ;
  assign n10429 = n9401 ^ n9371 ;
  assign n10430 = n10429 ^ n9361 ;
  assign n10431 = n9361 ^ n9185 ;
  assign n10432 = n10431 ^ n9361 ;
  assign n10433 = n10430 & ~n10432 ;
  assign n10434 = n10433 ^ n9361 ;
  assign n10435 = n9354 & n10434 ;
  assign n10444 = n10443 ^ n10435 ;
  assign n10449 = n10448 ^ n10444 ;
  assign n10450 = n9367 ^ n9354 ;
  assign n10451 = n10450 ^ n9367 ;
  assign n10452 = ~n9185 & n9365 ;
  assign n10453 = n10452 ^ n9367 ;
  assign n10454 = ~n10451 & n10453 ;
  assign n10455 = n10454 ^ n9367 ;
  assign n10456 = ~n10449 & n10455 ;
  assign n10457 = n10456 ^ n10449 ;
  assign n10458 = n9372 ^ n9349 ;
  assign n10459 = n9349 ^ n9154 ;
  assign n10460 = n10459 ^ n9349 ;
  assign n10461 = ~n10458 & ~n10460 ;
  assign n10462 = n10461 ^ n9349 ;
  assign n10463 = n9185 & n10462 ;
  assign n10464 = ~n10457 & ~n10463 ;
  assign n9188 = n9187 ^ n9154 ;
  assign n9329 = n9188 & n9328 ;
  assign n10466 = n9188 & n9360 ;
  assign n10465 = ~n9348 & n10439 ;
  assign n10467 = n10466 ^ n10465 ;
  assign n10468 = ~n9329 & ~n10467 ;
  assign n10469 = n10464 & n10468 ;
  assign n10470 = n10469 ^ n6277 ;
  assign n10471 = n10470 ^ x122 ;
  assign n10508 = ~n9991 & ~n10471 ;
  assign n10509 = n10508 ^ n10471 ;
  assign n10510 = n10402 & ~n10509 ;
  assign n10059 = n10058 ^ n10029 ;
  assign n10407 = n10059 ^ n10057 ;
  assign n10421 = ~n10395 & ~n10407 ;
  assign n10501 = n10471 ^ n10421 ;
  assign n10502 = n10501 ^ n10421 ;
  assign n10417 = n10058 & n10386 ;
  assign n10412 = n10058 & n10392 ;
  assign n10396 = n10395 ^ n10205 ;
  assign n10399 = n10059 & n10396 ;
  assign n10389 = n10385 ^ n10205 ;
  assign n10390 = n10385 ^ n10059 ;
  assign n10391 = n10389 & ~n10390 ;
  assign n10393 = n10392 ^ n10391 ;
  assign n10400 = n10399 ^ n10393 ;
  assign n10413 = n10412 ^ n10400 ;
  assign n10405 = n10386 & n10397 ;
  assign n10416 = n10413 ^ n10405 ;
  assign n10418 = n10417 ^ n10416 ;
  assign n10408 = n10392 & ~n10407 ;
  assign n10411 = n10408 ^ n10392 ;
  assign n10414 = n10413 ^ n10411 ;
  assign n10387 = n10059 & n10386 ;
  assign n10415 = n10414 ^ n10387 ;
  assign n10419 = n10418 ^ n10415 ;
  assign n10410 = n10408 ^ n10205 ;
  assign n10420 = n10419 ^ n10410 ;
  assign n10422 = n10421 ^ n10420 ;
  assign n10503 = n10422 ^ n10421 ;
  assign n10504 = n10503 ^ n10421 ;
  assign n10505 = n10502 & n10504 ;
  assign n10506 = n10505 ^ n10421 ;
  assign n10507 = ~n9991 & n10506 ;
  assign n10511 = n10510 ^ n10507 ;
  assign n10495 = n10412 ^ n10399 ;
  assign n10496 = n10399 ^ n9991 ;
  assign n10497 = n10496 ^ n10399 ;
  assign n10498 = n10495 & n10497 ;
  assign n10499 = n10498 ^ n10399 ;
  assign n10500 = n10471 & n10499 ;
  assign n12517 = n10500 ^ n10415 ;
  assign n10529 = n10471 ^ n9991 ;
  assign n10426 = n10417 ^ n10402 ;
  assign n10427 = n10426 ^ n10420 ;
  assign n10530 = ~n9991 & n10427 ;
  assign n10531 = n10530 ^ n10420 ;
  assign n10485 = n10417 ^ n10400 ;
  assign n10409 = n10408 ^ n10407 ;
  assign n10423 = n10422 ^ n10409 ;
  assign n10398 = n10396 & n10397 ;
  assign n10401 = n10400 ^ n10398 ;
  assign n10403 = n10402 ^ n10401 ;
  assign n10388 = n10387 ^ n10059 ;
  assign n10394 = n10393 ^ n10388 ;
  assign n10404 = n10403 ^ n10394 ;
  assign n10406 = n10405 ^ n10404 ;
  assign n10424 = n10423 ^ n10406 ;
  assign n10425 = n10424 ^ n10390 ;
  assign n10428 = n10427 ^ n10425 ;
  assign n10486 = n10485 ^ n10428 ;
  assign n10484 = n10413 ^ n10058 ;
  assign n10487 = n10486 ^ n10484 ;
  assign n10532 = n10531 ^ n10487 ;
  assign n10533 = n10532 ^ n10531 ;
  assign n10534 = n10531 ^ n10471 ;
  assign n10535 = n10534 ^ n10531 ;
  assign n10536 = ~n10533 & n10535 ;
  assign n10537 = n10536 ^ n10531 ;
  assign n10538 = n10529 & n10537 ;
  assign n10539 = n10538 ^ n10531 ;
  assign n12518 = n12517 ^ n10539 ;
  assign n12519 = n12518 ^ n10428 ;
  assign n12252 = n10423 ^ n10394 ;
  assign n12520 = n12519 ^ n12252 ;
  assign n12510 = n10415 ^ n10401 ;
  assign n12511 = n12510 ^ n10419 ;
  assign n12514 = n10471 & n12511 ;
  assign n12515 = n12514 ^ n10419 ;
  assign n12516 = n10529 & n12515 ;
  assign n12521 = n12520 ^ n12516 ;
  assign n12508 = n10421 ^ n10399 ;
  assign n12509 = ~n10509 & n12508 ;
  assign n12522 = n12521 ^ n12509 ;
  assign n12500 = n10428 ^ n10398 ;
  assign n12501 = n12500 ^ n10487 ;
  assign n12502 = n12501 ^ n10428 ;
  assign n12503 = n10428 ^ n9991 ;
  assign n12504 = n12503 ^ n10428 ;
  assign n12505 = ~n12502 & n12504 ;
  assign n12506 = n12505 ^ n10428 ;
  assign n12507 = n10471 & ~n12506 ;
  assign n12523 = n12522 ^ n12507 ;
  assign n12492 = n12252 ^ n10412 ;
  assign n10520 = n10408 ^ n10405 ;
  assign n12493 = n12492 ^ n10520 ;
  assign n12494 = n12493 ^ n12252 ;
  assign n12495 = n12252 ^ n10471 ;
  assign n12496 = n12495 ^ n12252 ;
  assign n12497 = n12494 & n12496 ;
  assign n12498 = n12497 ^ n12252 ;
  assign n12499 = n10529 & ~n12498 ;
  assign n12524 = n12523 ^ n12499 ;
  assign n12525 = ~n10511 & ~n12524 ;
  assign n12526 = n12525 ^ n9764 ;
  assign n13145 = n12526 ^ x94 ;
  assign n10815 = n10052 ^ n9058 ;
  assign n10816 = ~n9109 & ~n10815 ;
  assign n10803 = n10050 ^ n9027 ;
  assign n10804 = n10803 ^ n10050 ;
  assign n10805 = n10050 ^ n9067 ;
  assign n10806 = n10805 ^ n10050 ;
  assign n10807 = n10804 & ~n10806 ;
  assign n10808 = n10807 ^ n10050 ;
  assign n10809 = n9109 & n10808 ;
  assign n10810 = n10809 ^ n10045 ;
  assign n10811 = n10810 ^ n9116 ;
  assign n9078 = n9073 ^ n9039 ;
  assign n9079 = n9078 ^ n9052 ;
  assign n10795 = n9079 ^ n9069 ;
  assign n9071 = n9070 ^ n9067 ;
  assign n10796 = n9071 ^ n9044 ;
  assign n10799 = ~n9069 & ~n10796 ;
  assign n10800 = n10799 ^ n9044 ;
  assign n10801 = ~n10795 & n10800 ;
  assign n10802 = n10801 ^ n9079 ;
  assign n10812 = n10811 ^ n10802 ;
  assign n10813 = n10812 ^ n7693 ;
  assign n10791 = n9048 ^ n9030 ;
  assign n10792 = n10791 ^ n9039 ;
  assign n10793 = n10792 ^ n9056 ;
  assign n10794 = n9068 & ~n10793 ;
  assign n10814 = n10813 ^ n10794 ;
  assign n10817 = n10816 ^ n10814 ;
  assign n10790 = ~n9070 & n9078 ;
  assign n10818 = n10817 ^ n10790 ;
  assign n10787 = ~n9055 & n9067 ;
  assign n10788 = n10787 ^ n9051 ;
  assign n10789 = n9109 & n10788 ;
  assign n10819 = n10818 ^ n10789 ;
  assign n11565 = n10819 ^ x107 ;
  assign n10856 = n10186 ^ n10131 ;
  assign n11596 = n10150 & n10856 ;
  assign n11579 = n10167 ^ n10162 ;
  assign n11111 = n10175 ^ n10159 ;
  assign n11580 = n11579 ^ n11111 ;
  assign n11581 = ~n10126 & n11580 ;
  assign n11592 = n11581 ^ n8959 ;
  assign n10857 = n10143 ^ n10130 ;
  assign n11124 = n10857 ^ n10145 ;
  assign n11125 = n10857 ^ n10131 ;
  assign n11126 = n11125 ^ n10857 ;
  assign n11127 = n11124 & ~n11126 ;
  assign n11128 = n11127 ^ n10857 ;
  assign n11129 = ~n10126 & n11128 ;
  assign n11593 = n11592 ^ n11129 ;
  assign n11582 = n10177 ^ n10166 ;
  assign n11583 = n11582 ^ n11581 ;
  assign n11566 = n10171 ^ n10161 ;
  assign n11584 = n11583 ^ n11566 ;
  assign n11585 = n11584 ^ n10166 ;
  assign n11586 = n11585 ^ n11583 ;
  assign n11587 = n11583 ^ n10126 ;
  assign n11588 = n11587 ^ n11583 ;
  assign n11589 = n11586 & n11588 ;
  assign n11590 = n11589 ^ n11583 ;
  assign n11591 = n10138 & n11590 ;
  assign n11594 = n11593 ^ n11591 ;
  assign n11575 = n10152 ^ n10144 ;
  assign n11578 = n10186 & ~n11575 ;
  assign n11595 = n11594 ^ n11578 ;
  assign n11597 = n11596 ^ n11595 ;
  assign n11576 = n10186 ^ n10126 ;
  assign n11577 = ~n11575 & n11576 ;
  assign n11598 = n11597 ^ n11577 ;
  assign n11107 = n10151 ^ n10141 ;
  assign n11568 = n11107 ^ n10130 ;
  assign n11567 = n11566 ^ n10167 ;
  assign n11569 = n11568 ^ n11567 ;
  assign n11570 = n11567 ^ n10126 ;
  assign n11571 = n11570 ^ n11567 ;
  assign n11572 = ~n11569 & ~n11571 ;
  assign n11573 = n11572 ^ n11567 ;
  assign n11574 = ~n10138 & n11573 ;
  assign n11599 = n11598 ^ n11574 ;
  assign n11600 = n11599 ^ x80 ;
  assign n11602 = n11565 & ~n11600 ;
  assign n11601 = n11600 ^ n11565 ;
  assign n11603 = n11602 ^ n11601 ;
  assign n7430 = n7429 ^ x73 ;
  assign n6859 = n6858 ^ x82 ;
  assign n7748 = n7747 ^ x88 ;
  assign n7951 = n7921 & ~n7932 ;
  assign n7945 = n7936 ^ n7925 ;
  assign n7946 = n7945 ^ n7907 ;
  assign n7947 = n7793 & n7946 ;
  assign n7943 = n7942 ^ n7919 ;
  assign n7937 = n7936 ^ n7881 ;
  assign n7938 = n7937 ^ n7875 ;
  assign n7939 = ~n7793 & n7938 ;
  assign n7944 = n7943 ^ n7939 ;
  assign n7948 = n7947 ^ n7944 ;
  assign n7949 = n7749 & n7948 ;
  assign n7935 = n7934 ^ n7917 ;
  assign n7940 = n7939 ^ n7935 ;
  assign n7950 = n7949 ^ n7940 ;
  assign n7952 = n7951 ^ n7950 ;
  assign n7906 = n7904 & n7905 ;
  assign n7953 = n7952 ^ n7906 ;
  assign n7894 = n7893 ^ n7883 ;
  assign n7899 = n7894 ^ n7749 ;
  assign n7900 = n7899 ^ n7894 ;
  assign n7901 = n7896 & ~n7900 ;
  assign n7902 = n7901 ^ n7894 ;
  assign n7903 = n7794 & ~n7902 ;
  assign n7954 = n7953 ^ n7903 ;
  assign n7957 = n7956 ^ n7954 ;
  assign n7958 = n7957 ^ n6507 ;
  assign n7959 = n7958 ^ x114 ;
  assign n8192 = n8118 ^ n8101 ;
  assign n8193 = n8192 ^ n8030 ;
  assign n8194 = n8193 ^ n8121 ;
  assign n8195 = n8150 & ~n8194 ;
  assign n8190 = n8189 ^ n8101 ;
  assign n8175 = n8174 ^ n8097 ;
  assign n8177 = n8176 ^ n8175 ;
  assign n8191 = n8190 ^ n8177 ;
  assign n8196 = n8195 ^ n8191 ;
  assign n8197 = ~n8166 & n8196 ;
  assign n8181 = n8180 ^ n8177 ;
  assign n8182 = n8181 ^ n8172 ;
  assign n8183 = n8182 ^ n8165 ;
  assign n8186 = n8185 ^ n8183 ;
  assign n8187 = n8186 ^ n6605 ;
  assign n8198 = n8197 ^ n8187 ;
  assign n8199 = n8198 ^ n8121 ;
  assign n8122 = n8121 ^ n8109 ;
  assign n8153 = n8122 ^ n8106 ;
  assign n8154 = n8153 ^ n8122 ;
  assign n8155 = ~n8150 & ~n8154 ;
  assign n8156 = n8155 ^ n8122 ;
  assign n8157 = n7982 & n8156 ;
  assign n8200 = n8199 ^ n8157 ;
  assign n8201 = n8200 ^ x107 ;
  assign n8202 = n7959 & n8201 ;
  assign n8203 = ~n7748 & n8202 ;
  assign n8383 = n8203 ^ n8202 ;
  assign n8364 = n8363 ^ x97 ;
  assign n8365 = ~n7748 & ~n8364 ;
  assign n8378 = n8201 & n8365 ;
  assign n8379 = n8378 ^ n8365 ;
  assign n8368 = ~n7748 & ~n8201 ;
  assign n8380 = n8379 ^ n8368 ;
  assign n8374 = n7959 & n8364 ;
  assign n8376 = n8374 ^ n8364 ;
  assign n8377 = n8368 & n8376 ;
  assign n8381 = n8380 ^ n8377 ;
  assign n8369 = n8368 ^ n8201 ;
  assign n8370 = ~n7959 & ~n8369 ;
  assign n8371 = n8370 ^ n8369 ;
  assign n8372 = n8364 & ~n8371 ;
  assign n8366 = n8202 & n8365 ;
  assign n8367 = n8366 ^ n8203 ;
  assign n8373 = n8372 ^ n8367 ;
  assign n8375 = n8374 ^ n8373 ;
  assign n8382 = n8381 ^ n8375 ;
  assign n8384 = n8383 ^ n8382 ;
  assign n8449 = n8384 ^ n8366 ;
  assign n8450 = n6859 & n8449 ;
  assign n8451 = n8450 ^ n8366 ;
  assign n10597 = ~n7430 & n8451 ;
  assign n8389 = n6859 & n7430 ;
  assign n8391 = n8389 ^ n6859 ;
  assign n8398 = ~n7748 & n8376 ;
  assign n8393 = n8372 ^ n8371 ;
  assign n8394 = n8393 ^ n8365 ;
  assign n8385 = n8369 ^ n7748 ;
  assign n8386 = ~n8364 & ~n8385 ;
  assign n8392 = n8386 ^ n8364 ;
  assign n8395 = n8394 ^ n8392 ;
  assign n8396 = n8395 ^ n8370 ;
  assign n8397 = n8396 ^ n8376 ;
  assign n8399 = n8398 ^ n8397 ;
  assign n8400 = n8399 ^ n8381 ;
  assign n8401 = ~n8391 & ~n8400 ;
  assign n8390 = n8389 ^ n7430 ;
  assign n10569 = ~n8377 & ~n8390 ;
  assign n10570 = ~n8401 & ~n10569 ;
  assign n8412 = n8391 ^ n7430 ;
  assign n10565 = n8396 & ~n8412 ;
  assign n8455 = n8398 ^ n8377 ;
  assign n10556 = n8455 ^ n8395 ;
  assign n8431 = ~n7959 & n8379 ;
  assign n8432 = n8431 ^ n8379 ;
  assign n8433 = n8432 ^ n8384 ;
  assign n10557 = n10556 ^ n8433 ;
  assign n10558 = n10557 ^ n8455 ;
  assign n10559 = n8455 ^ n6859 ;
  assign n10560 = n10559 ^ n8455 ;
  assign n10561 = n10558 & n10560 ;
  assign n7431 = n7430 ^ n6859 ;
  assign n8416 = n8378 ^ n8366 ;
  assign n10548 = n8416 ^ n8373 ;
  assign n10549 = n8416 ^ n7430 ;
  assign n10550 = n10549 ^ n8416 ;
  assign n10551 = n10548 & ~n10550 ;
  assign n10552 = n10551 ^ n8416 ;
  assign n10553 = ~n7431 & n10552 ;
  assign n10554 = n10553 ^ n8455 ;
  assign n10555 = n10554 ^ n10553 ;
  assign n10562 = n10561 ^ n10555 ;
  assign n10563 = n7430 & n10562 ;
  assign n10564 = n10563 ^ n10554 ;
  assign n10566 = n10565 ^ n10564 ;
  assign n10546 = n8396 ^ n8377 ;
  assign n10547 = n8389 & n10546 ;
  assign n10567 = n10566 ^ n10547 ;
  assign n8444 = n8395 ^ n8366 ;
  assign n10544 = n8444 ^ n8432 ;
  assign n10545 = n10544 ^ n8382 ;
  assign n10568 = n10567 ^ n10545 ;
  assign n10571 = n10570 ^ n10568 ;
  assign n8387 = n8386 ^ n8384 ;
  assign n8438 = n8387 ^ n8373 ;
  assign n8439 = n8373 ^ n7430 ;
  assign n8440 = n8439 ^ n8373 ;
  assign n8441 = n8438 & ~n8440 ;
  assign n8442 = n8441 ^ n8373 ;
  assign n8443 = ~n7431 & n8442 ;
  assign n10592 = n10571 ^ n8443 ;
  assign n10586 = n8393 ^ n8387 ;
  assign n10587 = n8393 ^ n7430 ;
  assign n10588 = n10587 ^ n8393 ;
  assign n10589 = ~n10586 & n10588 ;
  assign n10590 = n10589 ^ n8393 ;
  assign n10591 = ~n6859 & ~n10590 ;
  assign n10593 = n10592 ^ n10591 ;
  assign n8429 = n8399 ^ n7430 ;
  assign n8430 = n8429 ^ n8399 ;
  assign n10580 = n8455 ^ n8399 ;
  assign n10583 = n8430 & n10580 ;
  assign n10584 = n10583 ^ n8399 ;
  assign n10585 = n7431 & n10584 ;
  assign n10594 = n10593 ^ n10585 ;
  assign n10595 = n10594 ^ n7981 ;
  assign n10572 = n10571 ^ n10567 ;
  assign n10573 = n10572 ^ n8431 ;
  assign n10574 = n10573 ^ n10572 ;
  assign n10577 = ~n6859 & n10574 ;
  assign n10578 = n10577 ^ n10572 ;
  assign n10579 = ~n7431 & n10578 ;
  assign n10596 = n10595 ^ n10579 ;
  assign n10598 = n10597 ^ n10596 ;
  assign n11604 = n10598 ^ x90 ;
  assign n12207 = n11603 & n11604 ;
  assign n12214 = n12207 ^ n11602 ;
  assign n11608 = n10351 ^ n10331 ;
  assign n11632 = n11608 ^ n10348 ;
  assign n11311 = n10344 ^ n10314 ;
  assign n11312 = n10314 ^ n10294 ;
  assign n11313 = n11312 ^ n10314 ;
  assign n11314 = n11311 & n11313 ;
  assign n11315 = n11314 ^ n10314 ;
  assign n11316 = ~n10366 & n11315 ;
  assign n11633 = n11632 ^ n11316 ;
  assign n11634 = n11633 ^ n8921 ;
  assign n11635 = n11634 ^ n10321 ;
  assign n11150 = n10344 ^ n10336 ;
  assign n11151 = n11150 ^ n10291 ;
  assign n11152 = n11151 ^ n10347 ;
  assign n11624 = n11152 ^ n10348 ;
  assign n11625 = n11624 ^ n10305 ;
  assign n11626 = n11625 ^ n10348 ;
  assign n11627 = n10348 ^ n10294 ;
  assign n11628 = n11627 ^ n10348 ;
  assign n11629 = ~n11626 & n11628 ;
  assign n11630 = n11629 ^ n10348 ;
  assign n11631 = ~n10293 & n11630 ;
  assign n11636 = n11635 ^ n11631 ;
  assign n11303 = n11151 ^ n10344 ;
  assign n11618 = n11303 ^ n10342 ;
  assign n11619 = n10342 ^ n10293 ;
  assign n11620 = n11619 ^ n10342 ;
  assign n11621 = ~n11618 & n11620 ;
  assign n11622 = n11621 ^ n10342 ;
  assign n11623 = ~n10294 & n11622 ;
  assign n11637 = n11636 ^ n11623 ;
  assign n11613 = n10314 ^ n10306 ;
  assign n11614 = n11613 ^ n10318 ;
  assign n11615 = n10294 & n11614 ;
  assign n11610 = n10318 ^ n10305 ;
  assign n11611 = n11610 ^ n10299 ;
  assign n11609 = n11608 ^ n10339 ;
  assign n11612 = n11611 ^ n11609 ;
  assign n11616 = n11615 ^ n11612 ;
  assign n11617 = n10366 & n11616 ;
  assign n11638 = n11637 ^ n11617 ;
  assign n11639 = n11638 ^ x89 ;
  assign n11640 = n11604 & ~n11639 ;
  assign n11641 = n11640 ^ n11604 ;
  assign n11642 = n11641 ^ n11639 ;
  assign n12215 = n12214 ^ n11642 ;
  assign n12209 = n11604 ^ n11565 ;
  assign n11661 = n11604 ^ n11602 ;
  assign n11606 = ~n11600 & n11604 ;
  assign n11660 = n11606 ^ n11565 ;
  assign n11662 = n11661 ^ n11660 ;
  assign n11663 = n11639 & ~n11662 ;
  assign n11664 = n11663 ^ n11660 ;
  assign n12210 = n12209 ^ n11664 ;
  assign n11643 = ~n11602 & ~n11642 ;
  assign n11644 = n11643 ^ n11639 ;
  assign n12211 = n12210 ^ n11644 ;
  assign n11605 = n11604 ^ n11603 ;
  assign n11607 = n11606 ^ n11605 ;
  assign n12205 = n11607 ^ n11565 ;
  assign n11665 = n11639 ^ n11600 ;
  assign n11666 = n11639 ^ n11604 ;
  assign n11667 = n11600 & ~n11666 ;
  assign n11668 = n11667 ^ n11565 ;
  assign n11669 = ~n11665 & ~n11668 ;
  assign n12206 = n12205 ^ n11669 ;
  assign n12208 = n12207 ^ n12206 ;
  assign n12212 = n12211 ^ n12208 ;
  assign n12213 = n12212 ^ n11639 ;
  assign n12216 = n12215 ^ n12213 ;
  assign n9808 = n9807 ^ n9803 ;
  assign n9818 = n9817 ^ n9808 ;
  assign n9820 = n9819 ^ n9817 ;
  assign n9821 = n9820 ^ n9817 ;
  assign n9822 = ~n9818 & ~n9821 ;
  assign n9823 = n9822 ^ n9817 ;
  assign n9824 = n9721 & ~n9823 ;
  assign n10611 = n9841 ^ n9811 ;
  assign n10612 = n10611 ^ n10002 ;
  assign n10613 = n10612 ^ n9994 ;
  assign n10614 = n9721 & n10613 ;
  assign n10615 = n10614 ^ n9836 ;
  assign n10607 = n9801 ^ n9765 ;
  assign n10608 = n10607 ^ n9800 ;
  assign n10609 = n10608 ^ n9768 ;
  assign n10610 = ~n9721 & n10609 ;
  assign n10616 = n10615 ^ n10610 ;
  assign n10617 = ~n9992 & n10616 ;
  assign n10618 = n10617 ^ n10614 ;
  assign n9849 = n9839 ^ n9766 ;
  assign n9868 = n9849 ^ n9829 ;
  assign n9869 = n9868 ^ n9816 ;
  assign n9838 = n9837 ^ n9826 ;
  assign n9870 = n9869 ^ n9838 ;
  assign n10601 = n9870 ^ n9868 ;
  assign n10602 = n9868 ^ n9721 ;
  assign n10603 = n10602 ^ n9868 ;
  assign n10604 = n10601 & ~n10603 ;
  assign n10605 = n10604 ^ n9868 ;
  assign n10606 = n9819 & ~n10605 ;
  assign n10619 = n10618 ^ n10606 ;
  assign n10620 = ~n10018 & ~n10619 ;
  assign n10621 = ~n9824 & n10620 ;
  assign n10622 = n10621 ^ n8093 ;
  assign n11563 = n10622 ^ x112 ;
  assign n12222 = n12206 ^ n11640 ;
  assign n11645 = n11603 ^ n11600 ;
  assign n11646 = ~n11639 & ~n11645 ;
  assign n12221 = n11667 ^ n11646 ;
  assign n12223 = n12222 ^ n12221 ;
  assign n11647 = n11646 ^ n11600 ;
  assign n11648 = ~n11604 & ~n11647 ;
  assign n11649 = n11648 ^ n11644 ;
  assign n11650 = n11649 ^ n11642 ;
  assign n12220 = n11660 ^ n11650 ;
  assign n12224 = n12223 ^ n12220 ;
  assign n12225 = n11563 & n12224 ;
  assign n12226 = n12225 ^ n12223 ;
  assign n12217 = n12213 ^ n12211 ;
  assign n12218 = ~n11563 & n12217 ;
  assign n12219 = n12218 ^ n12211 ;
  assign n12227 = n12226 ^ n12219 ;
  assign n9663 = n9535 ^ n9533 ;
  assign n9664 = n9663 ^ n9535 ;
  assign n9665 = n9581 & n9664 ;
  assign n9666 = n9665 ^ n9535 ;
  assign n9667 = ~n9580 & n9666 ;
  assign n10949 = n9552 & n9608 ;
  assign n10946 = n9588 ^ n9540 ;
  assign n10947 = n10946 ^ n9614 ;
  assign n10948 = n10947 ^ n9583 ;
  assign n10950 = n10949 ^ n10948 ;
  assign n9615 = n9614 ^ n9534 ;
  assign n9616 = n9615 ^ n9540 ;
  assign n10951 = n10950 ^ n9616 ;
  assign n10952 = n10951 ^ n9533 ;
  assign n10953 = n10952 ^ n10950 ;
  assign n10954 = n10950 ^ n9580 ;
  assign n10955 = n10954 ^ n10950 ;
  assign n10956 = n10953 & ~n10955 ;
  assign n10957 = n10956 ^ n10950 ;
  assign n10958 = ~n9581 & n10957 ;
  assign n10959 = n10958 ^ n10950 ;
  assign n10967 = n10959 ^ n9546 ;
  assign n10960 = n9592 ^ n9581 ;
  assign n10961 = n10960 ^ n9592 ;
  assign n10962 = n9977 ^ n9609 ;
  assign n10963 = n10962 ^ n9592 ;
  assign n10964 = ~n10961 & n10963 ;
  assign n10965 = n10964 ^ n9592 ;
  assign n10966 = ~n10959 & n10965 ;
  assign n10968 = n10967 ^ n10966 ;
  assign n10969 = n9618 & ~n10968 ;
  assign n10970 = n10969 ^ n10967 ;
  assign n10973 = n9597 ^ n9548 ;
  assign n10974 = n10973 ^ n9537 ;
  assign n10975 = n9581 & ~n10974 ;
  assign n10976 = n10975 ^ n9537 ;
  assign n10977 = n9580 & n10976 ;
  assign n10978 = n10977 ^ n9537 ;
  assign n10979 = ~n10970 & ~n10978 ;
  assign n10980 = ~n9667 & n10979 ;
  assign n10981 = n10980 ^ n7533 ;
  assign n11562 = n10981 ^ x65 ;
  assign n12228 = n12226 ^ n11562 ;
  assign n12229 = n12228 ^ n12226 ;
  assign n12230 = n12227 & n12229 ;
  assign n12231 = n12230 ^ n12226 ;
  assign n12232 = ~n12216 & ~n12231 ;
  assign n12233 = n12232 ^ n9527 ;
  assign n13146 = n12233 ^ x108 ;
  assign n13147 = n13145 & ~n13146 ;
  assign n13148 = n13147 ^ n13145 ;
  assign n13149 = n13148 ^ n13146 ;
  assign n10838 = n10177 ^ n10167 ;
  assign n10833 = n10147 ^ n10125 ;
  assign n10839 = n10838 ^ n10833 ;
  assign n10840 = n10131 & n10839 ;
  assign n10841 = n10840 ^ n10838 ;
  assign n10844 = n10841 ^ n10161 ;
  assign n10845 = n10844 ^ n10841 ;
  assign n10846 = ~n10131 & n10845 ;
  assign n10847 = n10846 ^ n10841 ;
  assign n10848 = ~n10126 & n10847 ;
  assign n10849 = n10848 ^ n10841 ;
  assign n11130 = n11129 ^ n10849 ;
  assign n11108 = n10171 ^ n10163 ;
  assign n11109 = n11108 ^ n11107 ;
  assign n11110 = n11109 ^ n10196 ;
  assign n11112 = n11111 ^ n11110 ;
  assign n11113 = n11112 ^ n11107 ;
  assign n11114 = n10126 & n11113 ;
  assign n11115 = n11114 ^ n11109 ;
  assign n11131 = n11130 ^ n11115 ;
  assign n11132 = n11131 ^ n7865 ;
  assign n11116 = n10857 ^ n10160 ;
  assign n11117 = n11116 ^ n10180 ;
  assign n11105 = n10838 ^ n10125 ;
  assign n11106 = n11105 ^ n10152 ;
  assign n11120 = n11117 ^ n11106 ;
  assign n11121 = ~n10126 & ~n11120 ;
  assign n11118 = n11117 ^ n11115 ;
  assign n11122 = n11121 ^ n11118 ;
  assign n11123 = ~n10138 & ~n11122 ;
  assign n11133 = n11132 ^ n11123 ;
  assign n11134 = n11133 ^ x85 ;
  assign n8452 = n8451 ^ n8444 ;
  assign n8453 = ~n7430 & n8452 ;
  assign n8417 = n8416 ^ n8393 ;
  assign n8402 = n8401 ^ n8367 ;
  assign n8418 = n8417 ^ n8402 ;
  assign n8413 = n8374 ^ n8365 ;
  assign n8414 = n8413 ^ n7748 ;
  assign n8415 = ~n8412 & ~n8414 ;
  assign n8419 = n8418 ^ n8415 ;
  assign n8403 = n8402 ^ n8367 ;
  assign n8405 = n8396 ^ n8381 ;
  assign n8404 = n8382 ^ n8377 ;
  assign n8406 = n8405 ^ n8404 ;
  assign n8409 = ~n8403 & ~n8406 ;
  assign n8410 = n8409 ^ n8367 ;
  assign n8411 = ~n8390 & n8410 ;
  assign n8420 = n8419 ^ n8411 ;
  assign n8445 = n8444 ^ n8420 ;
  assign n8446 = n8445 ^ n8443 ;
  assign n8434 = n8433 ^ n8399 ;
  assign n8435 = ~n8430 & n8434 ;
  assign n8436 = n8435 ^ n8399 ;
  assign n8437 = ~n7431 & n8436 ;
  assign n8447 = n8446 ^ n8437 ;
  assign n8421 = n8420 ^ n8415 ;
  assign n8388 = n8387 ^ n8379 ;
  assign n8422 = n8421 ^ n8388 ;
  assign n8423 = n8422 ^ n8421 ;
  assign n8424 = n8421 ^ n6859 ;
  assign n8425 = n8424 ^ n8421 ;
  assign n8426 = n8423 & n8425 ;
  assign n8427 = n8426 ^ n8421 ;
  assign n8428 = ~n7431 & n8427 ;
  assign n8448 = n8447 ^ n8428 ;
  assign n8454 = n8453 ^ n8448 ;
  assign n8456 = n8455 ^ n8396 ;
  assign n8457 = n8396 ^ n7430 ;
  assign n8458 = n8457 ^ n8396 ;
  assign n8459 = n8456 & ~n8458 ;
  assign n8460 = n8459 ^ n8396 ;
  assign n8461 = n7431 & n8460 ;
  assign n8462 = ~n8454 & ~n8461 ;
  assign n8463 = n8462 ^ n7828 ;
  assign n11135 = n8463 ^ x100 ;
  assign n11136 = ~n11134 & n11135 ;
  assign n11178 = n11136 ^ n11135 ;
  assign n8762 = n8761 ^ x81 ;
  assign n8804 = n8803 ^ x99 ;
  assign n8726 = n8725 ^ x123 ;
  assign n8614 = n8613 ^ x106 ;
  assign n8814 = n8726 ^ n8614 ;
  assign n8690 = n8689 ^ n5863 ;
  assign n8683 = n8682 ^ n7617 ;
  assign n8684 = n7735 & ~n8683 ;
  assign n8665 = ~n7694 & ~n7718 ;
  assign n8666 = n8665 ^ n7717 ;
  assign n8660 = n7701 ^ n7614 ;
  assign n8661 = n8660 ^ n7694 ;
  assign n8662 = n7603 & n8661 ;
  assign n8663 = n8660 & n8662 ;
  assign n8664 = n8663 ^ n8661 ;
  assign n8667 = n8666 ^ n8664 ;
  assign n8675 = n8666 ^ n7432 ;
  assign n8672 = n7626 & ~n7694 ;
  assign n8673 = n8672 ^ n7605 ;
  assign n8674 = n7432 & n8673 ;
  assign n8676 = n8675 ^ n8674 ;
  assign n8677 = n8676 ^ n7694 ;
  assign n8678 = n8677 ^ n8664 ;
  assign n8679 = n8678 ^ n8674 ;
  assign n8680 = ~n8667 & ~n8679 ;
  assign n8681 = n8680 ^ n8676 ;
  assign n8687 = n8684 ^ n8681 ;
  assign n8688 = ~n8659 & ~n8687 ;
  assign n8691 = n8690 ^ n8688 ;
  assign n8692 = n8691 ^ x105 ;
  assign n8811 = n8692 ^ n8614 ;
  assign n8619 = n8307 ^ n8288 ;
  assign n8630 = n8619 ^ n8284 ;
  assign n8631 = n8630 ^ n8310 ;
  assign n8629 = n8279 ^ n8249 ;
  assign n8632 = n8631 ^ n8629 ;
  assign n8633 = n8632 ^ n8349 ;
  assign n8634 = ~n8205 & n8633 ;
  assign n8635 = n8634 ^ n8349 ;
  assign n8636 = n8204 & n8635 ;
  assign n8615 = n8306 ^ n8302 ;
  assign n8617 = n8616 ^ n8615 ;
  assign n8618 = ~n8204 & n8617 ;
  assign n8621 = n8618 ^ n8299 ;
  assign n8620 = n8619 ^ n8618 ;
  assign n8622 = n8621 ^ n8620 ;
  assign n8625 = ~n8204 & ~n8622 ;
  assign n8626 = n8625 ^ n8621 ;
  assign n8627 = n8205 & n8626 ;
  assign n8628 = n8627 ^ n8618 ;
  assign n8637 = n8636 ^ n8628 ;
  assign n8641 = n8205 & n8302 ;
  assign n8642 = n8641 ^ n8286 ;
  assign n8643 = n8638 & n8642 ;
  assign n8644 = n8643 ^ n8286 ;
  assign n8645 = ~n8637 & n8644 ;
  assign n8646 = n8645 ^ n8637 ;
  assign n8647 = ~n8361 & ~n8646 ;
  assign n8654 = n8647 & ~n8653 ;
  assign n8655 = n8654 ^ n5827 ;
  assign n8656 = n8655 ^ x96 ;
  assign n8815 = n8811 ^ n8656 ;
  assign n8816 = ~n8726 & ~n8815 ;
  assign n8657 = n8656 ^ n8614 ;
  assign n10873 = n8816 ^ n8657 ;
  assign n10874 = ~n8814 & n10873 ;
  assign n8820 = n8726 ^ n8692 ;
  assign n8821 = n8820 ^ n8726 ;
  assign n8812 = n8811 ^ n8726 ;
  assign n8822 = n8820 ^ n8812 ;
  assign n8823 = n8822 ^ n8820 ;
  assign n8824 = ~n8821 & n8823 ;
  assign n8825 = n8824 ^ n8820 ;
  assign n8826 = n8656 & n8825 ;
  assign n8827 = n8826 ^ n8812 ;
  assign n10872 = n8827 ^ n8815 ;
  assign n10875 = n10874 ^ n10872 ;
  assign n10876 = n8804 & ~n10875 ;
  assign n10877 = n10876 ^ n8827 ;
  assign n8828 = n8692 ^ n8656 ;
  assign n8806 = n8614 & n8692 ;
  assign n8829 = n8806 ^ n8726 ;
  assign n8830 = ~n8828 & ~n8829 ;
  assign n10870 = n8830 ^ n8657 ;
  assign n10865 = n8614 & ~n8656 ;
  assign n10866 = n10865 ^ n8692 ;
  assign n10867 = ~n8820 & ~n10866 ;
  assign n10868 = n10867 ^ n8692 ;
  assign n10869 = ~n8804 & n10868 ;
  assign n10871 = n10870 ^ n10869 ;
  assign n10879 = n10877 ^ n10871 ;
  assign n10880 = n8762 & ~n10879 ;
  assign n10881 = n10880 ^ n10877 ;
  assign n11137 = n10881 ^ n7870 ;
  assign n11138 = n11137 ^ x91 ;
  assign n11172 = n10321 ^ n7157 ;
  assign n11173 = n11172 ^ n10330 ;
  assign n11157 = n10310 ^ n10306 ;
  assign n11154 = n10369 ^ n10339 ;
  assign n11153 = n11152 ^ n10316 ;
  assign n11155 = n11154 ^ n11153 ;
  assign n11158 = n11157 ^ n11155 ;
  assign n11159 = n10293 & ~n11158 ;
  assign n11156 = n11155 ^ n10291 ;
  assign n11160 = n11159 ^ n11156 ;
  assign n11161 = ~n10294 & ~n11160 ;
  assign n11142 = n10309 ^ n10288 ;
  assign n11143 = n10309 ^ n10294 ;
  assign n11144 = n11143 ^ n10309 ;
  assign n11145 = n11142 & n11144 ;
  assign n11146 = n11145 ^ n10309 ;
  assign n11147 = n10366 & n11146 ;
  assign n11148 = n11147 ^ n10291 ;
  assign n11141 = ~n10293 & n10316 ;
  assign n11149 = n11148 ^ n11141 ;
  assign n11162 = n11161 ^ n11149 ;
  assign n11140 = n10295 & ~n10334 ;
  assign n11163 = n11162 ^ n11140 ;
  assign n11139 = n10294 & n10299 ;
  assign n11164 = n11163 ^ n11139 ;
  assign n11165 = n10339 ^ n10307 ;
  assign n11166 = n10339 ^ n10294 ;
  assign n11167 = n11166 ^ n10339 ;
  assign n11168 = n11165 & ~n11167 ;
  assign n11169 = n11168 ^ n10339 ;
  assign n11170 = ~n10366 & n11169 ;
  assign n11171 = ~n11164 & ~n11170 ;
  assign n11174 = n11173 ^ n11171 ;
  assign n11175 = n11174 ^ x78 ;
  assign n11176 = n11138 & ~n11175 ;
  assign n11189 = n11176 ^ n11175 ;
  assign n11190 = n11178 & ~n11189 ;
  assign n11195 = n11190 ^ n11189 ;
  assign n11179 = n11178 ^ n11134 ;
  assign n11193 = n11176 & n11179 ;
  assign n11177 = n11136 & n11176 ;
  assign n11194 = n11193 ^ n11177 ;
  assign n11196 = n11195 ^ n11194 ;
  assign n11187 = n11136 ^ n11134 ;
  assign n11188 = n11176 & ~n11187 ;
  assign n11191 = n11190 ^ n11188 ;
  assign n11192 = n11191 ^ n11175 ;
  assign n11197 = n11196 ^ n11192 ;
  assign n11198 = n11197 ^ n11188 ;
  assign n11096 = n9053 ^ n9049 ;
  assign n11097 = ~n9070 & ~n11096 ;
  assign n11087 = n9062 ^ n9037 ;
  assign n11088 = n11087 ^ n8893 ;
  assign n11089 = n11088 ^ n9062 ;
  assign n11092 = n9066 & ~n11089 ;
  assign n11093 = n11092 ^ n9062 ;
  assign n11094 = ~n9109 & n11093 ;
  assign n11085 = n9119 ^ n9047 ;
  assign n11086 = n11085 ^ n10802 ;
  assign n11095 = n11094 ^ n11086 ;
  assign n11098 = n11097 ^ n11095 ;
  assign n11082 = ~n9043 & n9067 ;
  assign n11083 = n11082 ^ n9042 ;
  assign n11084 = n9109 & ~n11083 ;
  assign n11099 = n11098 ^ n11084 ;
  assign n11100 = n11099 ^ n7003 ;
  assign n11078 = n9044 ^ n9039 ;
  assign n11079 = ~n9067 & n11078 ;
  assign n11101 = n11100 ^ n11079 ;
  assign n11102 = n11101 ^ x118 ;
  assign n9402 = n9187 & n9401 ;
  assign n9389 = n9368 ^ n9333 ;
  assign n9390 = ~n9188 & n9389 ;
  assign n9391 = n9390 ^ n9337 ;
  assign n9392 = n9373 ^ n9367 ;
  assign n9393 = n9188 & n9392 ;
  assign n9394 = n9393 ^ n9154 ;
  assign n9395 = ~n9391 & n9394 ;
  assign n9380 = n9366 ^ n9325 ;
  assign n9379 = n9378 ^ n9372 ;
  assign n9381 = n9380 ^ n9379 ;
  assign n9382 = n9381 ^ n9378 ;
  assign n9383 = n9378 ^ n9185 ;
  assign n9384 = n9383 ^ n9378 ;
  assign n9385 = ~n9382 & ~n9384 ;
  assign n9386 = n9385 ^ n9378 ;
  assign n9387 = ~n9354 & n9386 ;
  assign n9388 = n9387 ^ n9378 ;
  assign n9396 = n9395 ^ n9388 ;
  assign n9350 = n9349 ^ n9344 ;
  assign n9352 = n9351 ^ n9350 ;
  assign n9353 = ~n9348 & n9352 ;
  assign n9397 = n9396 ^ n9353 ;
  assign n9346 = n9345 ^ n9341 ;
  assign n9347 = n9186 & n9346 ;
  assign n9398 = n9397 ^ n9347 ;
  assign n9403 = n9402 ^ n9398 ;
  assign n9405 = n9340 ^ n9187 ;
  assign n9406 = n9378 ^ n9154 ;
  assign n9409 = ~n9340 & ~n9406 ;
  assign n9410 = n9409 ^ n9154 ;
  assign n9411 = n9405 & n9410 ;
  assign n9412 = n9411 ^ n9187 ;
  assign n9404 = n9186 & n9399 ;
  assign n9413 = n9412 ^ n9404 ;
  assign n9414 = ~n9403 & ~n9413 ;
  assign n9415 = ~n9329 & n9414 ;
  assign n9416 = n9374 ^ n9368 ;
  assign n9417 = n9374 ^ n9185 ;
  assign n9418 = n9417 ^ n9374 ;
  assign n9419 = n9416 & n9418 ;
  assign n9420 = n9419 ^ n9374 ;
  assign n9421 = ~n9154 & n9420 ;
  assign n9422 = n9415 & ~n9421 ;
  assign n9423 = n9422 ^ n7792 ;
  assign n11103 = n9423 ^ x109 ;
  assign n11238 = n11102 & ~n11103 ;
  assign n11811 = n11198 & n11238 ;
  assign n11995 = n11811 ^ n9579 ;
  assign n11217 = n11179 & ~n11189 ;
  assign n11212 = n11136 & ~n11189 ;
  assign n11218 = n11217 ^ n11212 ;
  assign n11219 = n11218 ^ n11195 ;
  assign n11220 = n11219 ^ n11191 ;
  assign n11208 = n11189 ^ n11138 ;
  assign n11209 = ~n11187 & n11208 ;
  assign n11180 = n11176 ^ n11138 ;
  assign n11199 = n11136 & n11180 ;
  assign n11200 = n11199 ^ n11198 ;
  assign n11183 = ~n11134 & ~n11175 ;
  assign n11184 = n11183 ^ n11135 ;
  assign n11185 = ~n11138 & n11184 ;
  assign n11186 = n11185 ^ n11184 ;
  assign n11201 = n11200 ^ n11186 ;
  assign n11210 = n11209 ^ n11201 ;
  assign n11213 = n11212 ^ n11210 ;
  assign n11214 = n11213 ^ n11193 ;
  assign n11211 = n11210 ^ n11200 ;
  assign n11215 = n11214 ^ n11211 ;
  assign n11207 = n11176 ^ n11136 ;
  assign n11216 = n11215 ^ n11207 ;
  assign n11221 = n11220 ^ n11216 ;
  assign n11206 = n11188 ^ n11185 ;
  assign n11222 = n11221 ^ n11206 ;
  assign n11181 = n11179 & n11180 ;
  assign n11203 = n11199 ^ n11181 ;
  assign n11202 = n11201 ^ n11180 ;
  assign n11204 = n11203 ^ n11202 ;
  assign n11262 = n11222 ^ n11204 ;
  assign n11263 = n11204 ^ n11102 ;
  assign n11264 = n11263 ^ n11204 ;
  assign n11265 = ~n11262 & ~n11264 ;
  assign n11266 = n11265 ^ n11204 ;
  assign n11267 = n11103 & n11266 ;
  assign n11996 = n11995 ^ n11267 ;
  assign n11786 = n11217 ^ n11102 ;
  assign n11787 = n11786 ^ n11217 ;
  assign n11788 = n11218 ^ n11217 ;
  assign n11789 = n11788 ^ n11217 ;
  assign n11790 = ~n11787 & n11789 ;
  assign n11791 = n11790 ^ n11217 ;
  assign n11792 = n11103 & n11791 ;
  assign n11240 = n11238 ^ n11102 ;
  assign n11239 = n11238 ^ n11103 ;
  assign n11241 = n11240 ^ n11239 ;
  assign n11991 = n11203 & n11241 ;
  assign n11987 = n11217 ^ n11210 ;
  assign n11988 = n11987 ^ n11190 ;
  assign n11989 = n11238 & n11988 ;
  assign n11223 = n11222 ^ n11194 ;
  assign n11224 = n11223 ^ n11210 ;
  assign n11976 = n11224 ^ n11197 ;
  assign n11974 = n11193 ^ n11191 ;
  assign n11975 = n11974 ^ n11209 ;
  assign n11977 = n11976 ^ n11975 ;
  assign n11978 = n11102 & ~n11977 ;
  assign n11979 = n11978 ^ n11975 ;
  assign n11990 = n11989 ^ n11979 ;
  assign n11992 = n11991 ^ n11990 ;
  assign n11225 = n11224 ^ n11212 ;
  assign n11228 = n11225 ^ n11191 ;
  assign n11982 = n11979 ^ n11228 ;
  assign n11983 = n11982 ^ n11979 ;
  assign n11984 = ~n11102 & n11983 ;
  assign n11985 = n11984 ^ n11979 ;
  assign n11986 = ~n11103 & n11985 ;
  assign n11993 = n11992 ^ n11986 ;
  assign n11994 = ~n11792 & ~n11993 ;
  assign n11997 = n11996 ^ n11994 ;
  assign n13150 = n11997 ^ x69 ;
  assign n10600 = n10384 ^ x121 ;
  assign n10623 = n10622 ^ x97 ;
  assign n10624 = n9990 ^ x88 ;
  assign n10625 = ~n10623 & n10624 ;
  assign n10626 = n10625 ^ n10624 ;
  assign n10627 = n10626 ^ n10623 ;
  assign n8727 = n8692 & ~n8726 ;
  assign n8728 = n8657 & n8727 ;
  assign n10643 = n8728 ^ n8002 ;
  assign n8833 = n8726 ^ n8656 ;
  assign n8831 = n8830 ^ n8827 ;
  assign n8817 = n8816 ^ n8692 ;
  assign n8818 = n8814 & n8817 ;
  assign n8819 = n8818 ^ n8815 ;
  assign n8832 = n8831 ^ n8819 ;
  assign n8834 = n8833 ^ n8832 ;
  assign n10644 = n10643 ^ n8834 ;
  assign n8842 = n8692 & n8815 ;
  assign n8843 = n8842 ^ n8656 ;
  assign n8844 = ~n8812 & n8843 ;
  assign n8845 = n8844 ^ n8726 ;
  assign n10636 = n8845 ^ n8834 ;
  assign n8835 = n8834 ^ n8819 ;
  assign n10637 = n10636 ^ n8835 ;
  assign n10638 = n8835 ^ n8762 ;
  assign n10639 = n10638 ^ n8835 ;
  assign n10640 = n10637 & n10639 ;
  assign n10641 = n10640 ^ n8835 ;
  assign n10642 = ~n8804 & n10641 ;
  assign n10645 = n10644 ^ n10642 ;
  assign n10628 = n8834 ^ n8728 ;
  assign n8807 = n8806 ^ n8692 ;
  assign n8808 = n8807 ^ n8727 ;
  assign n8809 = n8808 ^ n8726 ;
  assign n8810 = ~n8656 & n8809 ;
  assign n8813 = n8812 ^ n8810 ;
  assign n10629 = n10628 ^ n8813 ;
  assign n10630 = n10629 ^ n8728 ;
  assign n10633 = n8804 & ~n10630 ;
  assign n10634 = n10633 ^ n8728 ;
  assign n10635 = ~n8762 & n10634 ;
  assign n10646 = n10645 ^ n10635 ;
  assign n10647 = n10646 ^ x115 ;
  assign n10669 = n10466 ^ n9380 ;
  assign n10655 = n9390 ^ n9351 ;
  assign n10656 = ~n9345 & ~n10436 ;
  assign n10657 = n10655 & n10656 ;
  assign n10658 = n10657 ^ n10436 ;
  assign n10670 = n10669 ^ n10658 ;
  assign n10671 = n10670 ^ n9413 ;
  assign n10660 = n9356 ^ n9249 ;
  assign n10661 = n10660 ^ n9366 ;
  assign n10662 = n10661 ^ n10658 ;
  assign n10659 = n10658 ^ n9332 ;
  assign n10663 = n10662 ^ n10659 ;
  assign n10664 = n10662 ^ n9185 ;
  assign n10665 = n10664 ^ n10662 ;
  assign n10666 = ~n10663 & n10665 ;
  assign n10667 = n10666 ^ n10662 ;
  assign n10668 = ~n9154 & n10667 ;
  assign n10672 = n10671 ^ n10668 ;
  assign n10648 = n9380 ^ n9328 ;
  assign n10649 = n10648 ^ n9380 ;
  assign n10650 = n9380 ^ n9185 ;
  assign n10651 = n10650 ^ n9380 ;
  assign n10652 = n10649 & n10651 ;
  assign n10653 = n10652 ^ n9380 ;
  assign n10654 = ~n9354 & n10653 ;
  assign n10673 = n10672 ^ n10654 ;
  assign n10674 = ~n9329 & n10673 ;
  assign n10675 = ~n9421 & n10674 ;
  assign n10676 = n10675 ^ n8029 ;
  assign n10677 = n10676 ^ x114 ;
  assign n10678 = n10647 & n10677 ;
  assign n10691 = n10627 & n10678 ;
  assign n10692 = n10691 ^ n10624 ;
  assign n10686 = n10627 & ~n10677 ;
  assign n10682 = n10625 ^ n10623 ;
  assign n10687 = n10686 ^ n10682 ;
  assign n10693 = n10692 ^ n10687 ;
  assign n10688 = ~n10647 & ~n10687 ;
  assign n10689 = n10688 ^ n10682 ;
  assign n10683 = n10678 ^ n10647 ;
  assign n10684 = ~n10682 & n10683 ;
  assign n10679 = n10678 ^ n10677 ;
  assign n10680 = n10679 ^ n10647 ;
  assign n10681 = n10627 & ~n10680 ;
  assign n10685 = n10684 ^ n10681 ;
  assign n10690 = n10689 ^ n10685 ;
  assign n10694 = n10693 ^ n10690 ;
  assign n10749 = n10694 ^ n10678 ;
  assign n10714 = n10625 & n10679 ;
  assign n10707 = n10691 ^ n10684 ;
  assign n10708 = n10707 ^ n10681 ;
  assign n10704 = n10677 ^ n10647 ;
  assign n10705 = ~n10624 & ~n10704 ;
  assign n10706 = n10705 ^ n10682 ;
  assign n10709 = n10708 ^ n10706 ;
  assign n10699 = n10625 & ~n10680 ;
  assign n10710 = n10709 ^ n10699 ;
  assign n10711 = n10710 ^ n10680 ;
  assign n10712 = n10711 ^ n10688 ;
  assign n10715 = n10714 ^ n10712 ;
  assign n10716 = n10715 ^ n10699 ;
  assign n10695 = n10625 & n10678 ;
  assign n10717 = n10716 ^ n10695 ;
  assign n10713 = n10712 ^ n10625 ;
  assign n10718 = n10717 ^ n10713 ;
  assign n10703 = n10686 ^ n10681 ;
  assign n10719 = n10718 ^ n10703 ;
  assign n10702 = n10684 ^ n10683 ;
  assign n10720 = n10719 ^ n10702 ;
  assign n10701 = n10694 ^ n10681 ;
  assign n10721 = n10720 ^ n10701 ;
  assign n10700 = n10699 ^ n10681 ;
  assign n10722 = n10721 ^ n10700 ;
  assign n10723 = n10722 ^ n10624 ;
  assign n10724 = n10723 ^ n10706 ;
  assign n10697 = n10647 ^ n10623 ;
  assign n10698 = n10697 ^ n10677 ;
  assign n10725 = n10724 ^ n10698 ;
  assign n10696 = n10695 ^ n10694 ;
  assign n10726 = n10725 ^ n10696 ;
  assign n10727 = n10726 ^ n10691 ;
  assign n10750 = n10749 ^ n10727 ;
  assign n10766 = n10750 ^ n10725 ;
  assign n10767 = n10766 ^ n10690 ;
  assign n10768 = n10767 ^ n10699 ;
  assign n13159 = n10768 ^ n10715 ;
  assign n13163 = n13159 ^ n10694 ;
  assign n13164 = ~n10600 & n13163 ;
  assign n13165 = n13164 ^ n10694 ;
  assign n10746 = n10709 ^ n10681 ;
  assign n10747 = n10746 ^ n10688 ;
  assign n10748 = n10747 ^ n10693 ;
  assign n13154 = n10748 ^ n10721 ;
  assign n13155 = n10600 & n13154 ;
  assign n13156 = n13155 ^ n10721 ;
  assign n13172 = n13165 ^ n13156 ;
  assign n11767 = n10747 ^ n10703 ;
  assign n11768 = n11767 ^ n10720 ;
  assign n10599 = n10598 ^ x82 ;
  assign n11769 = n10720 ^ n10599 ;
  assign n11770 = n11769 ^ n10720 ;
  assign n11771 = ~n11768 & n11770 ;
  assign n11772 = n11771 ^ n10720 ;
  assign n11773 = n10600 & n11772 ;
  assign n13173 = n13172 ^ n11773 ;
  assign n13174 = n13173 ^ n10121 ;
  assign n11754 = n10718 ^ n10709 ;
  assign n13157 = n13156 ^ n11754 ;
  assign n13158 = n13157 ^ n13156 ;
  assign n13160 = n13159 ^ n13158 ;
  assign n13161 = n10600 & n13160 ;
  assign n13162 = n13161 ^ n13157 ;
  assign n13175 = n13174 ^ n13162 ;
  assign n10745 = n10600 ^ n10599 ;
  assign n13170 = n10703 ^ n10691 ;
  assign n13171 = n10745 & n13170 ;
  assign n13176 = n13175 ^ n13171 ;
  assign n13166 = n13165 ^ n10717 ;
  assign n13167 = n13166 ^ n13162 ;
  assign n13151 = n10717 ^ n10710 ;
  assign n13152 = n13151 ^ n10726 ;
  assign n13153 = n10600 & n13152 ;
  assign n13168 = n13167 ^ n13153 ;
  assign n13169 = ~n10599 & ~n13168 ;
  assign n13177 = n13176 ^ n13169 ;
  assign n13178 = n13177 ^ x125 ;
  assign n13179 = n13150 & ~n13178 ;
  assign n13220 = n13179 ^ n13178 ;
  assign n13223 = n13220 ^ n13150 ;
  assign n11292 = n10295 & n10305 ;
  assign n11287 = n10307 ^ n10302 ;
  assign n11288 = n11287 ^ n10307 ;
  assign n11289 = n10296 & n10343 ;
  assign n11290 = ~n11288 & n11289 ;
  assign n11291 = n11290 ^ n11287 ;
  assign n11293 = n11292 ^ n11291 ;
  assign n11317 = n11293 ^ n10290 ;
  assign n11318 = n11317 ^ n11170 ;
  assign n11319 = n11318 ^ n11316 ;
  assign n11320 = n11319 ^ n10364 ;
  assign n11302 = n10312 ^ n10290 ;
  assign n11304 = n11303 ^ n11154 ;
  assign n11305 = n11304 ^ n10296 ;
  assign n11306 = n10296 ^ n10290 ;
  assign n11307 = n11306 ^ n10296 ;
  assign n11308 = n11305 & ~n11307 ;
  assign n11309 = n11308 ^ n10296 ;
  assign n11310 = n11302 & ~n11309 ;
  assign n11321 = n11320 ^ n11310 ;
  assign n11294 = n11293 ^ n10336 ;
  assign n11295 = n11294 ^ n10346 ;
  assign n11296 = n11295 ^ n11293 ;
  assign n11297 = n11293 ^ n10294 ;
  assign n11298 = n11297 ^ n11293 ;
  assign n11299 = ~n11296 & ~n11298 ;
  assign n11300 = n11299 ^ n11293 ;
  assign n11301 = ~n10293 & n11300 ;
  assign n11322 = n11321 ^ n11301 ;
  assign n11286 = n10296 & ~n11150 ;
  assign n11323 = n11322 ^ n11286 ;
  assign n11280 = n10347 ^ n10299 ;
  assign n11281 = n10299 ^ n10294 ;
  assign n11282 = n11281 ^ n10299 ;
  assign n11283 = n11280 & n11282 ;
  assign n11284 = n11283 ^ n10299 ;
  assign n11285 = ~n10366 & n11284 ;
  assign n11324 = n11323 ^ n11285 ;
  assign n11325 = ~n10322 & ~n11324 ;
  assign n11326 = n11325 ^ n6477 ;
  assign n11327 = n11326 ^ x113 ;
  assign n8805 = n8804 ^ n8762 ;
  assign n8836 = ~n8762 & ~n8835 ;
  assign n8837 = n8836 ^ n8819 ;
  assign n8846 = n8845 ^ n8837 ;
  assign n8838 = n8837 ^ n8813 ;
  assign n8847 = n8846 ^ n8838 ;
  assign n8848 = ~n8762 & n8847 ;
  assign n8849 = n8848 ^ n8838 ;
  assign n8850 = ~n8805 & ~n8849 ;
  assign n8851 = n8850 ^ n8837 ;
  assign n8852 = ~n8728 & n8851 ;
  assign n8853 = n8852 ^ n6072 ;
  assign n11278 = n8853 ^ x104 ;
  assign n11279 = n10470 ^ x73 ;
  assign n11332 = n11278 & ~n11279 ;
  assign n11331 = n11279 ^ n11278 ;
  assign n11333 = n11332 ^ n11331 ;
  assign n11367 = n8372 ^ n8369 ;
  assign n11368 = n11367 ^ n8381 ;
  assign n11369 = n6859 & ~n11368 ;
  assign n11370 = n11369 ^ n8395 ;
  assign n11371 = ~n7431 & n11370 ;
  assign n11352 = n8431 ^ n8366 ;
  assign n11353 = n11352 ^ n8384 ;
  assign n11348 = n10553 ^ n8391 ;
  assign n11349 = n11348 ^ n10585 ;
  assign n11337 = n8396 ^ n8393 ;
  assign n11338 = ~n10569 & ~n11337 ;
  assign n11336 = n8391 ^ n8381 ;
  assign n11339 = n11338 ^ n11336 ;
  assign n11340 = n8377 ^ n8372 ;
  assign n11341 = n11340 ^ n10569 ;
  assign n11342 = n11341 ^ n11340 ;
  assign n11343 = n11340 ^ n8381 ;
  assign n11344 = n11343 ^ n11340 ;
  assign n11345 = n11342 & n11344 ;
  assign n11346 = n11345 ^ n11340 ;
  assign n11347 = n11339 & ~n11346 ;
  assign n11350 = n11349 ^ n11347 ;
  assign n11354 = n11353 ^ n11350 ;
  assign n11364 = n11354 ^ n10591 ;
  assign n11351 = n11350 ^ n10580 ;
  assign n11355 = n11354 ^ n11351 ;
  assign n11356 = n11355 ^ n10544 ;
  assign n11357 = n11356 ^ n10580 ;
  assign n11358 = n11357 ^ n11355 ;
  assign n11359 = n11355 ^ n6859 ;
  assign n11360 = n11359 ^ n11355 ;
  assign n11361 = n11358 & n11360 ;
  assign n11362 = n11361 ^ n11355 ;
  assign n11363 = ~n7431 & n11362 ;
  assign n11365 = n11364 ^ n11363 ;
  assign n11335 = n8391 & n8416 ;
  assign n11366 = n11365 ^ n11335 ;
  assign n11372 = n11371 ^ n11366 ;
  assign n11373 = ~n8437 & ~n11372 ;
  assign n11374 = n11373 ^ n6773 ;
  assign n11375 = n11374 ^ x123 ;
  assign n11379 = n11333 & n11375 ;
  assign n11389 = n11379 ^ n11375 ;
  assign n11385 = n11278 & n11375 ;
  assign n11390 = n11389 ^ n11385 ;
  assign n11391 = n11327 & n11390 ;
  assign n11376 = n11327 & ~n11375 ;
  assign n11377 = n11333 & n11376 ;
  assign n11328 = n11279 & ~n11327 ;
  assign n11329 = n11278 & n11328 ;
  assign n11330 = n11329 ^ n11328 ;
  assign n11334 = n11333 ^ n11330 ;
  assign n11378 = n11377 ^ n11334 ;
  assign n11392 = n11391 ^ n11378 ;
  assign n11387 = n11328 & n11385 ;
  assign n11383 = n11332 & ~n11375 ;
  assign n11384 = n11383 ^ n11332 ;
  assign n11386 = n11385 ^ n11384 ;
  assign n11388 = n11387 ^ n11386 ;
  assign n11393 = n11392 ^ n11388 ;
  assign n11382 = n11376 ^ n11327 ;
  assign n11394 = n11393 ^ n11382 ;
  assign n11410 = n11394 ^ n11384 ;
  assign n11411 = n11410 ^ n11387 ;
  assign n9857 = n9843 ^ n9829 ;
  assign n9858 = n9857 ^ n9804 ;
  assign n9859 = n9858 ^ n9808 ;
  assign n9860 = n9859 ^ n9800 ;
  assign n9840 = n9839 ^ n9838 ;
  assign n9845 = n9844 ^ n9840 ;
  assign n9863 = n9860 ^ n9845 ;
  assign n9864 = n9721 & ~n9863 ;
  assign n9847 = n9846 ^ n9831 ;
  assign n9850 = n9849 ^ n9848 ;
  assign n9851 = n9848 ^ n9846 ;
  assign n9852 = n9851 ^ n9848 ;
  assign n9853 = ~n9850 & ~n9852 ;
  assign n9854 = n9853 ^ n9848 ;
  assign n9855 = n9847 & n9854 ;
  assign n9856 = n9855 ^ n9831 ;
  assign n9861 = n9860 ^ n9856 ;
  assign n9865 = n9864 ^ n9861 ;
  assign n9872 = n9865 ^ n9856 ;
  assign n9871 = ~n9721 & ~n9870 ;
  assign n9873 = n9872 ^ n9871 ;
  assign n9874 = ~n9819 & ~n9873 ;
  assign n9833 = n9832 ^ n9824 ;
  assign n9866 = n9865 ^ n9833 ;
  assign n9867 = n9866 ^ n5785 ;
  assign n9875 = n9874 ^ n9867 ;
  assign n11275 = n9875 ^ x99 ;
  assign n11276 = n10204 ^ x106 ;
  assign n11401 = n11275 & ~n11276 ;
  assign n11402 = n11401 ^ n11275 ;
  assign n11403 = n11402 ^ n11276 ;
  assign n11835 = n11403 ^ n11275 ;
  assign n13213 = n11411 & ~n11835 ;
  assign n11420 = n11391 ^ n11390 ;
  assign n11406 = n11333 ^ n11278 ;
  assign n11407 = n11406 ^ n11390 ;
  assign n11414 = ~n11327 & ~n11407 ;
  assign n11415 = n11414 ^ n11407 ;
  assign n11416 = n11415 ^ n11377 ;
  assign n11421 = n11420 ^ n11416 ;
  assign n11424 = n11421 ^ n11378 ;
  assign n11412 = n11332 & n11376 ;
  assign n11413 = n11412 ^ n11376 ;
  assign n11417 = n11416 ^ n11413 ;
  assign n13206 = n11424 ^ n11417 ;
  assign n11380 = n11379 ^ n11378 ;
  assign n13192 = n11391 ^ n11380 ;
  assign n11442 = n11387 ^ n11329 ;
  assign n12663 = n11442 ^ n11414 ;
  assign n13193 = n13192 ^ n12663 ;
  assign n11381 = n11380 ^ n11330 ;
  assign n13190 = n11392 ^ n11381 ;
  assign n13191 = n13190 ^ n11420 ;
  assign n13194 = n13193 ^ n13191 ;
  assign n13195 = ~n11276 & n13194 ;
  assign n13196 = n13195 ^ n13191 ;
  assign n13207 = n13206 ^ n13196 ;
  assign n11461 = n11412 ^ n11383 ;
  assign n13203 = n11461 ^ n11424 ;
  assign n11446 = n11412 ^ n11387 ;
  assign n11819 = n11446 ^ n11410 ;
  assign n11820 = n11819 ^ n11388 ;
  assign n13204 = n13203 ^ n11820 ;
  assign n13205 = n11276 & ~n13204 ;
  assign n13208 = n13207 ^ n13205 ;
  assign n13209 = ~n11275 & n13208 ;
  assign n13201 = n11276 & n11461 ;
  assign n13180 = n11442 ^ n11394 ;
  assign n13197 = n13196 ^ n13180 ;
  assign n11277 = n11276 ^ n11275 ;
  assign n11845 = n11392 ^ n11276 ;
  assign n11846 = n11845 ^ n11392 ;
  assign n11847 = n11393 & ~n11846 ;
  assign n11848 = n11847 ^ n11392 ;
  assign n11849 = n11277 & n11848 ;
  assign n13198 = n13197 ^ n11849 ;
  assign n13199 = n13198 ^ n10085 ;
  assign n13200 = n13199 ^ n11417 ;
  assign n13202 = n13201 ^ n13200 ;
  assign n13210 = n13209 ^ n13202 ;
  assign n13188 = n11414 ^ n11377 ;
  assign n13189 = n11403 & n13188 ;
  assign n13211 = n13210 ^ n13189 ;
  assign n13181 = n13180 ^ n11446 ;
  assign n13182 = n13181 ^ n13180 ;
  assign n13183 = n13180 ^ n11275 ;
  assign n13184 = n13183 ^ n13180 ;
  assign n13185 = n13182 & n13184 ;
  assign n13186 = n13185 ^ n13180 ;
  assign n13187 = n11277 & n13186 ;
  assign n13212 = n13211 ^ n13187 ;
  assign n13214 = n13213 ^ n13212 ;
  assign n13215 = n13214 ^ x76 ;
  assign n10878 = n10877 ^ n8762 ;
  assign n10882 = n10881 ^ n10878 ;
  assign n10883 = n10882 ^ n10871 ;
  assign n10884 = n10883 ^ n7117 ;
  assign n12050 = n10884 ^ x69 ;
  assign n12069 = n9994 ^ n9849 ;
  assign n12068 = n9807 ^ n9802 ;
  assign n12070 = n12069 ^ n12068 ;
  assign n12071 = ~n9721 & n12070 ;
  assign n12072 = n12071 ^ n12068 ;
  assign n12080 = n12072 ^ n7054 ;
  assign n12081 = n12080 ^ n9824 ;
  assign n12082 = n12081 ^ n10026 ;
  assign n12074 = n9842 ^ n9831 ;
  assign n12075 = n12074 ^ n9837 ;
  assign n12076 = ~n10008 & n12075 ;
  assign n12073 = n12072 ^ n9813 ;
  assign n12077 = n12076 ^ n12073 ;
  assign n12065 = n9994 ^ n9814 ;
  assign n12066 = n12065 ^ n9829 ;
  assign n12067 = n9819 & ~n12066 ;
  assign n12078 = n12077 ^ n12067 ;
  assign n12079 = n9992 & n12078 ;
  assign n12083 = n12082 ^ n12079 ;
  assign n12064 = n9830 & ~n9857 ;
  assign n12084 = n12083 ^ n12064 ;
  assign n12057 = n9842 ^ n9828 ;
  assign n12056 = n9842 ^ n9817 ;
  assign n12058 = n12057 ^ n12056 ;
  assign n12059 = n12057 ^ n9721 ;
  assign n12060 = n12059 ^ n12057 ;
  assign n12061 = ~n12058 & ~n12060 ;
  assign n12062 = n12061 ^ n12057 ;
  assign n12063 = ~n9819 & n12062 ;
  assign n12088 = n12084 ^ n12063 ;
  assign n12089 = n12088 ^ x125 ;
  assign n12095 = ~n9580 & n9612 ;
  assign n12096 = n12095 ^ n9595 ;
  assign n9652 = n9588 & n9647 ;
  assign n9653 = n9652 ^ n9581 ;
  assign n9654 = ~n9614 & ~n9653 ;
  assign n9655 = n9654 ^ n9581 ;
  assign n12105 = n12096 ^ n9655 ;
  assign n9634 = n9580 ^ n9538 ;
  assign n9635 = n9634 ^ n9538 ;
  assign n9636 = n9598 & ~n9635 ;
  assign n9637 = n9636 ^ n9538 ;
  assign n9638 = n9581 & n9637 ;
  assign n12106 = n12105 ^ n9638 ;
  assign n9584 = n9552 & n9582 ;
  assign n9585 = n9584 ^ n9583 ;
  assign n12107 = n12106 ^ n9585 ;
  assign n12108 = n12107 ^ n9972 ;
  assign n12109 = n12108 ^ n7329 ;
  assign n12097 = n12096 ^ n10946 ;
  assign n9620 = n9590 ^ n9464 ;
  assign n9621 = n9542 ^ n9505 ;
  assign n9622 = n9621 ^ n9507 ;
  assign n9623 = n9620 & n9622 ;
  assign n12098 = n12097 ^ n9623 ;
  assign n12099 = n12098 ^ n12096 ;
  assign n12102 = n9580 & n12099 ;
  assign n12103 = n12102 ^ n12096 ;
  assign n12104 = n9581 & ~n12103 ;
  assign n12110 = n12109 ^ n12104 ;
  assign n12090 = n9592 ^ n9544 ;
  assign n12091 = n12090 ^ n9592 ;
  assign n12092 = n10961 & n12091 ;
  assign n12093 = n12092 ^ n9592 ;
  assign n12094 = ~n9580 & ~n12093 ;
  assign n12111 = n12110 ^ n12094 ;
  assign n12112 = n12111 ^ x110 ;
  assign n12113 = ~n12089 & ~n12112 ;
  assign n12119 = n12113 ^ n12089 ;
  assign n12052 = n11101 ^ x108 ;
  assign n10858 = n10856 & n10857 ;
  assign n10850 = n10849 ^ n10175 ;
  assign n10823 = n10177 ^ n10145 ;
  assign n10824 = n10823 ^ n10144 ;
  assign n10825 = n10824 ^ n10177 ;
  assign n10826 = ~n10126 & n10825 ;
  assign n10827 = n10826 ^ n10823 ;
  assign n10851 = n10850 ^ n10827 ;
  assign n10852 = n10851 ^ n10202 ;
  assign n10853 = n10852 ^ n7102 ;
  assign n10834 = n10833 ^ n10141 ;
  assign n10835 = ~n10126 & n10834 ;
  assign n10829 = n10827 ^ n10149 ;
  assign n10830 = n10829 ^ n10173 ;
  assign n10828 = n10827 ^ n10125 ;
  assign n10831 = n10830 ^ n10828 ;
  assign n10832 = n10831 ^ n10827 ;
  assign n10836 = n10835 ^ n10832 ;
  assign n10837 = n10138 & n10836 ;
  assign n10854 = n10853 ^ n10837 ;
  assign n10821 = n10175 ^ n10169 ;
  assign n10822 = n10126 & n10821 ;
  assign n10855 = n10854 ^ n10822 ;
  assign n10859 = n10858 ^ n10855 ;
  assign n12053 = n10859 ^ x83 ;
  assign n12054 = n12052 & n12053 ;
  assign n12055 = n12054 ^ n12053 ;
  assign n12126 = n12055 ^ n12052 ;
  assign n12127 = ~n12119 & ~n12126 ;
  assign n12116 = n12054 ^ n12052 ;
  assign n12117 = n12113 & n12116 ;
  assign n12443 = n12127 ^ n12117 ;
  assign n12114 = n12113 ^ n12112 ;
  assign n12131 = n12054 & ~n12114 ;
  assign n12115 = n12055 & ~n12114 ;
  assign n12145 = n12131 ^ n12115 ;
  assign n12143 = ~n12114 & ~n12126 ;
  assign n12144 = n12143 ^ n12114 ;
  assign n12146 = n12145 ^ n12144 ;
  assign n12133 = n12054 & n12113 ;
  assign n12120 = n12119 ^ n12112 ;
  assign n12128 = n12116 & ~n12120 ;
  assign n12129 = n12128 ^ n12127 ;
  assign n12134 = n12133 ^ n12129 ;
  assign n12122 = n12054 & ~n12119 ;
  assign n12121 = n12055 & ~n12120 ;
  assign n12123 = n12122 ^ n12121 ;
  assign n12135 = n12134 ^ n12123 ;
  assign n12132 = n12131 ^ n12121 ;
  assign n12136 = n12135 ^ n12132 ;
  assign n12130 = n12129 ^ n12054 ;
  assign n12137 = n12136 ^ n12130 ;
  assign n12141 = n12137 ^ n12121 ;
  assign n12140 = n12128 ^ n12120 ;
  assign n12142 = n12141 ^ n12140 ;
  assign n12153 = n12146 ^ n12142 ;
  assign n12147 = n12113 & ~n12126 ;
  assign n12148 = n12147 ^ n12146 ;
  assign n12149 = n12148 ^ n12142 ;
  assign n12150 = n12149 ^ n12117 ;
  assign n12151 = n12150 ^ n12133 ;
  assign n12152 = n12151 ^ n12113 ;
  assign n12154 = n12153 ^ n12152 ;
  assign n12444 = n12443 ^ n12154 ;
  assign n12049 = n11174 ^ x86 ;
  assign n12445 = n12154 ^ n12049 ;
  assign n12446 = n12445 ^ n12154 ;
  assign n12447 = n12444 & n12446 ;
  assign n12448 = n12447 ^ n12154 ;
  assign n12449 = ~n12050 & n12448 ;
  assign n12155 = n12154 ^ n12141 ;
  assign n12138 = n12137 ^ n12115 ;
  assign n12139 = n12138 ^ n12055 ;
  assign n12156 = n12155 ^ n12139 ;
  assign n12163 = n12156 ^ n12128 ;
  assign n12158 = n12147 ^ n12128 ;
  assign n12159 = n12158 ^ n12117 ;
  assign n12160 = n12159 ^ n12116 ;
  assign n12161 = n12160 ^ n12148 ;
  assign n12162 = n12161 ^ n12147 ;
  assign n12164 = n12163 ^ n12162 ;
  assign n12165 = ~n12049 & ~n12164 ;
  assign n12166 = n12165 ^ n12162 ;
  assign n12450 = n12449 ^ n12166 ;
  assign n12191 = n12049 & n12050 ;
  assign n12192 = n12191 ^ n12050 ;
  assign n12196 = n12192 ^ n12049 ;
  assign n12439 = n12161 ^ n12142 ;
  assign n12440 = ~n12196 & n12439 ;
  assign n12437 = n12196 ^ n12050 ;
  assign n12438 = n12138 & n12437 ;
  assign n12441 = n12440 ^ n12438 ;
  assign n12435 = n12156 & n12191 ;
  assign n12430 = n12131 ^ n12050 ;
  assign n12431 = n12430 ^ n12131 ;
  assign n12432 = n12145 & n12431 ;
  assign n12433 = n12432 ^ n12131 ;
  assign n12434 = ~n12049 & n12433 ;
  assign n12436 = n12435 ^ n12434 ;
  assign n12442 = n12441 ^ n12436 ;
  assign n12451 = n12450 ^ n12442 ;
  assign n12193 = n12153 & n12192 ;
  assign n12452 = n12451 ^ n12193 ;
  assign n12453 = n12452 ^ n9720 ;
  assign n12421 = n12143 ^ n12122 ;
  assign n12422 = n12421 ^ n12148 ;
  assign n12423 = n12148 ^ n12049 ;
  assign n12424 = n12423 ^ n12148 ;
  assign n12425 = ~n12422 & n12424 ;
  assign n12426 = n12425 ^ n12148 ;
  assign n12427 = ~n12050 & ~n12426 ;
  assign n12454 = n12453 ^ n12427 ;
  assign n12181 = n12154 ^ n12138 ;
  assign n12419 = n12181 ^ n12153 ;
  assign n12420 = n12191 & n12419 ;
  assign n12455 = n12454 ^ n12420 ;
  assign n12051 = n12050 ^ n12049 ;
  assign n12411 = n12166 ^ n12132 ;
  assign n12414 = n12411 ^ n12136 ;
  assign n12415 = n12414 ^ n12411 ;
  assign n12416 = ~n12049 & n12415 ;
  assign n12417 = n12416 ^ n12411 ;
  assign n12418 = n12051 & ~n12417 ;
  assign n12456 = n12455 ^ n12418 ;
  assign n13216 = n12456 ^ x126 ;
  assign n13217 = ~n13215 & n13216 ;
  assign n13218 = n13217 ^ n13215 ;
  assign n13228 = n13218 ^ n13216 ;
  assign n13233 = n13223 & n13228 ;
  assign n13231 = n13179 & n13228 ;
  assign n13224 = n13223 ^ n13178 ;
  assign n13225 = ~n13218 & n13224 ;
  assign n13226 = n13225 ^ n13218 ;
  assign n13221 = ~n13218 & ~n13220 ;
  assign n13219 = n13179 & ~n13218 ;
  assign n13222 = n13221 ^ n13219 ;
  assign n13227 = n13226 ^ n13222 ;
  assign n13232 = n13231 ^ n13227 ;
  assign n13234 = n13233 ^ n13232 ;
  assign n13230 = n13224 & n13228 ;
  assign n13235 = n13234 ^ n13230 ;
  assign n13229 = n13228 ^ n13227 ;
  assign n13236 = n13235 ^ n13229 ;
  assign n13237 = n13236 ^ n13230 ;
  assign n13238 = n13149 & n13237 ;
  assign n13262 = n13236 ^ n13231 ;
  assign n13263 = n13262 ^ n13219 ;
  assign n13264 = n13263 ^ n13233 ;
  assign n13249 = n13217 & n13224 ;
  assign n13239 = n13217 ^ n13216 ;
  assign n13246 = ~n13220 & n13239 ;
  assign n13247 = n13246 ^ n13237 ;
  assign n13244 = n13230 ^ n13221 ;
  assign n13245 = n13244 ^ n13220 ;
  assign n13248 = n13247 ^ n13245 ;
  assign n13250 = n13249 ^ n13248 ;
  assign n13240 = n13223 & n13239 ;
  assign n13241 = n13240 ^ n13231 ;
  assign n13242 = n13241 ^ n13223 ;
  assign n13243 = n13242 ^ n13234 ;
  assign n13251 = n13250 ^ n13243 ;
  assign n13265 = n13264 ^ n13251 ;
  assign n13258 = n13216 ^ n13150 ;
  assign n13259 = ~n13215 & ~n13258 ;
  assign n13260 = n13259 ^ n13224 ;
  assign n13261 = n13260 ^ n13239 ;
  assign n13266 = n13265 ^ n13261 ;
  assign n13290 = n13266 ^ n13246 ;
  assign n13291 = n13147 & ~n13290 ;
  assign n13252 = n13251 ^ n13217 ;
  assign n13253 = n13252 ^ n13243 ;
  assign n13286 = n13253 ^ n13225 ;
  assign n13287 = ~n13146 & ~n13286 ;
  assign n13267 = n13266 ^ n13250 ;
  assign n13281 = n13149 ^ n13145 ;
  assign n13282 = n13267 & ~n13281 ;
  assign n13275 = n13246 ^ n13225 ;
  assign n13276 = n13225 ^ n13145 ;
  assign n13277 = n13276 ^ n13225 ;
  assign n13278 = n13275 & n13277 ;
  assign n13279 = n13278 ^ n13225 ;
  assign n13280 = n13146 & n13279 ;
  assign n13283 = n13282 ^ n13280 ;
  assign n13257 = n13146 ^ n13145 ;
  assign n13269 = n13236 ^ n13219 ;
  assign n13272 = n13269 ^ n13221 ;
  assign n13268 = n13267 ^ n13232 ;
  assign n13270 = n13269 ^ n13268 ;
  assign n13271 = n13145 & ~n13270 ;
  assign n13273 = n13272 ^ n13271 ;
  assign n13274 = ~n13257 & n13273 ;
  assign n13284 = n13283 ^ n13274 ;
  assign n13255 = n13241 ^ n13219 ;
  assign n13256 = n13149 & n13255 ;
  assign n13285 = n13284 ^ n13256 ;
  assign n13288 = n13287 ^ n13285 ;
  assign n13254 = ~n13145 & ~n13253 ;
  assign n13289 = n13288 ^ n13254 ;
  assign n13292 = n13291 ^ n13289 ;
  assign n13293 = ~n13238 & ~n13292 ;
  assign n13294 = n13240 & ~n13281 ;
  assign n13295 = n13294 ^ n13145 ;
  assign n13296 = n13295 ^ n13294 ;
  assign n13297 = n13240 ^ n13239 ;
  assign n13298 = n13297 ^ n13290 ;
  assign n13299 = n13298 ^ n13250 ;
  assign n13300 = n13299 ^ n13234 ;
  assign n13301 = n13146 & ~n13300 ;
  assign n13302 = n13301 ^ n13234 ;
  assign n13305 = n13296 & ~n13302 ;
  assign n13306 = n13305 ^ n13294 ;
  assign n13307 = n13293 & ~n13306 ;
  assign n13308 = n13307 ^ n10859 ;
  assign n13309 = n13308 ^ x69 ;
  assign n10523 = n10420 ^ n10413 ;
  assign n10512 = ~n9991 & ~n10486 ;
  assign n10513 = n10512 ^ n10428 ;
  assign n10524 = n10523 ^ n10513 ;
  assign n10518 = n10400 ^ n10387 ;
  assign n10519 = n10518 ^ n10420 ;
  assign n10521 = n10520 ^ n10519 ;
  assign n10522 = n9991 & n10521 ;
  assign n10525 = n10524 ^ n10522 ;
  assign n10526 = ~n10471 & ~n10525 ;
  assign n10472 = ~n10424 & n10471 ;
  assign n10473 = n10472 ^ n10423 ;
  assign n10514 = n10513 ^ n10473 ;
  assign n10515 = n10514 ^ n10511 ;
  assign n10516 = n10515 ^ n10500 ;
  assign n10488 = n10487 ^ n10399 ;
  assign n10489 = n10488 ^ n10398 ;
  assign n10490 = n10398 ^ n9991 ;
  assign n10491 = n10490 ^ n10398 ;
  assign n10492 = ~n10489 & n10491 ;
  assign n10493 = n10492 ^ n10398 ;
  assign n10494 = ~n10471 & n10493 ;
  assign n10517 = n10516 ^ n10494 ;
  assign n10527 = n10526 ^ n10517 ;
  assign n10475 = n10421 ^ n10414 ;
  assign n10476 = n10475 ^ n10423 ;
  assign n10477 = n10476 ^ n10473 ;
  assign n10474 = n10473 ^ n10428 ;
  assign n10478 = n10477 ^ n10474 ;
  assign n10479 = n10477 ^ n10471 ;
  assign n10480 = n10479 ^ n10477 ;
  assign n10481 = n10478 & ~n10480 ;
  assign n10482 = n10481 ^ n10477 ;
  assign n10483 = ~n9991 & n10482 ;
  assign n10528 = n10527 ^ n10483 ;
  assign n10540 = ~n10528 & ~n10539 ;
  assign n10541 = n10540 ^ n8613 ;
  assign n12615 = n10541 ^ x74 ;
  assign n10820 = n10819 ^ x75 ;
  assign n10860 = n10859 ^ x93 ;
  assign n10861 = n10820 & ~n10860 ;
  assign n10862 = n10861 ^ n10820 ;
  assign n10931 = n9367 ^ n9343 ;
  assign n10932 = ~n9185 & n10931 ;
  assign n10928 = n9343 ^ n9324 ;
  assign n10929 = n10928 ^ n9337 ;
  assign n10922 = n9368 ^ n9185 ;
  assign n10923 = n10922 ^ n9368 ;
  assign n10924 = ~n9376 & n10923 ;
  assign n10925 = n10924 ^ n9368 ;
  assign n10926 = ~n9354 & n10925 ;
  assign n10927 = n10926 ^ n9368 ;
  assign n10930 = n10929 ^ n10927 ;
  assign n10933 = n10932 ^ n10930 ;
  assign n10934 = n10933 ^ n10927 ;
  assign n10937 = n10934 ^ n9358 ;
  assign n10938 = n10937 ^ n10934 ;
  assign n10939 = ~n9185 & n10938 ;
  assign n10940 = n10939 ^ n10934 ;
  assign n10941 = n9154 & n10940 ;
  assign n10942 = n10941 ^ n10933 ;
  assign n10943 = ~n10463 & ~n10942 ;
  assign n10919 = n10467 ^ n7488 ;
  assign n10920 = n10919 ^ n9388 ;
  assign n10944 = n10943 ^ n10920 ;
  assign n10945 = n10944 ^ x76 ;
  assign n10982 = n10981 ^ x117 ;
  assign n10983 = ~n10945 & n10982 ;
  assign n10984 = n10983 ^ n10945 ;
  assign n10985 = n10984 ^ n10982 ;
  assign n10885 = n10884 ^ x94 ;
  assign n10903 = n8388 ^ n8384 ;
  assign n10906 = n10903 ^ n8461 ;
  assign n10901 = n8377 ^ n8376 ;
  assign n10902 = n10901 ^ n8367 ;
  assign n10904 = n10903 ^ n10902 ;
  assign n10905 = n7430 & n10904 ;
  assign n10907 = n10906 ^ n10905 ;
  assign n10908 = n10907 ^ n8461 ;
  assign n10899 = n8395 ^ n8388 ;
  assign n10900 = ~n7430 & n10899 ;
  assign n10909 = n10908 ^ n10900 ;
  assign n10910 = ~n6859 & n10909 ;
  assign n10911 = n10910 ^ n10907 ;
  assign n10896 = ~n6859 & ~n8392 ;
  assign n10894 = n8393 ^ n8379 ;
  assign n10895 = n10894 ^ n8384 ;
  assign n10897 = n10896 ^ n10895 ;
  assign n10898 = n7430 & ~n10897 ;
  assign n10912 = n10911 ^ n10898 ;
  assign n10893 = n8374 & ~n8412 ;
  assign n10913 = n10912 ^ n10893 ;
  assign n10888 = n8405 ^ n6859 ;
  assign n10889 = n10888 ^ n8405 ;
  assign n10890 = n8406 & ~n10889 ;
  assign n10891 = n10890 ^ n8405 ;
  assign n10892 = n7431 & n10891 ;
  assign n10914 = n10913 ^ n10892 ;
  assign n10915 = ~n10585 & ~n10914 ;
  assign n10916 = n10915 ^ n7593 ;
  assign n10917 = n10916 ^ x124 ;
  assign n10918 = ~n10885 & n10917 ;
  assign n10987 = n10918 ^ n10885 ;
  assign n10993 = n10985 & ~n10987 ;
  assign n10986 = n10918 & n10985 ;
  assign n11024 = n10993 ^ n10986 ;
  assign n10988 = n10987 ^ n10917 ;
  assign n10989 = n10985 & n10988 ;
  assign n11023 = n10989 ^ n10985 ;
  assign n11025 = n11024 ^ n11023 ;
  assign n10997 = n10918 & n10983 ;
  assign n10991 = n10985 ^ n10945 ;
  assign n10992 = n10988 & n10991 ;
  assign n10994 = n10993 ^ n10992 ;
  assign n11016 = n10997 ^ n10994 ;
  assign n11010 = n10983 ^ n10917 ;
  assign n11013 = n10945 ^ n10917 ;
  assign n11011 = n10982 ^ n10885 ;
  assign n11012 = n11011 ^ n10917 ;
  assign n11014 = n11013 ^ n11012 ;
  assign n11015 = ~n11010 & n11014 ;
  assign n11017 = n11016 ^ n11015 ;
  assign n11018 = n11017 ^ n10986 ;
  assign n11007 = n10918 & n10991 ;
  assign n11008 = n11007 ^ n10992 ;
  assign n10999 = n10988 ^ n10885 ;
  assign n11005 = n10991 & n10999 ;
  assign n11006 = n11005 ^ n10991 ;
  assign n11009 = n11008 ^ n11006 ;
  assign n11019 = n11018 ^ n11009 ;
  assign n11020 = n11019 ^ n10917 ;
  assign n11000 = n10983 & n10999 ;
  assign n10995 = n10983 & ~n10987 ;
  assign n11001 = n11000 ^ n10995 ;
  assign n10998 = n10997 ^ n10983 ;
  assign n11002 = n11001 ^ n10998 ;
  assign n10996 = n10995 ^ n10994 ;
  assign n11003 = n11002 ^ n10996 ;
  assign n10990 = n10989 ^ n10986 ;
  assign n11004 = n11003 ^ n10990 ;
  assign n11021 = n11020 ^ n11004 ;
  assign n12044 = n11025 ^ n11021 ;
  assign n12045 = n10862 & ~n12044 ;
  assign n12742 = n12045 ^ n10989 ;
  assign n12725 = n11016 ^ n11005 ;
  assign n12732 = n12725 ^ n11018 ;
  assign n11535 = n11005 ^ n10995 ;
  assign n11536 = n11535 ^ n11009 ;
  assign n12726 = n11536 ^ n10992 ;
  assign n12727 = n12726 ^ n12725 ;
  assign n11527 = n10860 ^ n10820 ;
  assign n12728 = n12725 ^ n10860 ;
  assign n12729 = ~n11527 & n12728 ;
  assign n12730 = n12729 ^ n10860 ;
  assign n12731 = n12727 & n12730 ;
  assign n12733 = n12732 ^ n12731 ;
  assign n12743 = n12742 ^ n12733 ;
  assign n11026 = n11025 ^ n10999 ;
  assign n11022 = n11005 ^ n11000 ;
  assign n11027 = n11026 ^ n11022 ;
  assign n11521 = n11027 ^ n10997 ;
  assign n11522 = n10997 ^ n10860 ;
  assign n11523 = n11522 ^ n10997 ;
  assign n11524 = n11521 & ~n11523 ;
  assign n11525 = n11524 ^ n10997 ;
  assign n11526 = n10820 & n11525 ;
  assign n12744 = n12743 ^ n11526 ;
  assign n10863 = n10862 ^ n10860 ;
  assign n10864 = n10863 ^ n10861 ;
  assign n12018 = n10993 ^ n10860 ;
  assign n12019 = n12018 ^ n10993 ;
  assign n12020 = n10994 & n12019 ;
  assign n12021 = n12020 ^ n10993 ;
  assign n12022 = ~n10864 & n12021 ;
  assign n12745 = n12744 ^ n12022 ;
  assign n12736 = n11022 ^ n10984 ;
  assign n11028 = n11027 ^ n11021 ;
  assign n12737 = n12736 ^ n11028 ;
  assign n11051 = n11007 ^ n11002 ;
  assign n12738 = n12737 ^ n11051 ;
  assign n12739 = ~n10860 & n12738 ;
  assign n12734 = n12733 ^ n10984 ;
  assign n12735 = n12734 ^ n11028 ;
  assign n12740 = n12739 ^ n12735 ;
  assign n12741 = ~n10864 & n12740 ;
  assign n12746 = n12745 ^ n12741 ;
  assign n12719 = n10989 ^ n10860 ;
  assign n12720 = n12719 ^ n10989 ;
  assign n12722 = n11002 & n12720 ;
  assign n12723 = n12722 ^ n10989 ;
  assign n12724 = n10820 & n12723 ;
  assign n12747 = n12746 ^ n12724 ;
  assign n12748 = n12747 ^ n11000 ;
  assign n12749 = n12748 ^ n12747 ;
  assign n11035 = n11028 ^ n11018 ;
  assign n11036 = n11035 ^ n11024 ;
  assign n11034 = n10993 ^ n10984 ;
  assign n11037 = n11036 ^ n11034 ;
  assign n12750 = n12749 ^ n11037 ;
  assign n12751 = n10820 & n12750 ;
  assign n12752 = n12751 ^ n12748 ;
  assign n12760 = n12752 ^ n7747 ;
  assign n12753 = n12752 ^ n12747 ;
  assign n12754 = n12753 ^ n12752 ;
  assign n11029 = n11028 ^ n11009 ;
  assign n11030 = ~n10860 & ~n11029 ;
  assign n11031 = n11030 ^ n11009 ;
  assign n12755 = n12752 ^ n11031 ;
  assign n12756 = n12755 ^ n12752 ;
  assign n12757 = ~n12754 & ~n12756 ;
  assign n12758 = n12757 ^ n12752 ;
  assign n12759 = ~n11527 & ~n12758 ;
  assign n12761 = n12760 ^ n12759 ;
  assign n12762 = n12761 ^ x113 ;
  assign n12789 = ~n12615 & ~n12762 ;
  assign n12796 = n12789 ^ n12615 ;
  assign n11254 = n11222 ^ n11203 ;
  assign n11255 = n11254 ^ n11208 ;
  assign n11252 = n11209 ^ n11203 ;
  assign n11253 = n11252 ^ n11216 ;
  assign n11256 = n11255 ^ n11253 ;
  assign n11268 = n11240 & ~n11256 ;
  assign n11269 = ~n11267 & n11268 ;
  assign n11270 = n11269 ^ n11267 ;
  assign n11257 = n11256 ^ n11190 ;
  assign n11258 = ~n11239 & ~n11257 ;
  assign n11249 = n11239 ^ n11102 ;
  assign n11250 = n11219 ^ n11197 ;
  assign n11251 = n11249 & ~n11250 ;
  assign n11259 = n11258 ^ n11251 ;
  assign n11182 = n11181 ^ n11177 ;
  assign n11205 = n11204 ^ n11182 ;
  assign n11226 = n11225 ^ n11205 ;
  assign n11227 = n11103 & n11226 ;
  assign n11229 = n11228 ^ n11227 ;
  assign n11260 = n11259 ^ n11229 ;
  assign n11242 = n11191 ^ n11103 ;
  assign n11243 = n11242 ^ n11191 ;
  assign n11246 = ~n11220 & ~n11243 ;
  assign n11247 = n11246 ^ n11191 ;
  assign n11248 = ~n11241 & n11247 ;
  assign n11261 = n11260 ^ n11248 ;
  assign n11271 = n11270 ^ n11261 ;
  assign n11272 = n11271 ^ n8803 ;
  assign n11104 = n11103 ^ n11102 ;
  assign n11230 = n11229 ^ n11214 ;
  assign n11231 = n11230 ^ n11215 ;
  assign n11232 = n11231 ^ n11230 ;
  assign n11233 = n11230 ^ n11102 ;
  assign n11234 = n11233 ^ n11230 ;
  assign n11235 = n11232 & ~n11234 ;
  assign n11236 = n11235 ^ n11230 ;
  assign n11237 = ~n11104 & n11236 ;
  assign n11273 = n11272 ^ n11237 ;
  assign n12616 = n11273 ^ x89 ;
  assign n12652 = n12193 ^ n8891 ;
  assign n12653 = n12652 ^ n12438 ;
  assign n12630 = n12191 ^ n12141 ;
  assign n12633 = n12159 ^ n12050 ;
  assign n12634 = n12051 & n12633 ;
  assign n12635 = n12634 ^ n12050 ;
  assign n12636 = n12116 & n12635 ;
  assign n12631 = n12159 ^ n12143 ;
  assign n12637 = n12636 ^ n12631 ;
  assign n12640 = ~n12630 & ~n12637 ;
  assign n12641 = n12640 ^ n12191 ;
  assign n12617 = n12156 ^ n12133 ;
  assign n12644 = n12617 ^ n12049 ;
  assign n12642 = n12617 ^ n12192 ;
  assign n12643 = n12642 ^ n12637 ;
  assign n12645 = n12644 ^ n12643 ;
  assign n12646 = n12641 & ~n12645 ;
  assign n12647 = n12646 ^ n12644 ;
  assign n12648 = n12647 ^ n12449 ;
  assign n12618 = n12131 ^ n12123 ;
  assign n12619 = n12618 ^ n12162 ;
  assign n12620 = ~n12049 & n12619 ;
  assign n12621 = n12620 ^ n12123 ;
  assign n12649 = n12648 ^ n12621 ;
  assign n12623 = n12621 ^ n12439 ;
  assign n12622 = n12621 ^ n12617 ;
  assign n12624 = n12623 ^ n12622 ;
  assign n12627 = ~n12049 & n12624 ;
  assign n12628 = n12627 ^ n12623 ;
  assign n12629 = ~n12050 & n12628 ;
  assign n12650 = n12649 ^ n12629 ;
  assign n12651 = ~n12434 & n12650 ;
  assign n12654 = n12653 ^ n12651 ;
  assign n12655 = n12654 ^ x106 ;
  assign n12656 = n12616 & n12655 ;
  assign n12660 = n12226 ^ n9019 ;
  assign n12657 = n12226 ^ n12216 ;
  assign n12658 = n12657 ^ n12219 ;
  assign n12659 = ~n11562 & ~n12658 ;
  assign n12661 = n12660 ^ n12659 ;
  assign n12662 = n12661 ^ x107 ;
  assign n12689 = n11461 ^ n11421 ;
  assign n11443 = n11442 ^ n11410 ;
  assign n11444 = n11443 ^ n11388 ;
  assign n12673 = n11444 ^ n11417 ;
  assign n11432 = n11415 ^ n11380 ;
  assign n12680 = n12673 ^ n11432 ;
  assign n12674 = n11388 ^ n11277 ;
  assign n12675 = ~n12673 & ~n12674 ;
  assign n12679 = n11276 & n12675 ;
  assign n12681 = n12680 ^ n12679 ;
  assign n12690 = n12689 ^ n12681 ;
  assign n12685 = n11461 ^ n11414 ;
  assign n12686 = n12685 ^ n11421 ;
  assign n11447 = n11446 ^ n11420 ;
  assign n12687 = n12686 ^ n11447 ;
  assign n12688 = ~n11276 & ~n12687 ;
  assign n12691 = n12690 ^ n12688 ;
  assign n12692 = n11277 & ~n12691 ;
  assign n11404 = n11391 & n11403 ;
  assign n11395 = n11394 ^ n11381 ;
  assign n11396 = n11394 ^ n11276 ;
  assign n11397 = n11396 ^ n11394 ;
  assign n11398 = n11395 & n11397 ;
  assign n11399 = n11398 ^ n11394 ;
  assign n11400 = n11277 & n11399 ;
  assign n11405 = n11404 ^ n11400 ;
  assign n12676 = n12675 ^ n11405 ;
  assign n11851 = n11410 ^ n11381 ;
  assign n11852 = n11410 ^ n11276 ;
  assign n11853 = n11852 ^ n11410 ;
  assign n11854 = n11851 & ~n11853 ;
  assign n11855 = n11854 ^ n11410 ;
  assign n11856 = n11277 & n11855 ;
  assign n12677 = n12676 ^ n11856 ;
  assign n12678 = n12677 ^ n6858 ;
  assign n12682 = n12681 ^ n12678 ;
  assign n12667 = n11378 ^ n11276 ;
  assign n12668 = n12667 ^ n11378 ;
  assign n12669 = n11392 ^ n11378 ;
  assign n12670 = n12668 & n12669 ;
  assign n12671 = n12670 ^ n11378 ;
  assign n12672 = n11275 & n12671 ;
  assign n12683 = n12682 ^ n12672 ;
  assign n12664 = n12663 ^ n11417 ;
  assign n11827 = n11394 ^ n11387 ;
  assign n12665 = n12664 ^ n11827 ;
  assign n12666 = ~n11835 & ~n12665 ;
  assign n12684 = n12683 ^ n12666 ;
  assign n12693 = n12692 ^ n12684 ;
  assign n12694 = n12693 ^ x80 ;
  assign n12695 = n12662 & n12694 ;
  assign n12697 = n12695 ^ n12694 ;
  assign n12707 = n12697 ^ n12662 ;
  assign n12709 = n12656 & ~n12707 ;
  assign n12699 = n12656 ^ n12655 ;
  assign n12701 = n12699 ^ n12616 ;
  assign n12708 = ~n12701 & ~n12707 ;
  assign n12710 = n12709 ^ n12708 ;
  assign n12702 = n12697 & ~n12701 ;
  assign n12711 = n12710 ^ n12702 ;
  assign n12704 = n12655 ^ n12616 ;
  assign n12705 = ~n12662 & n12704 ;
  assign n12706 = n12705 ^ n12662 ;
  assign n12712 = n12711 ^ n12706 ;
  assign n12696 = n12656 & n12695 ;
  assign n12703 = n12702 ^ n12696 ;
  assign n12713 = n12712 ^ n12703 ;
  assign n12700 = n12697 & n12699 ;
  assign n12714 = n12713 ^ n12700 ;
  assign n13134 = n12714 ^ n12694 ;
  assign n13135 = ~n12796 & ~n13134 ;
  assign n12780 = n12705 ^ n12616 ;
  assign n12781 = ~n12694 & ~n12780 ;
  assign n12811 = n12796 ^ n12762 ;
  assign n13132 = n12781 & ~n12811 ;
  assign n12764 = n12656 ^ n12616 ;
  assign n12769 = ~n12707 & n12764 ;
  assign n12790 = n12769 ^ n12707 ;
  assign n12791 = n12790 ^ n12710 ;
  assign n12773 = n12695 & ~n12701 ;
  assign n12774 = n12773 ^ n12696 ;
  assign n12771 = n12695 & n12699 ;
  assign n12772 = n12771 ^ n12695 ;
  assign n12775 = n12774 ^ n12772 ;
  assign n12792 = n12791 ^ n12775 ;
  assign n12793 = n12792 ^ n12702 ;
  assign n12794 = ~n12789 & n12793 ;
  assign n13124 = n12794 ^ n12771 ;
  assign n13127 = n12762 ^ n12714 ;
  assign n13128 = n13127 ^ n12762 ;
  assign n13129 = n12789 & n13128 ;
  assign n13130 = n13129 ^ n12762 ;
  assign n13131 = ~n13124 & ~n13130 ;
  assign n13133 = n13132 ^ n13131 ;
  assign n13136 = n13135 ^ n13133 ;
  assign n13122 = n12774 ^ n12700 ;
  assign n13123 = ~n12811 & n13122 ;
  assign n13137 = n13136 ^ n13123 ;
  assign n13138 = n13137 ^ n12769 ;
  assign n12766 = n12695 ^ n12662 ;
  assign n12767 = n12699 & n12766 ;
  assign n12768 = n12767 ^ n12709 ;
  assign n12770 = n12769 ^ n12768 ;
  assign n12776 = n12775 ^ n12770 ;
  assign n12777 = n12776 ^ n12768 ;
  assign n12698 = n12697 ^ n12696 ;
  assign n12715 = n12714 ^ n12698 ;
  assign n12765 = n12764 ^ n12715 ;
  assign n12778 = n12777 ^ n12765 ;
  assign n13117 = n12769 ^ n12762 ;
  assign n13118 = n13117 ^ n12769 ;
  assign n13119 = ~n12778 & ~n13118 ;
  assign n13120 = n13119 ^ n12769 ;
  assign n13121 = n12615 & n13120 ;
  assign n13139 = n13138 ^ n13121 ;
  assign n13140 = n13139 ^ n12710 ;
  assign n12763 = n12762 ^ n12615 ;
  assign n12779 = n12778 ^ n12767 ;
  assign n13109 = n12779 ^ n12712 ;
  assign n13110 = ~n12615 & n13109 ;
  assign n13111 = n13110 ^ n12712 ;
  assign n12782 = n12781 ^ n12770 ;
  assign n12783 = n12782 ^ n12710 ;
  assign n12784 = n12783 ^ n12766 ;
  assign n12785 = n12784 ^ n12779 ;
  assign n13112 = n13111 ^ n12785 ;
  assign n13113 = ~n12763 & n13112 ;
  assign n13114 = n13113 ^ n12785 ;
  assign n13141 = n13140 ^ n13114 ;
  assign n13142 = n13141 ^ n10819 ;
  assign n13106 = ~n12762 & n12783 ;
  assign n13107 = n13106 ^ n12710 ;
  assign n13108 = ~n12763 & n13107 ;
  assign n13143 = n13142 ^ n13108 ;
  assign n13144 = n13143 ^ x118 ;
  assign n14958 = n13309 ^ n13144 ;
  assign n11556 = n10863 & n11037 ;
  assign n11543 = n11008 ^ n11001 ;
  assign n11544 = n11543 ^ n11021 ;
  assign n11545 = n11544 ^ n11017 ;
  assign n11537 = n11536 ^ n11000 ;
  assign n11538 = n11537 ^ n10860 ;
  assign n11539 = n11527 ^ n10860 ;
  assign n11540 = n11538 & n11539 ;
  assign n11541 = n11540 ^ n10860 ;
  assign n11542 = n10991 & ~n11541 ;
  assign n11546 = n11545 ^ n11542 ;
  assign n11552 = n11546 ^ n11004 ;
  assign n11548 = n11004 ^ n11000 ;
  assign n11549 = n11548 ^ n11051 ;
  assign n11038 = n11037 ^ n10989 ;
  assign n11039 = n11038 ^ n10993 ;
  assign n11040 = n11039 ^ n11025 ;
  assign n11550 = n11549 ^ n11040 ;
  assign n11551 = n10860 & n11550 ;
  assign n11553 = n11552 ^ n11551 ;
  assign n11554 = n10820 & ~n11553 ;
  assign n11547 = n11546 ^ n11025 ;
  assign n11555 = n11554 ^ n11547 ;
  assign n11557 = n11556 ^ n11555 ;
  assign n11530 = n11025 ^ n10860 ;
  assign n11531 = n11530 ^ n11025 ;
  assign n11532 = n11038 & ~n11531 ;
  assign n11533 = n11532 ^ n11025 ;
  assign n11534 = ~n11527 & n11533 ;
  assign n11558 = n11557 ^ n11534 ;
  assign n11559 = ~n11526 & n11558 ;
  assign n11560 = n11559 ^ n9184 ;
  assign n11561 = n11560 ^ x78 ;
  assign n9619 = n9592 ^ n9548 ;
  assign n9656 = n9655 ^ n9619 ;
  assign n9657 = n9656 ^ n9638 ;
  assign n9624 = n9623 ^ n9619 ;
  assign n9625 = n9624 ^ n9533 ;
  assign n9626 = n9625 ^ n9619 ;
  assign n9627 = n9619 ^ n9580 ;
  assign n9628 = n9627 ^ n9619 ;
  assign n9629 = n9626 & n9628 ;
  assign n9630 = n9629 ^ n9619 ;
  assign n9631 = n9618 & n9630 ;
  assign n9658 = n9657 ^ n9631 ;
  assign n9617 = n9608 & n9616 ;
  assign n9659 = n9658 ^ n9617 ;
  assign n9586 = n9550 ^ n9546 ;
  assign n9602 = n9601 ^ n9586 ;
  assign n9603 = n9601 ^ n9581 ;
  assign n9604 = n9603 ^ n9601 ;
  assign n9605 = n9602 & ~n9604 ;
  assign n9606 = n9605 ^ n9601 ;
  assign n9607 = ~n9580 & ~n9606 ;
  assign n9660 = n9659 ^ n9607 ;
  assign n9668 = n9660 & ~n9667 ;
  assign n9669 = ~n9585 & n9668 ;
  assign n9676 = n9669 & ~n9675 ;
  assign n9677 = n9676 ^ n8278 ;
  assign n9678 = n9677 ^ x84 ;
  assign n9876 = n9875 ^ x77 ;
  assign n9877 = ~n9678 & n9876 ;
  assign n9878 = n9877 ^ n9876 ;
  assign n9130 = n9068 & n9072 ;
  assign n9127 = n9126 ^ n9060 ;
  assign n9128 = n9069 & n9127 ;
  assign n9121 = n9120 ^ n8247 ;
  assign n9122 = n9121 ^ n9116 ;
  assign n9077 = n9053 ^ n9033 ;
  assign n9080 = n9079 ^ n9077 ;
  assign n9081 = n9080 ^ n9066 ;
  assign n9074 = n9073 ^ n9052 ;
  assign n9075 = n9074 ^ n9037 ;
  assign n9076 = n9070 & n9075 ;
  assign n9082 = n9081 ^ n9076 ;
  assign n9083 = n9082 ^ n9066 ;
  assign n9084 = n9083 ^ n9082 ;
  assign n9088 = n9084 & n9085 ;
  assign n9089 = n9088 ^ n9082 ;
  assign n9090 = n9067 & n9089 ;
  assign n9091 = n9090 ^ n9082 ;
  assign n9123 = n9122 ^ n9091 ;
  assign n9104 = n9100 ^ n9067 ;
  assign n9105 = n9104 ^ n9100 ;
  assign n9106 = ~n9101 & n9105 ;
  assign n9107 = n9106 ^ n9100 ;
  assign n9108 = ~n9066 & ~n9107 ;
  assign n9124 = n9123 ^ n9108 ;
  assign n9065 = n9064 ^ n9061 ;
  assign n9092 = n9071 & ~n9091 ;
  assign n9093 = ~n9065 & n9092 ;
  assign n9125 = n9124 ^ n9093 ;
  assign n9129 = n9128 ^ n9125 ;
  assign n9131 = n9130 ^ n9129 ;
  assign n9132 = n9131 ^ x70 ;
  assign n9424 = n9423 ^ x67 ;
  assign n9425 = ~n9132 & n9424 ;
  assign n9426 = n9425 ^ n9424 ;
  assign n9427 = n9426 ^ n9132 ;
  assign n9884 = n9427 ^ n9424 ;
  assign n9891 = n9878 & ~n9884 ;
  assign n9880 = n9877 ^ n9678 ;
  assign n9881 = n9427 & ~n9880 ;
  assign n9917 = n9891 ^ n9881 ;
  assign n9933 = n9917 ^ n9878 ;
  assign n9931 = n9425 & n9878 ;
  assign n9879 = n9427 & n9878 ;
  assign n9882 = n9881 ^ n9879 ;
  assign n9932 = n9931 ^ n9882 ;
  assign n9934 = n9933 ^ n9932 ;
  assign n9898 = n9426 & ~n9880 ;
  assign n9899 = n9898 ^ n9426 ;
  assign n9935 = n9934 ^ n9899 ;
  assign n9909 = n9425 & ~n9880 ;
  assign n11686 = n9935 ^ n9909 ;
  assign n8464 = n8463 ^ x102 ;
  assign n8854 = n8853 ^ x116 ;
  assign n9959 = ~n8464 & ~n8854 ;
  assign n9960 = n9959 ^ n8464 ;
  assign n9885 = ~n9880 & ~n9884 ;
  assign n9892 = n9885 ^ n9427 ;
  assign n9883 = n9427 & n9877 ;
  assign n9886 = n9885 ^ n9883 ;
  assign n9887 = n9886 ^ n9882 ;
  assign n9893 = n9892 ^ n9887 ;
  assign n9894 = n9893 ^ n9891 ;
  assign n9962 = n9894 & n9959 ;
  assign n9961 = n9934 & ~n9960 ;
  assign n9963 = n9962 ^ n9961 ;
  assign n11700 = n9931 ^ n8464 ;
  assign n9900 = n9426 & n9678 ;
  assign n9901 = n9900 ^ n9899 ;
  assign n9902 = n9901 ^ n9877 ;
  assign n9889 = ~n9876 & ~n9884 ;
  assign n9890 = n9889 ^ n9885 ;
  assign n9895 = n9894 ^ n9890 ;
  assign n9888 = n9887 ^ n9424 ;
  assign n9896 = n9895 ^ n9888 ;
  assign n9897 = n9896 ^ n9883 ;
  assign n9903 = n9902 ^ n9897 ;
  assign n11689 = n9903 ^ n9898 ;
  assign n11703 = n11689 ^ n9881 ;
  assign n9914 = n9880 ^ n9876 ;
  assign n9915 = n9425 & n9914 ;
  assign n9910 = n9909 ^ n9901 ;
  assign n11701 = n9915 ^ n9910 ;
  assign n11704 = n11703 ^ n11701 ;
  assign n11705 = n8854 & ~n11704 ;
  assign n11702 = n11701 ^ n9931 ;
  assign n11706 = n11705 ^ n11702 ;
  assign n11707 = n11700 & ~n11706 ;
  assign n11708 = n11707 ^ n8464 ;
  assign n11698 = n9959 ^ n8854 ;
  assign n11699 = n9887 & ~n11698 ;
  assign n11709 = n11708 ^ n11699 ;
  assign n11690 = n9934 ^ n9915 ;
  assign n11691 = n11690 ^ n11689 ;
  assign n11687 = n9897 ^ n9893 ;
  assign n11688 = n11687 ^ n9915 ;
  assign n11692 = n11691 ^ n11688 ;
  assign n11693 = n11688 ^ n8854 ;
  assign n11694 = n11693 ^ n11688 ;
  assign n11695 = n11692 & ~n11694 ;
  assign n11696 = n11695 ^ n11688 ;
  assign n11697 = ~n8464 & ~n11696 ;
  assign n11710 = n11709 ^ n11697 ;
  assign n11711 = n9959 ^ n9885 ;
  assign n11712 = n11711 ^ n11710 ;
  assign n11685 = n9960 ^ n8854 ;
  assign n11713 = n11685 ^ n9896 ;
  assign n11714 = ~n9959 & ~n11713 ;
  assign n11715 = n11714 ^ n9896 ;
  assign n11716 = n11712 & n11715 ;
  assign n11717 = n11716 ^ n9959 ;
  assign n11718 = ~n11710 & ~n11717 ;
  assign n11719 = ~n9963 & n11718 ;
  assign n11720 = ~n9960 & n11719 ;
  assign n11721 = n11686 & n11720 ;
  assign n11722 = n11721 ^ n11719 ;
  assign n11725 = n11722 ^ n9288 ;
  assign n9938 = n9890 ^ n9879 ;
  assign n11684 = n9938 ^ n9893 ;
  assign n11723 = ~n11685 & n11722 ;
  assign n11724 = n11684 & n11723 ;
  assign n11726 = n11725 ^ n11724 ;
  assign n11727 = n11726 ^ x75 ;
  assign n11758 = n10695 & n10745 ;
  assign n10739 = ~n10599 & n10600 ;
  assign n10740 = n10739 ^ n10600 ;
  assign n11755 = n10740 & ~n11754 ;
  assign n11751 = n10739 & ~n10767 ;
  assign n11744 = n10695 ^ n10600 ;
  assign n11745 = n11744 ^ n10695 ;
  assign n11748 = ~n10696 & ~n11745 ;
  assign n11749 = n11748 ^ n10695 ;
  assign n11750 = ~n10745 & n11749 ;
  assign n11752 = n11751 ^ n11750 ;
  assign n11729 = n10727 ^ n10600 ;
  assign n11730 = n11729 ^ n10727 ;
  assign n11731 = n10726 & ~n10768 ;
  assign n11732 = n11731 ^ n10727 ;
  assign n11733 = n11730 & ~n11732 ;
  assign n11734 = n11733 ^ n10727 ;
  assign n11735 = n10599 & ~n11734 ;
  assign n11736 = n11735 ^ n10726 ;
  assign n11739 = ~n10600 & ~n10724 ;
  assign n11740 = n11739 ^ n10706 ;
  assign n11741 = ~n10745 & ~n11740 ;
  assign n11742 = n11741 ^ n10706 ;
  assign n11743 = n11736 & n11742 ;
  assign n11753 = n11752 ^ n11743 ;
  assign n11756 = n11755 ^ n11753 ;
  assign n10741 = n10740 ^ n10599 ;
  assign n11728 = n10715 & n10741 ;
  assign n11757 = n11756 ^ n11728 ;
  assign n11759 = n11758 ^ n11757 ;
  assign n11760 = n10720 ^ n10718 ;
  assign n11761 = n10718 ^ n10599 ;
  assign n11762 = n11761 ^ n10718 ;
  assign n11763 = n11760 & n11762 ;
  assign n11764 = n11763 ^ n10718 ;
  assign n11765 = ~n10600 & n11764 ;
  assign n11766 = n11759 & ~n11765 ;
  assign n11774 = n11766 & ~n11773 ;
  assign n11775 = n11774 ^ n9215 ;
  assign n11776 = n11775 ^ x100 ;
  assign n11777 = n11727 & ~n11776 ;
  assign n11812 = n11811 ^ n9248 ;
  assign n11778 = ~n11222 & n11238 ;
  assign n11779 = n11778 ^ n11258 ;
  assign n11802 = n11209 ^ n11199 ;
  assign n11794 = n11212 ^ n11193 ;
  assign n11793 = n11254 ^ n11201 ;
  assign n11795 = n11794 ^ n11793 ;
  assign n11796 = n11103 & ~n11795 ;
  assign n11797 = n11796 ^ n11794 ;
  assign n11801 = n11797 ^ n11182 ;
  assign n11803 = n11802 ^ n11801 ;
  assign n11804 = n11803 ^ n11797 ;
  assign n11805 = ~n11103 & n11804 ;
  assign n11806 = n11805 ^ n11801 ;
  assign n11807 = n11102 & n11806 ;
  assign n11782 = n11204 ^ n11201 ;
  assign n11783 = n11782 ^ n11216 ;
  assign n11798 = n11797 ^ n11783 ;
  assign n11799 = n11798 ^ n11792 ;
  assign n11800 = n11799 ^ n11248 ;
  assign n11808 = n11807 ^ n11800 ;
  assign n11780 = n11256 ^ n11219 ;
  assign n11781 = n11780 ^ n11177 ;
  assign n11784 = n11783 ^ n11781 ;
  assign n11785 = n11241 & n11784 ;
  assign n11809 = n11808 ^ n11785 ;
  assign n11810 = ~n11779 & ~n11809 ;
  assign n11813 = n11812 ^ n11810 ;
  assign n11814 = n11813 ^ x117 ;
  assign n11408 = n11401 & ~n11407 ;
  assign n11840 = ~n11276 & n11414 ;
  assign n11836 = n11416 ^ n11391 ;
  assign n11837 = ~n11835 & ~n11836 ;
  assign n11830 = n11461 ^ n11417 ;
  assign n11817 = n11442 ^ n11378 ;
  assign n11818 = n11817 ^ n11384 ;
  assign n11821 = n11820 ^ n11818 ;
  assign n11822 = n11276 & n11821 ;
  assign n11823 = n11822 ^ n11820 ;
  assign n11831 = n11830 ^ n11823 ;
  assign n11826 = n11461 ^ n11415 ;
  assign n11828 = n11827 ^ n11826 ;
  assign n11829 = n11276 & ~n11828 ;
  assign n11832 = n11831 ^ n11829 ;
  assign n11833 = n11277 & ~n11832 ;
  assign n11434 = n11420 ^ n11377 ;
  assign n11435 = n11402 & n11434 ;
  assign n11824 = n11823 ^ n11435 ;
  assign n11825 = n11824 ^ n11400 ;
  assign n11834 = n11833 ^ n11825 ;
  assign n11838 = n11837 ^ n11834 ;
  assign n11815 = n11414 ^ n11380 ;
  assign n11816 = n11275 & n11815 ;
  assign n11839 = n11838 ^ n11816 ;
  assign n11841 = n11840 ^ n11839 ;
  assign n11842 = ~n11408 & ~n11841 ;
  assign n11850 = n11842 & ~n11849 ;
  assign n11857 = n11850 & ~n11856 ;
  assign n11858 = n11857 ^ n9321 ;
  assign n11859 = n11858 ^ x102 ;
  assign n11860 = n11814 & n11859 ;
  assign n11861 = n11860 ^ n11859 ;
  assign n11886 = n11861 ^ n11814 ;
  assign n11907 = n11777 & ~n11886 ;
  assign n11865 = n11777 ^ n11727 ;
  assign n11899 = n11860 & n11865 ;
  assign n11908 = n11907 ^ n11899 ;
  assign n11868 = n11777 ^ n11776 ;
  assign n11872 = n11860 & ~n11868 ;
  assign n11871 = n11861 & ~n11868 ;
  assign n11873 = n11872 ^ n11871 ;
  assign n11863 = n11860 ^ n11814 ;
  assign n11869 = n11863 & ~n11868 ;
  assign n11870 = n11869 ^ n11868 ;
  assign n11874 = n11873 ^ n11870 ;
  assign n11866 = n11865 ^ n11776 ;
  assign n11867 = n11861 & n11866 ;
  assign n11875 = n11874 ^ n11867 ;
  assign n11864 = n11777 & n11863 ;
  assign n11876 = n11875 ^ n11864 ;
  assign n11877 = n11876 ^ n11861 ;
  assign n11862 = ~n11777 & n11861 ;
  assign n11878 = n11877 ^ n11862 ;
  assign n11879 = n11878 ^ n11876 ;
  assign n11909 = n11908 ^ n11879 ;
  assign n11910 = n11909 ^ n11727 ;
  assign n11904 = n11863 & n11865 ;
  assign n11891 = n11863 & n11866 ;
  assign n11890 = n11872 ^ n11867 ;
  assign n11892 = n11891 ^ n11890 ;
  assign n11887 = n11866 & ~n11886 ;
  assign n11888 = n11887 ^ n11872 ;
  assign n11889 = n11888 ^ n11866 ;
  assign n11893 = n11892 ^ n11889 ;
  assign n11901 = n11893 ^ n11872 ;
  assign n11900 = n11899 ^ n11860 ;
  assign n11902 = n11901 ^ n11900 ;
  assign n11897 = n11871 ^ n11867 ;
  assign n11898 = n11897 ^ n11862 ;
  assign n11903 = n11902 ^ n11898 ;
  assign n11905 = n11904 ^ n11903 ;
  assign n11906 = n11905 ^ n11864 ;
  assign n11911 = n11910 ^ n11906 ;
  assign n13347 = n11911 ^ n11867 ;
  assign n11564 = n11563 ^ n11562 ;
  assign n11670 = n11669 ^ n11666 ;
  assign n11671 = n11670 ^ n11664 ;
  assign n11672 = ~n11563 & n11671 ;
  assign n11673 = n11672 ^ n11664 ;
  assign n11651 = n11650 ^ n11607 ;
  assign n11652 = n11651 ^ n11565 ;
  assign n11653 = n11652 ^ n11651 ;
  assign n11654 = n11651 ^ n11606 ;
  assign n11655 = n11654 ^ n11651 ;
  assign n11656 = ~n11653 & n11655 ;
  assign n11657 = n11656 ^ n11651 ;
  assign n11658 = n11563 & n11657 ;
  assign n11659 = n11658 ^ n11649 ;
  assign n11674 = n11673 ^ n11659 ;
  assign n11675 = ~n11564 & ~n11674 ;
  assign n11676 = n11675 ^ n11673 ;
  assign n11677 = n11676 ^ n9153 ;
  assign n11678 = n11677 ^ x124 ;
  assign n13333 = ~n11678 & n11899 ;
  assign n13348 = n13347 ^ n13333 ;
  assign n11931 = n11907 ^ n11904 ;
  assign n13344 = n11931 ^ n11867 ;
  assign n13345 = n13344 ^ n11879 ;
  assign n13346 = ~n11678 & n13345 ;
  assign n13349 = n13348 ^ n13346 ;
  assign n13350 = n11561 & n13349 ;
  assign n11679 = n11561 & ~n11678 ;
  assign n11680 = n11679 ^ n11678 ;
  assign n11681 = n11680 ^ n11561 ;
  assign n13340 = n11906 ^ n11875 ;
  assign n13341 = n11681 & n13340 ;
  assign n13335 = ~n11680 & n11864 ;
  assign n11894 = n11893 ^ n11869 ;
  assign n11895 = n11681 & n11894 ;
  assign n13336 = n13335 ^ n11895 ;
  assign n11682 = n11681 ^ n11678 ;
  assign n11942 = n11891 ^ n11874 ;
  assign n11943 = n11682 & ~n11942 ;
  assign n13330 = n11943 ^ n11903 ;
  assign n13322 = n11678 ^ n11561 ;
  assign n13323 = n11903 ^ n11678 ;
  assign n13324 = n13323 ^ n11903 ;
  assign n13325 = n11903 ^ n11888 ;
  assign n13326 = n13325 ^ n11903 ;
  assign n13327 = ~n13324 & n13326 ;
  assign n13328 = n13327 ^ n11903 ;
  assign n13329 = n13322 & n13328 ;
  assign n13331 = n13330 ^ n13329 ;
  assign n13332 = n13331 ^ n11894 ;
  assign n13334 = n13333 ^ n13332 ;
  assign n13337 = n13336 ^ n13334 ;
  assign n13338 = n13337 ^ n10944 ;
  assign n13315 = n11894 ^ n11678 ;
  assign n13316 = n13315 ^ n11894 ;
  assign n13319 = n11942 & ~n13316 ;
  assign n13320 = n13319 ^ n11894 ;
  assign n13321 = ~n11561 & ~n13320 ;
  assign n13339 = n13338 ^ n13321 ;
  assign n13342 = n13341 ^ n13339 ;
  assign n13313 = n11887 ^ n11871 ;
  assign n13314 = ~n11678 & n13313 ;
  assign n13343 = n13342 ^ n13314 ;
  assign n13351 = n13350 ^ n13343 ;
  assign n13352 = n13351 ^ x83 ;
  assign n11409 = ~n11405 & ~n11408 ;
  assign n11418 = n11417 ^ n11411 ;
  assign n11419 = n11418 ^ n11276 ;
  assign n11422 = n11421 ^ n11392 ;
  assign n11423 = n11422 ^ n11276 ;
  assign n11425 = n11424 ^ n11275 ;
  assign n11428 = ~n11422 & ~n11425 ;
  assign n11429 = n11428 ^ n11275 ;
  assign n11430 = n11423 & n11429 ;
  assign n11431 = n11430 ^ n11276 ;
  assign n11433 = n11432 ^ n11392 ;
  assign n11436 = n11435 ^ n11433 ;
  assign n11437 = ~n11431 & ~n11436 ;
  assign n11440 = ~n11419 & ~n11437 ;
  assign n11441 = n11440 ^ n11276 ;
  assign n11445 = n11444 ^ n11384 ;
  assign n11448 = n11447 ^ n11445 ;
  assign n11449 = n11448 ^ n11444 ;
  assign n11450 = n11444 ^ n11276 ;
  assign n11451 = n11450 ^ n11444 ;
  assign n11452 = n11449 & n11451 ;
  assign n11453 = n11452 ^ n11444 ;
  assign n11454 = ~n11275 & n11453 ;
  assign n11456 = n11454 ^ n11275 ;
  assign n11455 = n11454 ^ n11437 ;
  assign n11457 = n11456 ^ n11455 ;
  assign n11458 = ~n11441 & n11457 ;
  assign n11459 = n11458 ^ n11456 ;
  assign n11460 = n11459 ^ n11454 ;
  assign n11462 = ~n11277 & n11461 ;
  assign n11463 = ~n11460 & n11462 ;
  assign n11464 = n11463 ^ n11459 ;
  assign n11465 = n11409 & ~n11464 ;
  assign n11466 = n11465 ^ n8761 ;
  assign n11467 = n11466 ^ x122 ;
  assign n11274 = n11273 ^ x104 ;
  assign n10542 = n10541 ^ x82 ;
  assign n11054 = n11005 ^ n10820 ;
  assign n11055 = n11005 ^ n10860 ;
  assign n11056 = n11019 ^ n10860 ;
  assign n11057 = ~n11055 & ~n11056 ;
  assign n11058 = n11057 ^ n10860 ;
  assign n11059 = ~n11054 & n11058 ;
  assign n11052 = n10862 & n11051 ;
  assign n11043 = n11023 ^ n11017 ;
  assign n11044 = n10820 & n11043 ;
  assign n11041 = n10997 ^ n10993 ;
  assign n11042 = n11041 ^ n11040 ;
  assign n11045 = n11044 ^ n11042 ;
  assign n11047 = n11041 ^ n10860 ;
  assign n11046 = n11041 ^ n10820 ;
  assign n11048 = n11047 ^ n11046 ;
  assign n11049 = n11045 & n11048 ;
  assign n11050 = n11049 ^ n11046 ;
  assign n11053 = n11052 ^ n11050 ;
  assign n11060 = n11059 ^ n11053 ;
  assign n11061 = n11060 ^ n11001 ;
  assign n11032 = n11031 ^ n11001 ;
  assign n11033 = ~n10864 & n11032 ;
  assign n11062 = n11061 ^ n11033 ;
  assign n11063 = n11028 ^ n11002 ;
  assign n11064 = n10820 & ~n11063 ;
  assign n11065 = n11064 ^ n11002 ;
  assign n11066 = n11065 ^ n10860 ;
  assign n11067 = n11066 ^ n11065 ;
  assign n11068 = n10820 & n11008 ;
  assign n11069 = n11068 ^ n11065 ;
  assign n11070 = ~n11067 & n11069 ;
  assign n11071 = n11070 ^ n11065 ;
  assign n11072 = n11062 & ~n11071 ;
  assign n11073 = n11072 ^ n8691 ;
  assign n11074 = n11073 ^ x81 ;
  assign n9964 = n9963 ^ n8655 ;
  assign n9919 = n9909 ^ n9883 ;
  assign n9920 = n9919 ^ n9890 ;
  assign n9918 = n9917 ^ n9900 ;
  assign n9921 = n9920 ^ n9918 ;
  assign n9922 = n8464 & n9921 ;
  assign n9905 = n9896 ^ n9885 ;
  assign n9904 = n9903 ^ n9882 ;
  assign n9906 = n9905 ^ n9904 ;
  assign n9907 = ~n8464 & n9906 ;
  assign n9908 = n9907 ^ n9905 ;
  assign n9946 = n9922 ^ n9908 ;
  assign n9936 = n9935 ^ n9903 ;
  assign n9937 = n9936 ^ n9903 ;
  assign n9939 = n9938 ^ n9937 ;
  assign n9940 = n9939 ^ n9903 ;
  assign n9941 = n9903 ^ n8464 ;
  assign n9942 = n9941 ^ n9903 ;
  assign n9943 = ~n9940 & n9942 ;
  assign n9944 = n9943 ^ n9903 ;
  assign n9945 = n8854 & ~n9944 ;
  assign n9947 = n9946 ^ n9945 ;
  assign n8855 = n8854 ^ n8464 ;
  assign n9925 = n9910 ^ n9898 ;
  assign n9926 = n9898 ^ n8464 ;
  assign n9927 = n9926 ^ n9898 ;
  assign n9928 = n9925 & ~n9927 ;
  assign n9929 = n9928 ^ n9898 ;
  assign n9930 = ~n8855 & n9929 ;
  assign n9948 = n9947 ^ n9930 ;
  assign n9911 = n9910 ^ n9894 ;
  assign n9912 = ~n8464 & n9911 ;
  assign n9913 = n9912 ^ n9908 ;
  assign n9949 = n9948 ^ n9913 ;
  assign n9916 = n9915 ^ n9913 ;
  assign n9923 = n9922 ^ n9916 ;
  assign n9924 = ~n8855 & ~n9923 ;
  assign n9950 = n9949 ^ n9924 ;
  assign n9951 = n9882 ^ n8464 ;
  assign n9952 = n9951 ^ n9882 ;
  assign n9955 = n9932 & n9952 ;
  assign n9956 = n9955 ^ n9882 ;
  assign n9957 = n8855 & n9956 ;
  assign n9958 = ~n9950 & ~n9957 ;
  assign n9965 = n9964 ^ n9958 ;
  assign n9966 = n9965 ^ x72 ;
  assign n11469 = n11074 ^ n9966 ;
  assign n13354 = ~n10542 & n11469 ;
  assign n13371 = n13354 ^ n10542 ;
  assign n10728 = n10600 & ~n10727 ;
  assign n10729 = n10728 ^ n10691 ;
  assign n10731 = n10729 ^ n10718 ;
  assign n10730 = n10729 ^ n10703 ;
  assign n10732 = n10731 ^ n10730 ;
  assign n10735 = ~n10600 & n10732 ;
  assign n10736 = n10735 ^ n10731 ;
  assign n10737 = ~n10599 & n10736 ;
  assign n10738 = n10737 ^ n10729 ;
  assign n10759 = ~n10600 & ~n10689 ;
  assign n10751 = n10750 ^ n10703 ;
  assign n10752 = n10751 ^ n10623 ;
  assign n10753 = n10752 ^ n10703 ;
  assign n10754 = n10703 ^ n10600 ;
  assign n10755 = n10754 ^ n10703 ;
  assign n10756 = n10753 & n10755 ;
  assign n10757 = n10756 ^ n10703 ;
  assign n10758 = n10748 & ~n10757 ;
  assign n10760 = n10759 ^ n10758 ;
  assign n10761 = n10745 & ~n10760 ;
  assign n10762 = n10761 ^ n10759 ;
  assign n10742 = n10720 ^ n10695 ;
  assign n10743 = n10742 ^ n10710 ;
  assign n10744 = n10741 & ~n10743 ;
  assign n10763 = n10762 ^ n10744 ;
  assign n10764 = ~n10738 & ~n10763 ;
  assign n10765 = n10745 ^ n10714 ;
  assign n10771 = n10767 ^ n10747 ;
  assign n10770 = n10718 ^ n10689 ;
  assign n10772 = n10771 ^ n10770 ;
  assign n10775 = n10772 ^ n10714 ;
  assign n10769 = n10768 ^ n10726 ;
  assign n10773 = n10772 ^ n10769 ;
  assign n10774 = ~n10599 & ~n10773 ;
  assign n10776 = n10775 ^ n10774 ;
  assign n10777 = ~n10765 & ~n10776 ;
  assign n10778 = n10777 ^ n10714 ;
  assign n10779 = n10764 & ~n10778 ;
  assign n10780 = n10779 ^ n8725 ;
  assign n10781 = n10780 ^ x99 ;
  assign n11075 = n10781 & n11074 ;
  assign n11477 = n11075 ^ n10781 ;
  assign n11498 = n11477 ^ n9966 ;
  assign n11496 = ~n9966 & ~n10781 ;
  assign n11497 = n11496 ^ n11074 ;
  assign n11499 = n11498 ^ n11497 ;
  assign n11500 = ~n10542 & ~n11499 ;
  assign n13368 = n11500 ^ n11075 ;
  assign n11472 = n11074 ^ n10542 ;
  assign n11473 = n11472 ^ n10781 ;
  assign n11481 = n11075 & n11473 ;
  assign n13369 = n13368 ^ n11481 ;
  assign n11468 = n10781 ^ n9966 ;
  assign n13370 = n13369 ^ n11468 ;
  assign n13372 = n13371 ^ n13370 ;
  assign n11470 = n11469 ^ n10542 ;
  assign n11471 = n11470 ^ n10542 ;
  assign n11479 = n11472 ^ n9966 ;
  assign n11480 = n11473 ^ n11074 ;
  assign n11482 = n11481 ^ n11480 ;
  assign n11483 = n11479 & ~n11482 ;
  assign n11478 = n11477 ^ n11074 ;
  assign n11484 = n11483 ^ n11478 ;
  assign n11485 = n11484 ^ n11480 ;
  assign n11486 = n11485 ^ n11472 ;
  assign n11474 = n11074 & n11473 ;
  assign n11475 = n11474 ^ n11473 ;
  assign n10543 = n9966 & n10542 ;
  assign n11076 = n10543 & ~n11075 ;
  assign n11476 = n11475 ^ n11076 ;
  assign n11487 = n11486 ^ n11476 ;
  assign n11488 = n11487 ^ n9966 ;
  assign n11491 = ~n11471 & ~n11488 ;
  assign n11492 = n11491 ^ n10542 ;
  assign n11493 = n11468 & n11492 ;
  assign n11494 = n11493 ^ n11488 ;
  assign n13367 = n11494 ^ n11076 ;
  assign n13373 = n13372 ^ n13367 ;
  assign n13374 = ~n11274 & ~n13373 ;
  assign n13375 = n13374 ^ n13370 ;
  assign n13355 = n13354 ^ n11472 ;
  assign n11501 = n11500 ^ n11497 ;
  assign n13356 = n13355 ^ n11501 ;
  assign n13353 = n11468 ^ n11074 ;
  assign n13357 = n13356 ^ n13353 ;
  assign n13358 = n13357 ^ n11473 ;
  assign n13359 = n13358 ^ n10542 ;
  assign n13360 = n13359 ^ n11474 ;
  assign n13361 = n13360 ^ n13357 ;
  assign n13362 = ~n9966 & n13361 ;
  assign n13363 = n13362 ^ n13358 ;
  assign n13364 = n11274 & n13363 ;
  assign n13365 = n13364 ^ n13357 ;
  assign n13376 = n13375 ^ n13365 ;
  assign n13377 = ~n11467 & ~n13376 ;
  assign n13366 = n13365 ^ n11467 ;
  assign n13378 = n13377 ^ n13366 ;
  assign n13379 = n13378 ^ n10884 ;
  assign n13380 = n13379 ^ x70 ;
  assign n13381 = ~n13352 & n13380 ;
  assign n11969 = ~n8464 & ~n9936 ;
  assign n11970 = n11969 ^ n9903 ;
  assign n11971 = n8854 & ~n11970 ;
  assign n11961 = n9898 ^ n9889 ;
  assign n11953 = n9900 ^ n9888 ;
  assign n11948 = n9897 ^ n9888 ;
  assign n11949 = n9897 ^ n8464 ;
  assign n11950 = n8855 & ~n11949 ;
  assign n11951 = n11950 ^ n8464 ;
  assign n11952 = n11948 & ~n11951 ;
  assign n11954 = n11953 ^ n11952 ;
  assign n11965 = n11961 ^ n11954 ;
  assign n11962 = n11961 ^ n9931 ;
  assign n11963 = n11962 ^ n9920 ;
  assign n11964 = ~n8464 & n11963 ;
  assign n11966 = n11965 ^ n11964 ;
  assign n11967 = n8855 & ~n11966 ;
  assign n11957 = n11690 ^ n9897 ;
  assign n11958 = ~n11698 & ~n11957 ;
  assign n11947 = n9962 ^ n9930 ;
  assign n11955 = n11954 ^ n11947 ;
  assign n11956 = n11955 ^ n9957 ;
  assign n11959 = n11958 ^ n11956 ;
  assign n11960 = n11959 ^ n8363 ;
  assign n11968 = n11967 ^ n11960 ;
  assign n11972 = n11971 ^ n11968 ;
  assign n11973 = n11972 ^ x98 ;
  assign n11998 = n11997 ^ x120 ;
  assign n12200 = n12129 & n12191 ;
  assign n12197 = n12161 ^ n12143 ;
  assign n12198 = ~n12196 & ~n12197 ;
  assign n12170 = n12133 ^ n12054 ;
  assign n12171 = ~n12049 & n12170 ;
  assign n12172 = n12171 ^ n12155 ;
  assign n12188 = n12172 ^ n12166 ;
  assign n12182 = n12181 ^ n12133 ;
  assign n12183 = n12133 ^ n12049 ;
  assign n12184 = n12183 ^ n12133 ;
  assign n12185 = n12182 & ~n12184 ;
  assign n12186 = n12185 ^ n12133 ;
  assign n12187 = ~n12051 & n12186 ;
  assign n12189 = n12188 ^ n12187 ;
  assign n12173 = n12172 ^ n12133 ;
  assign n12174 = n12173 ^ n12151 ;
  assign n12175 = n12174 ^ n12173 ;
  assign n12178 = n12049 & n12175 ;
  assign n12179 = n12178 ^ n12173 ;
  assign n12180 = ~n12050 & n12179 ;
  assign n12190 = n12189 ^ n12180 ;
  assign n12194 = n12193 ^ n12190 ;
  assign n12195 = n12194 ^ n7429 ;
  assign n12199 = n12198 ^ n12195 ;
  assign n12201 = n12200 ^ n12199 ;
  assign n12157 = n12156 ^ n12117 ;
  assign n12167 = n12166 ^ n12157 ;
  assign n12118 = n12117 ^ n12115 ;
  assign n12124 = n12123 ^ n12118 ;
  assign n12125 = n12049 & n12124 ;
  assign n12168 = n12167 ^ n12125 ;
  assign n12169 = n12051 & ~n12168 ;
  assign n12202 = n12201 ^ n12169 ;
  assign n12203 = n12202 ^ x65 ;
  assign n12234 = n12233 ^ x96 ;
  assign n12299 = n12203 & ~n12234 ;
  assign n12339 = n12299 ^ n12203 ;
  assign n12046 = n12045 ^ n9463 ;
  assign n12008 = n11017 ^ n10989 ;
  assign n12009 = n12008 ^ n11025 ;
  assign n12007 = n11022 ^ n10997 ;
  assign n12010 = n12009 ^ n12007 ;
  assign n12011 = n12009 ^ n10860 ;
  assign n12012 = n12011 ^ n12009 ;
  assign n12013 = n12010 & n12012 ;
  assign n12014 = n12013 ^ n12009 ;
  assign n12015 = ~n10864 & n12014 ;
  assign n12023 = n12022 ^ n12015 ;
  assign n12004 = n10997 ^ n10989 ;
  assign n12001 = n11002 ^ n10989 ;
  assign n12002 = n12001 ^ n11535 ;
  assign n12003 = ~n10820 & n12002 ;
  assign n12005 = n12004 ^ n12003 ;
  assign n12006 = ~n10860 & n12005 ;
  assign n12024 = n12023 ^ n12006 ;
  assign n12025 = n10820 & ~n12024 ;
  assign n12026 = n11024 ^ n10860 ;
  assign n12027 = n12026 ^ n11024 ;
  assign n12030 = ~n11036 & ~n12027 ;
  assign n12031 = n12030 ^ n11024 ;
  assign n12032 = n12025 & n12031 ;
  assign n12033 = n12032 ^ n12024 ;
  assign n12034 = n11051 ^ n10863 ;
  assign n12035 = n11015 ^ n11013 ;
  assign n12036 = n12035 ^ n10861 ;
  assign n12039 = ~n11051 & ~n12036 ;
  assign n12040 = n12039 ^ n10861 ;
  assign n12041 = n12034 & n12040 ;
  assign n12042 = n12041 ^ n10863 ;
  assign n12043 = ~n12033 & ~n12042 ;
  assign n12047 = n12046 ^ n12043 ;
  assign n12048 = n12047 ^ x105 ;
  assign n12281 = n10417 ^ n10394 ;
  assign n12253 = n10411 ^ n10387 ;
  assign n12254 = n12253 ^ n10402 ;
  assign n12255 = n12254 ^ n12252 ;
  assign n12256 = n9991 & ~n12255 ;
  assign n12257 = n12256 ^ n10411 ;
  assign n12282 = n12281 ^ n12257 ;
  assign n12244 = n10509 ^ n9991 ;
  assign n12245 = n12244 ^ n10471 ;
  assign n12278 = n10423 ^ n10387 ;
  assign n12279 = ~n12245 & ~n12278 ;
  assign n12280 = n12279 ^ n10507 ;
  assign n12283 = n12282 ^ n12280 ;
  assign n12266 = n10420 ^ n10398 ;
  assign n12267 = ~n9991 & n12266 ;
  assign n12268 = n12267 ^ n10420 ;
  assign n12269 = n12268 ^ n10471 ;
  assign n12270 = n12269 ^ n12268 ;
  assign n12271 = n12268 ^ n10417 ;
  assign n12272 = n12271 ^ n10412 ;
  assign n12273 = n12272 ^ n12268 ;
  assign n12274 = n12270 & n12273 ;
  assign n12275 = n12274 ^ n12268 ;
  assign n12276 = ~n10529 & n12275 ;
  assign n12277 = n12276 ^ n12268 ;
  assign n12284 = n12283 ^ n12277 ;
  assign n12258 = n12257 ^ n10403 ;
  assign n12259 = n12258 ^ n10387 ;
  assign n12260 = n12259 ^ n12257 ;
  assign n12263 = n9991 & n12260 ;
  assign n12264 = n12263 ^ n12257 ;
  assign n12265 = ~n10471 & n12264 ;
  assign n12285 = n12284 ^ n12265 ;
  assign n12243 = n10508 ^ n10394 ;
  assign n12246 = n12245 ^ n10391 ;
  assign n12249 = ~n10508 & n12246 ;
  assign n12250 = n12249 ^ n10391 ;
  assign n12251 = n12243 & n12250 ;
  assign n12286 = n12285 ^ n12251 ;
  assign n12238 = n10417 ^ n9991 ;
  assign n12239 = n12238 ^ n10417 ;
  assign n12240 = n10520 & n12239 ;
  assign n12241 = n12240 ^ n10417 ;
  assign n12242 = n10471 & n12241 ;
  assign n12287 = n12286 ^ n12242 ;
  assign n12288 = ~n10494 & ~n12287 ;
  assign n12289 = n12288 ^ n9504 ;
  assign n12290 = n12289 ^ x115 ;
  assign n12300 = ~n12048 & ~n12290 ;
  assign n12306 = n12299 ^ n12234 ;
  assign n12320 = n12306 ^ n12203 ;
  assign n12321 = n12300 & n12320 ;
  assign n12331 = n12321 ^ n12300 ;
  assign n12301 = n12300 ^ n12290 ;
  assign n12302 = n12301 ^ n12048 ;
  assign n12315 = ~n12302 & ~n12306 ;
  assign n12307 = n12300 ^ n12048 ;
  assign n12308 = ~n12306 & ~n12307 ;
  assign n12303 = n12299 & ~n12302 ;
  assign n12311 = n12308 ^ n12303 ;
  assign n12310 = n12299 & n12300 ;
  assign n12312 = n12311 ^ n12310 ;
  assign n12313 = n12312 ^ n12299 ;
  assign n12305 = n12299 & ~n12301 ;
  assign n12309 = n12308 ^ n12305 ;
  assign n12314 = n12313 ^ n12309 ;
  assign n12316 = n12315 ^ n12314 ;
  assign n12204 = n12203 ^ n12048 ;
  assign n12295 = n12234 ^ n12048 ;
  assign n12296 = ~n12204 & ~n12295 ;
  assign n12297 = n12296 ^ n12234 ;
  assign n12298 = n12290 & ~n12297 ;
  assign n12304 = n12303 ^ n12298 ;
  assign n12317 = n12316 ^ n12304 ;
  assign n12325 = n12321 ^ n12317 ;
  assign n12291 = n12290 ^ n12234 ;
  assign n12292 = ~n12204 & n12291 ;
  assign n12322 = n12321 ^ n12292 ;
  assign n12323 = n12322 ^ n12311 ;
  assign n12324 = n12323 ^ n12321 ;
  assign n12326 = n12325 ^ n12324 ;
  assign n12319 = n12308 ^ n12296 ;
  assign n12327 = n12326 ^ n12319 ;
  assign n12330 = n12327 ^ n12310 ;
  assign n12332 = n12331 ^ n12330 ;
  assign n12340 = n12339 ^ n12332 ;
  assign n12341 = n12340 ^ n12326 ;
  assign n12342 = n12341 ^ n12327 ;
  assign n12235 = n12234 ^ n12204 ;
  assign n12293 = n12292 ^ n12235 ;
  assign n12336 = n12290 ^ n12203 ;
  assign n12337 = ~n12293 & ~n12336 ;
  assign n12338 = n12337 ^ n12321 ;
  assign n12343 = n12342 ^ n12338 ;
  assign n13415 = n12343 ^ n12323 ;
  assign n13416 = n13415 ^ n12310 ;
  assign n13417 = ~n11998 & n13416 ;
  assign n13403 = n12330 ^ n12308 ;
  assign n13418 = n13417 ^ n13403 ;
  assign n13419 = ~n11973 & n13418 ;
  assign n11999 = n11973 & n11998 ;
  assign n12359 = n11999 ^ n11998 ;
  assign n13411 = n12316 ^ n12298 ;
  assign n12377 = ~n12301 & ~n12306 ;
  assign n13412 = n13411 ^ n12377 ;
  assign n13413 = n12359 & n13412 ;
  assign n12378 = n12377 ^ n12314 ;
  assign n13397 = n12378 ^ n12321 ;
  assign n13398 = n12321 ^ n11998 ;
  assign n13399 = n13398 ^ n12321 ;
  assign n13400 = n13397 & ~n13399 ;
  assign n13401 = n13400 ^ n12321 ;
  assign n13402 = ~n11973 & n13401 ;
  assign n13404 = n13403 ^ n13402 ;
  assign n12344 = n12343 ^ n12317 ;
  assign n12345 = n12344 ^ n12341 ;
  assign n12346 = n12341 ^ n11998 ;
  assign n12347 = n12346 ^ n12341 ;
  assign n12348 = n12345 & n12347 ;
  assign n12349 = n12348 ^ n12341 ;
  assign n12350 = n11973 & n12349 ;
  assign n13405 = n13404 ^ n12350 ;
  assign n12351 = n11998 ^ n11973 ;
  assign n12364 = n12308 ^ n11973 ;
  assign n12365 = n12364 ^ n12308 ;
  assign n13392 = n12309 ^ n12308 ;
  assign n13393 = n13392 ^ n12308 ;
  assign n13394 = n12365 & n13393 ;
  assign n13395 = n13394 ^ n12308 ;
  assign n13396 = ~n12351 & n13395 ;
  assign n13406 = n13405 ^ n13396 ;
  assign n12397 = n12302 ^ n12298 ;
  assign n12398 = n12397 ^ n12314 ;
  assign n12399 = n12359 ^ n11973 ;
  assign n12400 = ~n12398 & ~n12399 ;
  assign n12390 = n12327 ^ n11998 ;
  assign n12391 = n12390 ^ n12327 ;
  assign n12394 = n12342 & ~n12391 ;
  assign n12395 = n12394 ^ n12327 ;
  assign n12396 = ~n11973 & n12395 ;
  assign n12401 = n12400 ^ n12396 ;
  assign n13407 = n13406 ^ n12401 ;
  assign n12318 = n12317 ^ n12305 ;
  assign n12328 = n12327 ^ n12318 ;
  assign n12294 = n12293 ^ n12234 ;
  assign n12329 = n12328 ^ n12294 ;
  assign n12333 = n12332 ^ n12329 ;
  assign n12375 = ~n12333 & n12359 ;
  assign n12369 = n12323 ^ n12315 ;
  assign n12370 = n12315 ^ n11973 ;
  assign n12371 = n12370 ^ n12315 ;
  assign n12372 = n12369 & ~n12371 ;
  assign n12373 = n12372 ^ n12315 ;
  assign n12374 = n12351 & n12373 ;
  assign n12376 = n12375 ^ n12374 ;
  assign n13408 = n13407 ^ n12376 ;
  assign n13409 = n13408 ^ n10981 ;
  assign n13385 = n12343 ^ n12324 ;
  assign n13384 = n12398 ^ n12332 ;
  assign n13386 = n13385 ^ n13384 ;
  assign n13387 = n13385 ^ n11998 ;
  assign n13388 = n13387 ^ n13385 ;
  assign n13389 = ~n13386 & n13388 ;
  assign n13390 = n13389 ^ n13385 ;
  assign n13391 = n11973 & n13390 ;
  assign n13410 = n13409 ^ n13391 ;
  assign n13414 = n13413 ^ n13410 ;
  assign n13420 = n13419 ^ n13414 ;
  assign n13421 = n13420 ^ x93 ;
  assign n12863 = n11270 ^ n7958 ;
  assign n12864 = n12863 ^ n11779 ;
  assign n12839 = n11782 ^ n11197 ;
  assign n12840 = n11238 & n12839 ;
  assign n12833 = n11196 ^ n11102 ;
  assign n12834 = n12833 ^ n11196 ;
  assign n12835 = n11253 & ~n12834 ;
  assign n12836 = n12835 ^ n11196 ;
  assign n12837 = ~n11104 & ~n12836 ;
  assign n12838 = n12837 ^ n11195 ;
  assign n12841 = n12840 ^ n12838 ;
  assign n12842 = n12841 ^ n11188 ;
  assign n12843 = n12842 ^ n12841 ;
  assign n12844 = n12843 ^ n11206 ;
  assign n12845 = n11206 ^ n11102 ;
  assign n12846 = n12845 ^ n11206 ;
  assign n12847 = n12844 & ~n12846 ;
  assign n12848 = n12847 ^ n11206 ;
  assign n12849 = ~n11104 & n12848 ;
  assign n12850 = n12849 ^ n12842 ;
  assign n12851 = n12850 ^ n11213 ;
  assign n12853 = n12851 ^ n12850 ;
  assign n12854 = n12850 ^ n11249 ;
  assign n12855 = n12854 ^ n12850 ;
  assign n12856 = n12850 ^ n12841 ;
  assign n12857 = n12856 ^ n12850 ;
  assign n12858 = n12855 & n12857 ;
  assign n12859 = n12853 & n12858 ;
  assign n12860 = n12859 ^ n12853 ;
  assign n12861 = n12860 ^ n12851 ;
  assign n12862 = ~n11251 & n12861 ;
  assign n12865 = n12864 ^ n12862 ;
  assign n12866 = n12865 ^ x90 ;
  assign n12885 = n11751 ^ n10767 ;
  assign n12886 = n12885 ^ n11765 ;
  assign n12882 = n10709 ^ n10701 ;
  assign n12883 = n12882 ^ n10768 ;
  assign n12884 = n10745 & ~n12883 ;
  assign n12887 = n12886 ^ n12884 ;
  assign n12881 = ~n10600 & ~n10709 ;
  assign n12888 = n12887 ^ n12881 ;
  assign n12874 = n10767 ^ n10600 ;
  assign n12875 = n12874 ^ n10767 ;
  assign n12876 = n10767 ^ n10714 ;
  assign n12877 = n12876 ^ n10767 ;
  assign n12878 = ~n12875 & n12877 ;
  assign n12879 = n12878 ^ n10767 ;
  assign n12880 = n10599 & ~n12879 ;
  assign n12889 = n12888 ^ n12880 ;
  assign n12867 = n10715 ^ n10600 ;
  assign n12868 = n12867 ^ n10715 ;
  assign n12869 = n10715 ^ n10707 ;
  assign n12870 = n12869 ^ n10715 ;
  assign n12871 = n12868 & n12870 ;
  assign n12872 = n12871 ^ n10715 ;
  assign n12873 = ~n10745 & n12872 ;
  assign n12890 = n12889 ^ n12873 ;
  assign n12891 = ~n10738 & n12890 ;
  assign n12892 = ~n11750 & n12891 ;
  assign n12893 = ~n11773 & n12892 ;
  assign n12894 = n12893 ^ n8200 ;
  assign n12895 = n12894 ^ x112 ;
  assign n12896 = ~n12866 & n12895 ;
  assign n12897 = n12896 ^ n12895 ;
  assign n12898 = n12897 ^ n12866 ;
  assign n12827 = n11972 ^ x73 ;
  assign n12828 = n12761 ^ x64 ;
  assign n12829 = ~n12827 & ~n12828 ;
  assign n12830 = n12829 ^ n12828 ;
  assign n12908 = n12830 ^ n12827 ;
  assign n12912 = n12898 & ~n12908 ;
  assign n12915 = n12202 ^ x114 ;
  assign n12916 = n12693 ^ x123 ;
  assign n12917 = n12915 & ~n12916 ;
  assign n12982 = n12912 & n12917 ;
  assign n12901 = n12829 ^ n12827 ;
  assign n12920 = n12897 & ~n12901 ;
  assign n12899 = n12898 ^ n12895 ;
  assign n12900 = ~n12830 & ~n12899 ;
  assign n12976 = n12920 ^ n12900 ;
  assign n12977 = n12920 ^ n12916 ;
  assign n12978 = n12977 ^ n12920 ;
  assign n12979 = n12976 & ~n12978 ;
  assign n12980 = n12979 ^ n12920 ;
  assign n12981 = n12915 & n12980 ;
  assign n12983 = n12982 ^ n12981 ;
  assign n12933 = ~n12899 & ~n12901 ;
  assign n12906 = n12829 & ~n12899 ;
  assign n12904 = n12829 & n12866 ;
  assign n12905 = n12904 ^ n12829 ;
  assign n12907 = n12906 ^ n12905 ;
  assign n12934 = n12933 ^ n12907 ;
  assign n13422 = n12917 & n12934 ;
  assign n12921 = ~n12830 & n12898 ;
  assign n12918 = n12917 ^ n12915 ;
  assign n12952 = n12918 ^ n12916 ;
  assign n12953 = n12952 ^ n12915 ;
  assign n12984 = n12921 & ~n12953 ;
  assign n13423 = n13422 ^ n12984 ;
  assign n13424 = ~n12983 & ~n13423 ;
  assign n13425 = n12918 & n12933 ;
  assign n12966 = n12906 & n12918 ;
  assign n13426 = n13425 ^ n12966 ;
  assign n12919 = n12916 ^ n12915 ;
  assign n12909 = n12896 & ~n12908 ;
  assign n12954 = n12909 ^ n12908 ;
  assign n12928 = n12897 & ~n12908 ;
  assign n12929 = n12928 ^ n12912 ;
  assign n12955 = n12954 ^ n12929 ;
  assign n12958 = n12928 ^ n12916 ;
  assign n12959 = n12958 ^ n12928 ;
  assign n12962 = ~n12955 & n12959 ;
  assign n12963 = n12962 ^ n12928 ;
  assign n12964 = n12919 & n12963 ;
  assign n12965 = n12964 ^ n12928 ;
  assign n12910 = n12909 ^ n12907 ;
  assign n12902 = n12896 & ~n12901 ;
  assign n12903 = n12902 ^ n12896 ;
  assign n12911 = n12910 ^ n12903 ;
  assign n13449 = n12911 & n12952 ;
  assign n12989 = n12933 & ~n12953 ;
  assign n13437 = n12989 ^ n12907 ;
  assign n12992 = n12898 & ~n12901 ;
  assign n12936 = n12928 ^ n12921 ;
  assign n12937 = n12936 ^ n12911 ;
  assign n12938 = n12937 ^ n12902 ;
  assign n12932 = n12920 ^ n12912 ;
  assign n12935 = n12934 ^ n12932 ;
  assign n12939 = n12938 ^ n12935 ;
  assign n12931 = n12901 ^ n12898 ;
  assign n12940 = n12939 ^ n12931 ;
  assign n12930 = n12929 ^ n12906 ;
  assign n12941 = n12940 ^ n12930 ;
  assign n12913 = n12912 ^ n12911 ;
  assign n12927 = n12913 ^ n12829 ;
  assign n12942 = n12941 ^ n12927 ;
  assign n12993 = n12992 ^ n12942 ;
  assign n13438 = n13437 ^ n12993 ;
  assign n13436 = n12920 & n12952 ;
  assign n13439 = n13438 ^ n13436 ;
  assign n12943 = n12942 ^ n12936 ;
  assign n13445 = n13439 ^ n12943 ;
  assign n13441 = n12955 ^ n12897 ;
  assign n13442 = n13441 ^ n12920 ;
  assign n12971 = n12942 ^ n12904 ;
  assign n13443 = n13442 ^ n12971 ;
  assign n13444 = n12916 & n13443 ;
  assign n13446 = n13445 ^ n13444 ;
  assign n13447 = n12915 & n13446 ;
  assign n13433 = n12909 ^ n12900 ;
  assign n13434 = n12952 & n13433 ;
  assign n13427 = n12913 ^ n12902 ;
  assign n13428 = n12915 ^ n12902 ;
  assign n13429 = n13428 ^ n12902 ;
  assign n13430 = n13427 & ~n13429 ;
  assign n13431 = n13430 ^ n12902 ;
  assign n13432 = ~n12916 & n13431 ;
  assign n13435 = n13434 ^ n13432 ;
  assign n13440 = n13439 ^ n13435 ;
  assign n13448 = n13447 ^ n13440 ;
  assign n13450 = n13449 ^ n13448 ;
  assign n13451 = ~n12965 & n13450 ;
  assign n13452 = ~n13426 & n13451 ;
  assign n13453 = n13424 & n13452 ;
  assign n13454 = n13453 ^ n10916 ;
  assign n13455 = n13454 ^ x100 ;
  assign n13456 = n13421 & n13455 ;
  assign n13457 = n13456 ^ n13421 ;
  assign n13486 = n13381 & n13457 ;
  assign n13458 = n13457 ^ n13455 ;
  assign n13382 = n13381 ^ n13380 ;
  assign n13383 = n13382 ^ n13352 ;
  assign n13466 = n13383 ^ n13380 ;
  assign n13467 = ~n13458 & ~n13466 ;
  assign n13461 = n13382 & ~n13421 ;
  assign n13462 = n13455 & n13461 ;
  assign n13483 = n13467 ^ n13462 ;
  assign n13481 = n13456 & ~n13466 ;
  assign n13484 = n13483 ^ n13481 ;
  assign n13487 = n13486 ^ n13484 ;
  assign n13473 = n13383 & n13456 ;
  assign n13475 = n13473 ^ n13383 ;
  assign n13465 = n13381 & ~n13458 ;
  assign n13468 = n13467 ^ n13465 ;
  assign n13463 = n13462 ^ n13461 ;
  assign n13464 = n13463 ^ n13458 ;
  assign n13469 = n13468 ^ n13464 ;
  assign n13459 = n13458 ^ n13421 ;
  assign n13460 = n13383 & n13459 ;
  assign n13470 = n13469 ^ n13460 ;
  assign n13476 = n13475 ^ n13470 ;
  assign n13488 = n13487 ^ n13476 ;
  assign n13472 = n13382 & n13457 ;
  assign n13489 = n13488 ^ n13472 ;
  assign n13485 = n13484 ^ n13457 ;
  assign n13490 = n13489 ^ n13485 ;
  assign n13491 = n13490 ^ n13486 ;
  assign n13479 = n13352 & n13421 ;
  assign n13474 = n13473 ^ n13472 ;
  assign n13477 = n13476 ^ n13474 ;
  assign n13480 = n13479 ^ n13477 ;
  assign n13482 = n13481 ^ n13480 ;
  assign n13492 = n13491 ^ n13482 ;
  assign n13478 = n13477 ^ n13421 ;
  assign n13493 = n13492 ^ n13478 ;
  assign n13494 = n13493 ^ n13490 ;
  assign n13495 = n13494 ^ n13486 ;
  assign n13496 = n13495 ^ n13465 ;
  assign n13497 = n13496 ^ n13381 ;
  assign n13498 = n13497 ^ n13490 ;
  assign n13527 = n13498 ^ n13468 ;
  assign n13528 = n13527 ^ n13490 ;
  assign n13526 = n13494 ^ n13481 ;
  assign n13529 = n13528 ^ n13526 ;
  assign n13525 = n13491 ^ n13352 ;
  assign n13530 = n13529 ^ n13525 ;
  assign n14990 = n13530 ^ n13476 ;
  assign n14991 = n13309 & ~n14990 ;
  assign n14992 = n14991 ^ n13476 ;
  assign n14993 = n14958 & ~n14992 ;
  assign n15406 = n14993 ^ n14992 ;
  assign n15407 = n15406 ^ n11073 ;
  assign n14982 = n13468 ^ n13463 ;
  assign n14983 = n14982 ^ n13458 ;
  assign n14984 = n14983 ^ n13463 ;
  assign n14985 = n13463 ^ n13144 ;
  assign n14986 = n14985 ^ n13463 ;
  assign n14987 = ~n14984 & ~n14986 ;
  assign n14988 = n14987 ^ n13463 ;
  assign n14989 = ~n13309 & n14988 ;
  assign n15382 = n13460 & n14958 ;
  assign n13499 = n13498 ^ n13472 ;
  assign n15395 = n13530 ^ n13499 ;
  assign n14960 = n13465 ^ n13462 ;
  assign n15396 = n15395 ^ n14960 ;
  assign n15392 = n13468 ^ n13460 ;
  assign n14974 = n13493 ^ n13477 ;
  assign n15393 = n15392 ^ n14974 ;
  assign n15394 = n15393 ^ n13499 ;
  assign n15397 = n15396 ^ n15394 ;
  assign n15398 = ~n13309 & n15397 ;
  assign n15399 = n15398 ^ n15394 ;
  assign n15400 = ~n14958 & ~n15399 ;
  assign n15401 = n15400 ^ n13499 ;
  assign n13310 = n13144 & n13309 ;
  assign n13311 = n13310 ^ n13309 ;
  assign n13312 = n13311 ^ n13144 ;
  assign n13534 = n13312 ^ n13309 ;
  assign n15391 = n13492 & n13534 ;
  assign n15402 = n15401 ^ n15391 ;
  assign n15384 = n13494 ^ n13480 ;
  assign n15383 = n13487 ^ n13463 ;
  assign n15385 = n15384 ^ n15383 ;
  assign n15386 = n15384 ^ n13309 ;
  assign n15387 = n15386 ^ n15384 ;
  assign n15388 = ~n15385 & n15387 ;
  assign n15389 = n15388 ^ n15384 ;
  assign n15390 = ~n13144 & ~n15389 ;
  assign n15403 = n15402 ^ n15390 ;
  assign n15404 = ~n15382 & n15403 ;
  assign n15405 = ~n14989 & n15404 ;
  assign n15408 = n15407 ^ n15405 ;
  assign n15409 = n15408 ^ x114 ;
  assign n13709 = n11726 ^ x85 ;
  assign n13710 = n10780 ^ x67 ;
  assign n13711 = n13709 & ~n13710 ;
  assign n13701 = n11677 ^ x86 ;
  assign n13667 = n12441 ^ n10284 ;
  assign n13642 = n12156 ^ n12141 ;
  assign n13640 = n12145 ^ n12114 ;
  assign n13641 = n13640 ^ n12439 ;
  assign n13643 = n13642 ^ n13641 ;
  assign n13644 = n12049 & ~n13643 ;
  assign n13645 = n13644 ^ n13642 ;
  assign n13654 = n13645 ^ n12436 ;
  assign n13655 = n13654 ^ n12187 ;
  assign n13646 = n13645 ^ n12154 ;
  assign n13647 = n13646 ^ n12131 ;
  assign n13648 = n13647 ^ n13645 ;
  assign n13651 = n12049 & n13648 ;
  assign n13652 = n13651 ^ n13645 ;
  assign n13653 = ~n12051 & n13652 ;
  assign n13656 = n13655 ^ n13653 ;
  assign n13661 = n12148 ^ n12127 ;
  assign n13662 = n12050 & ~n13661 ;
  assign n13657 = n12143 ^ n12128 ;
  assign n13658 = n13657 ^ n12439 ;
  assign n13659 = n12050 & n13658 ;
  assign n13660 = n13659 ^ n12117 ;
  assign n13663 = n13662 ^ n13660 ;
  assign n13664 = ~n12049 & n13663 ;
  assign n13665 = n13664 ^ n13659 ;
  assign n13666 = ~n13656 & ~n13665 ;
  assign n13668 = n13667 ^ n13666 ;
  assign n13635 = n12122 ^ n12049 ;
  assign n13636 = n13635 ^ n12122 ;
  assign n13637 = n12154 & n13636 ;
  assign n13638 = n13637 ^ n12122 ;
  assign n13639 = ~n12050 & n13638 ;
  assign n13669 = n13668 ^ n13639 ;
  assign n13670 = n13669 ^ x68 ;
  assign n13698 = n10471 & ~n10513 ;
  assign n13690 = n12279 ^ n12245 ;
  assign n13687 = n10428 ^ n10394 ;
  assign n13688 = ~n10509 & ~n13687 ;
  assign n13685 = n10520 ^ n10400 ;
  assign n13686 = ~n10471 & n13685 ;
  assign n13689 = n13688 ^ n13686 ;
  assign n13691 = n13690 ^ n13689 ;
  assign n13692 = n13691 ^ n12277 ;
  assign n13693 = n13692 ^ n10494 ;
  assign n13694 = n13693 ^ n10539 ;
  assign n13695 = n13694 ^ n10246 ;
  assign n13677 = n10471 ^ n10402 ;
  assign n13678 = n13677 ^ n12244 ;
  assign n13679 = n12244 ^ n10408 ;
  assign n13680 = n10408 ^ n10402 ;
  assign n13681 = n13680 ^ n10408 ;
  assign n13682 = n13679 & n13681 ;
  assign n13683 = n13682 ^ n10408 ;
  assign n13684 = ~n13678 & ~n13683 ;
  assign n13696 = n13695 ^ n13684 ;
  assign n13671 = n12252 ^ n10476 ;
  assign n13672 = n10476 ^ n10471 ;
  assign n13673 = n13672 ^ n10476 ;
  assign n13674 = n13671 & ~n13673 ;
  assign n13675 = n13674 ^ n10476 ;
  assign n13676 = ~n10529 & ~n13675 ;
  assign n13697 = n13696 ^ n13676 ;
  assign n13699 = n13698 ^ n13697 ;
  assign n13700 = n13699 ^ x116 ;
  assign n13727 = n13670 & n13700 ;
  assign n13730 = n13727 ^ n13670 ;
  assign n13731 = n13701 & n13730 ;
  assign n13716 = ~n13670 & n13701 ;
  assign n13729 = n13716 ^ n13701 ;
  assign n13732 = n13731 ^ n13729 ;
  assign n13736 = n13732 ^ n13727 ;
  assign n13702 = n11466 ^ x109 ;
  assign n13703 = n13701 & ~n13702 ;
  assign n13704 = n13703 ^ n13702 ;
  assign n13705 = n13704 ^ n13701 ;
  assign n13706 = n13700 & n13705 ;
  assign n13707 = ~n13670 & n13706 ;
  assign n13708 = n13707 ^ n13706 ;
  assign n13737 = n13736 ^ n13708 ;
  assign n13721 = ~n13670 & ~n13704 ;
  assign n13735 = n13721 ^ n13704 ;
  assign n13738 = n13737 ^ n13735 ;
  assign n13896 = n13711 & ~n13738 ;
  assign n13712 = n13711 ^ n13710 ;
  assign n13722 = n13700 & n13721 ;
  assign n13723 = n13722 ^ n13721 ;
  assign n13724 = ~n13712 & n13723 ;
  assign n13897 = n13896 ^ n13724 ;
  assign n13713 = n13712 ^ n13709 ;
  assign n13714 = n13713 ^ n13710 ;
  assign n13717 = n13702 & n13716 ;
  assign n13751 = ~n13700 & n13717 ;
  assign n13921 = n13751 ^ n13707 ;
  assign n13755 = n13706 ^ n13705 ;
  assign n13734 = n13731 ^ n13730 ;
  assign n13739 = n13738 ^ n13734 ;
  assign n13756 = n13755 ^ n13739 ;
  assign n13757 = n13756 ^ n13751 ;
  assign n13728 = n13703 & n13727 ;
  assign n13733 = n13732 ^ n13728 ;
  assign n13740 = n13739 ^ n13733 ;
  assign n13758 = n13757 ^ n13740 ;
  assign n13752 = n13751 ^ n13717 ;
  assign n13753 = n13752 ^ n13706 ;
  assign n13754 = n13753 ^ n13702 ;
  assign n13759 = n13758 ^ n13754 ;
  assign n13922 = n13921 ^ n13759 ;
  assign n13923 = n13714 & n13922 ;
  assign n13718 = n13717 ^ n13716 ;
  assign n13719 = n13700 & n13718 ;
  assign n13747 = n13719 ^ n13718 ;
  assign n13786 = n13756 ^ n13747 ;
  assign n13787 = n13756 ^ n13709 ;
  assign n13788 = n13787 ^ n13756 ;
  assign n13789 = ~n13786 & ~n13788 ;
  assign n13790 = n13789 ^ n13756 ;
  assign n13791 = n13710 & ~n13790 ;
  assign n13924 = n13923 ^ n13791 ;
  assign n13904 = n13712 ^ n13706 ;
  assign n13905 = n13904 ^ n13759 ;
  assign n13906 = n13737 ^ n13712 ;
  assign n13794 = n13738 ^ n13728 ;
  assign n13795 = n13794 ^ n13719 ;
  assign n13907 = n13906 ^ n13795 ;
  assign n13908 = ~n13905 & n13907 ;
  assign n13909 = n13908 ^ n13712 ;
  assign n13911 = n13756 ^ n13733 ;
  assign n13912 = n13911 ^ n13752 ;
  assign n13771 = n13759 ^ n13731 ;
  assign n13772 = n13771 ^ n13722 ;
  assign n13773 = n13772 ^ n13708 ;
  assign n13774 = n13773 ^ n13723 ;
  assign n13913 = n13912 ^ n13774 ;
  assign n13748 = n13747 ^ n13738 ;
  assign n13749 = n13748 ^ n13737 ;
  assign n13910 = n13749 ^ n13733 ;
  assign n13914 = n13913 ^ n13910 ;
  assign n13915 = n13910 ^ n13710 ;
  assign n13916 = n13915 ^ n13910 ;
  assign n13917 = n13914 & ~n13916 ;
  assign n13918 = n13917 ^ n13910 ;
  assign n13919 = n13709 & ~n13918 ;
  assign n13920 = n13909 & ~n13919 ;
  assign n13925 = n13924 ^ n13920 ;
  assign n13776 = n13737 ^ n13722 ;
  assign n13901 = n13776 ^ n13728 ;
  assign n13898 = n13771 ^ n13737 ;
  assign n13899 = n13898 ^ n13700 ;
  assign n13760 = n13759 ^ n13752 ;
  assign n13761 = n13760 ^ n13756 ;
  assign n13762 = n13761 ^ n13707 ;
  assign n13750 = n13749 ^ n13723 ;
  assign n13763 = n13762 ^ n13750 ;
  assign n13900 = n13899 ^ n13763 ;
  assign n13902 = n13901 ^ n13900 ;
  assign n13903 = n13713 & ~n13902 ;
  assign n13926 = n13925 ^ n13903 ;
  assign n13927 = ~n13897 & n13926 ;
  assign n13928 = n13927 ^ n10384 ;
  assign n13929 = n13928 ^ x97 ;
  assign n14046 = n11973 & n12315 ;
  assign n14031 = n12398 ^ n12311 ;
  assign n14032 = n14031 ^ n12378 ;
  assign n14033 = ~n11973 & ~n14032 ;
  assign n14043 = n14033 ^ n12396 ;
  assign n14036 = n12298 ^ n12235 ;
  assign n14034 = n12344 ^ n12330 ;
  assign n14035 = n14034 ^ n14033 ;
  assign n14037 = n14036 ^ n14035 ;
  assign n14038 = n14035 ^ n11973 ;
  assign n14039 = n14038 ^ n14035 ;
  assign n14040 = n14037 & n14039 ;
  assign n14041 = n14040 ^ n14035 ;
  assign n14042 = ~n11998 & n14041 ;
  assign n14044 = n14043 ^ n14042 ;
  assign n14028 = n12341 ^ n12324 ;
  assign n14029 = n14028 ^ n12317 ;
  assign n14030 = n11999 & n14029 ;
  assign n14045 = n14044 ^ n14030 ;
  assign n14047 = n14046 ^ n14045 ;
  assign n14048 = ~n13396 & ~n14047 ;
  assign n14026 = n12305 & ~n12399 ;
  assign n12363 = n12343 ^ n12308 ;
  assign n12366 = n12363 & ~n12365 ;
  assign n12367 = n12366 ^ n12308 ;
  assign n12368 = n11998 & n12367 ;
  assign n14027 = n14026 ^ n12368 ;
  assign n14049 = n14048 ^ n14027 ;
  assign n14050 = ~n12332 & n14049 ;
  assign n14051 = n14050 ^ n9990 ;
  assign n14052 = n14051 ^ x64 ;
  assign n11507 = n11474 ^ n10542 ;
  assign n11508 = n9966 & n11507 ;
  assign n11509 = n11508 ^ n11473 ;
  assign n14055 = n11509 ^ n11501 ;
  assign n14056 = ~n11274 & ~n14055 ;
  assign n14057 = n14056 ^ n11501 ;
  assign n14061 = n14057 ^ n10646 ;
  assign n14058 = n14057 ^ n13367 ;
  assign n11505 = n11486 ^ n9966 ;
  assign n10782 = n10543 & ~n10781 ;
  assign n11495 = n11494 ^ n10782 ;
  assign n14053 = n11505 ^ n11495 ;
  assign n14054 = ~n11274 & ~n14053 ;
  assign n14059 = n14058 ^ n14054 ;
  assign n14060 = n11467 & n14059 ;
  assign n14062 = n14061 ^ n14060 ;
  assign n14063 = n14062 ^ x120 ;
  assign n14064 = ~n14052 & ~n14063 ;
  assign n13985 = n11908 ^ n11864 ;
  assign n13986 = n13985 ^ n11911 ;
  assign n13987 = n11682 & n13986 ;
  assign n13973 = n11931 ^ n11862 ;
  assign n13976 = n13973 ^ n11901 ;
  assign n13977 = n13976 ^ n11903 ;
  assign n13978 = n13977 ^ n11911 ;
  assign n13979 = n13978 ^ n13973 ;
  assign n13980 = ~n11561 & n13979 ;
  assign n13981 = n13980 ^ n13976 ;
  assign n13982 = n11678 & n13981 ;
  assign n13983 = n13982 ^ n11891 ;
  assign n13974 = n13973 ^ n11891 ;
  assign n13975 = ~n11679 & n13974 ;
  assign n13984 = n13983 ^ n13975 ;
  assign n13988 = n13987 ^ n13984 ;
  assign n11932 = n11931 ^ n11903 ;
  assign n13966 = n13313 ^ n11932 ;
  assign n13967 = n13966 ^ n13313 ;
  assign n13968 = n13313 ^ n11678 ;
  assign n13969 = n13968 ^ n13313 ;
  assign n13970 = n13967 & ~n13969 ;
  assign n13971 = n13970 ^ n13313 ;
  assign n13972 = n13322 & n13971 ;
  assign n13989 = n13988 ^ n13972 ;
  assign n13965 = ~n11680 & n11888 ;
  assign n13990 = n13989 ^ n13965 ;
  assign n11683 = n11682 ^ n11680 ;
  assign n11880 = n11879 ^ n11869 ;
  assign n11881 = n11869 ^ n11561 ;
  assign n11882 = n11881 ^ n11869 ;
  assign n11883 = n11880 & ~n11882 ;
  assign n11884 = n11883 ^ n11869 ;
  assign n11885 = n11683 & n11884 ;
  assign n13991 = n13990 ^ n11885 ;
  assign n13992 = n13991 ^ n13336 ;
  assign n13993 = n13992 ^ n11943 ;
  assign n13994 = n13993 ^ n10676 ;
  assign n13995 = n13994 ^ x90 ;
  assign n12457 = n12456 ^ x101 ;
  assign n12458 = n11775 ^ x110 ;
  assign n12459 = ~n12457 & n12458 ;
  assign n12460 = n12459 ^ n12458 ;
  assign n12461 = n12460 ^ n12457 ;
  assign n12527 = n12526 ^ x92 ;
  assign n12485 = n9898 ^ n9896 ;
  assign n12486 = n12485 ^ n11684 ;
  assign n12487 = ~n8464 & ~n12486 ;
  assign n12479 = n9917 ^ n9909 ;
  assign n12488 = n12487 ^ n12479 ;
  assign n12489 = n8855 & n12488 ;
  assign n12480 = n12479 ^ n9945 ;
  assign n12481 = n12480 ^ n11970 ;
  assign n12482 = n12481 ^ n11958 ;
  assign n12483 = n12482 ^ n9799 ;
  assign n12470 = n9931 ^ n9886 ;
  assign n12471 = n12470 ^ n11690 ;
  assign n12472 = n12471 ^ n11970 ;
  assign n12469 = n9911 ^ n9903 ;
  assign n12473 = n12472 ^ n12469 ;
  assign n12474 = n12472 ^ n8464 ;
  assign n12475 = n12474 ^ n12472 ;
  assign n12476 = n12473 & n12475 ;
  assign n12477 = n12476 ^ n12472 ;
  assign n12478 = ~n8854 & ~n12477 ;
  assign n12484 = n12483 ^ n12478 ;
  assign n12490 = n12489 ^ n12484 ;
  assign n12491 = n12490 ^ x77 ;
  assign n12558 = n12527 ^ n12491 ;
  assign n12462 = n11560 ^ x70 ;
  assign n12559 = n12558 ^ n12462 ;
  assign n12463 = n11659 ^ n11562 ;
  assign n12464 = n12463 ^ n11675 ;
  assign n12465 = n12464 ^ n9722 ;
  assign n12466 = n12465 ^ x83 ;
  assign n12533 = n12527 ^ n12462 ;
  assign n12534 = n12466 & n12533 ;
  assign n12535 = n12534 ^ n12527 ;
  assign n12552 = n12491 ^ n12466 ;
  assign n12557 = n12535 & ~n12552 ;
  assign n12560 = n12559 ^ n12557 ;
  assign n12597 = n12560 ^ n12462 ;
  assign n12528 = ~n12491 & n12527 ;
  assign n12467 = n12462 & ~n12466 ;
  assign n12468 = n12467 ^ n12462 ;
  assign n12536 = n12468 ^ n12466 ;
  assign n12565 = n12528 & n12536 ;
  assign n12553 = ~n12462 & ~n12552 ;
  assign n12561 = n12558 ^ n12553 ;
  assign n12562 = n12561 ^ n12560 ;
  assign n12555 = n12552 ^ n12462 ;
  assign n12531 = n12528 ^ n12491 ;
  assign n12542 = n12467 & ~n12531 ;
  assign n12556 = n12555 ^ n12542 ;
  assign n12563 = n12562 ^ n12556 ;
  assign n12546 = n12467 ^ n12466 ;
  assign n12529 = n12528 ^ n12527 ;
  assign n12547 = n12529 ^ n12491 ;
  assign n12548 = ~n12546 & n12547 ;
  assign n12564 = n12563 ^ n12548 ;
  assign n12566 = n12565 ^ n12564 ;
  assign n12567 = n12566 ^ n12536 ;
  assign n12550 = ~n12531 & ~n12546 ;
  assign n12551 = n12550 ^ n12548 ;
  assign n12554 = n12553 ^ n12551 ;
  assign n12568 = n12567 ^ n12554 ;
  assign n12569 = n12568 ^ n12564 ;
  assign n12537 = n12529 & n12536 ;
  assign n12570 = n12569 ^ n12537 ;
  assign n12571 = n12570 ^ n12567 ;
  assign n12572 = n12571 ^ n12565 ;
  assign n12541 = n12467 & n12529 ;
  assign n12543 = n12542 ^ n12541 ;
  assign n12539 = n12467 & n12528 ;
  assign n12540 = n12539 ^ n12467 ;
  assign n12544 = n12543 ^ n12540 ;
  assign n12530 = n12468 & n12529 ;
  assign n12545 = n12544 ^ n12530 ;
  assign n12549 = n12548 ^ n12545 ;
  assign n12573 = n12572 ^ n12549 ;
  assign n12598 = n12597 ^ n12573 ;
  assign n13996 = n12461 & ~n12598 ;
  assign n12580 = n12565 ^ n12550 ;
  assign n12608 = n12580 ^ n12462 ;
  assign n12609 = n12608 ^ n12567 ;
  assign n12610 = n12609 ^ n12571 ;
  assign n12611 = n12461 & ~n12610 ;
  assign n12538 = n12537 ^ n12535 ;
  assign n12574 = n12573 ^ n12538 ;
  assign n12532 = n12531 ^ n12530 ;
  assign n12575 = n12574 ^ n12532 ;
  assign n12599 = n12598 ^ n12575 ;
  assign n12596 = n12530 ^ n12468 ;
  assign n12600 = n12599 ^ n12596 ;
  assign n12601 = n12600 ^ n12566 ;
  assign n12602 = n12566 ^ n12458 ;
  assign n12603 = n12602 ^ n12566 ;
  assign n12604 = ~n12601 & ~n12603 ;
  assign n12605 = n12604 ^ n12566 ;
  assign n12606 = n12457 & ~n12605 ;
  assign n14009 = n12539 ^ n12537 ;
  assign n14010 = n12458 & n14009 ;
  assign n14011 = n14010 ^ n12539 ;
  assign n14005 = ~n12458 & ~n12562 ;
  assign n14006 = n14005 ^ n12560 ;
  assign n14012 = n14011 ^ n14006 ;
  assign n14013 = n14012 ^ n14006 ;
  assign n14008 = n12575 ^ n12541 ;
  assign n14014 = n14013 ^ n14008 ;
  assign n14001 = n12542 ^ n12539 ;
  assign n14002 = n14001 ^ n12600 ;
  assign n14003 = n12458 & n14002 ;
  assign n14004 = n14003 ^ n12542 ;
  assign n14007 = n14006 ^ n14004 ;
  assign n14015 = n14014 ^ n14007 ;
  assign n13997 = n12563 ^ n12541 ;
  assign n13998 = n13997 ^ n12544 ;
  assign n13999 = n13998 ^ n12575 ;
  assign n14000 = ~n12458 & n13999 ;
  assign n14016 = n14015 ^ n14000 ;
  assign n14017 = n12457 & n14016 ;
  assign n14018 = n14017 ^ n14006 ;
  assign n14019 = ~n12606 & n14018 ;
  assign n14020 = ~n12611 & n14019 ;
  assign n14021 = ~n13996 & n14020 ;
  assign n14022 = n14021 ^ n10622 ;
  assign n14023 = n14022 ^ x73 ;
  assign n14024 = ~n13995 & ~n14023 ;
  assign n14069 = n14024 ^ n14023 ;
  assign n14085 = n14069 ^ n13995 ;
  assign n14086 = n14064 & ~n14085 ;
  assign n14073 = n14024 & n14064 ;
  assign n14087 = n14086 ^ n14073 ;
  assign n14025 = n14024 ^ n13995 ;
  assign n14083 = ~n14025 & n14064 ;
  assign n14084 = n14083 ^ n14064 ;
  assign n14088 = n14087 ^ n14084 ;
  assign n14065 = n14064 ^ n14063 ;
  assign n14066 = n14065 ^ n14052 ;
  assign n14071 = n14066 ^ n14063 ;
  assign n14080 = n14024 & ~n14071 ;
  assign n14108 = n14088 ^ n14080 ;
  assign n14109 = n14108 ^ n14083 ;
  assign n14072 = ~n14025 & ~n14071 ;
  assign n14074 = n14073 ^ n14072 ;
  assign n14110 = n14109 ^ n14074 ;
  assign n14091 = ~n14069 & ~n14071 ;
  assign n14104 = n14091 ^ n14086 ;
  assign n14107 = n14104 ^ n14052 ;
  assign n14111 = n14110 ^ n14107 ;
  assign n14093 = ~n14066 & ~n14085 ;
  assign n14115 = n14111 ^ n14093 ;
  assign n13930 = ~n12966 & ~n13423 ;
  assign n13931 = n12917 & n12928 ;
  assign n13932 = n13931 ^ n12989 ;
  assign n12956 = ~n12953 & ~n12955 ;
  assign n12922 = n12921 ^ n12920 ;
  assign n12944 = n12922 ^ n12897 ;
  assign n12945 = n12944 ^ n12943 ;
  assign n12948 = ~n12916 & ~n12945 ;
  assign n12923 = ~n12916 & n12922 ;
  assign n12924 = n12923 ^ n12921 ;
  assign n12949 = n12948 ^ n12924 ;
  assign n12950 = ~n12919 & n12949 ;
  assign n12951 = n12950 ^ n12924 ;
  assign n12957 = n12956 ^ n12951 ;
  assign n13950 = n12918 & n12992 ;
  assign n12994 = n12993 ^ n12906 ;
  assign n13942 = n12994 ^ n12928 ;
  assign n13939 = n12971 ^ n12945 ;
  assign n13940 = n13939 ^ n12909 ;
  assign n13943 = n13942 ^ n13940 ;
  assign n13944 = n12916 & ~n13943 ;
  assign n13941 = n13940 ^ n12907 ;
  assign n13945 = n13944 ^ n13941 ;
  assign n13946 = n12919 & n13945 ;
  assign n13937 = n13434 ^ n12907 ;
  assign n13938 = n13937 ^ n12981 ;
  assign n13947 = n13946 ^ n13938 ;
  assign n13934 = n12955 ^ n12921 ;
  assign n13935 = n13934 ^ n12913 ;
  assign n13936 = n12918 & ~n13935 ;
  assign n13948 = n13947 ^ n13936 ;
  assign n13933 = n12932 & ~n12953 ;
  assign n13949 = n13948 ^ n13933 ;
  assign n13951 = n13950 ^ n13949 ;
  assign n13952 = n12906 ^ n12902 ;
  assign n13955 = n12916 & n13952 ;
  assign n13956 = n13955 ^ n12906 ;
  assign n13957 = ~n12915 & n13956 ;
  assign n13958 = ~n13951 & ~n13957 ;
  assign n13959 = ~n12957 & n13958 ;
  assign n13960 = ~n13932 & n13959 ;
  assign n13961 = n13930 & n13960 ;
  assign n13962 = n13961 ^ n10598 ;
  assign n13963 = n13962 ^ x123 ;
  assign n14766 = n14111 ^ n13963 ;
  assign n14767 = n14766 ^ n14111 ;
  assign n14768 = ~n14115 & n14767 ;
  assign n14769 = n14768 ^ n14111 ;
  assign n14770 = ~n13929 & ~n14769 ;
  assign n13964 = n13963 ^ n13929 ;
  assign n14070 = ~n14065 & ~n14069 ;
  assign n14089 = n14088 ^ n14070 ;
  assign n14090 = n14089 ^ n14069 ;
  assign n14092 = n14091 ^ n14090 ;
  assign n14094 = n14093 ^ n14092 ;
  assign n14067 = ~n14025 & ~n14066 ;
  assign n14082 = n14067 ^ n14066 ;
  assign n14095 = n14094 ^ n14082 ;
  assign n14096 = n14095 ^ n14073 ;
  assign n15187 = n14096 ^ n14083 ;
  assign n14081 = n14080 ^ n14024 ;
  assign n14097 = n14096 ^ n14081 ;
  assign n14754 = n14097 ^ n14092 ;
  assign n14114 = n14086 ^ n14085 ;
  assign n14116 = n14115 ^ n14114 ;
  assign n14755 = n14754 ^ n14116 ;
  assign n14756 = n14755 ^ n14094 ;
  assign n15188 = n15187 ^ n14756 ;
  assign n15189 = ~n13929 & n15188 ;
  assign n15183 = n14087 ^ n14070 ;
  assign n15184 = n15183 ^ n14091 ;
  assign n15185 = n15184 ^ n14080 ;
  assign n15186 = n15185 ^ n14756 ;
  assign n15190 = n15189 ^ n15186 ;
  assign n15191 = n13964 & n15190 ;
  assign n15181 = ~n13963 & n14083 ;
  assign n15175 = n14754 ^ n14088 ;
  assign n14117 = n14116 ^ n14097 ;
  assign n14113 = n14070 ^ n14065 ;
  assign n14118 = n14117 ^ n14113 ;
  assign n14119 = n14118 ^ n14092 ;
  assign n15173 = n14119 ^ n14095 ;
  assign n15176 = n15175 ^ n15173 ;
  assign n15177 = n13929 & ~n15176 ;
  assign n15174 = n15173 ^ n14067 ;
  assign n15178 = n15177 ^ n15174 ;
  assign n15179 = ~n13964 & n15178 ;
  assign n14733 = n13929 & n13963 ;
  assign n15169 = n14111 ^ n14072 ;
  assign n15170 = n14733 & ~n15169 ;
  assign n15171 = n15170 ^ n14087 ;
  assign n14122 = n14116 ^ n14072 ;
  assign n14123 = n14072 ^ n13929 ;
  assign n14124 = n14123 ^ n14072 ;
  assign n14125 = n14122 & ~n14124 ;
  assign n14126 = n14125 ^ n14072 ;
  assign n14127 = n13964 & n14126 ;
  assign n15172 = n15171 ^ n14127 ;
  assign n15180 = n15179 ^ n15172 ;
  assign n15182 = n15181 ^ n15180 ;
  assign n15192 = n15191 ^ n15182 ;
  assign n15193 = ~n14770 & ~n15192 ;
  assign n15194 = n15193 ^ n10780 ;
  assign n15195 = n15194 ^ x96 ;
  assign n15196 = n14051 ^ x107 ;
  assign n11912 = n11911 ^ n11890 ;
  assign n11913 = n11890 ^ n11561 ;
  assign n11914 = n11913 ^ n11890 ;
  assign n11915 = n11912 & ~n11914 ;
  assign n11916 = n11915 ^ n11890 ;
  assign n11917 = n11683 & n11916 ;
  assign n14203 = n11890 ^ n11869 ;
  assign n14204 = n11681 & n14203 ;
  assign n14199 = n11887 ^ n11869 ;
  assign n14200 = n11682 & n14199 ;
  assign n14191 = n11875 ^ n11871 ;
  assign n14192 = n14191 ^ n11878 ;
  assign n14193 = n14192 ^ n11907 ;
  assign n14194 = n11561 & n14193 ;
  assign n14190 = n11909 ^ n11898 ;
  assign n14195 = n14194 ^ n14190 ;
  assign n14196 = n14195 ^ n11893 ;
  assign n14197 = n14196 ^ n11874 ;
  assign n14201 = n14200 ^ n14197 ;
  assign n14187 = n11911 ^ n11871 ;
  assign n14188 = n14187 ^ n11902 ;
  assign n14189 = n14188 ^ n11904 ;
  assign n14198 = n14197 ^ n14189 ;
  assign n14202 = n14201 ^ n14198 ;
  assign n14205 = n14204 ^ n14202 ;
  assign n14206 = n11942 ^ n11931 ;
  assign n14207 = n11942 ^ n11561 ;
  assign n14208 = n14207 ^ n11942 ;
  assign n14209 = ~n14206 & ~n14208 ;
  assign n14210 = n14209 ^ n11942 ;
  assign n14211 = ~n14205 & n14210 ;
  assign n14212 = n14211 ^ n14201 ;
  assign n14213 = n11683 & n14212 ;
  assign n14214 = n14213 ^ n14201 ;
  assign n14215 = ~n13965 & n14214 ;
  assign n14216 = ~n11917 & n14215 ;
  assign n14217 = n14216 ^ n10470 ;
  assign n15197 = n14217 ^ x98 ;
  assign n15198 = n15196 & n15197 ;
  assign n15199 = n15198 ^ n15196 ;
  assign n12812 = n12778 ^ n12708 ;
  assign n12813 = ~n12811 & ~n12812 ;
  assign n15239 = n12783 ^ n12771 ;
  assign n15237 = n12774 ^ n12709 ;
  assign n15240 = n15239 ^ n15237 ;
  assign n15241 = n12615 & n15240 ;
  assign n12716 = n12715 ^ n12700 ;
  assign n15236 = n12770 ^ n12716 ;
  assign n15238 = n15237 ^ n15236 ;
  assign n15242 = n15241 ^ n15238 ;
  assign n15243 = ~n12763 & ~n15242 ;
  assign n15244 = n15243 ^ n12770 ;
  assign n15235 = ~n12615 & ~n12791 ;
  assign n15245 = n15244 ^ n15235 ;
  assign n13125 = n12789 ^ n12762 ;
  assign n15233 = n12775 ^ n12700 ;
  assign n15234 = ~n13125 & n15233 ;
  assign n15246 = n15245 ^ n15234 ;
  assign n15232 = n12703 & n12763 ;
  assign n15247 = n15246 ^ n15232 ;
  assign n15248 = n12785 ^ n12615 ;
  assign n15249 = n15248 ^ n12785 ;
  assign n13567 = n12775 ^ n12773 ;
  assign n15250 = n12762 & n13567 ;
  assign n15251 = n15250 ^ n12785 ;
  assign n15252 = ~n15249 & ~n15251 ;
  assign n15253 = n15252 ^ n12785 ;
  assign n15254 = ~n15247 & ~n15253 ;
  assign n15255 = n15254 ^ n15247 ;
  assign n15256 = ~n12813 & ~n15255 ;
  assign n15258 = ~n12763 & ~n13111 ;
  assign n15259 = n15256 & n15258 ;
  assign n15257 = n15256 ^ n10056 ;
  assign n15260 = n15259 ^ n15257 ;
  assign n15261 = n15260 ^ x96 ;
  assign n14283 = n13302 ^ n13221 ;
  assign n14280 = n13260 ^ n13235 ;
  assign n14281 = ~n13146 & ~n14280 ;
  assign n14282 = n14281 ^ n13235 ;
  assign n14284 = n14283 ^ n14282 ;
  assign n14285 = n14284 ^ n13240 ;
  assign n14286 = n14285 ^ n13221 ;
  assign n14287 = n14286 ^ n14284 ;
  assign n14290 = n13146 & n14287 ;
  assign n14291 = n14290 ^ n14284 ;
  assign n14292 = n13145 & n14291 ;
  assign n14293 = n14292 ^ n14282 ;
  assign n13615 = n13237 ^ n13145 ;
  assign n13616 = n13615 ^ n13237 ;
  assign n13619 = n13247 & ~n13616 ;
  assign n13620 = n13619 ^ n13237 ;
  assign n13621 = ~n13257 & n13620 ;
  assign n14306 = n14293 ^ n13621 ;
  assign n14301 = n13246 ^ n13146 ;
  assign n14302 = n14301 ^ n13246 ;
  assign n14303 = n13299 & ~n14302 ;
  assign n14304 = n14303 ^ n13246 ;
  assign n14305 = n13257 & n14304 ;
  assign n14307 = n14306 ^ n14305 ;
  assign n13608 = n13298 ^ n13253 ;
  assign n14278 = n13608 ^ n13145 ;
  assign n14279 = n14278 ^ n13608 ;
  assign n14294 = n13222 & n14293 ;
  assign n14295 = n14294 ^ n13608 ;
  assign n14296 = n14279 & n14295 ;
  assign n14297 = n14296 ^ n13608 ;
  assign n14298 = n13146 & n14297 ;
  assign n14308 = n14307 ^ n14298 ;
  assign n14309 = n14308 ^ n13294 ;
  assign n14310 = n14309 ^ n10204 ;
  assign n15262 = n14310 ^ x122 ;
  assign n15263 = n15261 & ~n15262 ;
  assign n15264 = n15263 ^ n15261 ;
  assign n15265 = n15264 ^ n15262 ;
  assign n15266 = n15265 ^ n15261 ;
  assign n15200 = n13928 ^ x113 ;
  assign n12576 = n12461 & ~n12575 ;
  assign n15219 = n12459 ^ n12457 ;
  assign n14401 = n12609 ^ n12568 ;
  assign n15220 = n14401 ^ n12580 ;
  assign n14392 = n12600 ^ n12541 ;
  assign n15215 = n14392 ^ n12542 ;
  assign n15221 = n15220 ^ n15215 ;
  assign n15222 = ~n15219 & ~n15221 ;
  assign n15216 = n15215 ^ n12598 ;
  assign n15217 = n12460 & ~n15216 ;
  assign n15210 = n12564 ^ n12545 ;
  assign n15211 = n15210 ^ n12599 ;
  assign n15212 = n12459 & ~n15211 ;
  assign n15209 = n12458 & ~n12571 ;
  assign n15213 = n15212 ^ n15209 ;
  assign n15202 = n12568 ^ n12563 ;
  assign n15203 = n15202 ^ n12573 ;
  assign n15204 = n12573 ^ n12458 ;
  assign n15205 = n15204 ^ n12573 ;
  assign n15206 = ~n15203 & n15205 ;
  assign n15207 = n15206 ^ n12573 ;
  assign n15208 = n12457 & ~n15207 ;
  assign n15214 = n15213 ^ n15208 ;
  assign n15218 = n15217 ^ n15214 ;
  assign n15223 = n15222 ^ n15218 ;
  assign n14384 = n14010 ^ n12537 ;
  assign n15224 = n15223 ^ n14384 ;
  assign n15225 = n15224 ^ n13996 ;
  assign n15201 = n12457 & n14009 ;
  assign n15226 = n15225 ^ n15201 ;
  assign n15227 = ~n12576 & ~n15226 ;
  assign n15228 = n15227 ^ n10028 ;
  assign n15229 = n15228 ^ x74 ;
  assign n15230 = ~n15200 & ~n15229 ;
  assign n15273 = n15230 ^ n15200 ;
  assign n15282 = ~n15266 & ~n15273 ;
  assign n15279 = n15230 & n15264 ;
  assign n15276 = n15265 & ~n15273 ;
  assign n15274 = n15273 ^ n15229 ;
  assign n15275 = n15265 & ~n15274 ;
  assign n15277 = n15276 ^ n15275 ;
  assign n15231 = n15230 ^ n15229 ;
  assign n15271 = ~n15231 & n15265 ;
  assign n15272 = n15271 ^ n15265 ;
  assign n15278 = n15277 ^ n15272 ;
  assign n15280 = n15279 ^ n15278 ;
  assign n15269 = n15230 & n15263 ;
  assign n15270 = n15269 ^ n15230 ;
  assign n15281 = n15280 ^ n15270 ;
  assign n15283 = n15282 ^ n15281 ;
  assign n15267 = ~n15231 & ~n15266 ;
  assign n15268 = n15267 ^ n15266 ;
  assign n15284 = n15283 ^ n15268 ;
  assign n15285 = n15199 & ~n15284 ;
  assign n15346 = n15199 ^ n15197 ;
  assign n15347 = n15346 ^ n15196 ;
  assign n15288 = n15263 & ~n15274 ;
  assign n15311 = n15288 ^ n15279 ;
  assign n15287 = ~n15231 & n15263 ;
  assign n15312 = n15311 ^ n15287 ;
  assign n15309 = n15262 ^ n15200 ;
  assign n15310 = n15261 & n15309 ;
  assign n15313 = n15312 ^ n15310 ;
  assign n15306 = n15282 ^ n15271 ;
  assign n15307 = n15306 ^ n15231 ;
  assign n15304 = n15287 ^ n15282 ;
  assign n15305 = n15304 ^ n15267 ;
  assign n15308 = n15307 ^ n15305 ;
  assign n15314 = n15313 ^ n15308 ;
  assign n15374 = n15314 ^ n15275 ;
  assign n15375 = n15347 & ~n15374 ;
  assign n15368 = n15284 ^ n15267 ;
  assign n15369 = n15267 ^ n15197 ;
  assign n15370 = n15369 ^ n15267 ;
  assign n15371 = ~n15368 & n15370 ;
  assign n15372 = n15371 ^ n15267 ;
  assign n15373 = n15196 & n15372 ;
  assign n15376 = n15375 ^ n15373 ;
  assign n15365 = ~n15284 & ~n15346 ;
  assign n15354 = n15313 ^ n15271 ;
  assign n15357 = n15197 & n15354 ;
  assign n15349 = n15278 ^ n15267 ;
  assign n15350 = ~n15197 & n15349 ;
  assign n15351 = n15350 ^ n15267 ;
  assign n15358 = n15357 ^ n15351 ;
  assign n15359 = n15196 & n15358 ;
  assign n15360 = n15359 ^ n15351 ;
  assign n15348 = n15269 & n15347 ;
  assign n15361 = n15360 ^ n15348 ;
  assign n15344 = n15199 & n15276 ;
  assign n15334 = n15311 ^ n15271 ;
  assign n15335 = n15334 ^ n15314 ;
  assign n15336 = n15335 ^ n15334 ;
  assign n15337 = n15334 ^ n15196 ;
  assign n15338 = n15337 ^ n15334 ;
  assign n15339 = ~n15336 & ~n15338 ;
  assign n15340 = n15339 ^ n15334 ;
  assign n15341 = ~n15197 & n15340 ;
  assign n15342 = n15341 ^ n15288 ;
  assign n15286 = n15197 ^ n15196 ;
  assign n15326 = n15308 ^ n15276 ;
  assign n15327 = n15326 ^ n15288 ;
  assign n15328 = n15327 ^ n15279 ;
  assign n15329 = n15279 ^ n15197 ;
  assign n15330 = n15329 ^ n15279 ;
  assign n15331 = ~n15328 & n15330 ;
  assign n15332 = n15331 ^ n15279 ;
  assign n15333 = ~n15286 & n15332 ;
  assign n15343 = n15342 ^ n15333 ;
  assign n15345 = n15344 ^ n15343 ;
  assign n15362 = n15361 ^ n15345 ;
  assign n15317 = n15269 ^ n15263 ;
  assign n15289 = n15288 ^ n15287 ;
  assign n15318 = n15317 ^ n15289 ;
  assign n15315 = n15314 ^ n15279 ;
  assign n15316 = n15315 ^ n15264 ;
  assign n15319 = n15318 ^ n15316 ;
  assign n15320 = n15318 ^ n15197 ;
  assign n15321 = n15320 ^ n15318 ;
  assign n15322 = ~n15319 & ~n15321 ;
  assign n15323 = n15322 ^ n15318 ;
  assign n15324 = n15286 & n15323 ;
  assign n15363 = n15362 ^ n15324 ;
  assign n15364 = n15363 ^ n15283 ;
  assign n15366 = n15365 ^ n15364 ;
  assign n15299 = n15288 ^ n15197 ;
  assign n15300 = n15299 ^ n15288 ;
  assign n15301 = n15289 & n15300 ;
  assign n15302 = n15301 ^ n15288 ;
  assign n15303 = ~n15286 & n15302 ;
  assign n15367 = n15366 ^ n15303 ;
  assign n15377 = n15376 ^ n15367 ;
  assign n15291 = n15283 ^ n15278 ;
  assign n15290 = n15289 ^ n15263 ;
  assign n15292 = n15291 ^ n15290 ;
  assign n15293 = n15292 ^ n15283 ;
  assign n15294 = ~n15197 & n15293 ;
  assign n15295 = n15294 ^ n15291 ;
  assign n15296 = n15286 & n15295 ;
  assign n15378 = n15377 ^ n15296 ;
  assign n15379 = ~n15285 & ~n15378 ;
  assign n15380 = n15379 ^ n10541 ;
  assign n15381 = n15380 ^ x115 ;
  assign n15468 = ~n15195 & ~n15381 ;
  assign n11077 = n11076 ^ n10782 ;
  assign n11502 = n11501 ^ n11495 ;
  assign n11503 = ~n11467 & ~n11502 ;
  assign n11504 = n11503 ^ n11501 ;
  assign n11510 = n11509 ^ n11504 ;
  assign n11506 = n11505 ^ n11504 ;
  assign n11511 = n11510 ^ n11506 ;
  assign n11512 = n11510 ^ n11467 ;
  assign n11513 = n11512 ^ n11510 ;
  assign n11514 = ~n11511 & ~n11513 ;
  assign n11515 = n11514 ^ n11510 ;
  assign n11516 = ~n11274 & ~n11515 ;
  assign n11517 = n11516 ^ n11504 ;
  assign n11518 = ~n11077 & n11517 ;
  assign n11519 = n11518 ^ n8853 ;
  assign n11520 = n11519 ^ x92 ;
  assign n12972 = n12971 ^ n12902 ;
  assign n12985 = n12984 ^ n12972 ;
  assign n12986 = n12985 ^ n12983 ;
  assign n12973 = n12972 ^ n12910 ;
  assign n12967 = n12895 ^ n12827 ;
  assign n12968 = n12967 ^ n12910 ;
  assign n12969 = n12968 ^ n12940 ;
  assign n12970 = ~n12915 & n12969 ;
  assign n12974 = n12973 ^ n12970 ;
  assign n12975 = n12919 & ~n12974 ;
  assign n12987 = n12986 ^ n12975 ;
  assign n12988 = n12987 ^ n12966 ;
  assign n12990 = n12989 ^ n12988 ;
  assign n12991 = ~n12916 & n12990 ;
  assign n12995 = n12994 ^ n12911 ;
  assign n12998 = n12915 & ~n12995 ;
  assign n12999 = n12998 ^ n12911 ;
  assign n13000 = n12991 & n12999 ;
  assign n13001 = n13000 ^ n12990 ;
  assign n13002 = ~n12965 & n13001 ;
  assign n13003 = ~n12957 & n13002 ;
  assign n13006 = n13003 ^ n8463 ;
  assign n12914 = n12913 ^ n12900 ;
  assign n13004 = n12918 & n13003 ;
  assign n13005 = n12914 & n13004 ;
  assign n13007 = n13006 ^ n13005 ;
  assign n13008 = n13007 ^ x78 ;
  assign n13017 = n11520 & n13008 ;
  assign n13056 = n13017 ^ n11520 ;
  assign n13057 = n13056 ^ n13008 ;
  assign n13058 = n13057 ^ n11520 ;
  assign n11919 = n11814 ^ n11727 ;
  assign n11920 = n11919 ^ n11871 ;
  assign n11921 = n11920 ^ n11878 ;
  assign n11922 = n11561 & n11921 ;
  assign n11923 = n11922 ^ n11871 ;
  assign n11924 = n11683 & n11923 ;
  assign n11925 = n11924 ^ n11871 ;
  assign n11933 = n11894 ^ n11874 ;
  assign n11934 = n11933 ^ n11932 ;
  assign n11935 = ~n11561 & ~n11934 ;
  assign n11926 = n11892 ^ n11864 ;
  assign n11927 = n11926 ^ n11905 ;
  assign n11930 = n11927 ^ n11905 ;
  assign n11936 = n11935 ^ n11930 ;
  assign n11928 = n11927 ^ n11908 ;
  assign n11929 = n11561 & n11928 ;
  assign n11937 = n11936 ^ n11929 ;
  assign n11938 = n11678 & n11937 ;
  assign n11939 = n11938 ^ n11935 ;
  assign n11940 = ~n11925 & ~n11939 ;
  assign n11896 = n11895 ^ n11885 ;
  assign n11918 = n11917 ^ n11896 ;
  assign n11941 = n11940 ^ n11918 ;
  assign n11944 = n11943 ^ n11941 ;
  assign n11945 = n11944 ^ n9423 ;
  assign n11946 = n11945 ^ x110 ;
  assign n12382 = n12314 ^ n12303 ;
  assign n12383 = n12382 ^ n12327 ;
  assign n12384 = ~n11973 & n12383 ;
  assign n12379 = n12378 ^ n12310 ;
  assign n12380 = n12379 ^ n12376 ;
  assign n12381 = n12380 ^ n12368 ;
  assign n12385 = n12384 ^ n12381 ;
  assign n12402 = n12401 ^ n12385 ;
  assign n12386 = n12385 ^ n12376 ;
  assign n12387 = n12386 ^ n12368 ;
  assign n12362 = n11973 & n12328 ;
  assign n12388 = n12387 ^ n12362 ;
  assign n12389 = n12351 & n12388 ;
  assign n12403 = n12402 ^ n12389 ;
  assign n12360 = n12316 ^ n12310 ;
  assign n12361 = n12359 & n12360 ;
  assign n12404 = n12403 ^ n12361 ;
  assign n12354 = n12324 ^ n11998 ;
  assign n12355 = n12354 ^ n12324 ;
  assign n12356 = n12326 & ~n12355 ;
  assign n12357 = n12356 ^ n12324 ;
  assign n12358 = ~n12351 & n12357 ;
  assign n12405 = n12404 ^ n12358 ;
  assign n12406 = n12405 ^ n12350 ;
  assign n12407 = n12406 ^ n9677 ;
  assign n12000 = n11999 ^ n11973 ;
  assign n12334 = n12333 ^ n12323 ;
  assign n12335 = n12000 & ~n12334 ;
  assign n12408 = n12407 ^ n12335 ;
  assign n12409 = n12408 ^ x91 ;
  assign n12410 = ~n11946 & ~n12409 ;
  assign n13018 = n12410 ^ n12409 ;
  assign n12612 = n12611 ^ n9875 ;
  assign n12578 = n12458 ^ n12457 ;
  assign n12581 = n12580 ^ n12541 ;
  assign n12582 = n12581 ^ n12539 ;
  assign n12579 = n12574 ^ n12555 ;
  assign n12583 = n12582 ^ n12579 ;
  assign n12584 = n12458 & n12583 ;
  assign n12585 = n12584 ^ n12582 ;
  assign n12586 = n12585 ^ n12560 ;
  assign n12587 = n12586 ^ n12571 ;
  assign n12588 = n12587 ^ n12543 ;
  assign n12589 = n12588 ^ n12585 ;
  assign n12590 = n12458 & n12589 ;
  assign n12591 = n12590 ^ n12586 ;
  assign n12592 = ~n12578 & ~n12591 ;
  assign n12593 = n12592 ^ n12585 ;
  assign n12577 = n12458 & n12545 ;
  assign n12594 = n12593 ^ n12577 ;
  assign n12595 = ~n12576 & ~n12594 ;
  assign n12607 = n12595 & ~n12606 ;
  assign n12613 = n12612 ^ n12607 ;
  assign n12614 = n12613 ^ x116 ;
  assign n12717 = n12716 ^ n12703 ;
  assign n12718 = n12615 & ~n12717 ;
  assign n12801 = ~n12615 & n12777 ;
  assign n12802 = n12801 ^ n12768 ;
  assign n12814 = n12802 ^ n9131 ;
  assign n12815 = n12814 ^ n12813 ;
  assign n12804 = n12802 ^ n12710 ;
  assign n12800 = n12791 ^ n12773 ;
  assign n12803 = n12802 ^ n12800 ;
  assign n12805 = n12804 ^ n12803 ;
  assign n12806 = n12804 ^ n12615 ;
  assign n12807 = n12806 ^ n12804 ;
  assign n12808 = ~n12805 & n12807 ;
  assign n12809 = n12808 ^ n12804 ;
  assign n12810 = n12763 & n12809 ;
  assign n12816 = n12815 ^ n12810 ;
  assign n12797 = n12794 ^ n12712 ;
  assign n12817 = n12816 ^ n12797 ;
  assign n12788 = n12771 ^ n12697 ;
  assign n12795 = n12794 ^ n12788 ;
  assign n12798 = n12796 & n12797 ;
  assign n12799 = ~n12795 & n12798 ;
  assign n12818 = n12817 ^ n12799 ;
  assign n12786 = n12785 ^ n12778 ;
  assign n12787 = n12763 & n12786 ;
  assign n12819 = n12818 ^ n12787 ;
  assign n12820 = n12819 ^ n12816 ;
  assign n12821 = n12718 & ~n12820 ;
  assign n12822 = n12821 ^ n12819 ;
  assign n12823 = n12822 ^ x109 ;
  assign n12824 = n12614 & ~n12823 ;
  assign n13041 = n12824 ^ n12823 ;
  assign n13042 = ~n13018 & ~n13041 ;
  assign n13009 = n12824 ^ n12614 ;
  assign n13019 = n13009 & ~n13018 ;
  assign n13043 = n13042 ^ n13019 ;
  assign n13035 = n12824 & ~n13018 ;
  assign n13011 = n12410 ^ n11946 ;
  assign n13021 = n12824 & ~n13011 ;
  assign n13012 = n13009 ^ n12823 ;
  assign n13013 = ~n13011 & n13012 ;
  assign n13034 = n13021 ^ n13013 ;
  assign n13036 = n13035 ^ n13034 ;
  assign n12825 = n12410 & n12824 ;
  assign n13032 = n13013 ^ n12825 ;
  assign n13033 = n13032 ^ n12824 ;
  assign n13037 = n13036 ^ n13033 ;
  assign n13030 = n13011 ^ n12409 ;
  assign n13031 = n13012 & ~n13030 ;
  assign n13038 = n13037 ^ n13031 ;
  assign n13025 = n13013 ^ n13011 ;
  assign n13022 = ~n12823 & ~n13011 ;
  assign n13026 = n13025 ^ n13022 ;
  assign n13023 = n13022 ^ n13021 ;
  assign n13010 = n12410 & n13009 ;
  assign n13024 = n13023 ^ n13010 ;
  assign n13027 = n13026 ^ n13024 ;
  assign n13028 = n13027 ^ n13023 ;
  assign n13020 = n13019 ^ n13009 ;
  assign n13029 = n13028 ^ n13020 ;
  assign n13039 = n13038 ^ n13029 ;
  assign n13040 = n13039 ^ n13030 ;
  assign n13044 = n13043 ^ n13040 ;
  assign n13075 = n13044 ^ n13035 ;
  assign n13074 = n13039 ^ n11946 ;
  assign n13076 = n13075 ^ n13074 ;
  assign n14713 = n13058 & ~n13076 ;
  assign n13049 = n12823 ^ n12614 ;
  assign n13050 = n11946 & ~n13049 ;
  assign n13051 = n13050 ^ n12614 ;
  assign n13052 = n13051 ^ n12823 ;
  assign n13053 = n13052 ^ n13027 ;
  assign n15423 = n13053 ^ n13026 ;
  assign n15424 = n15423 ^ n11520 ;
  assign n15426 = n15423 ^ n13022 ;
  assign n15425 = n15423 ^ n13032 ;
  assign n15427 = n15426 ^ n15425 ;
  assign n15428 = n15426 ^ n13008 ;
  assign n15429 = n15428 ^ n15426 ;
  assign n15430 = n15427 & n15429 ;
  assign n15431 = n15430 ^ n15426 ;
  assign n15432 = n15424 & n15431 ;
  assign n15433 = n15432 ^ n11520 ;
  assign n13047 = n13008 ^ n11520 ;
  assign n15422 = n13031 & ~n13047 ;
  assign n15434 = n15433 ^ n15422 ;
  assign n15414 = n13076 ^ n13035 ;
  assign n15415 = n15414 ^ n13019 ;
  assign n15416 = n15415 ^ n13037 ;
  assign n15413 = n12823 ^ n11946 ;
  assign n15417 = n15416 ^ n15413 ;
  assign n15412 = n12409 & n13051 ;
  assign n15418 = n15417 ^ n15412 ;
  assign n15419 = n13008 & ~n15418 ;
  assign n15420 = n15419 ^ n15416 ;
  assign n15421 = n11520 & ~n15420 ;
  assign n15435 = n15434 ^ n15421 ;
  assign n15436 = ~n14713 & n15435 ;
  assign n15437 = n13037 ^ n13029 ;
  assign n15438 = ~n11520 & ~n15437 ;
  assign n15439 = n15438 ^ n13040 ;
  assign n15441 = n15439 ^ n15426 ;
  assign n15440 = n15439 ^ n15415 ;
  assign n15442 = n15441 ^ n15440 ;
  assign n15445 = ~n11520 & n15442 ;
  assign n15446 = n15445 ^ n15441 ;
  assign n15447 = ~n13008 & ~n15446 ;
  assign n15448 = n15447 ^ n15439 ;
  assign n15449 = n15436 & ~n15448 ;
  assign n15450 = n15449 ^ n9965 ;
  assign n15451 = n15450 ^ x105 ;
  assign n15458 = ~n15195 & ~n15451 ;
  assign n15469 = n15468 ^ n15458 ;
  assign n15473 = ~n15409 & n15469 ;
  assign n13577 = n11945 ^ x85 ;
  assign n13572 = ~n12716 & ~n13125 ;
  assign n13568 = n13567 ^ n12711 ;
  assign n13569 = n12789 & n13568 ;
  assign n13560 = n12771 ^ n12703 ;
  assign n13561 = n13560 ^ n12800 ;
  assign n13562 = n12615 & ~n13561 ;
  assign n13556 = n12791 ^ n12783 ;
  assign n13557 = n13556 ^ n12769 ;
  assign n13564 = n13562 ^ n13557 ;
  assign n13565 = ~n12763 & ~n13564 ;
  assign n13558 = n13557 ^ n13114 ;
  assign n13555 = n12813 ^ n11101 ;
  assign n13559 = n13558 ^ n13555 ;
  assign n13566 = n13565 ^ n13559 ;
  assign n13570 = n13569 ^ n13566 ;
  assign n13553 = n12774 ^ n12695 ;
  assign n13554 = n12763 & n13553 ;
  assign n13571 = n13570 ^ n13554 ;
  assign n13573 = n13572 ^ n13571 ;
  assign n13551 = n12712 ^ n12696 ;
  assign n13552 = ~n12615 & ~n13551 ;
  assign n13574 = n13573 ^ n13552 ;
  assign n13550 = n12696 & n12789 ;
  assign n13575 = n13574 ^ n13550 ;
  assign n13576 = n13575 ^ x94 ;
  assign n13578 = n13577 ^ n13576 ;
  assign n13579 = n13007 ^ x76 ;
  assign n13626 = n13377 ^ n13375 ;
  assign n13627 = n13626 ^ n11137 ;
  assign n13628 = n13627 ^ x67 ;
  assign n13630 = ~n13579 & n13628 ;
  assign n13613 = ~n13232 & ~n13257 ;
  assign n13609 = n13608 ^ n13248 ;
  assign n13610 = n13148 & ~n13609 ;
  assign n13596 = ~n13146 & n13233 ;
  assign n13597 = n13596 ^ n13238 ;
  assign n13598 = n13597 ^ n13282 ;
  assign n13581 = n13257 ^ n13219 ;
  assign n13583 = n13233 ^ n13146 ;
  assign n13582 = n13257 ^ n13225 ;
  assign n13584 = n13583 ^ n13582 ;
  assign n13585 = n13225 ^ n13146 ;
  assign n13586 = n13585 ^ n13583 ;
  assign n13587 = n13584 & ~n13586 ;
  assign n13588 = n13587 ^ n13583 ;
  assign n13589 = n13581 & ~n13588 ;
  assign n13590 = n13589 ^ n13219 ;
  assign n13599 = n13598 ^ n13590 ;
  assign n13600 = n13599 ^ n13257 ;
  assign n13592 = ~n13149 & ~n13249 ;
  assign n13593 = n13592 ^ n13290 ;
  assign n13594 = ~n13240 & n13257 ;
  assign n13595 = ~n13593 & n13594 ;
  assign n13601 = n13600 ^ n13595 ;
  assign n13602 = n13601 ^ n13238 ;
  assign n13603 = n13602 ^ n13590 ;
  assign n13604 = n13299 ^ n13243 ;
  assign n13605 = n13146 & n13604 ;
  assign n13606 = n13603 & n13605 ;
  assign n13607 = n13606 ^ n13601 ;
  assign n13611 = n13610 ^ n13607 ;
  assign n13580 = ~n13146 & n13221 ;
  assign n13612 = n13611 ^ n13580 ;
  assign n13614 = n13613 ^ n13612 ;
  assign n13622 = ~n13614 & ~n13621 ;
  assign n13623 = n13622 ^ n11133 ;
  assign n13624 = n13623 ^ x124 ;
  assign n13715 = n13708 & n13714 ;
  assign n13720 = n13714 & n13719 ;
  assign n13725 = n13724 ^ n13720 ;
  assign n13726 = n13710 ^ n13709 ;
  assign n13783 = n13726 & n13751 ;
  assign n13765 = n13753 ^ n13723 ;
  assign n13764 = n13763 ^ n13700 ;
  assign n13766 = n13765 ^ n13764 ;
  assign n13767 = ~n13709 & ~n13766 ;
  assign n13768 = n13767 ^ n13765 ;
  assign n13779 = n13774 ^ n13768 ;
  assign n13770 = n13759 ^ n13740 ;
  assign n13775 = n13774 ^ n13770 ;
  assign n13777 = n13776 ^ n13775 ;
  assign n13778 = n13709 & ~n13777 ;
  assign n13780 = n13779 ^ n13778 ;
  assign n13781 = n13710 & n13780 ;
  assign n13741 = n13740 ^ n13719 ;
  assign n13742 = n13719 ^ n13709 ;
  assign n13743 = n13742 ^ n13719 ;
  assign n13744 = ~n13741 & ~n13743 ;
  assign n13745 = n13744 ^ n13719 ;
  assign n13746 = n13726 & n13745 ;
  assign n13769 = n13768 ^ n13746 ;
  assign n13782 = n13781 ^ n13769 ;
  assign n13784 = n13783 ^ n13782 ;
  assign n13785 = ~n13725 & ~n13784 ;
  assign n13792 = n13785 & ~n13791 ;
  assign n13793 = ~n13715 & n13792 ;
  assign n13798 = n13743 & ~n13795 ;
  assign n13799 = n13798 ^ n13719 ;
  assign n13800 = ~n13710 & n13799 ;
  assign n13801 = n13793 & ~n13800 ;
  assign n13802 = n13801 ^ n11174 ;
  assign n13803 = n13802 ^ x117 ;
  assign n13804 = ~n13624 & n13803 ;
  assign n13805 = n13804 ^ n13624 ;
  assign n13806 = n13805 ^ n13803 ;
  assign n13820 = n13630 & n13806 ;
  assign n13843 = n13820 ^ n13806 ;
  assign n13631 = n13630 ^ n13628 ;
  assign n13823 = n13631 ^ n13579 ;
  assign n13840 = n13823 ^ n13628 ;
  assign n13841 = n13806 & ~n13840 ;
  assign n13810 = n13631 & n13806 ;
  assign n13842 = n13841 ^ n13810 ;
  assign n13844 = n13843 ^ n13842 ;
  assign n13835 = n13804 & n13823 ;
  assign n13809 = n13630 & ~n13805 ;
  assign n13811 = n13810 ^ n13809 ;
  assign n13807 = n13806 ^ n13624 ;
  assign n13808 = n13631 & n13807 ;
  assign n13812 = n13811 ^ n13808 ;
  assign n13629 = ~n13624 & n13628 ;
  assign n13632 = n13631 ^ n13629 ;
  assign n13813 = n13812 ^ n13632 ;
  assign n13814 = n13813 ^ n13808 ;
  assign n13836 = n13835 ^ n13814 ;
  assign n13625 = ~n13579 & ~n13624 ;
  assign n13831 = n13628 ^ n13625 ;
  assign n13832 = n13803 & ~n13831 ;
  assign n13833 = n13832 ^ n13803 ;
  assign n13834 = n13833 ^ n13804 ;
  assign n13837 = n13836 ^ n13834 ;
  assign n13838 = n13837 ^ n13808 ;
  assign n13824 = ~n13805 & n13823 ;
  assign n13825 = n13824 ^ n13820 ;
  assign n13826 = n13825 ^ n13809 ;
  assign n13819 = n13631 & ~n13805 ;
  assign n13821 = n13820 ^ n13819 ;
  assign n13822 = n13821 ^ n13805 ;
  assign n13827 = n13826 ^ n13822 ;
  assign n13816 = n13624 ^ n13579 ;
  assign n13817 = n13803 ^ n13629 ;
  assign n13818 = ~n13816 & n13817 ;
  assign n13828 = n13827 ^ n13818 ;
  assign n13815 = n13814 ^ n13625 ;
  assign n13829 = n13828 ^ n13815 ;
  assign n13830 = n13829 ^ n13807 ;
  assign n13839 = n13838 ^ n13830 ;
  assign n13845 = n13844 ^ n13839 ;
  assign n13846 = n13844 ^ n13577 ;
  assign n13847 = n13846 ^ n13844 ;
  assign n13848 = ~n13845 & ~n13847 ;
  assign n13849 = n13848 ^ n13844 ;
  assign n13850 = n13578 & n13849 ;
  assign n15165 = n13850 ^ n11273 ;
  assign n13864 = n13827 ^ n13577 ;
  assign n13865 = n13864 ^ n13827 ;
  assign n13885 = n13631 & n13804 ;
  assign n13886 = n13885 ^ n13838 ;
  assign n13887 = n13886 ^ n13833 ;
  assign n13888 = n13887 ^ n13885 ;
  assign n13889 = n13888 ^ n13827 ;
  assign n13890 = ~n13865 & ~n13889 ;
  assign n13891 = n13890 ^ n13827 ;
  assign n13892 = n13576 & ~n13891 ;
  assign n13852 = n13576 & n13577 ;
  assign n13853 = n13852 ^ n13576 ;
  assign n13854 = n13844 & n13853 ;
  assign n15149 = n13844 ^ n13818 ;
  assign n15148 = n13825 ^ n13819 ;
  assign n15150 = n15149 ^ n15148 ;
  assign n15147 = n13839 ^ n13826 ;
  assign n15151 = n15150 ^ n15147 ;
  assign n15152 = n13577 & n15151 ;
  assign n15153 = n15152 ^ n15150 ;
  assign n15159 = n15153 ^ n13812 ;
  assign n15156 = n13844 ^ n13814 ;
  assign n15157 = n15156 ^ n13819 ;
  assign n15158 = n13577 & n15157 ;
  assign n15160 = n15159 ^ n15158 ;
  assign n15161 = n13576 & ~n15160 ;
  assign n15140 = n13837 ^ n13829 ;
  assign n15141 = n15140 ^ n13887 ;
  assign n15142 = n13887 ^ n13576 ;
  assign n15143 = n15142 ^ n13887 ;
  assign n15144 = ~n15141 & n15143 ;
  assign n15145 = n15144 ^ n13887 ;
  assign n15146 = n13577 & n15145 ;
  assign n15154 = n15153 ^ n15146 ;
  assign n14817 = n13827 ^ n13814 ;
  assign n14818 = n13814 ^ n13577 ;
  assign n14819 = n14818 ^ n13814 ;
  assign n14820 = ~n14817 & ~n14819 ;
  assign n14821 = n14820 ^ n13814 ;
  assign n14822 = n13578 & n14821 ;
  assign n15155 = n15154 ^ n14822 ;
  assign n15162 = n15161 ^ n15155 ;
  assign n15163 = ~n13854 & n15162 ;
  assign n15164 = ~n13892 & n15163 ;
  assign n15166 = n15165 ^ n15164 ;
  assign n15167 = n15166 ^ x72 ;
  assign n15410 = n15409 ^ n15381 ;
  assign n15411 = n15410 ^ n15195 ;
  assign n15452 = n15451 ^ n15381 ;
  assign n15453 = n15381 ^ n15195 ;
  assign n15454 = ~n15452 & ~n15453 ;
  assign n15455 = n15454 ^ n15381 ;
  assign n15456 = n15411 & ~n15455 ;
  assign n15459 = n15458 ^ n15381 ;
  assign n15460 = ~n15411 & n15459 ;
  assign n15461 = n15460 ^ n15452 ;
  assign n15471 = ~n15456 & n15461 ;
  assign n14163 = n12613 ^ x104 ;
  assign n14311 = n14310 ^ x82 ;
  assign n14164 = ~n12951 & ~n13426 ;
  assign n14176 = n12909 ^ n12904 ;
  assign n14177 = n14176 ^ n12939 ;
  assign n14178 = ~n12915 & n14177 ;
  assign n14179 = n14178 ^ n12938 ;
  assign n14180 = ~n12916 & n14179 ;
  assign n14173 = n12915 & n12939 ;
  assign n14171 = n13435 ^ n12935 ;
  assign n14172 = n14171 ^ n13957 ;
  assign n14174 = n14173 ^ n14172 ;
  assign n14181 = n14180 ^ n14174 ;
  assign n14165 = n12993 ^ n12941 ;
  assign n14166 = n12941 ^ n12916 ;
  assign n14167 = n14166 ^ n12941 ;
  assign n14168 = n14165 & n14167 ;
  assign n14169 = n14168 ^ n12941 ;
  assign n14170 = n12915 & ~n14169 ;
  assign n14182 = n14181 ^ n14170 ;
  assign n14183 = ~n13932 & ~n14182 ;
  assign n14184 = n14164 & n14183 ;
  assign n14185 = n14184 ^ n11374 ;
  assign n14186 = n14185 ^ x99 ;
  assign n14218 = n14217 ^ x114 ;
  assign n14219 = n14186 & ~n14218 ;
  assign n14327 = n14219 ^ n14186 ;
  assign n14229 = n13710 ^ n13706 ;
  assign n14230 = n13740 ^ n13710 ;
  assign n14231 = n14230 ^ n13758 ;
  assign n14232 = n14231 ^ n14230 ;
  assign n14233 = n14230 ^ n13709 ;
  assign n14234 = n14233 ^ n14230 ;
  assign n14235 = n14232 & ~n14234 ;
  assign n14236 = n14235 ^ n14230 ;
  assign n14237 = ~n14229 & ~n14236 ;
  assign n14238 = n14237 ^ n13706 ;
  assign n14224 = n13762 ^ n13709 ;
  assign n14225 = n14224 ^ n13762 ;
  assign n14226 = n13763 & ~n14225 ;
  assign n14227 = n14226 ^ n13762 ;
  assign n14228 = n13710 & ~n14227 ;
  assign n14239 = n14238 ^ n14228 ;
  assign n14221 = n13713 & n13760 ;
  assign n14240 = n14239 ^ n14221 ;
  assign n14241 = n13772 ^ n13710 ;
  assign n14242 = n14241 ^ n13709 ;
  assign n14243 = ~n14240 & ~n14242 ;
  assign n14244 = n14243 ^ n14240 ;
  assign n14245 = n14244 ^ n13728 ;
  assign n14246 = n14245 ^ n14244 ;
  assign n14251 = ~n13710 & n14243 ;
  assign n14252 = n14246 & n14251 ;
  assign n14253 = n14252 ^ n14246 ;
  assign n14254 = n14253 ^ n14245 ;
  assign n14255 = ~n13726 & ~n14254 ;
  assign n14256 = n14255 ^ n14240 ;
  assign n14257 = n13709 & ~n14256 ;
  assign n14258 = n13747 ^ n13710 ;
  assign n14259 = n14258 ^ n13747 ;
  assign n14260 = n13747 ^ n13722 ;
  assign n14261 = n14260 ^ n13747 ;
  assign n14262 = ~n14259 & n14261 ;
  assign n14263 = n14262 ^ n13747 ;
  assign n14264 = n14257 & n14263 ;
  assign n14265 = n14264 ^ n14256 ;
  assign n14266 = ~n13746 & ~n14265 ;
  assign n14267 = ~n13715 & ~n13897 ;
  assign n14268 = n14266 & n14267 ;
  assign n14269 = n14268 ^ n11326 ;
  assign n14270 = n14269 ^ x89 ;
  assign n14271 = n11519 ^ x80 ;
  assign n14272 = n14270 & n14271 ;
  assign n14334 = n14272 ^ n14271 ;
  assign n14335 = n14327 & n14334 ;
  assign n14220 = n14219 ^ n14218 ;
  assign n14318 = n14220 ^ n14186 ;
  assign n14330 = n14272 & n14318 ;
  assign n15133 = n14335 ^ n14330 ;
  assign n14339 = n14318 & n14334 ;
  assign n14338 = n14219 & n14334 ;
  assign n14340 = n14339 ^ n14338 ;
  assign n14328 = n14272 & n14327 ;
  assign n14341 = n14340 ^ n14328 ;
  assign n14329 = n14328 ^ n14272 ;
  assign n14336 = n14335 ^ n14329 ;
  assign n14337 = n14336 ^ n14271 ;
  assign n14342 = n14341 ^ n14337 ;
  assign n14371 = n14342 ^ n14328 ;
  assign n14372 = n14371 ^ n14338 ;
  assign n15134 = n15133 ^ n14372 ;
  assign n15135 = n14311 & n15134 ;
  assign n14273 = n14272 ^ n14270 ;
  assign n14274 = n14273 ^ n14271 ;
  assign n14275 = ~n14220 & ~n14274 ;
  assign n15136 = n15135 ^ n14275 ;
  assign n15137 = ~n14163 & n15136 ;
  assign n14317 = n14219 & ~n14274 ;
  assign n14651 = ~n14163 & n14311 ;
  assign n14653 = n14651 ^ n14311 ;
  assign n14682 = n14653 ^ n14163 ;
  assign n15131 = n14317 & n14682 ;
  assign n15124 = n14651 ^ n14163 ;
  assign n14320 = n14219 & n14273 ;
  assign n14319 = n14273 & n14318 ;
  assign n14321 = n14320 ^ n14319 ;
  assign n14357 = n14321 ^ n14273 ;
  assign n14343 = n14342 ^ n14220 ;
  assign n14276 = n14219 & n14272 ;
  assign n14331 = n14330 ^ n14276 ;
  assign n14332 = n14331 ^ n14329 ;
  assign n14333 = n14332 ^ n14275 ;
  assign n14344 = n14343 ^ n14333 ;
  assign n14358 = n14357 ^ n14344 ;
  assign n14324 = ~n14274 & n14318 ;
  assign n14325 = n14324 ^ n14274 ;
  assign n15125 = n14358 ^ n14325 ;
  assign n15126 = ~n15124 & n15125 ;
  assign n14323 = n14317 ^ n14275 ;
  assign n14326 = n14325 ^ n14323 ;
  assign n15119 = n14326 ^ n14320 ;
  assign n15120 = n15119 ^ n14324 ;
  assign n15121 = n15120 ^ n14332 ;
  assign n15122 = n14653 & ~n15121 ;
  assign n14368 = n14311 ^ n14163 ;
  assign n15103 = n14328 ^ n14276 ;
  assign n15104 = n15103 ^ n14336 ;
  assign n15105 = n14311 & n15104 ;
  assign n15106 = n15105 ^ n14336 ;
  assign n15107 = n15106 ^ n14163 ;
  assign n15108 = n15107 ^ n15106 ;
  assign n15109 = n15107 ^ n14276 ;
  assign n15110 = n15109 ^ n15107 ;
  assign n15111 = n15107 ^ n14341 ;
  assign n15112 = n15111 ^ n15107 ;
  assign n15113 = ~n15110 & ~n15112 ;
  assign n15114 = n15108 & n15113 ;
  assign n15115 = n15114 ^ n15108 ;
  assign n15116 = n15115 ^ n15106 ;
  assign n15117 = n14368 & n15116 ;
  assign n15118 = n15117 ^ n15106 ;
  assign n15123 = n15122 ^ n15118 ;
  assign n15127 = n15126 ^ n15123 ;
  assign n15128 = n15127 ^ n14275 ;
  assign n14345 = n14344 ^ n14326 ;
  assign n14346 = n14345 ^ n14339 ;
  assign n14347 = ~n14311 & n14346 ;
  assign n14348 = n14347 ^ n14339 ;
  assign n14322 = n14321 ^ n14317 ;
  assign n14349 = n14348 ^ n14322 ;
  assign n14350 = n14349 ^ n14348 ;
  assign n14353 = n14311 & n14350 ;
  assign n14354 = n14353 ^ n14348 ;
  assign n14355 = ~n14163 & n14354 ;
  assign n14356 = n14355 ^ n14348 ;
  assign n15129 = n15128 ^ n14356 ;
  assign n15130 = n15129 ^ n11466 ;
  assign n15132 = n15131 ^ n15130 ;
  assign n15138 = n15137 ^ n15132 ;
  assign n15139 = n15138 ^ x90 ;
  assign n16924 = n15471 ^ n15139 ;
  assign n15463 = n15451 ^ n15195 ;
  assign n15465 = n15463 ^ n15381 ;
  assign n15466 = n15410 & ~n15465 ;
  assign n15467 = n15466 ^ n15409 ;
  assign n15475 = n15451 ^ n15409 ;
  assign n15476 = ~n15467 & ~n15475 ;
  assign n16920 = n15476 ^ n15463 ;
  assign n16921 = n16920 ^ n15471 ;
  assign n16922 = n15139 & n16921 ;
  assign n16923 = n16922 ^ n16920 ;
  assign n16925 = n16924 ^ n16923 ;
  assign n16926 = n16925 ^ n16920 ;
  assign n16928 = n16926 ^ n15461 ;
  assign n15457 = n15456 ^ n15195 ;
  assign n16927 = n16926 ^ n15457 ;
  assign n16929 = n16928 ^ n16927 ;
  assign n16930 = n16928 ^ n15139 ;
  assign n16931 = n16930 ^ n16928 ;
  assign n16932 = ~n16929 & n16931 ;
  assign n16933 = n16932 ^ n16928 ;
  assign n16934 = n15167 & ~n16933 ;
  assign n16935 = n16934 ^ n16926 ;
  assign n16936 = ~n15473 & ~n16935 ;
  assign n16937 = n16936 ^ n11519 ;
  assign n16938 = n16937 ^ x113 ;
  assign n14837 = n14022 ^ x88 ;
  assign n14876 = ~n13294 & ~n13597 ;
  assign n14891 = n13266 ^ n13252 ;
  assign n14892 = n14891 ^ n13281 ;
  assign n14893 = n14892 ^ n13248 ;
  assign n14894 = ~n13592 & ~n14893 ;
  assign n14895 = n14894 ^ n13298 ;
  assign n14903 = n14895 ^ n13280 ;
  assign n14896 = n14895 ^ n13265 ;
  assign n14897 = n14896 ^ n13243 ;
  assign n14898 = n14897 ^ n13267 ;
  assign n14899 = n14898 ^ n14895 ;
  assign n14900 = ~n13146 & ~n14899 ;
  assign n14901 = n14900 ^ n14896 ;
  assign n14902 = n13145 & ~n14901 ;
  assign n14904 = n14903 ^ n14902 ;
  assign n14883 = n13246 ^ n13219 ;
  assign n14884 = n14883 ^ n13244 ;
  assign n14885 = n14884 ^ n13219 ;
  assign n14886 = n13219 ^ n13145 ;
  assign n14887 = n14886 ^ n13219 ;
  assign n14888 = n14885 & ~n14887 ;
  assign n14889 = n14888 ^ n13219 ;
  assign n14890 = ~n13146 & n14889 ;
  assign n14905 = n14904 ^ n14890 ;
  assign n14877 = n13262 ^ n13227 ;
  assign n14878 = n13227 ^ n13146 ;
  assign n14879 = n14878 ^ n13227 ;
  assign n14880 = ~n14877 & ~n14879 ;
  assign n14881 = n14880 ^ n13227 ;
  assign n14882 = n13257 & ~n14881 ;
  assign n14906 = n14905 ^ n14882 ;
  assign n14907 = n14876 & n14906 ;
  assign n14908 = n14907 ^ n11599 ;
  assign n14909 = n14908 ^ x121 ;
  assign n14838 = n13143 ^ x112 ;
  assign n14933 = n14909 ^ n14838 ;
  assign n14839 = n13962 ^ x66 ;
  assign n14946 = ~n14839 & n14909 ;
  assign n14948 = n14933 & ~n14946 ;
  assign n14863 = n13923 ^ n13715 ;
  assign n14852 = n13728 ^ n13704 ;
  assign n14853 = ~n13709 & ~n14852 ;
  assign n14851 = n13898 ^ n13723 ;
  assign n14854 = n14853 ^ n14851 ;
  assign n14864 = n14863 ^ n14854 ;
  assign n14855 = n14854 ^ n13762 ;
  assign n14858 = n14855 ^ n13702 ;
  assign n14859 = n14858 ^ n14855 ;
  assign n14860 = ~n13709 & n14859 ;
  assign n14861 = n14860 ^ n14855 ;
  assign n14862 = ~n13710 & ~n14861 ;
  assign n14865 = n14864 ^ n14862 ;
  assign n14849 = n13738 ^ n13722 ;
  assign n14850 = ~n13712 & ~n14849 ;
  assign n14866 = n14865 ^ n14850 ;
  assign n14867 = n14866 ^ n13747 ;
  assign n14848 = n13711 & n13733 ;
  assign n14868 = n14867 ^ n14848 ;
  assign n14841 = n13747 ^ n13713 ;
  assign n14842 = n13912 ^ n13711 ;
  assign n14845 = ~n13747 & n14842 ;
  assign n14846 = n14845 ^ n13711 ;
  assign n14847 = n14841 & ~n14846 ;
  assign n14869 = n14868 ^ n14847 ;
  assign n14870 = ~n13725 & ~n14869 ;
  assign n14871 = ~n13800 & n14870 ;
  assign n14872 = n14871 ^ n11638 ;
  assign n14873 = n14872 ^ x65 ;
  assign n14914 = n14873 ^ n14838 ;
  assign n14917 = n14914 ^ n14839 ;
  assign n14840 = n14839 ^ n14838 ;
  assign n14874 = ~n14840 & ~n14873 ;
  assign n14875 = n14874 ^ n14839 ;
  assign n14918 = n14917 ^ n14875 ;
  assign n14919 = n14909 & ~n14918 ;
  assign n14910 = n14909 ^ n14873 ;
  assign n14920 = n14910 ^ n14838 ;
  assign n14921 = ~n14840 & ~n14920 ;
  assign n14922 = n14839 & ~n14921 ;
  assign n14923 = n14921 ^ n14873 ;
  assign n14924 = n14923 ^ n14838 ;
  assign n14925 = n14922 & n14924 ;
  assign n14926 = n14925 ^ n14923 ;
  assign n14927 = ~n14919 & ~n14926 ;
  assign n14945 = n14927 ^ n14839 ;
  assign n14947 = n14946 ^ n14945 ;
  assign n14949 = n14948 ^ n14947 ;
  assign n14950 = n14837 & ~n14949 ;
  assign n14931 = n14873 ^ n14839 ;
  assign n14911 = ~n14839 & n14910 ;
  assign n14929 = n14911 ^ n14873 ;
  assign n14930 = n14929 ^ n14927 ;
  assign n14932 = n14931 ^ n14930 ;
  assign n14951 = n14950 ^ n14932 ;
  assign n14836 = n13420 ^ x106 ;
  assign n14954 = n14951 ^ n14836 ;
  assign n14934 = n14933 ^ n14932 ;
  assign n14915 = n14914 ^ n14909 ;
  assign n14912 = n14911 ^ n14909 ;
  assign n14913 = n14840 & n14912 ;
  assign n14916 = n14915 ^ n14913 ;
  assign n14928 = n14927 ^ n14916 ;
  assign n14935 = n14934 ^ n14928 ;
  assign n14936 = n14935 ^ n14917 ;
  assign n14937 = n14936 ^ n14875 ;
  assign n14938 = n14937 ^ n14936 ;
  assign n14941 = ~n14909 & n14938 ;
  assign n14942 = n14941 ^ n14936 ;
  assign n14943 = n14837 & n14942 ;
  assign n14944 = n14943 ^ n14935 ;
  assign n14952 = n14951 ^ n14944 ;
  assign n14953 = n14836 & n14952 ;
  assign n14955 = n14954 ^ n14953 ;
  assign n14956 = n14955 ^ n11677 ;
  assign n14957 = n14956 ^ x92 ;
  assign n14961 = n13460 ^ n13383 ;
  assign n13543 = n13495 ^ n13473 ;
  assign n14962 = n14961 ^ n13543 ;
  assign n14963 = n14962 ^ n14960 ;
  assign n14964 = n13309 & n14963 ;
  assign n14959 = n13470 ^ n13383 ;
  assign n14965 = n14964 ^ n14959 ;
  assign n14994 = n14993 ^ n14965 ;
  assign n14995 = n14994 ^ n14989 ;
  assign n13531 = n13144 & n13530 ;
  assign n14996 = n14995 ^ n13531 ;
  assign n13535 = n13460 & n13534 ;
  assign n14997 = n14996 ^ n13535 ;
  assign n13507 = n13498 ^ n13482 ;
  assign n13508 = n13482 ^ n13309 ;
  assign n13509 = n13508 ^ n13482 ;
  assign n13510 = n13507 & n13509 ;
  assign n13511 = n13510 ^ n13482 ;
  assign n13512 = ~n13144 & ~n13511 ;
  assign n14998 = n14997 ^ n13512 ;
  assign n14999 = n14998 ^ n11560 ;
  assign n14975 = n14974 ^ n13483 ;
  assign n14973 = n13472 ^ n13468 ;
  assign n14976 = n14975 ^ n14973 ;
  assign n14977 = n14973 ^ n13309 ;
  assign n14978 = n14977 ^ n14973 ;
  assign n14979 = n14976 & n14978 ;
  assign n14980 = n14979 ^ n14973 ;
  assign n14981 = ~n13144 & n14980 ;
  assign n15000 = n14999 ^ n14981 ;
  assign n14966 = n14965 ^ n13496 ;
  assign n14967 = n14966 ^ n14965 ;
  assign n14970 = ~n13309 & n14967 ;
  assign n14971 = n14970 ^ n14965 ;
  assign n14972 = n14958 & ~n14971 ;
  assign n15001 = n15000 ^ n14972 ;
  assign n15002 = n15001 ^ x109 ;
  assign n15003 = ~n14957 & ~n15002 ;
  assign n15004 = n15003 ^ n14957 ;
  assign n14277 = n14276 ^ n14275 ;
  assign n14314 = n14277 & ~n14311 ;
  assign n14315 = n14314 ^ n14276 ;
  assign n14316 = ~n14163 & n14315 ;
  assign n14687 = n14316 ^ n11858 ;
  assign n14685 = n14682 ^ n14358 ;
  assign n14657 = n14371 ^ n14335 ;
  assign n14658 = n14657 ^ n14276 ;
  assign n14664 = n14658 ^ n14324 ;
  assign n14655 = n14331 ^ n14326 ;
  assign n14656 = n14655 ^ n14338 ;
  assign n14659 = n14658 ^ n14656 ;
  assign n14660 = n14656 ^ n14163 ;
  assign n14661 = n14368 & n14660 ;
  assign n14662 = n14661 ^ n14163 ;
  assign n14663 = ~n14659 & n14662 ;
  assign n14665 = n14664 ^ n14663 ;
  assign n14686 = n14685 ^ n14665 ;
  assign n14688 = n14687 ^ n14686 ;
  assign n14676 = n14358 ^ n14219 ;
  assign n14677 = n14676 ^ n14320 ;
  assign n14674 = n14271 ^ n14270 ;
  assign n14675 = n14674 ^ n14218 ;
  assign n14678 = n14677 ^ n14675 ;
  assign n14679 = n14678 ^ n14368 ;
  assign n14680 = n14344 & n14679 ;
  assign n14681 = n14680 ^ n14368 ;
  assign n14683 = n14682 ^ n14344 ;
  assign n14684 = ~n14681 & ~n14683 ;
  assign n14689 = n14688 ^ n14684 ;
  assign n14666 = n14665 ^ n14319 ;
  assign n14667 = n14666 ^ n14325 ;
  assign n14668 = n14667 ^ n14665 ;
  assign n14669 = n14665 ^ n14311 ;
  assign n14670 = n14669 ^ n14665 ;
  assign n14671 = ~n14668 & n14670 ;
  assign n14672 = n14671 ^ n14665 ;
  assign n14673 = n14368 & n14672 ;
  assign n14690 = n14689 ^ n14673 ;
  assign n14654 = n14320 & n14653 ;
  assign n14691 = n14690 ^ n14654 ;
  assign n14652 = n14341 & n14651 ;
  assign n14692 = n14691 ^ n14652 ;
  assign n14644 = n14358 ^ n14317 ;
  assign n14645 = n14644 ^ n14358 ;
  assign n14646 = n14358 ^ n14311 ;
  assign n14647 = n14646 ^ n14358 ;
  assign n14648 = n14645 & ~n14647 ;
  assign n14649 = n14648 ^ n14358 ;
  assign n14650 = ~n14163 & ~n14649 ;
  assign n14693 = n14692 ^ n14650 ;
  assign n14694 = n14693 ^ x70 ;
  assign n13054 = n13053 ^ n12825 ;
  assign n13048 = n13010 ^ n12410 ;
  assign n13055 = n13054 ^ n13048 ;
  assign n14725 = n13055 ^ n13043 ;
  assign n14723 = n13038 ^ n12825 ;
  assign n13064 = n13053 ^ n13029 ;
  assign n14724 = n14723 ^ n13064 ;
  assign n14726 = n14725 ^ n14724 ;
  assign n14727 = n13056 & ~n14726 ;
  assign n14716 = n13064 ^ n13043 ;
  assign n14714 = n13024 & n13056 ;
  assign n14715 = n14714 ^ n14713 ;
  assign n14717 = n14716 ^ n14715 ;
  assign n14710 = n13035 ^ n13029 ;
  assign n14711 = n14710 ^ n13043 ;
  assign n14712 = n13058 & ~n14711 ;
  assign n14718 = n14717 ^ n14712 ;
  assign n14702 = n13064 ^ n13031 ;
  assign n14703 = n14702 ^ n13008 ;
  assign n14704 = n14703 ^ n14702 ;
  assign n14705 = n14702 ^ n13037 ;
  assign n14706 = n14705 ^ n14702 ;
  assign n14707 = ~n14704 & n14706 ;
  assign n14708 = n14707 ^ n14702 ;
  assign n14709 = ~n11520 & ~n14708 ;
  assign n14719 = n14718 ^ n14709 ;
  assign n14720 = n14719 ^ n13055 ;
  assign n13089 = ~n13008 & ~n13028 ;
  assign n13090 = n13089 ^ n13023 ;
  assign n13077 = n13076 ^ n13040 ;
  assign n13078 = n13077 ^ n13035 ;
  assign n13091 = n13090 ^ n13078 ;
  assign n13092 = n13091 ^ n13090 ;
  assign n13093 = n13090 ^ n11520 ;
  assign n13094 = n13093 ^ n13090 ;
  assign n13095 = ~n13092 & n13094 ;
  assign n13096 = n13095 ^ n13090 ;
  assign n13097 = n13047 & n13096 ;
  assign n13098 = n13097 ^ n13090 ;
  assign n14721 = n14720 ^ n13098 ;
  assign n14722 = n14721 ^ n11726 ;
  assign n14728 = n14727 ^ n14722 ;
  assign n14695 = n13054 ^ n13021 ;
  assign n14696 = n14695 ^ n13034 ;
  assign n14697 = n13034 ^ n11520 ;
  assign n14698 = n14697 ^ n13034 ;
  assign n14699 = n14696 & ~n14698 ;
  assign n14700 = n14699 ^ n13034 ;
  assign n14701 = n13008 & n14700 ;
  assign n14729 = n14728 ^ n14701 ;
  assign n14730 = n14729 ^ x110 ;
  assign n14731 = ~n14694 & n14730 ;
  assign n14098 = n13929 & n14074 ;
  assign n14776 = n14109 ^ n14098 ;
  assign n14777 = ~n13964 & n14776 ;
  assign n14075 = n14074 ^ n14070 ;
  assign n14076 = n13929 & n14075 ;
  assign n14077 = n14076 ^ n14074 ;
  assign n14078 = n13963 & n14077 ;
  assign n14068 = ~n13964 & n14067 ;
  assign n14079 = n14078 ^ n14068 ;
  assign n14773 = n14079 ^ n11775 ;
  assign n14153 = n14111 ^ n14104 ;
  assign n14154 = n13963 & ~n14153 ;
  assign n14155 = n14154 ^ n14104 ;
  assign n14752 = n14155 ^ n14074 ;
  assign n14771 = n14770 ^ n14752 ;
  assign n14744 = n14116 ^ n13929 ;
  assign n14772 = n14771 ^ n14744 ;
  assign n14774 = n14773 ^ n14772 ;
  assign n14761 = n13963 & n14756 ;
  assign n14753 = n14752 ^ n14094 ;
  assign n14762 = n14761 ^ n14753 ;
  assign n14763 = ~n13929 & ~n14762 ;
  assign n14775 = n14774 ^ n14763 ;
  assign n14778 = n14777 ^ n14775 ;
  assign n14749 = n14733 ^ n13929 ;
  assign n14750 = n14097 ^ n14067 ;
  assign n14751 = n14749 & n14750 ;
  assign n14779 = n14778 ^ n14751 ;
  assign n14745 = n14744 ^ n14116 ;
  assign n14746 = n14119 & n14745 ;
  assign n14747 = n14746 ^ n14116 ;
  assign n14748 = n13963 & ~n14747 ;
  assign n14780 = n14779 ^ n14748 ;
  assign n14145 = n14088 ^ n13963 ;
  assign n14734 = n14733 ^ n13964 ;
  assign n14735 = n14734 ^ n14088 ;
  assign n14736 = n14735 ^ n13964 ;
  assign n14739 = ~n14145 & n14736 ;
  assign n14740 = n14739 ^ n13964 ;
  assign n14741 = ~n14095 & n14740 ;
  assign n14781 = n14780 ^ n14741 ;
  assign n14782 = n14781 ^ x68 ;
  assign n14783 = n13852 ^ n13577 ;
  assign n14784 = n14783 ^ n13576 ;
  assign n14785 = n13888 ^ n13839 ;
  assign n14798 = n13810 ^ n13805 ;
  assign n14799 = n14798 ^ n13836 ;
  assign n14800 = n14799 ^ n13824 ;
  assign n14801 = ~n13576 & ~n14800 ;
  assign n14802 = n14801 ^ n13836 ;
  assign n14803 = ~n13577 & n14802 ;
  assign n14796 = n13852 & n13886 ;
  assign n14786 = n13819 ^ n13577 ;
  assign n14791 = n13819 ^ n13809 ;
  assign n14792 = n14791 ^ n13841 ;
  assign n14787 = n13841 ^ n13805 ;
  assign n14788 = n14787 ^ n13819 ;
  assign n14789 = n14788 ^ n13839 ;
  assign n14790 = n13576 & n14789 ;
  assign n14793 = n14792 ^ n14790 ;
  assign n14794 = n14786 & ~n14793 ;
  assign n14795 = n14794 ^ n13577 ;
  assign n14797 = n14796 ^ n14795 ;
  assign n14804 = n14803 ^ n14797 ;
  assign n14805 = ~n13850 & ~n14804 ;
  assign n14806 = ~n14785 & n14805 ;
  assign n14807 = ~n14784 & n14806 ;
  assign n14808 = n14807 ^ n14805 ;
  assign n14809 = n13829 ^ n13578 ;
  assign n14810 = n14809 ^ n13829 ;
  assign n14811 = n13576 & n13825 ;
  assign n14812 = n14811 ^ n13829 ;
  assign n14813 = n14810 & ~n14812 ;
  assign n14814 = n14813 ^ n13829 ;
  assign n14815 = n14808 & ~n14814 ;
  assign n14816 = n14815 ^ n14808 ;
  assign n14823 = n14816 & ~n14822 ;
  assign n14824 = ~n13854 & n14823 ;
  assign n13858 = n13837 ^ n13835 ;
  assign n14826 = n13858 & n14783 ;
  assign n14827 = n14824 & n14826 ;
  assign n14825 = n14824 ^ n11813 ;
  assign n14828 = n14827 ^ n14825 ;
  assign n14829 = n14828 ^ x85 ;
  assign n14830 = ~n14782 & ~n14829 ;
  assign n14832 = n14830 ^ n14829 ;
  assign n14833 = n14832 ^ n14782 ;
  assign n15034 = n14731 & ~n14833 ;
  assign n15035 = n15034 ^ n14731 ;
  assign n14732 = n14731 ^ n14694 ;
  assign n15018 = n14732 ^ n14730 ;
  assign n15019 = n14830 & n15018 ;
  assign n15013 = n14830 ^ n14782 ;
  assign n15014 = ~n14732 & ~n15013 ;
  assign n15015 = n15014 ^ n14732 ;
  assign n14834 = ~n14732 & ~n14833 ;
  assign n14831 = ~n14732 & n14830 ;
  assign n14835 = n14834 ^ n14831 ;
  assign n15016 = n15015 ^ n14835 ;
  assign n15020 = n15019 ^ n15016 ;
  assign n15021 = n15020 ^ n14834 ;
  assign n15022 = n15021 ^ n15014 ;
  assign n15011 = n14829 ^ n14694 ;
  assign n15012 = ~n14730 & n15011 ;
  assign n15017 = n15016 ^ n15012 ;
  assign n15023 = n15022 ^ n15017 ;
  assign n15024 = n15023 ^ n15016 ;
  assign n15008 = n14731 ^ n14730 ;
  assign n15009 = ~n14832 & n15008 ;
  assign n15010 = n15009 ^ n14832 ;
  assign n15025 = n15024 ^ n15010 ;
  assign n15007 = n14731 & n14830 ;
  assign n15026 = n15025 ^ n15007 ;
  assign n15036 = n15035 ^ n15026 ;
  assign n16970 = ~n15004 & n15036 ;
  assign n15005 = n15004 ^ n15002 ;
  assign n15044 = n15008 & ~n15013 ;
  assign n16967 = n15044 ^ n15025 ;
  assign n16968 = ~n15005 & n16967 ;
  assign n16324 = n15002 ^ n14957 ;
  assign n15050 = n15023 ^ n15020 ;
  assign n15051 = n15050 ^ n14831 ;
  assign n15052 = n15051 ^ n15025 ;
  assign n15048 = n15009 ^ n15007 ;
  assign n15049 = n15048 ^ n14829 ;
  assign n15053 = n15052 ^ n15049 ;
  assign n15054 = n15053 ^ n15008 ;
  assign n15045 = n15044 ^ n15009 ;
  assign n15055 = n15054 ^ n15045 ;
  assign n15056 = n15055 ^ n15034 ;
  assign n15057 = n15056 ^ n14833 ;
  assign n15058 = n15057 ^ n15022 ;
  assign n15059 = n15058 ^ n15019 ;
  assign n15047 = n15016 ^ n15014 ;
  assign n15060 = n15059 ^ n15047 ;
  assign n16952 = n15060 ^ n15053 ;
  assign n16954 = n16952 ^ n15024 ;
  assign n16955 = n16954 ^ n15053 ;
  assign n16956 = n16954 ^ n15002 ;
  assign n16957 = n16956 ^ n16954 ;
  assign n16958 = n16955 & n16957 ;
  assign n16959 = n16958 ^ n16954 ;
  assign n16960 = n16324 & n16959 ;
  assign n16961 = n16960 ^ n16952 ;
  assign n16943 = n15018 ^ n14831 ;
  assign n16944 = n16943 ^ n15059 ;
  assign n16945 = ~n14957 & n16944 ;
  assign n16946 = n16945 ^ n15022 ;
  assign n16962 = n16961 ^ n16946 ;
  assign n15061 = n15060 ^ n15024 ;
  assign n15062 = n15061 ^ n15018 ;
  assign n15063 = n15062 ^ n15020 ;
  assign n15070 = n15005 ^ n14957 ;
  assign n15097 = ~n15063 & ~n15070 ;
  assign n16963 = n16962 ^ n15097 ;
  assign n16340 = n15044 ^ n15034 ;
  assign n16341 = n16340 ^ n15048 ;
  assign n16342 = n15048 ^ n15002 ;
  assign n16343 = n16342 ^ n15048 ;
  assign n16344 = n16341 & ~n16343 ;
  assign n16345 = n16344 ^ n15048 ;
  assign n16346 = ~n14957 & n16345 ;
  assign n16964 = n16963 ^ n16346 ;
  assign n16965 = n16964 ^ n14217 ;
  assign n16948 = n15060 ^ n15055 ;
  assign n16947 = n16946 ^ n15012 ;
  assign n16949 = n16948 ^ n16947 ;
  assign n16939 = n14832 ^ n14731 ;
  assign n16940 = n16939 ^ n15022 ;
  assign n16941 = n16940 ^ n15055 ;
  assign n16942 = n14957 & n16941 ;
  assign n16950 = n16949 ^ n16942 ;
  assign n16951 = ~n15002 & n16950 ;
  assign n16966 = n16965 ^ n16951 ;
  assign n16969 = n16968 ^ n16966 ;
  assign n16971 = n16970 ^ n16969 ;
  assign n16972 = n16971 ^ x82 ;
  assign n16973 = n16938 & n16972 ;
  assign n16974 = n16973 ^ n16938 ;
  assign n16975 = n16974 ^ n16972 ;
  assign n13099 = n13098 ^ n11972 ;
  assign n13014 = n13013 ^ n13010 ;
  assign n13015 = n13008 & n13014 ;
  assign n12826 = ~n11520 & n12825 ;
  assign n13016 = n13015 ^ n12826 ;
  assign n13062 = n13042 ^ n13039 ;
  assign n13059 = n13055 & n13058 ;
  assign n13067 = n13062 ^ n13059 ;
  assign n13061 = n13034 ^ n12825 ;
  assign n13063 = n13062 ^ n13061 ;
  assign n13065 = n13064 ^ n13063 ;
  assign n13066 = ~n13008 & n13065 ;
  assign n13068 = n13067 ^ n13066 ;
  assign n13060 = n13059 ^ n13037 ;
  assign n13069 = n13068 ^ n13060 ;
  assign n13070 = n13069 ^ n13037 ;
  assign n13071 = n13070 ^ n13069 ;
  assign n13072 = n13069 ^ n13008 ;
  assign n13073 = n13072 ^ n13069 ;
  assign n13079 = n13078 ^ n13069 ;
  assign n13080 = n13079 ^ n13069 ;
  assign n13081 = ~n13073 & ~n13080 ;
  assign n13082 = ~n13071 & n13081 ;
  assign n13083 = n13082 ^ n13071 ;
  assign n13084 = n13083 ^ n13070 ;
  assign n13085 = ~n13047 & ~n13084 ;
  assign n13086 = n13085 ^ n13068 ;
  assign n13045 = n13044 ^ n13026 ;
  assign n13046 = n13017 & ~n13045 ;
  assign n13087 = n13086 ^ n13046 ;
  assign n13088 = ~n13016 & n13087 ;
  assign n13100 = n13099 ^ n13088 ;
  assign n13101 = n13100 ^ x106 ;
  assign n13542 = n13467 ^ n13463 ;
  assign n13544 = n13543 ^ n13542 ;
  assign n13545 = n13311 & n13544 ;
  assign n13540 = ~n13489 & n13534 ;
  assign n13518 = n13476 ^ n13469 ;
  assign n13519 = n13469 ^ n13144 ;
  assign n13520 = n13519 ^ n13469 ;
  assign n13521 = n13518 & n13520 ;
  assign n13522 = n13521 ^ n13469 ;
  assign n13523 = n13309 & ~n13522 ;
  assign n13524 = n13523 ^ n13470 ;
  assign n13532 = n13531 ^ n13524 ;
  assign n13513 = n13479 ^ n13455 ;
  assign n13514 = n13310 & ~n13513 ;
  assign n13515 = n13421 ^ n13380 ;
  assign n13516 = n13515 ^ n13479 ;
  assign n13517 = n13514 & n13516 ;
  assign n13533 = n13532 ^ n13517 ;
  assign n13536 = n13535 ^ n13533 ;
  assign n13537 = n13536 ^ n13512 ;
  assign n13538 = n13537 ^ n12761 ;
  assign n13471 = n13470 ^ n13312 ;
  assign n13500 = n13499 ^ n13494 ;
  assign n13501 = n13500 ^ n13310 ;
  assign n13504 = ~n13312 & n13501 ;
  assign n13505 = n13504 ^ n13310 ;
  assign n13506 = n13471 & ~n13505 ;
  assign n13539 = n13538 ^ n13506 ;
  assign n13541 = n13540 ^ n13539 ;
  assign n13546 = n13545 ^ n13541 ;
  assign n13547 = n13546 ^ x97 ;
  assign n13548 = n13101 & n13547 ;
  assign n13549 = n13548 ^ n13101 ;
  assign n13871 = n13829 ^ n13814 ;
  assign n13872 = n13871 ^ n13809 ;
  assign n13873 = n13872 ^ n13832 ;
  assign n13874 = n13832 ^ n13577 ;
  assign n13875 = n13874 ^ n13832 ;
  assign n13876 = ~n13873 & ~n13875 ;
  assign n13877 = n13876 ^ n13832 ;
  assign n13878 = ~n13576 & n13877 ;
  assign n13879 = n13878 ^ n13827 ;
  assign n13870 = n13578 & n13821 ;
  assign n13880 = n13879 ^ n13870 ;
  assign n13866 = n13828 ^ n13827 ;
  assign n13867 = n13865 & n13866 ;
  assign n13868 = n13867 ^ n13827 ;
  assign n13869 = n13576 & ~n13868 ;
  assign n13881 = n13880 ^ n13869 ;
  assign n13855 = n13842 ^ n13824 ;
  assign n13882 = n13881 ^ n13855 ;
  assign n13856 = n13855 ^ n13576 ;
  assign n13857 = n13856 ^ n13855 ;
  assign n13861 = n13857 & n13858 ;
  assign n13862 = n13861 ^ n13855 ;
  assign n13863 = n13578 & n13862 ;
  assign n13883 = n13882 ^ n13863 ;
  assign n13884 = ~n13854 & n13883 ;
  assign n13893 = n13884 & ~n13892 ;
  assign n13851 = n13850 ^ n12865 ;
  assign n13894 = n13893 ^ n13851 ;
  assign n13895 = n13894 ^ x123 ;
  assign n14099 = n14098 ^ n14074 ;
  assign n14100 = n14099 ^ n14097 ;
  assign n14101 = n14100 ^ n14077 ;
  assign n14102 = n13964 & n14101 ;
  assign n14103 = n14102 ^ n14097 ;
  assign n14128 = n14118 ^ n14093 ;
  assign n14129 = n14128 ^ n14088 ;
  assign n14132 = n14095 ^ n13929 ;
  assign n14133 = n14132 ^ n14095 ;
  assign n14134 = ~n14129 & n14133 ;
  assign n14135 = n14134 ^ n14095 ;
  assign n14136 = ~n13963 & n14135 ;
  assign n14137 = n14136 ^ n14127 ;
  assign n14112 = n14111 ^ n14080 ;
  assign n14120 = n14119 ^ n14112 ;
  assign n14121 = ~n13929 & ~n14120 ;
  assign n14138 = n14137 ^ n14121 ;
  assign n14105 = n14104 ^ n14083 ;
  assign n14106 = n14105 ^ n14093 ;
  assign n14139 = n14138 ^ n14106 ;
  assign n14140 = n14139 ^ n14136 ;
  assign n14141 = ~n13964 & n14140 ;
  assign n14142 = n14141 ^ n14138 ;
  assign n14146 = n14145 ^ n14088 ;
  assign n14147 = n14089 & n14146 ;
  assign n14148 = n14147 ^ n14088 ;
  assign n14149 = ~n13929 & n14148 ;
  assign n14150 = ~n14142 & ~n14149 ;
  assign n14151 = ~n14103 & n14150 ;
  assign n14152 = ~n14079 & n14151 ;
  assign n14158 = n14152 ^ n12894 ;
  assign n14156 = n13929 & n14155 ;
  assign n14157 = n14152 & n14156 ;
  assign n14159 = n14158 ^ n14157 ;
  assign n14160 = n14159 ^ x80 ;
  assign n14161 = ~n13895 & n14160 ;
  assign n14162 = n14161 ^ n13895 ;
  assign n14362 = n14331 ^ n14325 ;
  assign n14360 = n14344 ^ n14330 ;
  assign n14361 = n14360 ^ n14341 ;
  assign n14363 = n14362 ^ n14361 ;
  assign n14364 = n14311 & n14363 ;
  assign n14365 = n14364 ^ n14361 ;
  assign n14375 = n14365 ^ n14358 ;
  assign n14373 = n14372 ^ n14321 ;
  assign n14374 = ~n14311 & n14373 ;
  assign n14376 = n14375 ^ n14374 ;
  assign n14369 = n14333 ^ n14324 ;
  assign n14370 = ~n14163 & n14369 ;
  assign n14377 = n14376 ^ n14370 ;
  assign n14378 = n14368 & n14377 ;
  assign n14359 = n14358 ^ n14356 ;
  assign n14366 = n14365 ^ n14359 ;
  assign n14367 = n14366 ^ n14316 ;
  assign n14379 = n14378 ^ n14367 ;
  assign n14380 = n14379 ^ n14335 ;
  assign n14381 = n14380 ^ n12693 ;
  assign n14382 = n14381 ^ x120 ;
  assign n14459 = n13379 ^ x108 ;
  assign n14383 = n13575 ^ x84 ;
  assign n14410 = n12598 ^ n12544 ;
  assign n14411 = ~n12457 & ~n14410 ;
  assign n14387 = ~n12457 & n12570 ;
  assign n14388 = n14387 ^ n12537 ;
  assign n14409 = n14388 ^ n12542 ;
  assign n14412 = n14411 ^ n14409 ;
  assign n14413 = n12458 & n14412 ;
  assign n14407 = n12460 & n12530 ;
  assign n14393 = n14392 ^ n12599 ;
  assign n14390 = n12565 ^ n12553 ;
  assign n14391 = n14390 ^ n12563 ;
  assign n14394 = n14393 ^ n14391 ;
  assign n14395 = n12458 & ~n14394 ;
  assign n14396 = n14395 ^ n14393 ;
  assign n14398 = n14396 ^ n12551 ;
  assign n14399 = n14398 ^ n12564 ;
  assign n14400 = n14399 ^ n14396 ;
  assign n14402 = n14401 ^ n14400 ;
  assign n14403 = n12458 & n14402 ;
  assign n14404 = n14403 ^ n14398 ;
  assign n14405 = n12457 & n14404 ;
  assign n14389 = n14388 ^ n12611 ;
  assign n14397 = n14396 ^ n14389 ;
  assign n14406 = n14405 ^ n14397 ;
  assign n14408 = n14407 ^ n14406 ;
  assign n14414 = n14413 ^ n14408 ;
  assign n14415 = n14414 ^ n14384 ;
  assign n14385 = n14384 ^ n14004 ;
  assign n14386 = n12457 & n14385 ;
  assign n14416 = n14415 ^ n14386 ;
  assign n14417 = ~n12576 & ~n13996 ;
  assign n14418 = ~n14416 & n14417 ;
  assign n14419 = n14418 ^ n12088 ;
  assign n14420 = n14419 ^ x101 ;
  assign n14421 = ~n14383 & n14420 ;
  assign n14422 = n14421 ^ n14420 ;
  assign n14441 = n12315 & ~n12399 ;
  assign n14437 = n12337 ^ n12235 ;
  assign n14438 = n14437 ^ n12341 ;
  assign n14439 = n12000 & ~n14438 ;
  assign n14433 = n13402 ^ n12374 ;
  assign n14428 = n12344 ^ n12311 ;
  assign n14429 = n14428 ^ n12321 ;
  assign n14430 = ~n12399 & ~n14429 ;
  assign n14431 = n14430 ^ n12312 ;
  assign n14432 = ~n11973 & ~n14431 ;
  assign n14434 = n14433 ^ n14432 ;
  assign n14427 = ~n12342 & n12359 ;
  assign n14435 = n14434 ^ n14427 ;
  assign n14423 = n12343 ^ n12327 ;
  assign n14424 = n14423 ^ n12316 ;
  assign n14425 = n14424 ^ n12334 ;
  assign n14426 = n11999 & ~n14425 ;
  assign n14436 = n14435 ^ n14426 ;
  assign n14440 = n14439 ^ n14436 ;
  assign n14442 = n14441 ^ n14440 ;
  assign n14443 = ~n14027 & ~n14442 ;
  assign n14444 = n14443 ^ n12111 ;
  assign n14445 = n14444 ^ x86 ;
  assign n14446 = n13308 ^ x126 ;
  assign n14447 = ~n14445 & ~n14446 ;
  assign n14449 = n14447 ^ n14446 ;
  assign n14482 = n14449 ^ n14445 ;
  assign n14483 = n14422 & ~n14482 ;
  assign n14506 = n14483 ^ n14482 ;
  assign n14454 = n14422 ^ n14383 ;
  assign n14496 = n14454 & ~n14482 ;
  assign n14495 = n14421 & ~n14482 ;
  assign n14497 = n14496 ^ n14495 ;
  assign n14507 = n14506 ^ n14497 ;
  assign n14450 = n14421 ^ n14383 ;
  assign n14522 = n14507 ^ n14450 ;
  assign n14465 = n14447 & ~n14450 ;
  assign n14451 = ~n14449 & ~n14450 ;
  assign n14521 = n14465 ^ n14451 ;
  assign n14523 = n14522 ^ n14521 ;
  assign n14524 = n14523 ^ n14497 ;
  assign n14531 = n14524 ^ n14446 ;
  assign n14504 = n14483 ^ n14422 ;
  assign n14455 = ~n14449 & n14454 ;
  assign n14453 = n14421 & ~n14449 ;
  assign n14456 = n14455 ^ n14453 ;
  assign n14452 = n14451 ^ n14449 ;
  assign n14457 = n14456 ^ n14452 ;
  assign n14448 = n14422 & n14447 ;
  assign n14458 = n14457 ^ n14448 ;
  assign n14505 = n14504 ^ n14458 ;
  assign n14508 = n14507 ^ n14505 ;
  assign n14500 = n14482 ^ n14446 ;
  assign n14501 = n14421 & ~n14500 ;
  assign n14502 = n14501 ^ n14483 ;
  assign n14530 = n14508 ^ n14502 ;
  assign n14532 = n14531 ^ n14530 ;
  assign n14533 = n14459 & n14532 ;
  assign n14460 = n13802 ^ x125 ;
  assign n14461 = ~n14459 & n14460 ;
  assign n14515 = n14508 ^ n14501 ;
  assign n14516 = n14515 ^ n14496 ;
  assign n14517 = n14461 & n14516 ;
  assign n14464 = n14461 ^ n14459 ;
  assign n14518 = n14517 ^ n14464 ;
  assign n14525 = n14524 ^ n14505 ;
  assign n14519 = n14507 ^ n14501 ;
  assign n14520 = n14461 & ~n14519 ;
  assign n14526 = n14525 ^ n14520 ;
  assign n14527 = ~n14518 & ~n14526 ;
  assign n14503 = n14502 ^ n14453 ;
  assign n14509 = n14508 ^ n14503 ;
  assign n14498 = n14497 ^ n14455 ;
  assign n14470 = n14421 & n14447 ;
  assign n14479 = n14470 ^ n14448 ;
  assign n14480 = n14479 ^ n14465 ;
  assign n14499 = n14498 ^ n14480 ;
  assign n14510 = n14509 ^ n14499 ;
  assign n14511 = n14460 & n14510 ;
  assign n14512 = n14511 ^ n14509 ;
  assign n14513 = n14459 & n14512 ;
  assign n14463 = n14460 ^ n14459 ;
  assign n14485 = n14483 ^ n14453 ;
  assign n14481 = n14480 ^ n14447 ;
  assign n14484 = n14483 ^ n14481 ;
  assign n14486 = n14485 ^ n14484 ;
  assign n14487 = n14485 ^ n14460 ;
  assign n14488 = n14487 ^ n14485 ;
  assign n14489 = n14486 & ~n14488 ;
  assign n14490 = n14489 ^ n14485 ;
  assign n14491 = n14463 & n14490 ;
  assign n14492 = n14491 ^ n14483 ;
  assign n14466 = n14465 ^ n14455 ;
  assign n14467 = ~n14464 & n14466 ;
  assign n14468 = n14467 ^ n14451 ;
  assign n14469 = n14468 ^ n14467 ;
  assign n14471 = n14470 ^ n14469 ;
  assign n14472 = n14471 ^ n14469 ;
  assign n14473 = n14469 ^ n14460 ;
  assign n14474 = n14473 ^ n14469 ;
  assign n14475 = n14472 & ~n14474 ;
  assign n14476 = n14475 ^ n14469 ;
  assign n14477 = ~n14463 & n14476 ;
  assign n14478 = n14477 ^ n14468 ;
  assign n14493 = n14492 ^ n14478 ;
  assign n14494 = n14493 ^ n12202 ;
  assign n14514 = n14513 ^ n14494 ;
  assign n14528 = n14527 ^ n14514 ;
  assign n14462 = ~n14458 & n14461 ;
  assign n14529 = n14528 ^ n14462 ;
  assign n14534 = n14533 ^ n14529 ;
  assign n14535 = n14534 ^ x82 ;
  assign n14537 = n14382 & n14535 ;
  assign n14536 = n14535 ^ n14382 ;
  assign n14538 = n14537 ^ n14536 ;
  assign n14539 = n14538 ^ n14535 ;
  assign n14540 = ~n14162 & n14539 ;
  assign n14541 = n13549 & n14540 ;
  assign n16877 = n14541 ^ n14185 ;
  assign n14561 = n13549 & n14161 ;
  assign n14557 = n13548 & n14161 ;
  assign n14602 = n14561 ^ n14557 ;
  assign n14542 = n13548 ^ n13547 ;
  assign n14575 = n14161 & n14542 ;
  assign n14601 = n14575 ^ n14161 ;
  assign n14603 = n14602 ^ n14601 ;
  assign n14544 = n14162 ^ n14160 ;
  assign n14545 = n14544 ^ n13895 ;
  assign n14577 = n14542 & n14545 ;
  assign n14543 = ~n14162 & n14542 ;
  assign n14578 = n14577 ^ n14543 ;
  assign n14576 = n14575 ^ n14542 ;
  assign n14579 = n14578 ^ n14576 ;
  assign n14604 = n14603 ^ n14579 ;
  assign n14581 = n14542 ^ n13101 ;
  assign n14582 = n14545 & ~n14581 ;
  assign n14605 = n14604 ^ n14582 ;
  assign n14593 = ~n14162 & ~n14581 ;
  assign n14594 = n14593 ^ n14579 ;
  assign n14600 = n14594 ^ n14581 ;
  assign n14606 = n14605 ^ n14600 ;
  assign n14609 = ~n14535 & ~n14606 ;
  assign n14595 = n14594 ^ n14582 ;
  assign n14596 = n14535 & n14595 ;
  assign n14597 = n14596 ^ n14582 ;
  assign n14610 = n14609 ^ n14597 ;
  assign n14611 = n14382 & n14610 ;
  assign n14612 = n14611 ^ n14597 ;
  assign n14632 = n14593 ^ n14577 ;
  assign n14633 = n14632 ^ n14575 ;
  assign n16867 = n14633 ^ n14579 ;
  assign n14547 = n13548 & n14544 ;
  assign n14562 = n14561 ^ n14547 ;
  assign n16865 = n14575 ^ n14562 ;
  assign n14565 = n13549 & n14544 ;
  assign n14555 = n13548 & ~n14162 ;
  assign n16864 = n14565 ^ n14555 ;
  assign n16866 = n16865 ^ n16864 ;
  assign n16868 = n16867 ^ n16866 ;
  assign n16869 = n16866 ^ n14535 ;
  assign n16870 = n16869 ^ n16866 ;
  assign n16871 = n16868 & ~n16870 ;
  assign n16872 = n16871 ^ n16866 ;
  assign n16873 = n14382 & n16872 ;
  assign n16850 = n14606 ^ n14602 ;
  assign n14546 = n13549 & n14545 ;
  assign n14556 = n14555 ^ n14546 ;
  assign n14558 = n14557 ^ n14556 ;
  assign n14559 = n14558 ^ n13548 ;
  assign n14548 = n14547 ^ n14546 ;
  assign n14560 = n14559 ^ n14548 ;
  assign n14615 = n14565 ^ n14560 ;
  assign n16851 = n16850 ^ n14615 ;
  assign n14566 = n14565 ^ n14558 ;
  assign n14563 = n14562 ^ n14560 ;
  assign n14564 = n14563 ^ n13101 ;
  assign n14567 = n14566 ^ n14564 ;
  assign n16847 = n14567 ^ n14557 ;
  assign n16848 = n16847 ^ n14606 ;
  assign n16849 = n16848 ^ n14547 ;
  assign n16852 = n16851 ^ n16849 ;
  assign n16853 = n14535 & n16852 ;
  assign n16854 = n16853 ^ n16849 ;
  assign n16855 = ~n14382 & ~n16854 ;
  assign n16856 = n16855 ^ n14582 ;
  assign n16840 = n14582 ^ n14382 ;
  assign n16841 = n16840 ^ n14582 ;
  assign n16842 = n14582 ^ n14562 ;
  assign n16843 = n16842 ^ n14582 ;
  assign n16844 = n16841 & n16843 ;
  assign n16845 = n16844 ^ n14582 ;
  assign n16846 = ~n14535 & n16845 ;
  assign n16857 = n16856 ^ n16846 ;
  assign n16859 = ~n14536 & n14578 ;
  assign n16860 = ~n16857 & n16859 ;
  assign n16861 = n16860 ^ n16857 ;
  assign n16874 = n16873 ^ n16861 ;
  assign n16858 = n16857 ^ n14538 ;
  assign n16863 = n14603 & ~n16858 ;
  assign n16875 = n16874 ^ n16863 ;
  assign n16876 = ~n14612 & ~n16875 ;
  assign n16878 = n16877 ^ n16876 ;
  assign n16879 = n16878 ^ x96 ;
  assign n16395 = n15194 ^ x102 ;
  assign n16396 = n14729 ^ x116 ;
  assign n16518 = n16395 & ~n16396 ;
  assign n16519 = n16518 ^ n16395 ;
  assign n16520 = n16519 ^ n16396 ;
  assign n16397 = n14956 ^ x117 ;
  assign n15502 = n15279 ^ n15196 ;
  assign n15503 = n15502 ^ n15279 ;
  assign n15504 = n15280 & n15503 ;
  assign n15505 = n15504 ^ n15279 ;
  assign n15506 = n15197 & n15505 ;
  assign n16420 = n15199 & n15287 ;
  assign n16412 = n15304 ^ n15198 ;
  assign n16413 = n16412 ^ n15316 ;
  assign n16414 = n16413 ^ n15326 ;
  assign n16415 = ~n15346 & ~n16414 ;
  assign n16416 = n16415 ^ n15198 ;
  assign n16417 = n15346 ^ n15318 ;
  assign n16418 = ~n16416 & ~n16417 ;
  assign n15729 = n15288 ^ n15281 ;
  assign n16408 = n15729 ^ n15275 ;
  assign n16409 = n15198 & n16408 ;
  assign n15759 = n15316 ^ n15282 ;
  assign n15760 = n15347 & ~n15759 ;
  assign n15761 = n15760 ^ n15344 ;
  assign n16405 = n15761 ^ n15360 ;
  assign n16406 = n16405 ^ n15324 ;
  assign n16398 = n15284 ^ n15278 ;
  assign n16399 = n16398 ^ n15314 ;
  assign n16400 = n15314 ^ n15197 ;
  assign n16401 = n16400 ^ n15314 ;
  assign n16402 = n16399 & n16401 ;
  assign n16403 = n16402 ^ n15314 ;
  assign n16404 = n15286 & ~n16403 ;
  assign n16407 = n16406 ^ n16404 ;
  assign n16410 = n16409 ^ n16407 ;
  assign n16411 = n16410 ^ n15318 ;
  assign n16419 = n16418 ^ n16411 ;
  assign n16421 = n16420 ^ n16419 ;
  assign n16422 = ~n15373 & ~n16421 ;
  assign n16423 = ~n15506 & n16422 ;
  assign n15751 = n15280 ^ n15230 ;
  assign n15752 = n15199 & n15751 ;
  assign n15755 = ~n15308 & n15347 ;
  assign n15756 = n15755 ^ n15365 ;
  assign n16424 = ~n15752 & ~n15756 ;
  assign n16425 = n16423 & n16424 ;
  assign n16426 = n16425 ^ n13699 ;
  assign n16427 = n16426 ^ x84 ;
  assign n16428 = n16397 & ~n16427 ;
  assign n16431 = n15138 ^ x77 ;
  assign n15817 = n14464 ^ n14460 ;
  assign n16450 = n14532 ^ n14505 ;
  assign n16451 = n16450 ^ n14465 ;
  assign n16452 = n15817 & ~n16451 ;
  assign n16445 = n14495 ^ n14465 ;
  assign n16446 = n16445 ^ n14505 ;
  assign n15769 = n14532 ^ n14507 ;
  assign n16436 = n15769 ^ n14483 ;
  assign n16435 = n14496 ^ n14480 ;
  assign n16437 = n16436 ^ n16435 ;
  assign n16433 = n14523 ^ n14505 ;
  assign n16434 = n16433 ^ n14451 ;
  assign n16438 = n16437 ^ n16434 ;
  assign n16439 = n14460 & n16438 ;
  assign n16440 = n16439 ^ n16437 ;
  assign n16447 = n16446 ^ n16440 ;
  assign n16448 = n14459 & n16447 ;
  assign n16013 = n14481 ^ n14470 ;
  assign n16014 = n14470 ^ n14460 ;
  assign n16015 = n16014 ^ n14470 ;
  assign n16016 = n16013 & n16015 ;
  assign n16017 = n16016 ^ n14470 ;
  assign n16018 = n14463 & n16017 ;
  assign n15778 = n14457 ^ n14456 ;
  assign n15777 = n14481 ^ n14456 ;
  assign n15779 = n15778 ^ n15777 ;
  assign n15780 = n15778 ^ n14460 ;
  assign n15781 = n15780 ^ n15778 ;
  assign n15782 = ~n15779 & n15781 ;
  assign n15783 = n15782 ^ n15778 ;
  assign n15784 = ~n14463 & ~n15783 ;
  assign n15785 = n15784 ^ n14456 ;
  assign n16432 = n16018 ^ n15785 ;
  assign n16441 = n16440 ^ n16432 ;
  assign n16033 = n14460 & n14530 ;
  assign n16034 = n16033 ^ n14508 ;
  assign n16037 = n16034 ^ n14456 ;
  assign n16038 = n16037 ^ n16034 ;
  assign n16039 = n14460 & n16038 ;
  assign n16040 = n16039 ^ n16034 ;
  assign n16041 = ~n14463 & n16040 ;
  assign n16042 = n16041 ^ n16034 ;
  assign n16442 = n16441 ^ n16042 ;
  assign n15825 = n15769 ^ n14523 ;
  assign n15826 = n14523 ^ n14460 ;
  assign n15827 = n15826 ^ n14523 ;
  assign n15828 = ~n15825 & n15827 ;
  assign n15829 = n15828 ^ n14523 ;
  assign n15830 = n14459 & n15829 ;
  assign n16443 = n16442 ^ n15830 ;
  assign n16444 = n16443 ^ n13669 ;
  assign n16449 = n16448 ^ n16444 ;
  assign n16453 = n16452 ^ n16449 ;
  assign n16454 = n16453 ^ x67 ;
  assign n16455 = ~n16431 & n16454 ;
  assign n16458 = n16455 ^ n16454 ;
  assign n16462 = n16458 ^ n16431 ;
  assign n16466 = n16462 ^ n16454 ;
  assign n16478 = n16428 & ~n16466 ;
  assign n16429 = n16428 ^ n16397 ;
  assign n16430 = n16429 ^ n16427 ;
  assign n16463 = n16430 ^ n16397 ;
  assign n16472 = n16455 & ~n16463 ;
  assign n16533 = n16478 ^ n16472 ;
  assign n16534 = n16520 & n16533 ;
  assign n16474 = n16458 & ~n16463 ;
  assign n16459 = n16428 & n16458 ;
  assign n16485 = n16474 ^ n16459 ;
  assign n16526 = n16485 ^ n16474 ;
  assign n16527 = n16526 ^ n16474 ;
  assign n16528 = n16474 ^ n16395 ;
  assign n16529 = n16528 ^ n16474 ;
  assign n16530 = n16527 & ~n16529 ;
  assign n16531 = n16530 ^ n16474 ;
  assign n16532 = ~n16396 & n16531 ;
  assign n16535 = n16534 ^ n16532 ;
  assign n16464 = n16462 & ~n16463 ;
  assign n16475 = n16474 ^ n16464 ;
  assign n16473 = n16472 ^ n16463 ;
  assign n16476 = n16475 ^ n16473 ;
  assign n16467 = n16429 & ~n16466 ;
  assign n16477 = n16476 ^ n16467 ;
  assign n16479 = n16478 ^ n16477 ;
  assign n16480 = n16479 ^ n16466 ;
  assign n16880 = n16480 ^ n16396 ;
  assign n16881 = n16880 ^ n16480 ;
  assign n16469 = n16430 & n16462 ;
  assign n16481 = n16480 ^ n16469 ;
  assign n16882 = n16481 ^ n16480 ;
  assign n16883 = ~n16881 & n16882 ;
  assign n16884 = n16883 ^ n16480 ;
  assign n16885 = ~n16395 & n16884 ;
  assign n16886 = n16885 ^ n16480 ;
  assign n16887 = ~n16535 & ~n16886 ;
  assign n16456 = n16430 & n16455 ;
  assign n16888 = n16456 & n16520 ;
  assign n16900 = n16479 ^ n16456 ;
  assign n16482 = n16481 ^ n16430 ;
  assign n16483 = n16482 ^ n16456 ;
  assign n16484 = n16483 ^ n16458 ;
  assign n16486 = n16485 ^ n16484 ;
  assign n16487 = n16486 ^ n16469 ;
  assign n16471 = n16429 & n16462 ;
  assign n16488 = n16487 ^ n16471 ;
  assign n16489 = n16488 ^ n16464 ;
  assign n16465 = n16464 ^ n16459 ;
  assign n16468 = n16467 ^ n16465 ;
  assign n16470 = n16469 ^ n16468 ;
  assign n16490 = n16489 ^ n16470 ;
  assign n16460 = n16459 ^ n16428 ;
  assign n16461 = n16460 ^ n16397 ;
  assign n16491 = n16490 ^ n16461 ;
  assign n16901 = n16900 ^ n16491 ;
  assign n16902 = n16901 ^ n16459 ;
  assign n16903 = n16902 ^ n16479 ;
  assign n16904 = n16903 ^ n16901 ;
  assign n16905 = n16901 ^ n16396 ;
  assign n16906 = n16905 ^ n16901 ;
  assign n16907 = ~n16904 & n16906 ;
  assign n16908 = n16907 ^ n16901 ;
  assign n16909 = ~n16395 & ~n16908 ;
  assign n16910 = n16909 ^ n16456 ;
  assign n16897 = n16486 ^ n16483 ;
  assign n16896 = n16477 ^ n16465 ;
  assign n16898 = n16897 ^ n16896 ;
  assign n16899 = n16519 & ~n16898 ;
  assign n16911 = n16910 ^ n16899 ;
  assign n16511 = n16396 ^ n16395 ;
  assign n16492 = n16491 ^ n16472 ;
  assign n16457 = n16456 ^ n16455 ;
  assign n16493 = n16492 ^ n16457 ;
  assign n16500 = n16493 ^ n16478 ;
  assign n16501 = n16500 ^ n16460 ;
  assign n16522 = n16501 ^ n16483 ;
  assign n16895 = n16511 & n16522 ;
  assign n16912 = n16911 ^ n16895 ;
  assign n16889 = n16475 ^ n16472 ;
  assign n16890 = n16889 ^ n16471 ;
  assign n16891 = n16890 ^ n16493 ;
  assign n16892 = n16395 & n16891 ;
  assign n16893 = n16892 ^ n16475 ;
  assign n16894 = ~n16396 & n16893 ;
  assign n16913 = n16912 ^ n16894 ;
  assign n16521 = n16480 & n16520 ;
  assign n16914 = n16913 ^ n16521 ;
  assign n16915 = ~n16888 & ~n16914 ;
  assign n16916 = n16887 & n16915 ;
  assign n16917 = n16916 ^ n14269 ;
  assign n16918 = n16917 ^ x122 ;
  assign n16919 = n16879 & ~n16918 ;
  assign n16991 = n16919 ^ n16879 ;
  assign n17009 = ~n16975 & n16991 ;
  assign n16987 = n16975 ^ n16938 ;
  assign n16992 = n16987 & n16991 ;
  assign n17010 = n17009 ^ n16992 ;
  assign n16994 = n16973 & n16991 ;
  assign n17008 = n16994 ^ n16991 ;
  assign n17011 = n17010 ^ n17008 ;
  assign n15818 = n15817 ^ n14459 ;
  assign n15819 = n14470 ^ n14457 ;
  assign n15820 = n15818 & ~n15819 ;
  assign n15821 = n15820 ^ n14467 ;
  assign n15793 = n14465 ^ n14460 ;
  assign n15794 = n15793 ^ n14465 ;
  assign n15810 = n14523 ^ n14465 ;
  assign n15811 = n15794 & n15810 ;
  assign n15812 = n15811 ^ n14465 ;
  assign n15813 = n14459 & n15812 ;
  assign n15800 = n14458 ^ n14422 ;
  assign n15801 = n15800 ^ n14460 ;
  assign n15802 = n15801 ^ n15800 ;
  assign n15803 = n15800 ^ n14501 ;
  assign n15804 = n15803 ^ n14451 ;
  assign n15805 = n15804 ^ n15800 ;
  assign n15806 = ~n15802 & n15805 ;
  assign n15807 = n15806 ^ n15800 ;
  assign n15808 = ~n14463 & ~n15807 ;
  assign n15809 = n15808 ^ n15800 ;
  assign n15814 = n15813 ^ n15809 ;
  assign n15815 = n15814 ^ n14497 ;
  assign n15795 = n14521 & ~n15794 ;
  assign n15796 = n15795 ^ n14465 ;
  assign n15797 = n14463 & n15796 ;
  assign n15798 = n15797 ^ n14448 ;
  assign n15790 = ~n14460 & n14532 ;
  assign n15791 = n15790 ^ n14448 ;
  assign n15792 = ~n14463 & n15791 ;
  assign n15799 = n15798 ^ n15792 ;
  assign n15816 = n15815 ^ n15799 ;
  assign n15822 = n15821 ^ n15816 ;
  assign n15823 = n15822 ^ n15785 ;
  assign n15772 = n14497 ^ n14460 ;
  assign n15773 = n15772 ^ n14497 ;
  assign n15774 = ~n15769 & n15773 ;
  assign n15775 = n15774 ^ n14497 ;
  assign n15776 = n14463 & n15775 ;
  assign n15824 = n15823 ^ n15776 ;
  assign n15831 = n15824 & ~n15830 ;
  assign n15832 = n15831 ^ n12456 ;
  assign n16656 = n15832 ^ x69 ;
  assign n16657 = n14781 ^ x78 ;
  assign n16658 = n16656 & ~n16657 ;
  assign n16659 = n16658 ^ n16656 ;
  assign n16677 = n13078 ^ n13019 ;
  assign n16678 = n13017 & ~n16677 ;
  assign n16667 = n13058 ^ n13055 ;
  assign n16668 = n16667 ^ n13059 ;
  assign n16669 = n13057 ^ n13034 ;
  assign n16670 = n16669 ^ n13027 ;
  assign n16671 = n16668 & n16670 ;
  assign n16672 = n16671 ^ n13034 ;
  assign n16673 = n16672 ^ n12825 ;
  assign n16665 = n15423 ^ n12825 ;
  assign n16666 = n11520 & ~n16665 ;
  assign n16674 = n16673 ^ n16666 ;
  assign n16663 = n15423 ^ n13034 ;
  assign n16664 = ~n13008 & ~n16663 ;
  assign n16675 = n16674 ^ n16664 ;
  assign n16662 = n13056 & n13075 ;
  assign n16676 = n16675 ^ n16662 ;
  assign n16679 = n16678 ^ n16676 ;
  assign n16680 = n13075 ^ n11946 ;
  assign n16681 = n16680 ^ n13038 ;
  assign n16682 = n13038 ^ n13008 ;
  assign n16683 = n16682 ^ n13038 ;
  assign n16684 = n16681 & ~n16683 ;
  assign n16685 = n16684 ^ n13038 ;
  assign n16686 = ~n11520 & n16685 ;
  assign n16687 = ~n16679 & ~n16686 ;
  assign n16688 = n13047 & n16687 ;
  assign n16689 = n13035 ^ n13008 ;
  assign n16690 = n16689 ^ n13035 ;
  assign n16691 = n13036 & ~n16690 ;
  assign n16692 = n16691 ^ n13035 ;
  assign n16693 = n16688 & n16692 ;
  assign n16694 = n16693 ^ n16687 ;
  assign n16695 = ~n14715 & n16694 ;
  assign n16696 = n16695 ^ n12490 ;
  assign n16697 = n16696 ^ x108 ;
  assign n16700 = n14953 ^ n14944 ;
  assign n16701 = n16700 ^ n12465 ;
  assign n16702 = n16701 ^ x118 ;
  assign n16705 = ~n16697 & n16702 ;
  assign n16660 = n15001 ^ x101 ;
  assign n15748 = n15289 ^ n15231 ;
  assign n15749 = n15748 ^ n15349 ;
  assign n15750 = n15199 & ~n15749 ;
  assign n15753 = n15752 ^ n15750 ;
  assign n15736 = n15287 ^ n15275 ;
  assign n15509 = n15318 ^ n15279 ;
  assign n15737 = n15736 ^ n15509 ;
  assign n15730 = n15729 ^ n15287 ;
  assign n15731 = n15287 ^ n15196 ;
  assign n15732 = n15731 ^ n15287 ;
  assign n15733 = n15730 & ~n15732 ;
  assign n15734 = n15733 ^ n15287 ;
  assign n15735 = ~n15286 & n15734 ;
  assign n15738 = n15737 ^ n15735 ;
  assign n15728 = n15198 & n15305 ;
  assign n15739 = n15738 ^ n15728 ;
  assign n15754 = n15753 ^ n15739 ;
  assign n15757 = n15756 ^ n15754 ;
  assign n15758 = n15757 ^ n15361 ;
  assign n15762 = n15761 ^ n15758 ;
  assign n15763 = n15762 ^ n15285 ;
  assign n15764 = n15763 ^ n12526 ;
  assign n15740 = n15739 ^ n15276 ;
  assign n15741 = n15740 ^ n15354 ;
  assign n15742 = n15741 ^ n15739 ;
  assign n15743 = n15739 ^ n15197 ;
  assign n15744 = n15743 ^ n15739 ;
  assign n15745 = n15742 & n15744 ;
  assign n15746 = n15745 ^ n15739 ;
  assign n15747 = n15286 & n15746 ;
  assign n15765 = n15764 ^ n15747 ;
  assign n16661 = n15765 ^ x91 ;
  assign n16708 = n16660 & ~n16661 ;
  assign n16713 = n16705 & n16708 ;
  assign n16706 = n16705 ^ n16702 ;
  assign n16711 = n16706 ^ n16697 ;
  assign n16712 = n16708 & n16711 ;
  assign n16714 = n16713 ^ n16712 ;
  assign n16709 = n16706 & n16708 ;
  assign n16710 = n16709 ^ n16708 ;
  assign n16715 = n16714 ^ n16710 ;
  assign n16707 = n16660 & n16706 ;
  assign n16716 = n16715 ^ n16707 ;
  assign n16698 = n16697 ^ n16661 ;
  assign n16699 = ~n16661 & ~n16698 ;
  assign n16703 = n16702 ^ n16699 ;
  assign n16704 = n16660 & n16703 ;
  assign n16717 = n16716 ^ n16704 ;
  assign n16718 = n16659 & n16717 ;
  assign n16720 = n16708 ^ n16661 ;
  assign n16721 = n16720 ^ n16660 ;
  assign n16734 = n16711 & n16721 ;
  assign n16732 = n16708 ^ n16660 ;
  assign n16733 = n16711 & n16732 ;
  assign n16735 = n16734 ^ n16733 ;
  assign n16731 = n16712 ^ n16711 ;
  assign n16736 = n16735 ^ n16731 ;
  assign n16722 = n16711 ^ n16702 ;
  assign n16723 = n16721 & ~n16722 ;
  assign n16749 = n16736 ^ n16723 ;
  assign n16729 = n16715 ^ n16713 ;
  assign n16728 = n16720 ^ n16699 ;
  assign n16730 = n16729 ^ n16728 ;
  assign n16737 = n16736 ^ n16730 ;
  assign n16719 = n16707 ^ n16706 ;
  assign n16745 = n16737 ^ n16719 ;
  assign n16750 = n16749 ^ n16745 ;
  assign n16793 = n16659 & ~n16750 ;
  assign n16741 = n16705 & n16721 ;
  assign n16742 = n16741 ^ n16736 ;
  assign n16740 = n16717 ^ n16714 ;
  assign n16743 = n16742 ^ n16740 ;
  assign n16725 = n16702 ^ n16698 ;
  assign n16726 = n16725 ^ n16661 ;
  assign n16739 = n16735 ^ n16726 ;
  assign n16744 = n16743 ^ n16739 ;
  assign n16746 = n16745 ^ n16744 ;
  assign n16738 = n16737 ^ n16723 ;
  assign n16747 = n16746 ^ n16738 ;
  assign n16748 = n16747 ^ n16720 ;
  assign n16751 = n16750 ^ n16748 ;
  assign n16727 = n16726 ^ n16716 ;
  assign n16752 = n16751 ^ n16727 ;
  assign n16724 = n16723 ^ n16719 ;
  assign n16753 = n16752 ^ n16724 ;
  assign n16754 = n16753 ^ n16712 ;
  assign n16755 = n16658 & ~n16754 ;
  assign n16789 = n16751 ^ n16734 ;
  assign n16790 = n16658 & n16789 ;
  assign n16784 = n16709 ^ n16707 ;
  assign n16785 = n16784 ^ n16715 ;
  assign n16786 = n16659 & n16785 ;
  assign n16767 = n16735 ^ n16716 ;
  assign n16768 = n16767 ^ n16749 ;
  assign n16764 = n16733 ^ n16709 ;
  assign n16765 = n16764 ^ n16746 ;
  assign n16756 = n16657 ^ n16656 ;
  assign n16757 = n16744 ^ n16657 ;
  assign n16758 = n16757 ^ n16744 ;
  assign n16759 = n16744 ^ n16712 ;
  assign n16760 = n16759 ^ n16744 ;
  assign n16761 = n16758 & n16760 ;
  assign n16762 = n16761 ^ n16744 ;
  assign n16763 = ~n16756 & n16762 ;
  assign n16766 = n16765 ^ n16763 ;
  assign n16769 = n16768 ^ n16766 ;
  assign n16770 = n16769 ^ n16763 ;
  assign n16771 = ~n16656 & ~n16770 ;
  assign n16772 = n16771 ^ n16766 ;
  assign n16787 = n16786 ^ n16772 ;
  assign n16776 = n16702 ^ n16660 ;
  assign n16777 = n16776 ^ n16661 ;
  assign n16778 = n16777 ^ n16752 ;
  assign n16781 = ~n16656 & n16778 ;
  assign n16773 = n16772 ^ n16763 ;
  assign n16782 = n16781 ^ n16773 ;
  assign n16783 = n16657 & ~n16782 ;
  assign n16788 = n16787 ^ n16783 ;
  assign n16791 = n16790 ^ n16788 ;
  assign n16792 = ~n16755 & n16791 ;
  assign n16794 = n16793 ^ n16792 ;
  assign n16795 = ~n16718 & n16794 ;
  assign n16796 = n16795 ^ n12613 ;
  assign n16797 = n16796 ^ x72 ;
  assign n15593 = n13888 ^ n13809 ;
  assign n15594 = n15593 ^ n13844 ;
  assign n15600 = n15594 ^ n13871 ;
  assign n15601 = n15600 ^ n13821 ;
  assign n15602 = n15601 ^ n15594 ;
  assign n15603 = n15594 ^ n13576 ;
  assign n15604 = n15603 ^ n15594 ;
  assign n15605 = ~n15602 & ~n15604 ;
  assign n15606 = n15605 ^ n15594 ;
  assign n15607 = n13578 & n15606 ;
  assign n15608 = n15607 ^ n15594 ;
  assign n15591 = n15150 ^ n13577 ;
  assign n15592 = n15591 ^ n15150 ;
  assign n15596 = n15150 ^ n13825 ;
  assign n15597 = n15592 & ~n15596 ;
  assign n15598 = n15597 ^ n15150 ;
  assign n15599 = n13576 & ~n15598 ;
  assign n15609 = n15608 ^ n15599 ;
  assign n15618 = n15609 ^ n11997 ;
  assign n15619 = n15618 ^ n15146 ;
  assign n15610 = ~n13576 & ~n15609 ;
  assign n15611 = n13842 ^ n13577 ;
  assign n15612 = n15611 ^ n13842 ;
  assign n15613 = n13842 ^ n13838 ;
  assign n15614 = n15613 ^ n13842 ;
  assign n15615 = ~n15612 & n15614 ;
  assign n15616 = n15615 ^ n13842 ;
  assign n15617 = n15610 & n15616 ;
  assign n15620 = n15619 ^ n15617 ;
  assign n15768 = n15620 ^ x100 ;
  assign n15833 = n15832 ^ x94 ;
  assign n15834 = n15768 & n15833 ;
  assign n15835 = n15834 ^ n15833 ;
  assign n15836 = n15835 ^ n15768 ;
  assign n15841 = n14326 ^ n14322 ;
  assign n15840 = n14330 ^ n14273 ;
  assign n15842 = n15841 ^ n15840 ;
  assign n15843 = n15842 ^ n14322 ;
  assign n15844 = ~n14311 & ~n15843 ;
  assign n15845 = n15844 ^ n15841 ;
  assign n15854 = n15845 ^ n14316 ;
  assign n15847 = n15845 ^ n14657 ;
  assign n15846 = n15845 ^ n15120 ;
  assign n15848 = n15847 ^ n15846 ;
  assign n15851 = ~n14311 & ~n15848 ;
  assign n15852 = n15851 ^ n15847 ;
  assign n15853 = ~n14163 & ~n15852 ;
  assign n15855 = n15854 ^ n15853 ;
  assign n15838 = n14338 ^ n14330 ;
  assign n15839 = ~n14368 & n15838 ;
  assign n15856 = n15855 ^ n15839 ;
  assign n15837 = n14657 & n14682 ;
  assign n15857 = n15856 ^ n15837 ;
  assign n15865 = n14332 ^ n14324 ;
  assign n15866 = n15865 ^ n14317 ;
  assign n15867 = n15866 ^ n14345 ;
  assign n15868 = ~n14163 & n15867 ;
  assign n15869 = n15868 ^ n14332 ;
  assign n15870 = n14311 & n15869 ;
  assign n15871 = n15870 ^ n14339 ;
  assign n15860 = n14339 ^ n14311 ;
  assign n15861 = n15860 ^ n14339 ;
  assign n15862 = n15103 & ~n15861 ;
  assign n15863 = n15862 ^ n14339 ;
  assign n15864 = ~n14163 & n15863 ;
  assign n15872 = n15871 ^ n15864 ;
  assign n15873 = n15857 & ~n15872 ;
  assign n15874 = n15873 ^ n13214 ;
  assign n15875 = n15874 ^ x75 ;
  assign n15899 = n15170 ^ n14103 ;
  assign n15891 = n14116 ^ n14067 ;
  assign n15890 = n14086 ^ n14074 ;
  assign n15892 = n15891 ^ n15890 ;
  assign n15893 = n15892 ^ n14754 ;
  assign n15894 = ~n13929 & ~n15893 ;
  assign n15895 = n15894 ^ n14754 ;
  assign n15896 = ~n13963 & ~n15895 ;
  assign n15888 = n13964 & ~n14118 ;
  assign n15883 = n14104 ^ n14097 ;
  assign n15884 = n13963 & n15883 ;
  assign n14130 = n14129 ^ n14095 ;
  assign n15876 = n14149 ^ n14130 ;
  assign n15877 = n15876 ^ n14067 ;
  assign n15878 = n15877 ^ n14105 ;
  assign n15879 = n15878 ^ n14149 ;
  assign n15880 = ~n13963 & ~n15879 ;
  assign n15881 = n15880 ^ n15876 ;
  assign n15882 = n15881 ^ n14149 ;
  assign n15885 = n15884 ^ n15882 ;
  assign n15886 = ~n13929 & ~n15885 ;
  assign n15887 = n15886 ^ n15881 ;
  assign n15889 = n15888 ^ n15887 ;
  assign n15897 = n15896 ^ n15889 ;
  assign n15898 = ~n14078 & n15897 ;
  assign n15900 = n15899 ^ n15898 ;
  assign n15901 = ~n14770 & n15900 ;
  assign n15902 = n15901 ^ n13177 ;
  assign n15903 = n15902 ^ x93 ;
  assign n15904 = n15875 & ~n15903 ;
  assign n15916 = n15904 ^ n15903 ;
  assign n15917 = ~n15836 & ~n15916 ;
  assign n15766 = n15765 ^ x125 ;
  assign n15540 = n14927 ^ n14926 ;
  assign n15541 = n14837 ^ n14836 ;
  assign n15548 = n14919 ^ n14917 ;
  assign n15542 = ~n14839 & ~n14915 ;
  assign n15543 = n15542 ^ n14948 ;
  assign n15544 = n15543 ^ n14916 ;
  assign n15545 = n14836 & ~n15544 ;
  assign n15546 = n15545 ^ n15543 ;
  assign n15549 = n15548 ^ n15546 ;
  assign n15547 = n15546 ^ n14926 ;
  assign n15550 = n15549 ^ n15547 ;
  assign n15551 = n15549 ^ n14836 ;
  assign n15552 = n15551 ^ n15549 ;
  assign n15553 = ~n15550 & ~n15552 ;
  assign n15554 = n15553 ^ n15549 ;
  assign n15555 = n15541 & ~n15554 ;
  assign n15556 = n15555 ^ n15546 ;
  assign n15557 = n15540 & ~n15556 ;
  assign n15558 = n15557 ^ n12233 ;
  assign n15767 = n15558 ^ x76 ;
  assign n15933 = n15766 & n15767 ;
  assign n16836 = n15917 & n15933 ;
  assign n15905 = ~n15836 & n15904 ;
  assign n15976 = n15905 ^ n15836 ;
  assign n15906 = n15904 ^ n15875 ;
  assign n15949 = ~n15836 & n15906 ;
  assign n15961 = n15949 ^ n15917 ;
  assign n15977 = n15976 ^ n15961 ;
  assign n15914 = n15836 ^ n15833 ;
  assign n15956 = n15914 & ~n15916 ;
  assign n15978 = n15977 ^ n15956 ;
  assign n16830 = n15978 ^ n15905 ;
  assign n15926 = n15834 & n15904 ;
  assign n16815 = n15926 ^ n15835 ;
  assign n15946 = n15834 & ~n15916 ;
  assign n16816 = n16815 ^ n15946 ;
  assign n15907 = n15906 ^ n15903 ;
  assign n15925 = n15834 & n15907 ;
  assign n16817 = n16816 ^ n15925 ;
  assign n16818 = n15766 & n16817 ;
  assign n15939 = n15835 & n15904 ;
  assign n15908 = n15835 & n15907 ;
  assign n15943 = n15939 ^ n15908 ;
  assign n15927 = n15835 & n15906 ;
  assign n15942 = n15927 ^ n15835 ;
  assign n15944 = n15943 ^ n15942 ;
  assign n15928 = n15927 ^ n15926 ;
  assign n15945 = n15944 ^ n15928 ;
  assign n16819 = n16818 ^ n15945 ;
  assign n16831 = n16830 ^ n16819 ;
  assign n15947 = n15946 ^ n15928 ;
  assign n15948 = n15947 ^ n15945 ;
  assign n16826 = n15948 ^ n15905 ;
  assign n15938 = n15834 & n15906 ;
  assign n15940 = n15939 ^ n15938 ;
  assign n16827 = n16826 ^ n15940 ;
  assign n16828 = n16827 ^ n15978 ;
  assign n16829 = n15766 & ~n16828 ;
  assign n16832 = n16831 ^ n16829 ;
  assign n16833 = n15767 & ~n16832 ;
  assign n15974 = n15907 & n15914 ;
  assign n16820 = n16819 ^ n15974 ;
  assign n15915 = n15906 & n15914 ;
  assign n16806 = n15977 ^ n15915 ;
  assign n16821 = n16820 ^ n16806 ;
  assign n15934 = n15933 ^ n15767 ;
  assign n15935 = n15934 ^ n15766 ;
  assign n15970 = ~n15935 & n15946 ;
  assign n15955 = n15904 & n15914 ;
  assign n15969 = n15934 & n15955 ;
  assign n15971 = n15970 ^ n15969 ;
  assign n16822 = n16821 ^ n15971 ;
  assign n16823 = n16822 ^ n14310 ;
  assign n16807 = n16806 ^ n15955 ;
  assign n15918 = n15917 ^ n15915 ;
  assign n16808 = n16807 ^ n15918 ;
  assign n16809 = n16808 ^ n16806 ;
  assign n16810 = n16806 ^ n15767 ;
  assign n16811 = n16810 ^ n16806 ;
  assign n16812 = n16809 & ~n16811 ;
  assign n16813 = n16812 ^ n16806 ;
  assign n16814 = ~n15766 & ~n16813 ;
  assign n16824 = n16823 ^ n16814 ;
  assign n16800 = n15767 ^ n15766 ;
  assign n16354 = n15974 ^ n15767 ;
  assign n16355 = n16354 ^ n15974 ;
  assign n16362 = n15955 ^ n15949 ;
  assign n16803 = ~n16355 & n16362 ;
  assign n16804 = n16803 ^ n15974 ;
  assign n16805 = n16800 & n16804 ;
  assign n16825 = n16824 ^ n16805 ;
  assign n16834 = n16833 ^ n16825 ;
  assign n16370 = n15944 ^ n15926 ;
  assign n16363 = n15927 ^ n15925 ;
  assign n16798 = n16370 ^ n16363 ;
  assign n16799 = n15934 & n16798 ;
  assign n16835 = n16834 ^ n16799 ;
  assign n16837 = n16836 ^ n16835 ;
  assign n16838 = n16837 ^ x115 ;
  assign n17001 = ~n16797 & ~n16838 ;
  assign n17002 = n17001 ^ n16838 ;
  assign n16977 = n16919 ^ n16918 ;
  assign n16986 = n16977 ^ n16879 ;
  assign n17012 = n16973 & n16986 ;
  assign n19062 = n17012 ^ n17009 ;
  assign n16976 = n16919 & ~n16975 ;
  assign n17048 = n16976 ^ n16919 ;
  assign n17006 = n16919 & n16974 ;
  assign n16995 = n16919 & n16973 ;
  assign n17047 = n17006 ^ n16995 ;
  assign n17049 = n17048 ^ n17047 ;
  assign n16981 = ~n16975 & ~n16977 ;
  assign n18544 = n17049 ^ n16981 ;
  assign n19063 = n19062 ^ n18544 ;
  assign n19064 = ~n17002 & n19063 ;
  assign n16980 = n16974 & ~n16977 ;
  assign n16982 = n16981 ^ n16980 ;
  assign n17018 = n16981 ^ n16797 ;
  assign n17019 = n17018 ^ n16981 ;
  assign n17020 = n16982 & n17019 ;
  assign n17021 = n17020 ^ n16981 ;
  assign n17022 = n16838 & n17021 ;
  assign n19055 = n17022 ^ n17006 ;
  assign n16997 = n16974 & n16986 ;
  assign n19053 = n16997 ^ n16994 ;
  assign n19054 = n17001 & n19053 ;
  assign n19056 = n19055 ^ n19054 ;
  assign n19057 = n19056 ^ n17022 ;
  assign n19051 = n16997 ^ n16995 ;
  assign n19052 = n16797 & n19051 ;
  assign n19058 = n19057 ^ n19052 ;
  assign n19059 = n16838 & n19058 ;
  assign n19060 = n19059 ^ n19056 ;
  assign n16989 = ~n16975 & n16986 ;
  assign n17050 = n17049 ^ n16989 ;
  assign n16988 = n16986 & n16987 ;
  assign n17051 = n17050 ^ n16988 ;
  assign n19049 = n17001 ^ n16797 ;
  assign n19050 = n17051 & ~n19049 ;
  assign n19061 = n19060 ^ n19050 ;
  assign n19065 = n19064 ^ n19061 ;
  assign n16839 = n16838 ^ n16797 ;
  assign n16978 = n16973 & ~n16977 ;
  assign n16979 = n16978 ^ n16977 ;
  assign n16983 = n16982 ^ n16979 ;
  assign n19043 = n16992 ^ n16983 ;
  assign n19044 = n16983 ^ n16838 ;
  assign n19045 = n19044 ^ n16983 ;
  assign n19046 = ~n19043 & n19045 ;
  assign n19047 = n19046 ^ n16983 ;
  assign n19048 = ~n16839 & ~n19047 ;
  assign n19066 = n19065 ^ n19048 ;
  assign n19067 = n19066 ^ n16976 ;
  assign n18570 = ~n16839 & n16988 ;
  assign n18564 = n16983 ^ n16980 ;
  assign n18565 = n16980 ^ n16797 ;
  assign n18566 = n18565 ^ n16980 ;
  assign n18567 = ~n18564 & n18566 ;
  assign n18568 = n18567 ^ n16980 ;
  assign n18569 = ~n16838 & n18568 ;
  assign n18571 = n18570 ^ n18569 ;
  assign n19068 = n19067 ^ n18571 ;
  assign n17042 = n16994 & ~n17002 ;
  assign n17037 = n17009 ^ n16797 ;
  assign n17038 = n17037 ^ n17009 ;
  assign n17039 = n17010 & ~n17038 ;
  assign n17040 = n17039 ^ n17009 ;
  assign n17041 = n16838 & n17040 ;
  assign n17043 = n17042 ^ n17041 ;
  assign n19069 = n19068 ^ n17043 ;
  assign n18528 = n16995 ^ n16978 ;
  assign n19038 = n16976 ^ n16838 ;
  assign n19039 = n19038 ^ n16976 ;
  assign n19040 = n18528 & n19039 ;
  assign n19041 = n19040 ^ n16976 ;
  assign n19042 = n16839 & n19041 ;
  assign n19070 = n19069 ^ n19042 ;
  assign n19071 = ~n17011 & ~n19070 ;
  assign n19072 = n19071 ^ n14381 ;
  assign n19073 = n19072 ^ x88 ;
  assign n15988 = n13546 ^ x81 ;
  assign n16056 = n15380 ^ x107 ;
  assign n16149 = n15988 & ~n16056 ;
  assign n16005 = n14381 ^ x113 ;
  assign n16019 = n14453 ^ n14448 ;
  assign n16020 = n16019 ^ n14523 ;
  assign n16021 = n16020 ^ n15818 ;
  assign n16022 = ~n14464 & ~n16021 ;
  assign n16023 = n16022 ^ n15818 ;
  assign n16026 = n15799 ^ n14459 ;
  assign n16024 = n14501 ^ n14461 ;
  assign n16025 = n16024 ^ n15799 ;
  assign n16027 = n16026 ^ n16025 ;
  assign n16028 = n16023 & ~n16027 ;
  assign n16029 = n16028 ^ n16026 ;
  assign n16030 = n16029 ^ n14492 ;
  assign n16031 = n16030 ^ n16018 ;
  assign n16032 = n16031 ^ n15821 ;
  assign n16043 = n16042 ^ n16032 ;
  assign n16044 = n16043 ^ n15830 ;
  assign n16045 = n16044 ^ n12654 ;
  assign n16006 = n14496 ^ n14461 ;
  assign n16007 = n15817 ^ n14495 ;
  assign n16008 = n14495 ^ n14461 ;
  assign n16009 = n16008 ^ n14495 ;
  assign n16010 = ~n16007 & ~n16009 ;
  assign n16011 = n16010 ^ n14495 ;
  assign n16012 = n16006 & ~n16011 ;
  assign n16046 = n16045 ^ n16012 ;
  assign n16047 = n16046 ^ x74 ;
  assign n16048 = n16005 & n16047 ;
  assign n15989 = n15166 ^ x122 ;
  assign n15990 = n15548 ^ n15543 ;
  assign n15991 = ~n14836 & n15990 ;
  assign n15992 = n15991 ^ n15543 ;
  assign n16001 = n15992 ^ n12661 ;
  assign n15994 = n15992 ^ n14927 ;
  assign n15993 = n15992 ^ n14916 ;
  assign n15995 = n15994 ^ n15993 ;
  assign n15998 = ~n14836 & ~n15995 ;
  assign n15999 = n15998 ^ n15994 ;
  assign n16000 = n14837 & ~n15999 ;
  assign n16002 = n16001 ^ n16000 ;
  assign n16003 = n16002 ^ x104 ;
  assign n16004 = n15989 & ~n16003 ;
  assign n16071 = n16004 ^ n15989 ;
  assign n16072 = n16071 ^ n16003 ;
  assign n16105 = n16072 ^ n15989 ;
  assign n16106 = n16048 & ~n16105 ;
  assign n16049 = n16048 ^ n16047 ;
  assign n16081 = n16004 & n16049 ;
  assign n16050 = n16049 ^ n16005 ;
  assign n16073 = ~n16050 & n16072 ;
  assign n16095 = n16081 ^ n16073 ;
  assign n16094 = n16048 & n16072 ;
  assign n16096 = n16095 ^ n16094 ;
  assign n16053 = ~n16003 & ~n16050 ;
  assign n16054 = ~n15989 & n16053 ;
  assign n16069 = n16054 ^ n16053 ;
  assign n16063 = n16047 ^ n15989 ;
  assign n16064 = ~n16005 & n16063 ;
  assign n16078 = n16069 ^ n16064 ;
  assign n16074 = n16073 ^ n16050 ;
  assign n16075 = n16074 ^ n16053 ;
  assign n16065 = n16047 ^ n16003 ;
  assign n16066 = n16065 ^ n15989 ;
  assign n16067 = n16066 ^ n16005 ;
  assign n16068 = n16064 & n16067 ;
  assign n16070 = n16069 ^ n16068 ;
  assign n16076 = n16075 ^ n16070 ;
  assign n16079 = n16078 ^ n16076 ;
  assign n16080 = n16079 ^ n16075 ;
  assign n16082 = n16081 ^ n16080 ;
  assign n16097 = n16096 ^ n16082 ;
  assign n16093 = n16075 ^ n16072 ;
  assign n16098 = n16097 ^ n16093 ;
  assign n16089 = ~n16003 & ~n16063 ;
  assign n16090 = n16089 ^ n15989 ;
  assign n16091 = n16005 & ~n16090 ;
  assign n16092 = n16091 ^ n16048 ;
  assign n16099 = n16098 ^ n16092 ;
  assign n16107 = n16106 ^ n16099 ;
  assign n16297 = n16107 ^ n16081 ;
  assign n16298 = n16297 ^ n16049 ;
  assign n16299 = n16149 & ~n16298 ;
  assign n16062 = n16056 ^ n15988 ;
  assign n16051 = n16050 ^ n16047 ;
  assign n16052 = n16004 & n16051 ;
  assign n16121 = n16098 ^ n16052 ;
  assign n16289 = ~n16121 & n16149 ;
  assign n16150 = n16149 ^ n16056 ;
  assign n16151 = n16150 ^ n15988 ;
  assign n16157 = n16069 & n16151 ;
  assign n16290 = n16289 ^ n16157 ;
  assign n16286 = n16054 ^ n16050 ;
  assign n16287 = n16286 ^ n16068 ;
  assign n16288 = ~n15988 & ~n16287 ;
  assign n16291 = n16290 ^ n16288 ;
  assign n16285 = n16068 ^ n16067 ;
  assign n16292 = n16291 ^ n16285 ;
  assign n16293 = n16292 ^ n16289 ;
  assign n16294 = n16293 ^ n16157 ;
  assign n16295 = ~n16062 & n16294 ;
  assign n16296 = n16295 ^ n16291 ;
  assign n16300 = n16299 ^ n16296 ;
  assign n16301 = n16300 ^ n16069 ;
  assign n16279 = n16107 ^ n16054 ;
  assign n16280 = n16054 ^ n15988 ;
  assign n16281 = n16280 ^ n16054 ;
  assign n16282 = ~n16279 & ~n16281 ;
  assign n16283 = n16282 ^ n16054 ;
  assign n16284 = n16056 & n16283 ;
  assign n16302 = n16301 ^ n16284 ;
  assign n16303 = n16302 ^ n13575 ;
  assign n16077 = n16076 ^ n16049 ;
  assign n16083 = n16082 ^ n16077 ;
  assign n16084 = n16083 ^ n16079 ;
  assign n16100 = n16099 ^ n16084 ;
  assign n16101 = n16100 ^ n16071 ;
  assign n16102 = n16101 ^ n16080 ;
  assign n16122 = n16102 ^ n16051 ;
  assign n16123 = n16122 ^ n16121 ;
  assign n16271 = n16123 ^ n16079 ;
  assign n16274 = n16069 ^ n15988 ;
  assign n16275 = n16274 ^ n16069 ;
  assign n16276 = ~n16271 & ~n16275 ;
  assign n16277 = n16276 ^ n16069 ;
  assign n16278 = n16056 & n16277 ;
  assign n16304 = n16303 ^ n16278 ;
  assign n16265 = n16081 ^ n16075 ;
  assign n16266 = n16081 ^ n15988 ;
  assign n16267 = n16266 ^ n16081 ;
  assign n16268 = ~n16265 & ~n16267 ;
  assign n16269 = n16268 ^ n16081 ;
  assign n16270 = ~n16062 & n16269 ;
  assign n16305 = n16304 ^ n16270 ;
  assign n16306 = n16305 ^ x125 ;
  assign n15006 = n14835 & ~n15005 ;
  assign n16325 = n15060 ^ n15007 ;
  assign n16326 = ~n16324 & ~n16325 ;
  assign n16317 = n15021 ^ n15009 ;
  assign n16318 = n16317 ^ n15052 ;
  assign n16319 = n15052 ^ n14957 ;
  assign n16320 = n16319 ^ n15052 ;
  assign n16321 = n16318 & ~n16320 ;
  assign n16322 = n16321 ^ n15052 ;
  assign n16323 = ~n15002 & n16322 ;
  assign n16327 = n16326 ^ n16323 ;
  assign n16309 = n15053 ^ n15002 ;
  assign n16310 = n15045 ^ n15008 ;
  assign n16311 = n16310 ^ n15053 ;
  assign n16312 = n16311 ^ n15045 ;
  assign n16313 = n16312 ^ n15034 ;
  assign n16314 = n14957 & n16313 ;
  assign n16315 = n16314 ^ n16310 ;
  assign n16316 = n16309 & ~n16315 ;
  assign n16328 = n16327 ^ n16316 ;
  assign n16307 = n15063 ^ n15023 ;
  assign n16308 = ~n15004 & ~n16307 ;
  assign n16329 = n16328 ^ n16308 ;
  assign n16330 = n15055 ^ n15036 ;
  assign n16331 = n16330 ^ n15047 ;
  assign n16332 = n15047 ^ n15002 ;
  assign n16333 = n16332 ^ n15047 ;
  assign n16334 = ~n16331 & ~n16333 ;
  assign n16335 = n16334 ^ n15047 ;
  assign n16336 = n16324 & ~n16335 ;
  assign n16337 = n16329 & ~n16336 ;
  assign n16338 = ~n15006 & n16337 ;
  assign n16339 = ~n15097 & n16338 ;
  assign n16347 = n16339 & ~n16346 ;
  assign n16348 = n16347 ^ n11945 ;
  assign n16349 = n16348 ^ x116 ;
  assign n16350 = n16306 & n16349 ;
  assign n16351 = n16350 ^ n16306 ;
  assign n15936 = n15935 ^ n15767 ;
  assign n15937 = n15936 ^ n15934 ;
  assign n15975 = n15974 ^ n15908 ;
  assign n15979 = n15978 ^ n15975 ;
  assign n15980 = n15978 ^ n15766 ;
  assign n15981 = n15980 ^ n15978 ;
  assign n15982 = ~n15979 & ~n15981 ;
  assign n15983 = n15982 ^ n15978 ;
  assign n15984 = ~n15937 & ~n15983 ;
  assign n15921 = n15767 & n15918 ;
  assign n15909 = n15908 ^ n15905 ;
  assign n15910 = n15767 & n15909 ;
  assign n15911 = n15910 ^ n15908 ;
  assign n15922 = n15921 ^ n15911 ;
  assign n15923 = ~n15766 & n15922 ;
  assign n15924 = n15923 ^ n15911 ;
  assign n16369 = n15978 ^ n15939 ;
  assign n16371 = n16370 ^ n16369 ;
  assign n16372 = n15767 & ~n16371 ;
  assign n16373 = n16372 ^ n15947 ;
  assign n16367 = n15946 ^ n15944 ;
  assign n16368 = n15767 & n16367 ;
  assign n16374 = n16373 ^ n16368 ;
  assign n16375 = n15766 & n16374 ;
  assign n16376 = n16375 ^ n16372 ;
  assign n16364 = n16363 ^ n15905 ;
  assign n16365 = n16364 ^ n16362 ;
  assign n16366 = ~n15935 & n16365 ;
  assign n16377 = n16376 ^ n16366 ;
  assign n16361 = n15933 & n15938 ;
  assign n16378 = n16377 ^ n16361 ;
  assign n16356 = n15974 ^ n15918 ;
  assign n16357 = n16356 ^ n15974 ;
  assign n16358 = ~n16355 & n16357 ;
  assign n16359 = n16358 ^ n15974 ;
  assign n16360 = n15766 & n16359 ;
  assign n16379 = n16378 ^ n16360 ;
  assign n16380 = n16379 ^ n15970 ;
  assign n16381 = n15955 ^ n15938 ;
  assign n16382 = n15955 ^ n15766 ;
  assign n16383 = n16382 ^ n15955 ;
  assign n16384 = n16381 & ~n16383 ;
  assign n16385 = n16384 ^ n15955 ;
  assign n16386 = n15937 & n16385 ;
  assign n16387 = ~n16380 & ~n16386 ;
  assign n16388 = ~n15924 & n16387 ;
  assign n16389 = ~n15984 & n16388 ;
  assign n16390 = n16389 ^ n13623 ;
  assign n16391 = n16390 ^ x92 ;
  assign n14580 = n14579 ^ n14557 ;
  assign n14583 = n14582 ^ n14580 ;
  assign n14584 = n14535 & n14583 ;
  assign n14585 = n14584 ^ n14579 ;
  assign n16569 = n14585 ^ n14563 ;
  assign n16570 = n16569 ^ n14577 ;
  assign n16571 = n16570 ^ n14605 ;
  assign n16572 = n16571 ^ n14585 ;
  assign n16573 = n14535 & n16572 ;
  assign n16574 = n16573 ^ n16569 ;
  assign n16575 = ~n14382 & n16574 ;
  assign n14613 = n14603 ^ n14543 ;
  assign n16562 = n14613 ^ n14577 ;
  assign n16551 = n14606 ^ n14575 ;
  assign n16560 = n16551 ^ n14566 ;
  assign n16561 = n16560 ^ n14561 ;
  assign n16563 = n16562 ^ n16561 ;
  assign n16564 = n16563 ^ n16551 ;
  assign n16565 = ~n14535 & n16564 ;
  assign n16566 = n16565 ^ n16560 ;
  assign n16567 = n14536 & ~n16566 ;
  assign n16555 = n14537 & n14556 ;
  assign n16554 = n14540 & ~n14581 ;
  assign n16556 = n16555 ^ n16554 ;
  assign n16552 = n16551 ^ n14585 ;
  assign n16545 = n14632 ^ n14615 ;
  assign n16546 = n14632 ^ n14382 ;
  assign n16547 = n16546 ^ n14632 ;
  assign n16548 = n16545 & n16547 ;
  assign n16549 = n16548 ^ n14632 ;
  assign n16550 = ~n14535 & n16549 ;
  assign n16553 = n16552 ^ n16550 ;
  assign n16557 = n16556 ^ n16553 ;
  assign n14568 = n14567 ^ n14535 ;
  assign n14569 = n14568 ^ n14567 ;
  assign n14570 = n14567 ^ n14547 ;
  assign n14571 = n14570 ^ n14567 ;
  assign n14572 = n14569 & n14571 ;
  assign n14573 = n14572 ^ n14567 ;
  assign n14574 = ~n14536 & n14573 ;
  assign n16558 = n16557 ^ n14574 ;
  assign n16559 = n16558 ^ n13007 ;
  assign n16568 = n16567 ^ n16559 ;
  assign n16576 = n16575 ^ n16568 ;
  assign n16577 = n16576 ^ x75 ;
  assign n16578 = ~n16391 & ~n16577 ;
  assign n16591 = n16578 ^ n16577 ;
  assign n15168 = n15167 ^ n15139 ;
  assign n15474 = n15473 ^ n15461 ;
  assign n15477 = n15476 ^ n15474 ;
  assign n15470 = n15469 ^ n15467 ;
  assign n15472 = n15471 ^ n15470 ;
  assign n15478 = n15477 ^ n15472 ;
  assign n15479 = n15478 ^ n15452 ;
  assign n15487 = n15479 ^ n15472 ;
  assign n15488 = ~n15167 & n15487 ;
  assign n15489 = n15488 ^ n15472 ;
  assign n15482 = n15458 ^ n15409 ;
  assign n15483 = ~n15381 & n15482 ;
  assign n15462 = n15461 ^ n15457 ;
  assign n15464 = n15463 ^ n15462 ;
  assign n15480 = n15479 ^ n15464 ;
  assign n15481 = n15480 ^ n15463 ;
  assign n15484 = n15483 ^ n15481 ;
  assign n15485 = n15167 & ~n15484 ;
  assign n15486 = n15485 ^ n15480 ;
  assign n15490 = n15489 ^ n15486 ;
  assign n15491 = ~n15168 & n15490 ;
  assign n16392 = n15491 ^ n15486 ;
  assign n16393 = n16392 ^ n13627 ;
  assign n16394 = n16393 ^ x102 ;
  assign n16523 = n16520 ^ n16395 ;
  assign n16524 = n16522 & ~n16523 ;
  assign n16525 = n16524 ^ n16521 ;
  assign n16536 = n16535 ^ n16525 ;
  assign n16537 = n16536 ^ n13802 ;
  assign n16502 = n16501 ^ n16487 ;
  assign n16498 = n16474 ^ n16462 ;
  assign n16499 = n16396 & n16498 ;
  assign n16503 = n16502 ^ n16499 ;
  assign n16496 = n16483 ^ n16467 ;
  assign n16497 = n16496 ^ n16487 ;
  assign n16504 = n16503 ^ n16497 ;
  assign n16494 = n16493 ^ n16477 ;
  assign n16495 = n16494 ^ n16474 ;
  assign n16505 = n16504 ^ n16495 ;
  assign n16506 = n16505 ^ n16503 ;
  assign n16507 = ~n16396 & ~n16506 ;
  assign n16508 = n16507 ^ n16504 ;
  assign n16509 = ~n16395 & n16508 ;
  assign n16510 = n16509 ^ n16503 ;
  assign n16538 = n16537 ^ n16510 ;
  assign n16515 = n16472 ^ n16431 ;
  assign n16516 = n16515 ^ n16479 ;
  assign n16517 = n16395 & n16516 ;
  assign n16539 = n16538 ^ n16517 ;
  assign n16514 = ~n16396 & n16480 ;
  assign n16540 = n16539 ^ n16514 ;
  assign n16512 = ~n16476 & n16511 ;
  assign n16513 = ~n16510 & n16512 ;
  assign n16541 = n16540 ^ n16513 ;
  assign n16542 = n16541 ^ x85 ;
  assign n16543 = n16394 & n16542 ;
  assign n16589 = n16543 ^ n16542 ;
  assign n16621 = n16589 ^ n16394 ;
  assign n16624 = ~n16591 & ~n16621 ;
  assign n16581 = n16578 ^ n16391 ;
  assign n16623 = ~n16581 & ~n16621 ;
  assign n16625 = n16624 ^ n16623 ;
  assign n16602 = n16542 & n16577 ;
  assign n16603 = n16602 ^ n16589 ;
  assign n16579 = n16543 ^ n16394 ;
  assign n16580 = n16578 & n16579 ;
  assign n16617 = n16603 ^ n16580 ;
  assign n16618 = n16617 ^ n16578 ;
  assign n16598 = n16589 & ~n16591 ;
  assign n16544 = ~n16391 & n16543 ;
  assign n16593 = n16544 ^ n16543 ;
  assign n16592 = n16543 & ~n16591 ;
  assign n16594 = n16593 ^ n16592 ;
  assign n16599 = n16598 ^ n16594 ;
  assign n16605 = n16599 ^ n16544 ;
  assign n16619 = n16618 ^ n16605 ;
  assign n16622 = n16621 ^ n16619 ;
  assign n16626 = n16625 ^ n16622 ;
  assign n19105 = n16351 & ~n16626 ;
  assign n16597 = ~n16581 & n16589 ;
  assign n16600 = n16599 ^ n16597 ;
  assign n16352 = n16350 ^ n16349 ;
  assign n16615 = n16352 ^ n16306 ;
  assign n19103 = n16600 & ~n16615 ;
  assign n19099 = n16306 & n16619 ;
  assign n16353 = n16352 ^ n16351 ;
  assign n19094 = n16625 ^ n16580 ;
  assign n16590 = n16578 & n16589 ;
  assign n16595 = n16594 ^ n16590 ;
  assign n16596 = n16595 ^ n16589 ;
  assign n16601 = n16600 ^ n16596 ;
  assign n18378 = n16601 ^ n16592 ;
  assign n19088 = n18378 ^ n16544 ;
  assign n19095 = n19094 ^ n19088 ;
  assign n16604 = n16603 ^ n16590 ;
  assign n16606 = n16605 ^ n16604 ;
  assign n19090 = n16606 ^ n16580 ;
  assign n19091 = n19090 ^ n16600 ;
  assign n19092 = n19091 ^ n16625 ;
  assign n19093 = n16349 & n19092 ;
  assign n19096 = n19095 ^ n19093 ;
  assign n19097 = ~n16353 & n19096 ;
  assign n16582 = n16581 ^ n16577 ;
  assign n16583 = n16579 & ~n16582 ;
  assign n19089 = n19088 ^ n16583 ;
  assign n19098 = n19097 ^ n19089 ;
  assign n19100 = n19099 ^ n19098 ;
  assign n16630 = n16349 ^ n16306 ;
  assign n16585 = n16579 & ~n16581 ;
  assign n19081 = n16585 ^ n16349 ;
  assign n19082 = n19081 ^ n16585 ;
  assign n19083 = n16585 ^ n16583 ;
  assign n19084 = n19083 ^ n16585 ;
  assign n19085 = ~n19082 & n19084 ;
  assign n19086 = n19085 ^ n16585 ;
  assign n19087 = ~n16630 & n19086 ;
  assign n19101 = n19100 ^ n19087 ;
  assign n19102 = n19101 ^ n16590 ;
  assign n19104 = n19103 ^ n19102 ;
  assign n19106 = n19105 ^ n19104 ;
  assign n19074 = n16590 ^ n16352 ;
  assign n18368 = n16626 ^ n16580 ;
  assign n19075 = n18368 ^ n16351 ;
  assign n19078 = ~n16590 & n19075 ;
  assign n19079 = n19078 ^ n16351 ;
  assign n19080 = n19074 & ~n19079 ;
  assign n19107 = n19106 ^ n19080 ;
  assign n16586 = n16585 ^ n16579 ;
  assign n16584 = n16583 ^ n16580 ;
  assign n16587 = n16586 ^ n16584 ;
  assign n18593 = ~n16353 & n16587 ;
  assign n19108 = n19107 ^ n18593 ;
  assign n19109 = n19108 ^ n13894 ;
  assign n19110 = n19109 ^ x120 ;
  assign n15985 = n15984 ^ n13308 ;
  assign n15957 = n15956 ^ n15905 ;
  assign n15958 = n15957 ^ n15917 ;
  assign n15959 = n15958 ^ n15955 ;
  assign n15960 = ~n15767 & n15959 ;
  assign n15962 = n15961 ^ n15960 ;
  assign n15950 = n15918 ^ n15908 ;
  assign n15951 = n15950 ^ n15949 ;
  assign n15954 = n15951 ^ n15908 ;
  assign n15963 = n15962 ^ n15954 ;
  assign n15952 = n15951 ^ n15948 ;
  assign n15953 = n15767 & n15952 ;
  assign n15964 = n15963 ^ n15953 ;
  assign n15965 = ~n15766 & n15964 ;
  assign n15966 = n15965 ^ n15962 ;
  assign n15941 = ~n15937 & n15940 ;
  assign n15967 = n15966 ^ n15941 ;
  assign n15931 = n15767 & n15928 ;
  assign n15929 = n15928 ^ n15925 ;
  assign n15930 = n15766 & n15929 ;
  assign n15932 = n15931 ^ n15930 ;
  assign n15968 = n15967 ^ n15932 ;
  assign n15972 = ~n15968 & ~n15971 ;
  assign n15973 = ~n15924 & n15972 ;
  assign n15986 = n15985 ^ n15973 ;
  assign n15987 = n15986 ^ x100 ;
  assign n16158 = n16157 ^ n13143 ;
  assign n16103 = ~n16062 & ~n16102 ;
  assign n16055 = n16054 ^ n16052 ;
  assign n16057 = n16056 ^ n16054 ;
  assign n16058 = n16057 ^ n16054 ;
  assign n16059 = n16055 & ~n16058 ;
  assign n16060 = n16059 ^ n16054 ;
  assign n16061 = ~n15988 & n16060 ;
  assign n16104 = n16103 ^ n16061 ;
  assign n16152 = n16080 & n16151 ;
  assign n16137 = ~n15988 & ~n16100 ;
  assign n16138 = n16137 ^ n16099 ;
  assign n16141 = n16138 ^ n16052 ;
  assign n16142 = n16141 ^ n16138 ;
  assign n16143 = n15988 & n16142 ;
  assign n16144 = n16143 ^ n16138 ;
  assign n16145 = n16056 & ~n16144 ;
  assign n16146 = n16145 ^ n16138 ;
  assign n16120 = n16083 ^ n16070 ;
  assign n16124 = n16123 ^ n16120 ;
  assign n16125 = n16124 ^ n16073 ;
  assign n16118 = n16098 ^ n16076 ;
  assign n16117 = n16094 ^ n16053 ;
  assign n16119 = n16118 ^ n16117 ;
  assign n16126 = n16125 ^ n16119 ;
  assign n16127 = ~n16056 & ~n16126 ;
  assign n16128 = n16127 ^ n16125 ;
  assign n16147 = n16146 ^ n16128 ;
  assign n16130 = n16128 ^ n16095 ;
  assign n16129 = n16128 ^ n16091 ;
  assign n16131 = n16130 ^ n16129 ;
  assign n16134 = n16056 & n16131 ;
  assign n16135 = n16134 ^ n16130 ;
  assign n16136 = ~n15988 & ~n16135 ;
  assign n16148 = n16147 ^ n16136 ;
  assign n16153 = n16152 ^ n16148 ;
  assign n16114 = n16094 ^ n16048 ;
  assign n16115 = n16114 ^ n16107 ;
  assign n16116 = ~n16056 & ~n16115 ;
  assign n16154 = n16153 ^ n16116 ;
  assign n16108 = n16107 ^ n16106 ;
  assign n16109 = n16106 ^ n15988 ;
  assign n16110 = n16109 ^ n16106 ;
  assign n16111 = ~n16108 & n16110 ;
  assign n16112 = n16111 ^ n16106 ;
  assign n16113 = ~n16062 & n16112 ;
  assign n16155 = n16154 ^ n16113 ;
  assign n16156 = ~n16104 & ~n16155 ;
  assign n16159 = n16158 ^ n16156 ;
  assign n16160 = n16159 ^ x86 ;
  assign n15492 = n15489 ^ n15139 ;
  assign n15493 = n15492 ^ n15491 ;
  assign n15494 = n15493 ^ n13379 ;
  assign n15495 = n15494 ^ x101 ;
  assign n15621 = n15620 ^ x88 ;
  assign n15590 = n13100 ^ x66 ;
  assign n15646 = n15621 ^ n15590 ;
  assign n15559 = n15558 ^ x64 ;
  assign n15507 = ~n15197 & n15277 ;
  assign n15508 = n15507 ^ n15276 ;
  assign n15529 = n15508 ^ n15315 ;
  assign n15530 = n15529 ^ n15304 ;
  assign n15531 = n15530 ^ n15318 ;
  assign n15532 = n15531 ^ n15508 ;
  assign n15533 = n15197 & ~n15532 ;
  assign n15534 = n15533 ^ n15529 ;
  assign n15535 = n15286 & ~n15534 ;
  assign n15520 = n15509 ^ n15304 ;
  assign n15521 = n15197 & n15520 ;
  assign n15517 = n15376 ^ n15304 ;
  assign n15518 = n15517 ^ n15303 ;
  assign n15519 = n15518 ^ n15285 ;
  assign n15522 = n15521 ^ n15519 ;
  assign n15510 = n15509 ^ n15271 ;
  assign n15511 = n15510 ^ n15287 ;
  assign n15512 = n15287 ^ n15197 ;
  assign n15513 = n15512 ^ n15287 ;
  assign n15514 = n15511 & n15513 ;
  assign n15515 = n15514 ^ n15287 ;
  assign n15516 = n15286 & n15515 ;
  assign n15523 = n15522 ^ n15516 ;
  assign n15524 = n15523 ^ n15508 ;
  assign n15525 = n15524 ^ n15506 ;
  assign n15526 = n15525 ^ n12289 ;
  assign n15498 = n15316 ^ n15271 ;
  assign n15499 = ~n15286 & ~n15498 ;
  assign n15527 = n15526 ^ n15499 ;
  assign n15496 = n15278 ^ n15269 ;
  assign n15497 = ~n15197 & n15496 ;
  assign n15528 = n15527 ^ n15497 ;
  assign n15536 = n15535 ^ n15528 ;
  assign n15537 = n15536 ^ x112 ;
  assign n15538 = n14534 ^ x98 ;
  assign n15539 = n15537 & ~n15538 ;
  assign n15649 = n15539 ^ n15538 ;
  assign n15650 = n15649 ^ n15537 ;
  assign n15651 = n15650 ^ n15538 ;
  assign n15576 = n13486 ^ n13480 ;
  assign n15577 = n13311 & ~n15576 ;
  assign n15570 = n13483 ^ n13463 ;
  assign n15571 = n15570 ^ n13474 ;
  assign n15572 = n15571 ^ n14992 ;
  assign n15568 = n13498 ^ n13463 ;
  assign n15569 = ~n13309 & ~n15568 ;
  assign n15573 = n15572 ^ n15569 ;
  assign n15574 = ~n14958 & ~n15573 ;
  assign n15575 = n15574 ^ n13474 ;
  assign n15578 = n15577 ^ n15575 ;
  assign n15584 = ~n13312 & ~n13491 ;
  assign n15585 = ~n15578 & n15584 ;
  assign n15579 = n15578 ^ n13523 ;
  assign n15567 = n15382 ^ n14993 ;
  assign n15580 = n15579 ^ n15567 ;
  assign n15581 = n15580 ^ n13512 ;
  assign n15582 = n15581 ^ n12047 ;
  assign n15562 = n13526 ^ n13309 ;
  assign n15563 = n15562 ^ n13526 ;
  assign n15564 = n13529 & ~n15563 ;
  assign n15565 = n15564 ^ n13526 ;
  assign n15566 = n13144 & n15565 ;
  assign n15583 = n15582 ^ n15566 ;
  assign n15586 = n15585 ^ n15583 ;
  assign n15587 = n15586 ^ x73 ;
  assign n15652 = n15651 ^ n15587 ;
  assign n15657 = ~n15559 & ~n15652 ;
  assign n15588 = n15559 & n15587 ;
  assign n15633 = n15588 ^ n15559 ;
  assign n15635 = n15539 & n15633 ;
  assign n15634 = ~n15537 & n15633 ;
  assign n15636 = n15635 ^ n15634 ;
  assign n15656 = n15652 ^ n15636 ;
  assign n15658 = n15657 ^ n15656 ;
  assign n15626 = n15538 ^ n15537 ;
  assign n15638 = n15626 & n15633 ;
  assign n15639 = n15638 ^ n15636 ;
  assign n15659 = n15658 ^ n15639 ;
  assign n15629 = n15587 ^ n15559 ;
  assign n15630 = n15629 ^ n15537 ;
  assign n15631 = n15630 ^ n15538 ;
  assign n15653 = ~n15631 & n15652 ;
  assign n15654 = n15653 ^ n15636 ;
  assign n15655 = n15654 ^ n15631 ;
  assign n15660 = n15659 ^ n15655 ;
  assign n15627 = n15626 ^ n15587 ;
  assign n15628 = ~n15559 & n15627 ;
  assign n15671 = n15660 ^ n15628 ;
  assign n15672 = n15671 ^ n15657 ;
  assign n15647 = n15633 ^ n15587 ;
  assign n15664 = ~n15647 & n15651 ;
  assign n15665 = n15664 ^ n15647 ;
  assign n15666 = n15665 ^ n15657 ;
  assign n15673 = n15672 ^ n15666 ;
  assign n15668 = n15647 ^ n15559 ;
  assign n15669 = n15539 & n15668 ;
  assign n15670 = n15669 ^ n15668 ;
  assign n15674 = n15673 ^ n15670 ;
  assign n15648 = n15539 & ~n15647 ;
  assign n15661 = n15660 ^ n15648 ;
  assign n15662 = n15661 ^ n15657 ;
  assign n15663 = n15590 & n15662 ;
  assign n15667 = n15666 ^ n15663 ;
  assign n15677 = n15667 ^ n15621 ;
  assign n15678 = n15677 ^ n15667 ;
  assign n15679 = ~n15674 & n15678 ;
  assign n15680 = n15679 ^ n15667 ;
  assign n15681 = ~n15646 & ~n15680 ;
  assign n15682 = n15681 ^ n15667 ;
  assign n15685 = n15665 ^ n15661 ;
  assign n15686 = n15621 & ~n15685 ;
  assign n15683 = n15664 ^ n15648 ;
  assign n15684 = n15590 & n15683 ;
  assign n15687 = n15686 ^ n15684 ;
  assign n15622 = n15590 & n15621 ;
  assign n15637 = n15636 ^ n15633 ;
  assign n15640 = n15639 ^ n15637 ;
  assign n15718 = n15622 & n15640 ;
  assign n15706 = n15658 ^ n15621 ;
  assign n17139 = n15706 ^ n15658 ;
  assign n15709 = n17139 ^ n15590 ;
  assign n15713 = ~n15590 & n15706 ;
  assign n15691 = n15653 ^ n15559 ;
  assign n15692 = n15691 ^ n15671 ;
  assign n15625 = n15622 ^ n15621 ;
  assign n15589 = n15539 & n15588 ;
  assign n15641 = n15640 ^ n15589 ;
  assign n15632 = n15631 ^ n15628 ;
  assign n15642 = n15641 ^ n15632 ;
  assign n15710 = n15642 ^ n15635 ;
  assign n15711 = ~n15625 & ~n15710 ;
  assign n15712 = n15692 & n15711 ;
  assign n15714 = n15713 ^ n15712 ;
  assign n15715 = n15709 & n15714 ;
  assign n15716 = n15715 ^ n15713 ;
  assign n15717 = n15716 ^ n15706 ;
  assign n15719 = n15718 ^ n15717 ;
  assign n15703 = n15661 ^ n15589 ;
  assign n15704 = n15625 & n15703 ;
  assign n15720 = n15719 ^ n15704 ;
  assign n15693 = n15692 ^ n15637 ;
  assign n15689 = n15638 ^ n15589 ;
  assign n15688 = n15673 ^ n15664 ;
  assign n15690 = n15689 ^ n15688 ;
  assign n15694 = n15693 ^ n15690 ;
  assign n15695 = n15694 ^ n15669 ;
  assign n15698 = n15669 ^ n15590 ;
  assign n15699 = n15698 ^ n15669 ;
  assign n15700 = n15695 & ~n15699 ;
  assign n15701 = n15700 ^ n15669 ;
  assign n15702 = ~n15621 & n15701 ;
  assign n15721 = n15720 ^ n15702 ;
  assign n15722 = ~n15687 & ~n15721 ;
  assign n15723 = n15682 & n15722 ;
  assign n15643 = n15642 ^ n15639 ;
  assign n15644 = n15625 & n15643 ;
  assign n15623 = n15589 & n15622 ;
  assign n15624 = n15623 ^ n13420 ;
  assign n15645 = n15644 ^ n15624 ;
  assign n15724 = n15723 ^ n15645 ;
  assign n15725 = n15724 ^ x124 ;
  assign n15726 = n15495 & n15725 ;
  assign n15727 = n15726 ^ n15495 ;
  assign n14630 = n14602 ^ n14560 ;
  assign n14636 = n14630 ^ n14613 ;
  assign n14631 = n14630 ^ n14558 ;
  assign n14634 = n14633 ^ n14631 ;
  assign n14635 = ~n14382 & n14634 ;
  assign n14637 = n14636 ^ n14635 ;
  assign n14638 = ~n14535 & n14637 ;
  assign n14616 = n14615 ^ n14582 ;
  assign n14617 = ~n14382 & n14616 ;
  assign n14618 = n14617 ^ n14582 ;
  assign n14621 = n14618 ^ n14561 ;
  assign n14622 = n14621 ^ n14618 ;
  assign n14623 = n14382 & n14622 ;
  assign n14624 = n14623 ^ n14618 ;
  assign n14625 = ~n14536 & n14624 ;
  assign n14626 = n14625 ^ n14618 ;
  assign n14614 = n14613 ^ n14612 ;
  assign n14627 = n14626 ^ n14614 ;
  assign n14588 = n14579 ^ n14535 ;
  assign n14589 = n14588 ^ n14579 ;
  assign n14590 = n14585 & n14589 ;
  assign n14591 = n14590 ^ n14579 ;
  assign n14592 = n14382 & n14591 ;
  assign n14628 = n14627 ^ n14592 ;
  assign n14629 = n14628 ^ n14574 ;
  assign n14639 = n14638 ^ n14629 ;
  assign n14549 = n14548 ^ n14543 ;
  assign n14550 = n14548 ^ n14382 ;
  assign n14551 = n14550 ^ n14548 ;
  assign n14552 = n14549 & n14551 ;
  assign n14553 = n14552 ^ n14548 ;
  assign n14554 = n14536 & n14553 ;
  assign n14640 = n14639 ^ n14554 ;
  assign n14641 = ~n14541 & ~n14640 ;
  assign n14642 = n14641 ^ n13454 ;
  assign n14643 = n14642 ^ x68 ;
  assign n15098 = n15097 ^ n13351 ;
  assign n15093 = n15053 ^ n15025 ;
  assign n15094 = n15003 & n15093 ;
  assign n15090 = n15056 ^ n15007 ;
  assign n15091 = ~n15004 & n15090 ;
  assign n15087 = n15026 ^ n15020 ;
  assign n15088 = ~n15002 & ~n15087 ;
  assign n15082 = n15036 ^ n15005 ;
  assign n15072 = n15060 ^ n15003 ;
  assign n15073 = n15014 ^ n14957 ;
  assign n15074 = n15060 ^ n14957 ;
  assign n15075 = n15074 ^ n14957 ;
  assign n15076 = n15073 & n15075 ;
  assign n15077 = n15076 ^ n14957 ;
  assign n15078 = ~n15072 & ~n15077 ;
  assign n15079 = n15078 ^ n15003 ;
  assign n15071 = n15045 & ~n15070 ;
  assign n15080 = n15079 ^ n15071 ;
  assign n15081 = n15080 ^ n15020 ;
  assign n15083 = n15082 ^ n15081 ;
  assign n15046 = n15045 ^ n15005 ;
  assign n15064 = n15063 ^ n15003 ;
  assign n15065 = n15045 ^ n15003 ;
  assign n15066 = n15065 ^ n15003 ;
  assign n15067 = n15064 & ~n15066 ;
  assign n15068 = n15067 ^ n15003 ;
  assign n15069 = ~n15046 & n15068 ;
  assign n15084 = n15083 ^ n15069 ;
  assign n15037 = n15036 ^ n14957 ;
  assign n15038 = n15037 ^ n15036 ;
  assign n15039 = n15036 ^ n15021 ;
  assign n15040 = n15039 ^ n15036 ;
  assign n15041 = n15038 & ~n15040 ;
  assign n15042 = n15041 ^ n15036 ;
  assign n15043 = ~n15002 & n15042 ;
  assign n15085 = n15084 ^ n15043 ;
  assign n15027 = n15026 ^ n14835 ;
  assign n15028 = n15027 ^ n15023 ;
  assign n15029 = n15023 ^ n15002 ;
  assign n15030 = n15029 ^ n15023 ;
  assign n15031 = n15028 & ~n15030 ;
  assign n15032 = n15031 ^ n15023 ;
  assign n15033 = ~n14957 & n15032 ;
  assign n15086 = n15085 ^ n15033 ;
  assign n15089 = n15088 ^ n15086 ;
  assign n15092 = n15091 ^ n15089 ;
  assign n15095 = n15094 ^ n15092 ;
  assign n15096 = ~n15006 & ~n15095 ;
  assign n15099 = n15098 ^ n15096 ;
  assign n15100 = n15099 ^ x118 ;
  assign n15101 = ~n14643 & n15100 ;
  assign n15102 = n15101 ^ n14643 ;
  assign n16172 = n15102 ^ n15100 ;
  assign n16208 = n15727 & n16172 ;
  assign n16165 = n15100 ^ n14643 ;
  assign n16166 = n15727 & n16165 ;
  assign n16164 = n15101 & ~n15725 ;
  assign n16167 = n16166 ^ n16164 ;
  assign n16209 = n16208 ^ n16167 ;
  assign n16182 = n15727 ^ n15725 ;
  assign n16210 = n16209 ^ n16182 ;
  assign n16206 = n16172 & ~n16182 ;
  assign n16187 = ~n15102 & ~n16182 ;
  assign n16207 = n16206 ^ n16187 ;
  assign n16211 = n16210 ^ n16207 ;
  assign n16173 = n16172 ^ n14643 ;
  assign n16205 = n15727 & n16173 ;
  assign n16212 = n16211 ^ n16205 ;
  assign n16174 = n15726 & n16173 ;
  assign n16204 = n16174 ^ n16173 ;
  assign n16213 = n16212 ^ n16204 ;
  assign n16254 = n16213 ^ n16211 ;
  assign n16255 = n16254 ^ n16206 ;
  assign n16189 = n15101 & n15726 ;
  assign n16214 = n16213 ^ n16189 ;
  assign n16190 = n16189 ^ n15101 ;
  assign n16191 = n16190 ^ n16164 ;
  assign n16215 = n16214 ^ n16191 ;
  assign n16199 = n15726 & n16172 ;
  assign n16183 = n16182 ^ n15495 ;
  assign n16184 = n16172 & n16183 ;
  assign n16193 = n16189 ^ n16184 ;
  assign n16203 = n16199 ^ n16193 ;
  assign n16216 = n16215 ^ n16203 ;
  assign n16202 = n16199 ^ n16183 ;
  assign n16217 = n16216 ^ n16202 ;
  assign n16256 = n16255 ^ n16217 ;
  assign n16257 = ~n16160 & ~n16256 ;
  assign n16258 = n16257 ^ n16213 ;
  assign n16259 = ~n15987 & ~n16258 ;
  assign n16161 = ~n15987 & ~n16160 ;
  assign n18727 = n16161 & ~n16214 ;
  assign n16245 = n16211 ^ n16160 ;
  assign n16246 = n16245 ^ n16211 ;
  assign n16249 = ~n16212 & n16246 ;
  assign n16250 = n16249 ^ n16211 ;
  assign n16251 = n15987 & ~n16250 ;
  assign n18728 = n18727 ^ n16251 ;
  assign n19138 = ~n16259 & ~n18728 ;
  assign n16168 = n16161 ^ n16160 ;
  assign n16169 = n16168 ^ n15987 ;
  assign n18220 = ~n16169 & n16187 ;
  assign n18215 = n15987 ^ n14643 ;
  assign n18216 = n15727 & n18215 ;
  assign n18217 = n16160 ^ n15100 ;
  assign n18218 = ~n16165 & ~n18217 ;
  assign n18219 = n18216 & n18218 ;
  assign n18221 = n18220 ^ n18219 ;
  assign n16185 = n16161 ^ n15987 ;
  assign n19151 = n16174 & ~n16185 ;
  assign n19149 = ~n16168 & ~n16217 ;
  assign n19147 = n16207 ^ n16191 ;
  assign n19148 = n19147 ^ n16199 ;
  assign n19150 = n19149 ^ n19148 ;
  assign n19152 = n19151 ^ n19150 ;
  assign n18224 = n16160 ^ n15987 ;
  assign n16197 = n16189 ^ n16174 ;
  assign n16198 = n16197 ^ n15726 ;
  assign n16200 = n16199 ^ n16198 ;
  assign n18720 = n16200 ^ n14643 ;
  assign n16201 = n16200 ^ n16184 ;
  assign n16218 = n16217 ^ n16201 ;
  assign n16219 = n16218 ^ n16164 ;
  assign n16220 = n16219 ^ n16174 ;
  assign n16221 = n16220 ^ n16187 ;
  assign n18721 = n18720 ^ n16221 ;
  assign n16192 = n16191 ^ n16174 ;
  assign n16194 = n16193 ^ n16192 ;
  assign n18722 = n18721 ^ n16194 ;
  assign n18723 = n15987 & n18722 ;
  assign n18724 = n18723 ^ n16200 ;
  assign n18725 = ~n18224 & n18724 ;
  assign n19154 = n18725 ^ n16207 ;
  assign n19153 = n18725 ^ n18224 ;
  assign n19155 = n19154 ^ n19153 ;
  assign n19156 = n19152 & n19155 ;
  assign n19157 = n19156 ^ n19154 ;
  assign n19158 = n19157 ^ n18725 ;
  assign n19159 = n16209 ^ n16194 ;
  assign n19160 = ~n16169 & n19159 ;
  assign n19161 = ~n19158 & n19160 ;
  assign n19162 = n19161 ^ n19157 ;
  assign n19145 = n16209 ^ n16164 ;
  assign n19146 = ~n16168 & n19145 ;
  assign n19165 = n19162 ^ n19146 ;
  assign n19139 = n16200 ^ n16167 ;
  assign n19140 = n16167 ^ n16160 ;
  assign n19141 = n19140 ^ n16167 ;
  assign n19142 = n19139 & n19141 ;
  assign n19143 = n19142 ^ n16167 ;
  assign n19144 = ~n15987 & n19143 ;
  assign n19166 = n19165 ^ n19144 ;
  assign n19167 = ~n18221 & ~n19166 ;
  assign n19168 = n19138 & n19167 ;
  assign n19169 = n19168 ^ n13546 ;
  assign n19170 = n19169 ^ x65 ;
  assign n19185 = n19110 & n19170 ;
  assign n19224 = n19185 ^ n19170 ;
  assign n19247 = n19224 ^ n19110 ;
  assign n17398 = n13548 & n14540 ;
  assign n17380 = n14602 ^ n14548 ;
  assign n17381 = n17380 ^ n14604 ;
  assign n17379 = n16848 ^ n16562 ;
  assign n17382 = n17381 ^ n17379 ;
  assign n17383 = ~n14535 & ~n17382 ;
  assign n17384 = n17383 ^ n17379 ;
  assign n17393 = n17384 ^ n16550 ;
  assign n17394 = n17393 ^ n14626 ;
  assign n17395 = n17394 ^ n16556 ;
  assign n17396 = n17395 ^ n14592 ;
  assign n17386 = n17384 ^ n14575 ;
  assign n17385 = n17384 ^ n14632 ;
  assign n17387 = n17386 ^ n17385 ;
  assign n17390 = n14535 & n17387 ;
  assign n17391 = n17390 ^ n17386 ;
  assign n17392 = n14382 & ~n17391 ;
  assign n17397 = n17396 ^ n17392 ;
  assign n17399 = n17398 ^ n17397 ;
  assign n17400 = ~n14541 & n17399 ;
  assign n17401 = n17400 ^ n13962 ;
  assign n17402 = n17401 ^ x120 ;
  assign n17138 = n15658 ^ n15648 ;
  assign n17140 = ~n17138 & n17139 ;
  assign n17141 = n17140 ^ n15658 ;
  assign n17142 = ~n15590 & ~n17141 ;
  assign n17247 = n15664 ^ n15539 ;
  assign n17248 = n17247 ^ n15692 ;
  assign n17249 = n17248 ^ n15695 ;
  assign n17250 = n15621 & ~n17249 ;
  assign n17251 = n17250 ^ n15664 ;
  assign n17252 = n15590 & n17251 ;
  assign n17253 = n17252 ^ n15664 ;
  assign n17112 = n15622 ^ n15590 ;
  assign n17268 = n15641 & n17112 ;
  assign n17257 = n15674 ^ n15659 ;
  assign n17254 = n15654 ^ n15648 ;
  assign n17255 = n17254 ^ n15641 ;
  assign n17256 = ~n15621 & ~n17255 ;
  assign n17258 = n17257 ^ n17256 ;
  assign n17259 = ~n15590 & n17258 ;
  assign n17260 = n17259 ^ n15674 ;
  assign n17261 = n17112 ^ n15625 ;
  assign n17262 = n17261 ^ n15692 ;
  assign n17263 = n15685 ^ n15669 ;
  assign n17264 = n17263 ^ n15692 ;
  assign n17265 = ~n17262 & n17264 ;
  assign n17266 = n17265 ^ n15692 ;
  assign n17267 = n17260 & n17266 ;
  assign n17269 = n17268 ^ n17267 ;
  assign n17270 = ~n17253 & n17269 ;
  assign n17271 = n17270 ^ n15623 ;
  assign n17272 = ~n15635 & n17271 ;
  assign n17273 = ~n17142 & n17272 ;
  assign n17274 = n17273 ^ n14051 ;
  assign n17275 = n17274 ^ x97 ;
  assign n17301 = n15019 ^ n15002 ;
  assign n17302 = n17301 ^ n15019 ;
  assign n17303 = ~n15059 & ~n17302 ;
  assign n17304 = n17303 ^ n15019 ;
  assign n17305 = n14957 & n17304 ;
  assign n17283 = n15093 ^ n14731 ;
  assign n17284 = n15002 & ~n17283 ;
  assign n17285 = n17284 ^ n15026 ;
  assign n17289 = n17285 ^ n14831 ;
  assign n17290 = n17289 ^ n16340 ;
  assign n17291 = n17290 ^ n17285 ;
  assign n17294 = n15002 & ~n17291 ;
  assign n17286 = n17285 ^ n15080 ;
  assign n17287 = n17286 ^ n16336 ;
  assign n17288 = n17287 ^ n15080 ;
  assign n17295 = n17294 ^ n17288 ;
  assign n17296 = n17295 ^ n16336 ;
  assign n17297 = n16324 & n17296 ;
  assign n17298 = n17297 ^ n17287 ;
  assign n17306 = n17305 ^ n17298 ;
  assign n17276 = n15023 ^ n15003 ;
  assign n17277 = n15063 ^ n15005 ;
  assign n17280 = ~n15023 & ~n17277 ;
  assign n17281 = n17280 ^ n15005 ;
  assign n17282 = n17276 & ~n17281 ;
  assign n17307 = n17306 ^ n17282 ;
  assign n17308 = ~n15006 & n17307 ;
  assign n17309 = ~n16346 & n17308 ;
  assign n17310 = n17309 ^ n13994 ;
  assign n17311 = n17310 ^ x123 ;
  assign n17312 = ~n17275 & n17311 ;
  assign n17313 = n16659 & n16713 ;
  assign n17320 = n16742 ^ n16717 ;
  assign n17321 = n17320 ^ n16751 ;
  assign n17322 = n17321 ^ n16776 ;
  assign n17323 = ~n16657 & n17322 ;
  assign n17318 = n16751 ^ n16745 ;
  assign n17316 = n16753 ^ n16733 ;
  assign n17317 = n17316 ^ n16736 ;
  assign n17319 = n17318 ^ n17317 ;
  assign n17324 = n17323 ^ n17319 ;
  assign n17341 = n17324 ^ n16786 ;
  assign n17337 = n16784 ^ n16744 ;
  assign n17338 = ~n16758 & n17337 ;
  assign n17339 = n17338 ^ n16744 ;
  assign n17340 = n16756 & n17339 ;
  assign n17342 = n17341 ^ n17340 ;
  assign n17331 = n16789 ^ n16784 ;
  assign n17332 = n16789 ^ n16657 ;
  assign n17333 = n17332 ^ n16789 ;
  assign n17334 = n17331 & n17333 ;
  assign n17335 = n17334 ^ n16789 ;
  assign n17336 = n16756 & n17335 ;
  assign n17343 = n17342 ^ n17336 ;
  assign n17325 = n17324 ^ n16778 ;
  assign n17314 = n16735 ^ n16729 ;
  assign n17315 = n17314 ^ n16738 ;
  assign n17326 = n17325 ^ n17315 ;
  assign n17327 = n17326 ^ n17324 ;
  assign n17328 = n16657 & ~n17327 ;
  assign n17329 = n17328 ^ n17325 ;
  assign n17330 = ~n16656 & n17329 ;
  assign n17344 = n17343 ^ n17330 ;
  assign n17345 = ~n17313 & ~n17344 ;
  assign n17346 = n17345 ^ n14022 ;
  assign n17347 = n17346 ^ x106 ;
  assign n17351 = n15457 ^ n14062 ;
  assign n17349 = n15474 ^ n15457 ;
  assign n17350 = n15139 & n17349 ;
  assign n17352 = n17351 ^ n17350 ;
  assign n17353 = n17352 ^ n14062 ;
  assign n17354 = n17353 ^ n16923 ;
  assign n17355 = ~n15167 & ~n17354 ;
  assign n17356 = n17355 ^ n17352 ;
  assign n17348 = ~n15139 & n15473 ;
  assign n17357 = n17356 ^ n17348 ;
  assign n17358 = n17357 ^ x88 ;
  assign n17359 = ~n17347 & n17358 ;
  assign n17364 = n17359 ^ n17347 ;
  assign n17445 = n17364 ^ n17358 ;
  assign n17450 = n17312 & n17445 ;
  assign n17366 = ~n17275 & ~n17347 ;
  assign n17361 = n17312 ^ n17275 ;
  assign n17365 = ~n17361 & ~n17364 ;
  assign n17367 = n17366 ^ n17365 ;
  assign n17451 = n17450 ^ n17367 ;
  assign n17362 = n17359 & ~n17361 ;
  assign n17449 = n17362 ^ n17312 ;
  assign n17452 = n17451 ^ n17449 ;
  assign n17446 = ~n17361 & n17445 ;
  assign n17447 = n17446 ^ n17362 ;
  assign n17444 = n17365 ^ n17361 ;
  assign n17448 = n17447 ^ n17444 ;
  assign n17453 = n17452 ^ n17448 ;
  assign n17370 = n17361 ^ n17311 ;
  assign n17441 = n17359 ^ n17358 ;
  assign n17442 = n17370 & n17441 ;
  assign n17443 = n17442 ^ n17441 ;
  assign n17454 = n17453 ^ n17443 ;
  assign n17423 = n16478 ^ n16456 ;
  assign n17424 = n16518 & n17423 ;
  assign n17411 = n16475 ^ n16467 ;
  assign n17412 = n17411 ^ n16522 ;
  assign n17413 = n16396 & n17412 ;
  assign n17414 = n17413 ^ n16470 ;
  assign n17415 = n17414 ^ n16490 ;
  assign n17416 = n17415 ^ n17414 ;
  assign n17419 = ~n16396 & n17416 ;
  assign n17420 = n17419 ^ n17414 ;
  assign n17421 = n16511 & n17420 ;
  assign n17422 = n17421 ^ n17413 ;
  assign n17425 = n17424 ^ n17422 ;
  assign n17405 = n16476 ^ n16456 ;
  assign n17406 = n17405 ^ n16483 ;
  assign n17407 = n17406 ^ n16491 ;
  assign n17408 = ~n16396 & ~n17407 ;
  assign n17409 = n17408 ^ n16493 ;
  assign n17410 = ~n16395 & n17409 ;
  assign n17426 = n17425 ^ n17410 ;
  assign n17427 = ~n16886 & ~n17426 ;
  assign n17428 = n16492 ^ n16471 ;
  assign n17429 = n16471 ^ n16396 ;
  assign n17430 = n17429 ^ n16471 ;
  assign n17431 = n17428 & n17430 ;
  assign n17432 = n17431 ^ n16471 ;
  assign n17433 = ~n16511 & n17432 ;
  assign n17434 = n17427 & ~n17433 ;
  assign n17403 = n16535 ^ n13928 ;
  assign n17404 = n17403 ^ n16888 ;
  assign n17435 = n17434 ^ n17404 ;
  assign n17436 = n17435 ^ x65 ;
  assign n17455 = n17454 ^ n17436 ;
  assign n17456 = n17455 ^ n17454 ;
  assign n17371 = n17370 ^ n17275 ;
  assign n17460 = n17371 & n17445 ;
  assign n17374 = n17359 & n17370 ;
  assign n17461 = n17460 ^ n17374 ;
  assign n17462 = n17461 ^ n17454 ;
  assign n17360 = n17312 & n17359 ;
  assign n17363 = n17362 ^ n17360 ;
  assign n17373 = n17363 ^ n17359 ;
  assign n17375 = n17374 ^ n17373 ;
  assign n17463 = n17462 ^ n17375 ;
  assign n17372 = ~n17347 & n17371 ;
  assign n17376 = n17375 ^ n17372 ;
  assign n17457 = n17442 ^ n17376 ;
  assign n17377 = n17376 ^ n17365 ;
  assign n17368 = n17367 ^ n17363 ;
  assign n17369 = n17368 ^ n17364 ;
  assign n17378 = n17377 ^ n17369 ;
  assign n17458 = n17457 ^ n17378 ;
  assign n17459 = n17458 ^ n17275 ;
  assign n17464 = n17463 ^ n17459 ;
  assign n17465 = n17464 ^ n17454 ;
  assign n17468 = n17456 & ~n17465 ;
  assign n17469 = n17468 ^ n17454 ;
  assign n17470 = n17402 & ~n17469 ;
  assign n19135 = n17470 ^ n14159 ;
  assign n17437 = ~n17402 & n17436 ;
  assign n17438 = n17437 ^ n17402 ;
  assign n18633 = ~n17378 & ~n17438 ;
  assign n19127 = n17448 ^ n17360 ;
  assign n19128 = n19127 ^ n17461 ;
  assign n19129 = n17436 & ~n19128 ;
  assign n17485 = n17375 ^ n17365 ;
  assign n19130 = n19129 ^ n17485 ;
  assign n19131 = n17402 & n19130 ;
  assign n17439 = n17438 ^ n17436 ;
  assign n18609 = n17439 ^ n17437 ;
  assign n18618 = n17452 ^ n17378 ;
  assign n18621 = ~n17436 & ~n18618 ;
  assign n18622 = n18621 ^ n17378 ;
  assign n18623 = ~n18609 & ~n18622 ;
  assign n19122 = n18623 ^ n17485 ;
  assign n17500 = n17452 ^ n17368 ;
  assign n17501 = n17500 ^ n17448 ;
  assign n17502 = n17448 ^ n17436 ;
  assign n17503 = n17502 ^ n17448 ;
  assign n17504 = ~n17501 & n17503 ;
  assign n17505 = n17504 ^ n17448 ;
  assign n17506 = n17402 & ~n17505 ;
  assign n19123 = n19122 ^ n17506 ;
  assign n17472 = n17436 ^ n17402 ;
  assign n17507 = n17450 ^ n17447 ;
  assign n17508 = n17507 ^ n17450 ;
  assign n17509 = n17450 ^ n17436 ;
  assign n17510 = n17509 ^ n17450 ;
  assign n17511 = n17508 & ~n17510 ;
  assign n17512 = n17511 ^ n17450 ;
  assign n17513 = ~n17472 & n17512 ;
  assign n17514 = n17513 ^ n17450 ;
  assign n19124 = n19123 ^ n17514 ;
  assign n19117 = n17460 ^ n17442 ;
  assign n19115 = n17454 ^ n17442 ;
  assign n19116 = n19115 ^ n17376 ;
  assign n19118 = n19117 ^ n19116 ;
  assign n19119 = n17436 & ~n19118 ;
  assign n19120 = n19119 ^ n19117 ;
  assign n19121 = ~n17402 & n19120 ;
  assign n19125 = n19124 ^ n19121 ;
  assign n19114 = n17447 & n18609 ;
  assign n19126 = n19125 ^ n19114 ;
  assign n19132 = n19131 ^ n19126 ;
  assign n19113 = n17439 & ~n17458 ;
  assign n19133 = n19132 ^ n19113 ;
  assign n19134 = ~n18633 & ~n19133 ;
  assign n19136 = n19135 ^ n19134 ;
  assign n19137 = n19136 ^ x113 ;
  assign n19171 = n19137 & ~n19170 ;
  assign n19177 = ~n19110 & n19171 ;
  assign n19248 = n19247 ^ n19177 ;
  assign n17074 = n16937 ^ x91 ;
  assign n17075 = n16576 ^ x109 ;
  assign n17076 = ~n17074 & n17075 ;
  assign n17077 = n17076 ^ n17074 ;
  assign n17104 = n16115 ^ n16095 ;
  assign n17105 = n17104 ^ n16120 ;
  assign n17103 = n16271 ^ n16076 ;
  assign n17106 = n17105 ^ n17103 ;
  assign n17107 = ~n16056 & n17106 ;
  assign n17108 = n17107 ^ n17103 ;
  assign n17109 = n15988 & n17108 ;
  assign n17100 = n16124 ^ n16069 ;
  assign n17101 = ~n16150 & ~n17100 ;
  assign n17093 = n16054 & n16149 ;
  assign n17094 = n17093 ^ n16284 ;
  assign n17091 = n16099 ^ n16081 ;
  assign n17092 = n17091 ^ n16104 ;
  assign n17095 = n17094 ^ n17092 ;
  assign n17096 = n17095 ^ n16289 ;
  assign n17097 = n17096 ^ n12822 ;
  assign n17083 = n16099 ^ n16052 ;
  assign n17084 = n17083 ^ n16118 ;
  assign n17085 = n17084 ^ n16099 ;
  assign n17086 = n16099 ^ n16056 ;
  assign n17087 = n17086 ^ n16099 ;
  assign n17088 = n17085 & n17087 ;
  assign n17089 = n17088 ^ n16099 ;
  assign n17090 = n16062 & ~n17089 ;
  assign n17098 = n17097 ^ n17090 ;
  assign n17080 = n16106 & ~n16267 ;
  assign n17081 = n17080 ^ n16081 ;
  assign n17082 = ~n16056 & n17081 ;
  assign n17099 = n17098 ^ n17082 ;
  assign n17102 = n17101 ^ n17099 ;
  assign n17110 = n17109 ^ n17102 ;
  assign n17111 = n17110 ^ x77 ;
  assign n17148 = n15674 ^ n15660 ;
  assign n17149 = n15625 ^ n15590 ;
  assign n17150 = ~n17148 & ~n17149 ;
  assign n17145 = n17112 ^ n15644 ;
  assign n17126 = n15657 ^ n15647 ;
  assign n17127 = n17126 ^ n15671 ;
  assign n17128 = ~n15590 & ~n17127 ;
  assign n17129 = n17128 ^ n15657 ;
  assign n17143 = n17142 ^ n17129 ;
  assign n17131 = n17129 ^ n15654 ;
  assign n17130 = n17129 ^ n15689 ;
  assign n17132 = n17131 ^ n17130 ;
  assign n17135 = ~n15590 & n17132 ;
  assign n17136 = n17135 ^ n17131 ;
  assign n17137 = ~n15646 & n17136 ;
  assign n17144 = n17143 ^ n17137 ;
  assign n17146 = n17145 ^ n17144 ;
  assign n17120 = n15683 ^ n15658 ;
  assign n17121 = n15658 ^ n15590 ;
  assign n17122 = n17121 ^ n15658 ;
  assign n17123 = ~n17120 & ~n17122 ;
  assign n17124 = n17123 ^ n15658 ;
  assign n17125 = ~n15621 & ~n17124 ;
  assign n17147 = n17146 ^ n17125 ;
  assign n17151 = n17150 ^ n17147 ;
  assign n17113 = n17112 ^ n15693 ;
  assign n17114 = n15625 ^ n15589 ;
  assign n17115 = n17112 ^ n15589 ;
  assign n17116 = n17115 ^ n15589 ;
  assign n17117 = ~n17114 & ~n17116 ;
  assign n17118 = n17117 ^ n15589 ;
  assign n17119 = ~n17113 & ~n17118 ;
  assign n17152 = n17151 ^ n17119 ;
  assign n17153 = n17152 ^ n15623 ;
  assign n17154 = n17153 ^ n12408 ;
  assign n17155 = n17154 ^ x126 ;
  assign n17156 = n17111 & n17155 ;
  assign n17157 = n17156 ^ n17155 ;
  assign n17158 = n16796 ^ x84 ;
  assign n17159 = n16348 ^ x78 ;
  assign n17160 = n17158 & ~n17159 ;
  assign n17161 = n17160 ^ n17158 ;
  assign n17162 = n17157 & n17161 ;
  assign n17163 = ~n17077 & n17162 ;
  assign n17164 = n17077 ^ n17075 ;
  assign n17165 = n17164 ^ n17074 ;
  assign n17166 = n17160 ^ n17159 ;
  assign n17167 = n17166 ^ n17158 ;
  assign n17186 = n17157 & n17167 ;
  assign n17181 = n17156 & n17161 ;
  assign n17182 = n17181 ^ n17162 ;
  assign n17169 = n17157 ^ n17111 ;
  assign n17170 = n17161 & ~n17169 ;
  assign n17180 = n17170 ^ n17161 ;
  assign n17183 = n17182 ^ n17180 ;
  assign n17176 = n17156 & ~n17166 ;
  assign n17175 = n17111 & ~n17166 ;
  assign n17177 = n17176 ^ n17175 ;
  assign n17173 = n17156 ^ n17111 ;
  assign n17174 = n17160 & n17173 ;
  assign n17178 = n17177 ^ n17174 ;
  assign n17179 = n17178 ^ n17173 ;
  assign n17184 = n17183 ^ n17179 ;
  assign n17185 = n17184 ^ n17170 ;
  assign n17187 = n17186 ^ n17185 ;
  assign n17168 = n17156 & n17167 ;
  assign n17171 = n17170 ^ n17168 ;
  assign n17172 = n17171 ^ n17167 ;
  assign n17188 = n17187 ^ n17172 ;
  assign n17189 = n17165 & n17188 ;
  assign n17190 = ~n17163 & ~n17189 ;
  assign n17913 = n17156 & n17160 ;
  assign n17196 = n17186 ^ n17162 ;
  assign n17194 = n17157 & n17160 ;
  assign n17195 = n17194 ^ n17157 ;
  assign n17197 = n17196 ^ n17195 ;
  assign n17917 = n17913 ^ n17197 ;
  assign n18418 = n17176 ^ n17074 ;
  assign n18419 = n18418 ^ n17176 ;
  assign n18420 = n17917 & ~n18419 ;
  assign n18421 = n18420 ^ n17176 ;
  assign n18422 = ~n17075 & n18421 ;
  assign n18423 = n18422 ^ n17176 ;
  assign n18415 = n17076 & n17182 ;
  assign n18424 = n18423 ^ n18415 ;
  assign n17215 = n17188 ^ n17170 ;
  assign n17212 = n17197 ^ n17160 ;
  assign n17211 = n17175 ^ n17159 ;
  assign n17213 = n17212 ^ n17211 ;
  assign n17214 = n17213 ^ n17169 ;
  assign n17216 = n17215 ^ n17214 ;
  assign n18414 = n17216 ^ n17174 ;
  assign n18425 = n18424 ^ n18414 ;
  assign n17192 = n17075 ^ n17074 ;
  assign n17944 = n17174 ^ n17075 ;
  assign n17945 = n17944 ^ n17174 ;
  assign n17919 = n17194 ^ n17176 ;
  assign n17946 = n17919 ^ n17186 ;
  assign n17947 = n17946 ^ n17174 ;
  assign n17948 = ~n17945 & n17947 ;
  assign n17949 = n17948 ^ n17174 ;
  assign n17950 = n17192 & n17949 ;
  assign n18426 = n18425 ^ n17950 ;
  assign n17953 = n17165 & n17186 ;
  assign n17952 = n17165 & n17183 ;
  assign n17954 = n17953 ^ n17952 ;
  assign n18427 = n18426 ^ n17954 ;
  assign n18408 = n17213 ^ n17174 ;
  assign n18409 = n18408 ^ n17181 ;
  assign n18410 = n18409 ^ n17174 ;
  assign n18411 = ~n17945 & ~n18410 ;
  assign n18412 = n18411 ^ n17174 ;
  assign n18413 = n17192 & n18412 ;
  assign n18428 = n18427 ^ n18413 ;
  assign n17225 = n17216 ^ n17177 ;
  assign n17926 = n17225 ^ n17168 ;
  assign n18401 = n17926 ^ n17188 ;
  assign n18402 = n18401 ^ n17187 ;
  assign n18403 = n17187 ^ n17075 ;
  assign n18404 = n18403 ^ n17187 ;
  assign n18405 = n18402 & n18404 ;
  assign n18406 = n18405 ^ n17187 ;
  assign n18407 = ~n17074 & n18406 ;
  assign n18429 = n18428 ^ n18407 ;
  assign n17918 = n17917 ^ n17162 ;
  assign n18396 = n17216 ^ n17074 ;
  assign n18397 = n18396 ^ n17216 ;
  assign n18398 = n17918 & n18397 ;
  assign n18399 = n18398 ^ n17216 ;
  assign n18400 = n17075 & n18399 ;
  assign n18430 = n18429 ^ n18400 ;
  assign n17234 = n17164 & n17185 ;
  assign n18431 = n18430 ^ n17234 ;
  assign n18432 = n17190 & ~n18431 ;
  assign n18433 = n18432 ^ n13100 ;
  assign n19111 = n18433 ^ x74 ;
  assign n19181 = n19111 ^ n19110 ;
  assign n19182 = ~n19170 & ~n19181 ;
  assign n19178 = n19111 & n19177 ;
  assign n19179 = n19178 ^ n19177 ;
  assign n19112 = n19110 & n19111 ;
  assign n19173 = n19112 & ~n19170 ;
  assign n19180 = n19179 ^ n19173 ;
  assign n19183 = n19182 ^ n19180 ;
  assign n19249 = n19248 ^ n19183 ;
  assign n19206 = n19177 ^ n19171 ;
  assign n19172 = n19112 & n19171 ;
  assign n19212 = n19206 ^ n19172 ;
  assign n19270 = n19249 ^ n19212 ;
  assign n17735 = n15494 ^ x76 ;
  assign n17734 = n16541 ^ x93 ;
  assign n17824 = n17735 ^ n17734 ;
  assign n17737 = n15986 ^ x94 ;
  assign n17747 = n16753 ^ n16656 ;
  assign n17749 = n16753 ^ n16737 ;
  assign n17748 = n16753 ^ n16716 ;
  assign n17750 = n17749 ^ n17748 ;
  assign n17751 = n17749 ^ n16657 ;
  assign n17752 = n17751 ^ n17749 ;
  assign n17753 = ~n17750 & ~n17752 ;
  assign n17754 = n17753 ^ n17749 ;
  assign n17755 = ~n17747 & ~n17754 ;
  assign n17756 = n17755 ^ n16656 ;
  assign n17740 = n17316 ^ n16729 ;
  assign n17738 = n16741 ^ n16737 ;
  assign n17739 = n17738 ^ n16789 ;
  assign n17741 = n17740 ^ n17739 ;
  assign n17742 = n17739 ^ n16657 ;
  assign n17743 = n17742 ^ n17739 ;
  assign n17744 = n17741 & ~n17743 ;
  assign n17745 = n17744 ^ n17739 ;
  assign n17746 = ~n16656 & ~n17745 ;
  assign n17757 = n17756 ^ n17746 ;
  assign n17758 = n17757 ^ n16718 ;
  assign n17759 = ~n17313 & ~n17758 ;
  assign n17760 = n16657 & n16743 ;
  assign n17761 = n17760 ^ n16742 ;
  assign n17763 = n17761 ^ n16734 ;
  assign n17762 = n17761 ^ n16747 ;
  assign n17764 = n17763 ^ n17762 ;
  assign n17767 = ~n16657 & n17764 ;
  assign n17768 = n17767 ^ n17763 ;
  assign n17769 = ~n16756 & n17768 ;
  assign n17770 = n17769 ^ n17761 ;
  assign n17771 = n17759 & ~n17770 ;
  assign n17772 = ~n16793 & n17771 ;
  assign n17773 = ~n17336 & n17772 ;
  assign n17774 = n17773 ^ n14419 ;
  assign n17775 = n17774 ^ x69 ;
  assign n17776 = n17737 & ~n17775 ;
  assign n17777 = n17776 ^ n17737 ;
  assign n17778 = n17777 ^ n17775 ;
  assign n17780 = n16305 ^ x83 ;
  assign n17801 = n15590 & ~n17148 ;
  assign n17798 = n15641 & ~n17149 ;
  assign n17794 = n15685 ^ n15672 ;
  assign n17795 = ~n17261 & ~n17794 ;
  assign n17789 = n15693 ^ n15658 ;
  assign n17790 = ~n15622 & ~n17789 ;
  assign n17788 = ~n15640 & n15711 ;
  assign n17791 = n17790 ^ n17788 ;
  assign n17792 = n15621 & ~n17791 ;
  assign n17785 = n17125 ^ n15682 ;
  assign n17786 = n17785 ^ n17142 ;
  assign n17787 = n17786 ^ n14444 ;
  assign n17793 = n17792 ^ n17787 ;
  assign n17796 = n17795 ^ n17793 ;
  assign n17783 = n15689 ^ n15664 ;
  assign n17784 = n17112 & n17783 ;
  assign n17797 = n17796 ^ n17784 ;
  assign n17799 = n17798 ^ n17797 ;
  assign n17781 = n17148 ^ n15669 ;
  assign n17782 = n15621 & ~n17781 ;
  assign n17800 = n17799 ^ n17782 ;
  assign n17802 = n17801 ^ n17800 ;
  assign n17803 = n17802 ^ x117 ;
  assign n17804 = ~n17780 & n17803 ;
  assign n17805 = n17804 ^ n17780 ;
  assign n17815 = n17805 ^ n17803 ;
  assign n17851 = n17778 & n17815 ;
  assign n17779 = n17778 ^ n17737 ;
  assign n17831 = ~n17779 & n17804 ;
  assign n17832 = n17831 ^ n17804 ;
  assign n17829 = n17776 & n17804 ;
  assign n17817 = n17777 & n17804 ;
  assign n17830 = n17829 ^ n17817 ;
  assign n17833 = n17832 ^ n17830 ;
  assign n17852 = n17851 ^ n17833 ;
  assign n17807 = n17804 ^ n17803 ;
  assign n17827 = n17776 & n17807 ;
  assign n17893 = n17852 ^ n17827 ;
  assign n17894 = n17827 ^ n17734 ;
  assign n17895 = n17894 ^ n17827 ;
  assign n17896 = n17893 & n17895 ;
  assign n17897 = n17896 ^ n17827 ;
  assign n17898 = n17824 & n17897 ;
  assign n17808 = ~n17779 & n17807 ;
  assign n17806 = ~n17779 & ~n17805 ;
  assign n17809 = n17808 ^ n17806 ;
  assign n17838 = n17831 ^ n17809 ;
  assign n18320 = n17838 ^ n17829 ;
  assign n17839 = n17838 ^ n17779 ;
  assign n17840 = n17839 ^ n17806 ;
  assign n17834 = n17803 ^ n17775 ;
  assign n17835 = n17775 ^ n17737 ;
  assign n17836 = ~n17834 & ~n17835 ;
  assign n17837 = n17836 ^ n17817 ;
  assign n17841 = n17840 ^ n17837 ;
  assign n17842 = n17841 ^ n17777 ;
  assign n17816 = n17777 & n17815 ;
  assign n17818 = n17817 ^ n17816 ;
  assign n17843 = n17842 ^ n17818 ;
  assign n18319 = n17843 ^ n17817 ;
  assign n18321 = n18320 ^ n18319 ;
  assign n18322 = n18320 ^ n17735 ;
  assign n18323 = n18322 ^ n18320 ;
  assign n18324 = ~n18321 & n18323 ;
  assign n18325 = n18324 ^ n18320 ;
  assign n18326 = ~n17734 & n18325 ;
  assign n18327 = n18326 ^ n17829 ;
  assign n17812 = n17778 & n17807 ;
  assign n18318 = n17812 & ~n17824 ;
  assign n18328 = n18327 ^ n18318 ;
  assign n17825 = n17776 & n17815 ;
  assign n17846 = n17829 ^ n17825 ;
  assign n17845 = n17827 ^ n17776 ;
  assign n17847 = n17846 ^ n17845 ;
  assign n17864 = n17847 ^ n17816 ;
  assign n18340 = n17864 ^ n17817 ;
  assign n18337 = n17852 ^ n17840 ;
  assign n18341 = n18340 ^ n18337 ;
  assign n17736 = ~n17734 & n17735 ;
  assign n17884 = n17736 ^ n17734 ;
  assign n18339 = ~n17827 & n17884 ;
  assign n18342 = n18341 ^ n18339 ;
  assign n18343 = n17734 & n18342 ;
  assign n17844 = n17843 ^ n17841 ;
  assign n17848 = n17847 ^ n17844 ;
  assign n18333 = n17848 ^ n17825 ;
  assign n18332 = n17737 & ~n17834 ;
  assign n18334 = n18333 ^ n18332 ;
  assign n18335 = n17734 & n18334 ;
  assign n18336 = n18335 ^ n18332 ;
  assign n18338 = n18337 ^ n18336 ;
  assign n18344 = n18343 ^ n18338 ;
  assign n18345 = n17824 & ~n18344 ;
  assign n18346 = n18345 ^ n18336 ;
  assign n18329 = n17736 ^ n17735 ;
  assign n17900 = n17812 ^ n17778 ;
  assign n17901 = n17900 ^ n17852 ;
  assign n18330 = n17901 ^ n17808 ;
  assign n18331 = n18329 & n18330 ;
  assign n18347 = n18346 ^ n18331 ;
  assign n18348 = ~n18328 & ~n18347 ;
  assign n18349 = ~n17898 & n18348 ;
  assign n18353 = n18349 ^ n14534 ;
  assign n18350 = n17884 ^ n17735 ;
  assign n18351 = ~n17839 & n18350 ;
  assign n18352 = n18349 & n18351 ;
  assign n18354 = n18353 ^ n18352 ;
  assign n19035 = n18354 ^ x115 ;
  assign n19271 = n19249 ^ n19035 ;
  assign n19272 = n19271 ^ n19249 ;
  assign n19273 = ~n19270 & ~n19272 ;
  assign n19274 = n19273 ^ n19249 ;
  assign n19275 = n19073 & ~n19274 ;
  assign n19189 = n19182 ^ n19112 ;
  assign n19190 = n19189 ^ n19110 ;
  assign n19188 = n19173 ^ n19111 ;
  assign n19191 = n19190 ^ n19188 ;
  assign n19192 = n19137 & ~n19191 ;
  assign n19193 = n19192 ^ n19191 ;
  assign n19184 = ~n19111 & ~n19137 ;
  assign n19194 = n19193 ^ n19184 ;
  assign n19186 = n19184 & n19185 ;
  assign n19187 = n19186 ^ n19183 ;
  assign n19195 = n19194 ^ n19187 ;
  assign n19196 = n19195 ^ n19192 ;
  assign n19174 = n19173 ^ n19112 ;
  assign n19175 = n19174 ^ n19172 ;
  assign n19176 = n19175 ^ n19112 ;
  assign n19197 = n19196 ^ n19176 ;
  assign n19198 = n19073 & ~n19197 ;
  assign n19199 = n19198 ^ n19196 ;
  assign n19200 = ~n19035 & ~n19199 ;
  assign n19223 = ~n19137 & n19174 ;
  assign n20674 = n19223 ^ n19178 ;
  assign n20675 = n20674 ^ n19073 ;
  assign n20676 = n20675 ^ n20674 ;
  assign n20677 = n20674 ^ n19186 ;
  assign n20678 = n20677 ^ n20674 ;
  assign n20679 = n20676 & n20678 ;
  assign n20680 = n20679 ^ n20674 ;
  assign n20681 = n19035 & n20680 ;
  assign n19201 = n19073 ^ n19035 ;
  assign n19225 = n19224 ^ n19191 ;
  assign n19226 = n19137 & ~n19225 ;
  assign n19208 = n19186 ^ n19185 ;
  assign n19209 = n19208 ^ n19174 ;
  assign n19231 = n19226 ^ n19209 ;
  assign n20436 = n19231 ^ n19183 ;
  assign n19251 = n19223 ^ n19174 ;
  assign n19227 = n19226 ^ n19225 ;
  assign n20431 = n19251 ^ n19227 ;
  assign n19229 = n19193 ^ n19179 ;
  assign n20435 = n20431 ^ n19229 ;
  assign n20437 = n20436 ^ n20435 ;
  assign n20667 = n20437 ^ n20436 ;
  assign n20668 = n20436 ^ n19073 ;
  assign n20669 = n20668 ^ n20436 ;
  assign n20670 = n20667 & n20669 ;
  assign n20671 = n20670 ^ n20436 ;
  assign n20672 = n19201 & n20671 ;
  assign n20659 = n19227 ^ n19173 ;
  assign n20660 = n20659 ^ n19193 ;
  assign n20661 = n19193 ^ n19035 ;
  assign n20662 = n20661 ^ n19193 ;
  assign n20663 = n20660 & ~n20662 ;
  assign n20664 = n20663 ^ n19193 ;
  assign n20665 = ~n19073 & ~n20664 ;
  assign n19240 = n19035 & ~n19073 ;
  assign n19250 = n19249 ^ n19195 ;
  assign n19252 = n19251 ^ n19250 ;
  assign n19253 = n19240 & n19252 ;
  assign n20657 = n20436 ^ n19253 ;
  assign n20444 = n19196 ^ n19172 ;
  assign n20445 = n19035 & ~n20444 ;
  assign n20446 = n20445 ^ n19196 ;
  assign n19213 = n19212 ^ n19186 ;
  assign n20449 = n20446 ^ n19213 ;
  assign n20450 = n20449 ^ n20446 ;
  assign n20451 = n19035 & n20450 ;
  assign n20452 = n20451 ^ n20446 ;
  assign n20453 = ~n19073 & ~n20452 ;
  assign n20454 = n20453 ^ n20446 ;
  assign n20658 = n20657 ^ n20454 ;
  assign n20666 = n20665 ^ n20658 ;
  assign n20673 = n20672 ^ n20666 ;
  assign n20682 = n20681 ^ n20673 ;
  assign n20683 = ~n19200 & n20682 ;
  assign n20684 = ~n19275 & n20683 ;
  assign n20685 = n20684 ^ n16576 ;
  assign n20686 = n20685 ^ x77 ;
  assign n18026 = n17274 ^ x104 ;
  assign n18027 = n16971 ^ x66 ;
  assign n18028 = n18026 & n18027 ;
  assign n18029 = n18028 ^ n18026 ;
  assign n18030 = n18029 ^ n18027 ;
  assign n18020 = n17435 ^ x81 ;
  assign n17993 = ~n16718 & ~n16755 ;
  assign n18010 = n16764 ^ n16734 ;
  assign n18008 = n17738 ^ n17318 ;
  assign n18009 = ~n16657 & n18008 ;
  assign n18011 = n18010 ^ n18009 ;
  assign n18012 = n16756 & n18011 ;
  assign n18006 = n16659 & ~n16746 ;
  assign n17997 = n16729 ^ n16717 ;
  assign n17998 = n17997 ^ n17318 ;
  assign n17999 = ~n16656 & ~n17998 ;
  assign n18003 = n17999 ^ n16734 ;
  assign n18000 = n17999 ^ n16715 ;
  assign n17995 = n16704 ^ n16698 ;
  assign n17996 = ~n16656 & n17995 ;
  assign n18001 = n18000 ^ n17996 ;
  assign n18002 = n16657 & n18001 ;
  assign n18004 = n18003 ^ n18002 ;
  assign n18005 = n18004 ^ n16764 ;
  assign n18007 = n18006 ^ n18005 ;
  assign n18013 = n18012 ^ n18007 ;
  assign n17994 = n16658 & n16713 ;
  assign n18014 = n18013 ^ n17994 ;
  assign n18015 = ~n17340 & ~n18014 ;
  assign n18016 = ~n17313 & n18015 ;
  assign n18017 = n17993 & n18016 ;
  assign n18018 = n18017 ^ n15228 ;
  assign n18019 = n18018 ^ x107 ;
  assign n18073 = n18020 ^ n18019 ;
  assign n17971 = n16118 ^ n16115 ;
  assign n17981 = n17971 ^ n16123 ;
  assign n17980 = n16146 ^ n16061 ;
  assign n17982 = n17981 ^ n17980 ;
  assign n17983 = n17982 ^ n17094 ;
  assign n17972 = n17971 ^ n16082 ;
  assign n17975 = n17972 ^ n15988 ;
  assign n17976 = n17975 ^ n17972 ;
  assign n17977 = n16097 & ~n17976 ;
  assign n17978 = n17977 ^ n17972 ;
  assign n17979 = n16062 & ~n17978 ;
  assign n17984 = n17983 ^ n17979 ;
  assign n17963 = n16121 ^ n16051 ;
  assign n17964 = n17963 ^ n15988 ;
  assign n17965 = n17964 ^ n17963 ;
  assign n17966 = n17963 ^ n16083 ;
  assign n17967 = n17966 ^ n17963 ;
  assign n17968 = n17965 & ~n17967 ;
  assign n17969 = n17968 ^ n17963 ;
  assign n17970 = n16056 & ~n17969 ;
  assign n17985 = n17984 ^ n17970 ;
  assign n17986 = n17985 ^ n16157 ;
  assign n17987 = n17986 ^ n16289 ;
  assign n17988 = n17987 ^ n15260 ;
  assign n17989 = n17988 ^ x64 ;
  assign n18021 = ~n18019 & n18020 ;
  assign n18022 = n18021 ^ n18020 ;
  assign n18023 = n18022 ^ n18019 ;
  assign n18024 = n18023 ^ n18020 ;
  assign n17990 = n16837 ^ x90 ;
  assign n18069 = n18024 ^ n17990 ;
  assign n18070 = n17989 & n18069 ;
  assign n18074 = n18073 ^ n18070 ;
  assign n18075 = n18074 ^ n18022 ;
  assign n17991 = ~n17989 & n17990 ;
  assign n17992 = n17991 ^ n17989 ;
  assign n18034 = n17992 ^ n17990 ;
  assign n18043 = ~n18024 & n18034 ;
  assign n18050 = n18043 ^ n18034 ;
  assign n18047 = n18021 & n18034 ;
  assign n18039 = n18023 & n18034 ;
  assign n18048 = n18047 ^ n18039 ;
  assign n18051 = n18050 ^ n18048 ;
  assign n18052 = n18051 ^ n18043 ;
  assign n18025 = ~n17992 & ~n18024 ;
  assign n18053 = n18052 ^ n18025 ;
  assign n18054 = n18053 ^ n18048 ;
  assign n18076 = n18075 ^ n18054 ;
  assign n18273 = ~n18030 & ~n18076 ;
  assign n18031 = n18030 ^ n18026 ;
  assign n18044 = n18031 & n18043 ;
  assign n18274 = n18273 ^ n18044 ;
  assign n18063 = n18031 ^ n18029 ;
  assign n18067 = n17991 & n18022 ;
  assign n18033 = n17991 & n18023 ;
  assign n18072 = n18067 ^ n18033 ;
  assign n18077 = n18076 ^ n18072 ;
  assign n18078 = n18077 ^ n17991 ;
  assign n18071 = n18070 ^ n18050 ;
  assign n18079 = n18078 ^ n18071 ;
  assign n18080 = n18079 ^ n18072 ;
  assign n18064 = n18019 ^ n17989 ;
  assign n18065 = n18064 ^ n18020 ;
  assign n18066 = n17990 & n18065 ;
  assign n18068 = n18067 ^ n18066 ;
  assign n18081 = n18080 ^ n18068 ;
  assign n18095 = n18081 ^ n18071 ;
  assign n18035 = n18034 ^ n17989 ;
  assign n18036 = n18021 & n18035 ;
  assign n18094 = n18036 ^ n18035 ;
  assign n18096 = n18095 ^ n18094 ;
  assign n18045 = ~n17992 & n18022 ;
  assign n18695 = n18096 ^ n18045 ;
  assign n18696 = n18063 & ~n18695 ;
  assign n18040 = ~n17992 & n18021 ;
  assign n18086 = n18040 ^ n18025 ;
  assign n18085 = n18045 ^ n17992 ;
  assign n18087 = n18086 ^ n18085 ;
  assign n18266 = n18087 ^ n18051 ;
  assign n18263 = n18027 & n18086 ;
  assign n18264 = n18263 ^ n18025 ;
  assign n18265 = n18264 ^ n18096 ;
  assign n18267 = n18266 ^ n18265 ;
  assign n18268 = n18267 ^ n18264 ;
  assign n18269 = n18027 & n18268 ;
  assign n18270 = n18269 ^ n18265 ;
  assign n18271 = ~n18063 & ~n18270 ;
  assign n18272 = n18271 ^ n18264 ;
  assign n18690 = ~n18030 & n18067 ;
  assign n18691 = ~n18272 & n18690 ;
  assign n18692 = n18691 ^ n18272 ;
  assign n18088 = n18087 ^ n18047 ;
  assign n18688 = ~n18030 & ~n18088 ;
  assign n18037 = n18036 ^ n18033 ;
  assign n18038 = n18029 & n18037 ;
  assign n18689 = n18688 ^ n18038 ;
  assign n18693 = n18692 ^ n18689 ;
  assign n18681 = n18072 ^ n18036 ;
  assign n18682 = n18681 ^ n18066 ;
  assign n18683 = n18066 ^ n18026 ;
  assign n18684 = n18683 ^ n18066 ;
  assign n18685 = n18682 & ~n18684 ;
  assign n18686 = n18685 ^ n18066 ;
  assign n18687 = n18027 & n18686 ;
  assign n18694 = n18693 ^ n18687 ;
  assign n18697 = n18696 ^ n18694 ;
  assign n18680 = n18029 & ~n18078 ;
  assign n18698 = n18697 ^ n18680 ;
  assign n18673 = n18047 ^ n18025 ;
  assign n18672 = n18052 ^ n18036 ;
  assign n18674 = n18673 ^ n18672 ;
  assign n18675 = n18673 ^ n18026 ;
  assign n18676 = n18675 ^ n18673 ;
  assign n18677 = n18674 & ~n18676 ;
  assign n18678 = n18677 ^ n18673 ;
  assign n18679 = ~n18063 & n18678 ;
  assign n18699 = n18698 ^ n18679 ;
  assign n18700 = ~n18274 & ~n18699 ;
  assign n18032 = n18025 & n18031 ;
  assign n18041 = n18040 ^ n18039 ;
  assign n18042 = n18029 & n18041 ;
  assign n18701 = ~n18032 & ~n18042 ;
  assign n18702 = n18700 & n18701 ;
  assign n18703 = n18702 ^ n15380 ;
  assign n19695 = n18703 ^ x104 ;
  assign n19725 = n19072 ^ x81 ;
  assign n16647 = n16624 ^ n16583 ;
  assign n16648 = n16352 & n16647 ;
  assign n16607 = n16606 ^ n16601 ;
  assign n18587 = n16607 ^ n16595 ;
  assign n18588 = ~n16306 & n18587 ;
  assign n18389 = n18368 ^ n16619 ;
  assign n18390 = n16350 & ~n18389 ;
  assign n18589 = n18588 ^ n18390 ;
  assign n18585 = n18368 ^ n16623 ;
  assign n18586 = ~n16615 & ~n18585 ;
  assign n18590 = n18589 ^ n18586 ;
  assign n18359 = n16597 ^ n16583 ;
  assign n18381 = n18359 ^ n16603 ;
  assign n18382 = n18381 ^ n18368 ;
  assign n18584 = n16351 & n18382 ;
  assign n18591 = n18590 ^ n18584 ;
  assign n18577 = n16619 ^ n16597 ;
  assign n18578 = n18577 ^ n16603 ;
  assign n18579 = n16603 ^ n16306 ;
  assign n18580 = n18579 ^ n16603 ;
  assign n18581 = n18578 & ~n18580 ;
  assign n18582 = n18581 ^ n16603 ;
  assign n18583 = n16349 & n18582 ;
  assign n18592 = n18591 ^ n18583 ;
  assign n18594 = n18593 ^ n18592 ;
  assign n18595 = ~n16648 & ~n18594 ;
  assign n18596 = n18595 ^ n15166 ;
  assign n19698 = n18596 ^ x90 ;
  assign n18888 = n17833 ^ n17808 ;
  assign n18901 = n17736 & n18888 ;
  assign n19715 = n17846 ^ n17734 ;
  assign n19716 = n17735 & ~n19715 ;
  assign n17885 = n17851 ^ n17809 ;
  assign n17886 = ~n17884 & n17885 ;
  assign n17865 = n17864 ^ n17829 ;
  assign n17866 = n17735 & ~n17865 ;
  assign n17867 = n17866 ^ n17829 ;
  assign n17868 = n17867 ^ n17734 ;
  assign n17869 = n17868 ^ n17735 ;
  assign n17870 = n17869 ^ n17867 ;
  assign n17871 = n17843 ^ n17735 ;
  assign n17879 = ~n17841 & ~n17871 ;
  assign n17880 = n17879 ^ n17871 ;
  assign n17881 = n17880 ^ n17867 ;
  assign n17882 = n17870 & n17881 ;
  assign n17883 = n17882 ^ n17868 ;
  assign n17887 = n17886 ^ n17883 ;
  assign n17810 = n17809 ^ n17779 ;
  assign n17811 = n17736 & ~n17810 ;
  assign n19713 = n17887 ^ n17811 ;
  assign n19706 = n17901 ^ n17884 ;
  assign n17826 = n17825 ^ n17817 ;
  assign n17828 = n17827 ^ n17826 ;
  assign n19707 = n18329 ^ n17828 ;
  assign n19708 = n17901 ^ n17828 ;
  assign n19709 = n19708 ^ n17828 ;
  assign n19710 = ~n19707 & n19709 ;
  assign n19711 = n19710 ^ n17828 ;
  assign n19712 = ~n19706 & ~n19711 ;
  assign n19714 = n19713 ^ n19712 ;
  assign n19717 = n19716 ^ n19714 ;
  assign n17853 = n17852 ^ n17809 ;
  assign n19701 = n17853 ^ n17816 ;
  assign n19699 = n17836 ^ n17812 ;
  assign n19702 = n19701 ^ n19699 ;
  assign n19703 = ~n17735 & n19702 ;
  assign n19700 = n19699 ^ n17846 ;
  assign n19704 = n19703 ^ n19700 ;
  assign n19705 = n17734 & ~n19704 ;
  assign n19718 = n19717 ^ n19705 ;
  assign n19719 = ~n18901 & n19718 ;
  assign n19720 = n19719 ^ n16046 ;
  assign n19721 = n19720 ^ x107 ;
  assign n19722 = n19698 & n19721 ;
  assign n19770 = n19722 ^ n19721 ;
  assign n19771 = ~n19725 & n19770 ;
  assign n17660 = n15724 ^ x74 ;
  assign n17619 = n15984 ^ n14908 ;
  assign n17615 = ~n15766 & ~n15958 ;
  assign n17607 = n15948 ^ n15934 ;
  assign n17608 = n17607 ^ n15977 ;
  assign n17609 = n17608 ^ n16364 ;
  assign n17610 = n15936 & n17609 ;
  assign n17611 = n17610 ^ n15934 ;
  assign n17612 = n15974 ^ n15936 ;
  assign n17613 = n17611 & n17612 ;
  assign n17603 = n15949 ^ n15915 ;
  assign n17604 = n15767 & ~n17603 ;
  assign n17600 = n15938 ^ n15835 ;
  assign n17601 = ~n15766 & n17600 ;
  assign n17597 = n15942 ^ n15926 ;
  assign n17602 = n17601 ^ n17597 ;
  assign n17605 = n17604 ^ n17602 ;
  assign n17606 = ~n16800 & n17605 ;
  assign n17614 = n17613 ^ n17606 ;
  assign n17616 = n17615 ^ n17614 ;
  assign n17596 = n15934 & n15947 ;
  assign n17617 = n17616 ^ n17596 ;
  assign n17618 = ~n16386 & n17617 ;
  assign n17620 = n17619 ^ n17618 ;
  assign n17621 = n17620 ^ x89 ;
  assign n17538 = n16471 ^ n16465 ;
  assign n17574 = n17433 ^ n16525 ;
  assign n17541 = n16478 ^ n16466 ;
  assign n17542 = n17541 ^ n16493 ;
  assign n17559 = n17542 ^ n17423 ;
  assign n17543 = n17542 ^ n16395 ;
  assign n17544 = n17543 ^ n16466 ;
  assign n17551 = n16511 & ~n17544 ;
  assign n17539 = n16511 ^ n16478 ;
  assign n17540 = n17539 ^ n16493 ;
  assign n17552 = n17551 ^ n17540 ;
  assign n17553 = n16493 ^ n16466 ;
  assign n17547 = n16511 ^ n16466 ;
  assign n17554 = n17551 ^ n17547 ;
  assign n17555 = n17554 ^ n16466 ;
  assign n17556 = n17553 & n17555 ;
  assign n17557 = n17556 ^ n16466 ;
  assign n17558 = ~n17552 & ~n17557 ;
  assign n17560 = n17559 ^ n17558 ;
  assign n17561 = n17560 ^ n17423 ;
  assign n17562 = n16523 & ~n17561 ;
  assign n17563 = n17562 ^ n17423 ;
  assign n17564 = ~n16519 & n17563 ;
  assign n17565 = n17564 ^ n17423 ;
  assign n17566 = n16518 ^ n16464 ;
  assign n17567 = n17566 ^ n17565 ;
  assign n17568 = n16897 ^ n16523 ;
  assign n17569 = ~n16518 & n17568 ;
  assign n17570 = n17569 ^ n16897 ;
  assign n17571 = n17567 & ~n17570 ;
  assign n17572 = n17571 ^ n16518 ;
  assign n17573 = ~n17565 & ~n17572 ;
  assign n17575 = n17574 ^ n17573 ;
  assign n17576 = ~n16888 & n17575 ;
  assign n17577 = n16502 ^ n16474 ;
  assign n17578 = n17577 ^ n16492 ;
  assign n17579 = n16492 ^ n16396 ;
  assign n17580 = n17579 ^ n16492 ;
  assign n17581 = n17578 & n17580 ;
  assign n17582 = n17581 ^ n16492 ;
  assign n17583 = ~n16395 & n17582 ;
  assign n17584 = n17576 & ~n17583 ;
  assign n17585 = ~n16532 & n17584 ;
  assign n17586 = n16519 & n17585 ;
  assign n17587 = n17538 & n17586 ;
  assign n17588 = n17587 ^ n17585 ;
  assign n17590 = n16467 & ~n16511 ;
  assign n17591 = n17588 & n17590 ;
  assign n17589 = n17588 ^ n14872 ;
  assign n17592 = n17591 ^ n17589 ;
  assign n17593 = n17592 ^ x98 ;
  assign n17595 = n17401 ^ x99 ;
  assign n17537 = n16159 ^ x80 ;
  assign n17594 = n17593 ^ n17537 ;
  assign n17633 = n17595 ^ n17594 ;
  assign n17653 = ~n17593 & ~n17633 ;
  assign n17654 = n17653 ^ n17594 ;
  assign n17655 = n17621 & ~n17654 ;
  assign n17656 = n17655 ^ n17633 ;
  assign n17651 = n17621 ^ n17594 ;
  assign n17627 = n17595 ^ n17537 ;
  assign n17628 = n17621 ^ n17593 ;
  assign n17629 = n17595 & n17628 ;
  assign n17630 = n17629 ^ n17593 ;
  assign n17631 = n17627 & n17630 ;
  assign n17652 = n17651 ^ n17631 ;
  assign n17657 = n17656 ^ n17652 ;
  assign n18301 = n17657 ^ n17630 ;
  assign n17648 = n17595 ^ n17593 ;
  assign n17634 = n17621 ^ n17595 ;
  assign n17641 = n17537 & n17593 ;
  assign n17642 = n17634 & n17641 ;
  assign n17643 = n17642 ^ n17629 ;
  assign n17644 = n17643 ^ n17631 ;
  assign n17645 = n17644 ^ n17634 ;
  assign n17637 = n17627 & n17634 ;
  assign n17638 = n17637 ^ n17537 ;
  assign n17639 = n17633 & ~n17638 ;
  assign n17640 = n17639 ^ n17537 ;
  assign n17646 = n17645 ^ n17640 ;
  assign n17632 = n17631 ^ n17595 ;
  assign n17647 = n17646 ^ n17632 ;
  assign n17649 = n17648 ^ n17647 ;
  assign n18302 = n18301 ^ n17649 ;
  assign n19726 = n18302 ^ n17642 ;
  assign n17536 = n17346 ^ x121 ;
  assign n19727 = n19726 ^ n17536 ;
  assign n19728 = n19727 ^ n19726 ;
  assign n19729 = n19726 ^ n18302 ;
  assign n19730 = n17640 & ~n19729 ;
  assign n19731 = n19730 ^ n19726 ;
  assign n19732 = n19728 & ~n19731 ;
  assign n19733 = n19732 ^ n19726 ;
  assign n19734 = n17660 & ~n19733 ;
  assign n19735 = n19734 ^ n17660 ;
  assign n18298 = n17653 ^ n17595 ;
  assign n18299 = ~n17621 & n18298 ;
  assign n18300 = n18299 ^ n17633 ;
  assign n19736 = ~n17660 & n18300 ;
  assign n19737 = n19736 ^ n17642 ;
  assign n19738 = n19737 ^ n17660 ;
  assign n19739 = n19738 ^ n19736 ;
  assign n19740 = n19736 ^ n17645 ;
  assign n19741 = n19740 ^ n19736 ;
  assign n19742 = ~n19739 & n19741 ;
  assign n19743 = n19742 ^ n19736 ;
  assign n19744 = n17536 & n19743 ;
  assign n19745 = n19744 ^ n19736 ;
  assign n19746 = ~n19735 & ~n19745 ;
  assign n19747 = n19746 ^ n16002 ;
  assign n19748 = n19747 ^ x72 ;
  assign n19749 = ~n19725 & n19748 ;
  assign n19750 = n19749 ^ n19725 ;
  assign n19723 = n19722 ^ n19698 ;
  assign n19724 = n19723 ^ n19721 ;
  assign n19756 = n19724 ^ n19698 ;
  assign n19758 = ~n19750 & n19756 ;
  assign n19772 = n19771 ^ n19758 ;
  assign n19765 = n19722 & ~n19750 ;
  assign n19764 = n19722 & n19749 ;
  assign n19766 = n19765 ^ n19764 ;
  assign n19751 = n19750 ^ n19748 ;
  assign n19752 = ~n19724 & n19751 ;
  assign n19762 = n19752 ^ n19724 ;
  assign n19755 = n19749 ^ n19748 ;
  assign n19760 = ~n19724 & n19755 ;
  assign n19759 = ~n19724 & ~n19750 ;
  assign n19761 = n19760 ^ n19759 ;
  assign n19763 = n19762 ^ n19761 ;
  assign n19767 = n19766 ^ n19763 ;
  assign n19773 = n19772 ^ n19767 ;
  assign n19774 = n19773 ^ n19756 ;
  assign n19768 = n19767 ^ n19758 ;
  assign n19757 = n19755 & n19756 ;
  assign n19769 = n19768 ^ n19757 ;
  assign n19775 = n19774 ^ n19769 ;
  assign n19754 = n19723 & n19751 ;
  assign n19776 = n19775 ^ n19754 ;
  assign n19753 = n19752 ^ n19751 ;
  assign n19777 = n19776 ^ n19753 ;
  assign n20274 = n19777 ^ n19772 ;
  assign n19694 = n19169 ^ x114 ;
  assign n20275 = n19772 ^ n19694 ;
  assign n20276 = n20275 ^ n19772 ;
  assign n20277 = n20274 & ~n20276 ;
  assign n20278 = n20277 ^ n19772 ;
  assign n20279 = n19695 & n20278 ;
  assign n19696 = n19695 ^ n19694 ;
  assign n19835 = n19777 ^ n19757 ;
  assign n19836 = n19757 ^ n19694 ;
  assign n19837 = n19836 ^ n19757 ;
  assign n19838 = n19835 & n19837 ;
  assign n19839 = n19838 ^ n19757 ;
  assign n19840 = n19696 & n19839 ;
  assign n20725 = n20279 ^ n19840 ;
  assign n19824 = n19760 ^ n19754 ;
  assign n19825 = n19694 & n19824 ;
  assign n19786 = n19777 ^ n19722 ;
  assign n19787 = n19786 ^ n19766 ;
  assign n20717 = n19825 ^ n19787 ;
  assign n19782 = n19765 ^ n19750 ;
  assign n19809 = n19782 ^ n19725 ;
  assign n19810 = n19809 ^ n19773 ;
  assign n19811 = n19810 ^ n19772 ;
  assign n20696 = n19811 ^ n19758 ;
  assign n20706 = n20696 ^ n19763 ;
  assign n19781 = n19759 ^ n19758 ;
  assign n19783 = n19782 ^ n19781 ;
  assign n19784 = n19783 ^ n19764 ;
  assign n19785 = n19784 ^ n19763 ;
  assign n20694 = n19785 ^ n19757 ;
  assign n20695 = n20694 ^ n19763 ;
  assign n20697 = n20696 ^ n20695 ;
  assign n20700 = ~n20694 & n20697 ;
  assign n20707 = n20706 ^ n20700 ;
  assign n20698 = n20697 ^ n20696 ;
  assign n20702 = n20700 ^ n20698 ;
  assign n20703 = n19694 & ~n20702 ;
  assign n20704 = n20703 ^ n20696 ;
  assign n20705 = ~n19695 & ~n20704 ;
  assign n20708 = n20707 ^ n20705 ;
  assign n20718 = n20717 ^ n20708 ;
  assign n20026 = n19765 ^ n19763 ;
  assign n20711 = n20026 ^ n19811 ;
  assign n19788 = n19787 ^ n19761 ;
  assign n20709 = n19788 ^ n19759 ;
  assign n20710 = n20709 ^ n19776 ;
  assign n20712 = n20711 ^ n20710 ;
  assign n20713 = ~n19694 & n20712 ;
  assign n20714 = n20713 ^ n20710 ;
  assign n20715 = n19695 & n20714 ;
  assign n20716 = ~n20708 & n20715 ;
  assign n20719 = n20718 ^ n20716 ;
  assign n19697 = ~n19694 & n19695 ;
  assign n19794 = n19697 ^ n19696 ;
  assign n19832 = n19794 ^ n19695 ;
  assign n19789 = n19788 ^ n19785 ;
  assign n19790 = n19789 ^ n19769 ;
  assign n19780 = n19748 ^ n19725 ;
  assign n19791 = n19790 ^ n19780 ;
  assign n20022 = n19791 ^ n19775 ;
  assign n20692 = n20022 ^ n19783 ;
  assign n20693 = ~n19832 & ~n20692 ;
  assign n20720 = n20719 ^ n20693 ;
  assign n20726 = n20725 ^ n20720 ;
  assign n20727 = n20726 ^ n17110 ;
  assign n20688 = n19759 ^ n19754 ;
  assign n20687 = n20026 ^ n19810 ;
  assign n20689 = n20688 ^ n20687 ;
  assign n20690 = ~n19694 & n20689 ;
  assign n20691 = n20690 ^ n20687 ;
  assign n20721 = n20720 ^ n20717 ;
  assign n20722 = n20691 & ~n20721 ;
  assign n20723 = n20722 ^ n20717 ;
  assign n20724 = n19695 & n20723 ;
  assign n20728 = n20727 ^ n20724 ;
  assign n20729 = n20728 ^ x108 ;
  assign n18434 = n18433 ^ x99 ;
  assign n18388 = n16648 ^ n15620 ;
  assign n18391 = n18390 ^ n18388 ;
  assign n18367 = n16623 ^ n16351 ;
  assign n16640 = n16624 ^ n16595 ;
  assign n18369 = n18368 ^ n16640 ;
  assign n18370 = n18369 ^ n16352 ;
  assign n18373 = ~n16623 & n18370 ;
  assign n18374 = n18373 ^ n16352 ;
  assign n18375 = n18367 & n18374 ;
  assign n18376 = n18375 ^ n16351 ;
  assign n18360 = n18359 ^ n16598 ;
  assign n18361 = n18360 ^ n16617 ;
  assign n18362 = n16617 ^ n16306 ;
  assign n18363 = n18362 ^ n16617 ;
  assign n18364 = n18361 & n18363 ;
  assign n18365 = n18364 ^ n16617 ;
  assign n18366 = n16349 & n18365 ;
  assign n18377 = n18376 ^ n18366 ;
  assign n18379 = n18378 ^ n16306 ;
  assign n18380 = n18379 ^ n18378 ;
  assign n18383 = ~n16349 & n18382 ;
  assign n18384 = n18383 ^ n18378 ;
  assign n18385 = ~n18380 & n18384 ;
  assign n18386 = n18385 ^ n18378 ;
  assign n18387 = ~n18377 & ~n18386 ;
  assign n18392 = n18391 ^ n18387 ;
  assign n18393 = n18392 ^ x121 ;
  assign n18435 = n18434 ^ n18393 ;
  assign n18245 = n15987 & ~n16216 ;
  assign n18237 = n16183 ^ n16174 ;
  assign n18238 = n18237 ^ n16184 ;
  assign n18239 = n18238 ^ n16185 ;
  assign n18240 = ~n16167 & n18239 ;
  assign n18241 = n18240 ^ n16185 ;
  assign n18242 = n16168 ^ n16167 ;
  assign n18243 = n18241 & ~n18242 ;
  assign n16162 = n15727 & n16161 ;
  assign n18232 = n16162 & n16173 ;
  assign n18225 = n16206 ^ n16160 ;
  assign n18226 = n18225 ^ n16206 ;
  assign n18227 = n16206 ^ n16200 ;
  assign n18228 = n18227 ^ n16206 ;
  assign n18229 = n18226 & n18228 ;
  assign n18230 = n18229 ^ n16206 ;
  assign n18231 = ~n18224 & n18230 ;
  assign n18233 = n18232 ^ n18231 ;
  assign n16252 = ~n16169 & ~n16211 ;
  assign n16253 = n16252 ^ n16251 ;
  assign n18222 = n18221 ^ n16253 ;
  assign n18214 = n16215 ^ n16167 ;
  assign n18223 = n18222 ^ n18214 ;
  assign n18234 = n18233 ^ n18223 ;
  assign n16238 = n16216 ^ n16183 ;
  assign n16239 = n16238 ^ n16191 ;
  assign n16240 = n16191 ^ n16160 ;
  assign n16241 = n16240 ^ n16191 ;
  assign n16242 = ~n16239 & n16241 ;
  assign n16243 = n16242 ^ n16191 ;
  assign n16244 = ~n15987 & n16243 ;
  assign n18235 = n18234 ^ n16244 ;
  assign n18236 = n18235 ^ n15586 ;
  assign n18244 = n18243 ^ n18236 ;
  assign n18246 = n18245 ^ n18244 ;
  assign n18207 = n16219 ^ n16215 ;
  assign n18205 = n16216 ^ n16215 ;
  assign n18208 = n18207 ^ n18205 ;
  assign n18209 = n18205 ^ n15987 ;
  assign n18210 = n18209 ^ n18205 ;
  assign n18211 = n18208 & ~n18210 ;
  assign n18212 = n18211 ^ n18205 ;
  assign n18213 = ~n16160 & n18212 ;
  assign n18247 = n18246 ^ n18213 ;
  assign n18248 = n18247 ^ x106 ;
  assign n18291 = n18028 & ~n18086 ;
  assign n18256 = n18081 ^ n18047 ;
  assign n18286 = n18256 ^ n18041 ;
  assign n18276 = n18076 ^ n17990 ;
  assign n18277 = n18276 ^ n18067 ;
  assign n18278 = n18027 & ~n18277 ;
  assign n18279 = n18278 ^ n18080 ;
  assign n18287 = n18286 ^ n18279 ;
  assign n18282 = n18077 ^ n18041 ;
  assign n18283 = n18282 ^ n18071 ;
  assign n18284 = n18283 ^ n18256 ;
  assign n18285 = n18027 & n18284 ;
  assign n18288 = n18287 ^ n18285 ;
  assign n18289 = ~n18026 & ~n18288 ;
  assign n18275 = n18274 ^ n18272 ;
  assign n18280 = n18279 ^ n18275 ;
  assign n18281 = n18280 ^ n15536 ;
  assign n18290 = n18289 ^ n18281 ;
  assign n18292 = n18291 ^ n18290 ;
  assign n18255 = n18039 ^ n18029 ;
  assign n18257 = n18256 ^ n18031 ;
  assign n18260 = ~n18039 & n18257 ;
  assign n18261 = n18260 ^ n18031 ;
  assign n18262 = n18255 & n18261 ;
  assign n18293 = n18292 ^ n18262 ;
  assign n18249 = n18051 ^ n18037 ;
  assign n18250 = n18037 ^ n18027 ;
  assign n18251 = n18250 ^ n18037 ;
  assign n18252 = n18249 & n18251 ;
  assign n18253 = n18252 ^ n18037 ;
  assign n18254 = ~n18026 & n18253 ;
  assign n18294 = n18293 ^ n18254 ;
  assign n18295 = n18294 ^ x80 ;
  assign n18296 = n18248 & n18295 ;
  assign n18297 = n18296 ^ n18248 ;
  assign n18303 = n18302 ^ n18300 ;
  assign n18304 = n17660 & ~n18303 ;
  assign n18305 = n18304 ^ n18302 ;
  assign n18307 = n18305 ^ n17645 ;
  assign n18306 = n18305 ^ n17640 ;
  assign n18308 = n18307 ^ n18306 ;
  assign n18311 = ~n17660 & n18308 ;
  assign n18312 = n18311 ^ n18307 ;
  assign n18313 = n17536 & ~n18312 ;
  assign n18314 = n18313 ^ n18305 ;
  assign n18315 = ~n17642 & ~n18314 ;
  assign n18316 = n18315 ^ n15558 ;
  assign n18317 = n18316 ^ x97 ;
  assign n18355 = n18354 ^ x66 ;
  assign n18356 = n18317 & n18355 ;
  assign n18440 = n18356 ^ n18355 ;
  assign n18447 = n18297 & n18440 ;
  assign n18446 = n18296 & n18440 ;
  assign n18448 = n18447 ^ n18446 ;
  assign n18436 = n18297 ^ n18295 ;
  assign n18444 = ~n18436 & n18440 ;
  assign n18445 = n18444 ^ n18440 ;
  assign n18449 = n18448 ^ n18445 ;
  assign n18487 = n18449 ^ n18434 ;
  assign n18488 = n18487 ^ n18449 ;
  assign n18466 = n18356 & ~n18436 ;
  assign n18494 = n18466 ^ n18449 ;
  assign n18495 = ~n18488 & n18494 ;
  assign n18496 = n18495 ^ n18449 ;
  assign n18497 = ~n18435 & n18496 ;
  assign n18441 = n18440 ^ n18317 ;
  assign n18454 = n18297 & ~n18441 ;
  assign n20733 = n18454 ^ n18444 ;
  assign n18455 = n18454 ^ n18448 ;
  assign n18443 = n18296 & ~n18441 ;
  assign n18450 = n18449 ^ n18443 ;
  assign n18442 = ~n18436 & ~n18441 ;
  assign n18451 = n18450 ^ n18442 ;
  assign n18452 = n18451 ^ n18444 ;
  assign n18453 = n18452 ^ n18317 ;
  assign n18456 = n18455 ^ n18453 ;
  assign n20734 = n20733 ^ n18456 ;
  assign n18357 = n18356 ^ n18317 ;
  assign n18358 = n18297 & n18357 ;
  assign n18462 = n18455 ^ n18358 ;
  assign n18461 = n18446 ^ n18297 ;
  assign n18463 = n18462 ^ n18461 ;
  assign n18457 = n18456 ^ n18449 ;
  assign n18437 = n18436 ^ n18248 ;
  assign n18438 = n18357 & n18437 ;
  assign n18439 = n18438 ^ n18437 ;
  assign n18458 = n18457 ^ n18439 ;
  assign n18468 = n18463 ^ n18458 ;
  assign n18467 = n18466 ^ n18356 ;
  assign n18469 = n18468 ^ n18467 ;
  assign n19653 = n18469 ^ n18358 ;
  assign n18460 = n18357 & ~n18436 ;
  assign n19654 = n19653 ^ n18460 ;
  assign n20731 = n19654 ^ n18456 ;
  assign n20732 = ~n18393 & n20731 ;
  assign n20735 = n20734 ^ n20732 ;
  assign n20738 = ~n18434 & ~n20735 ;
  assign n20730 = n19654 ^ n18447 ;
  assign n20736 = n20735 ^ n20730 ;
  assign n20737 = ~n18393 & n20736 ;
  assign n20739 = n20738 ^ n20737 ;
  assign n20740 = n20739 ^ n18447 ;
  assign n20747 = n18468 ^ n18438 ;
  assign n18478 = n18469 ^ n18296 ;
  assign n18473 = n18446 ^ n18443 ;
  assign n18479 = n18478 ^ n18473 ;
  assign n18480 = n18479 ^ n18447 ;
  assign n18509 = n18393 & ~n18480 ;
  assign n18510 = n18509 ^ n18447 ;
  assign n18513 = n18510 ^ n18438 ;
  assign n18514 = n18513 ^ n18510 ;
  assign n18515 = ~n18393 & n18514 ;
  assign n18516 = n18515 ^ n18510 ;
  assign n18517 = n18434 & n18516 ;
  assign n18518 = n18517 ^ n18510 ;
  assign n18464 = n18463 ^ n18460 ;
  assign n18500 = n18393 & n18434 ;
  assign n18507 = n18500 ^ n18434 ;
  assign n18508 = n18464 & n18507 ;
  assign n18519 = n18518 ^ n18508 ;
  assign n20748 = n20747 ^ n18519 ;
  assign n20743 = n18454 ^ n18450 ;
  assign n20744 = n20743 ^ n18438 ;
  assign n20745 = n20744 ^ n18468 ;
  assign n20746 = ~n18393 & ~n20745 ;
  assign n20749 = n20748 ^ n20746 ;
  assign n19681 = n18479 ^ n18466 ;
  assign n19682 = n18466 ^ n18393 ;
  assign n19683 = n19682 ^ n18466 ;
  assign n19684 = ~n19681 & n19683 ;
  assign n19685 = n19684 ^ n18466 ;
  assign n19686 = n18434 & n19685 ;
  assign n20758 = n20749 ^ n19686 ;
  assign n20750 = n20749 ^ n18519 ;
  assign n20751 = n20750 ^ n19654 ;
  assign n20752 = n20751 ^ n20750 ;
  assign n20753 = n20750 ^ n18393 ;
  assign n20754 = n20753 ^ n20750 ;
  assign n20755 = ~n20752 & n20754 ;
  assign n20756 = n20755 ^ n20750 ;
  assign n20757 = n18434 & ~n20756 ;
  assign n20759 = n20758 ^ n20757 ;
  assign n20230 = n18442 ^ n18438 ;
  assign n20742 = n18500 & n20230 ;
  assign n20760 = n20759 ^ n20742 ;
  assign n20741 = n18473 & n18507 ;
  assign n20761 = n20760 ^ n20741 ;
  assign n20762 = ~n20740 & n20761 ;
  assign n20763 = ~n18497 & n20762 ;
  assign n20764 = n20763 ^ n17154 ;
  assign n20765 = n20764 ^ x94 ;
  assign n20766 = n20729 & n20765 ;
  assign n20767 = n20766 ^ n20765 ;
  assign n17849 = n17848 ^ n17833 ;
  assign n17850 = n17849 ^ n17829 ;
  assign n17854 = n17853 ^ n17850 ;
  assign n17855 = n17734 & n17854 ;
  assign n17856 = n17855 ^ n17849 ;
  assign n17888 = n17856 ^ n17812 ;
  assign n17889 = n17888 ^ n17887 ;
  assign n17857 = n17856 ^ n17828 ;
  assign n17858 = n17857 ^ n17856 ;
  assign n17859 = n17856 ^ n17735 ;
  assign n17860 = n17859 ^ n17856 ;
  assign n17861 = n17858 & ~n17860 ;
  assign n17862 = n17861 ^ n17856 ;
  assign n17863 = n17824 & n17862 ;
  assign n17890 = n17889 ^ n17863 ;
  assign n17813 = n17812 ^ n17735 ;
  assign n17814 = n17813 ^ n17812 ;
  assign n17821 = n17814 & n17818 ;
  assign n17822 = n17821 ^ n17812 ;
  assign n17823 = ~n17734 & n17822 ;
  assign n17891 = n17890 ^ n17823 ;
  assign n17892 = ~n17811 & ~n17891 ;
  assign n17899 = n17892 & ~n17898 ;
  assign n17902 = n17901 ^ n17831 ;
  assign n17903 = n17831 ^ n17734 ;
  assign n17904 = n17903 ^ n17831 ;
  assign n17905 = n17902 & ~n17904 ;
  assign n17906 = n17905 ^ n17831 ;
  assign n17907 = n17824 & n17906 ;
  assign n17908 = n17899 & ~n17907 ;
  assign n17909 = n17908 ^ n15832 ;
  assign n17910 = n17909 ^ x100 ;
  assign n17473 = n17465 ^ n17374 ;
  assign n17474 = n17473 ^ n17442 ;
  assign n17475 = n17474 ^ n17402 ;
  assign n17476 = ~n17472 & ~n17475 ;
  assign n17477 = n17476 ^ n17402 ;
  assign n17480 = n17461 ^ n17365 ;
  assign n17481 = n17480 ^ n17360 ;
  assign n17478 = n17365 ^ n17360 ;
  assign n17479 = n17478 ^ n17474 ;
  assign n17482 = n17481 ^ n17479 ;
  assign n17483 = ~n17477 & ~n17482 ;
  assign n17484 = n17483 ^ n17481 ;
  assign n17515 = n17514 ^ n17484 ;
  assign n17516 = n17515 ^ n17506 ;
  assign n17489 = n17358 ^ n17347 ;
  assign n17490 = n17489 ^ n17447 ;
  assign n17491 = n17490 ^ n17373 ;
  assign n17492 = n17491 ^ n17311 ;
  assign n17493 = n17492 ^ n17484 ;
  assign n17486 = n17485 ^ n17374 ;
  assign n17487 = n17486 ^ n17457 ;
  assign n17488 = n17487 ^ n17484 ;
  assign n17494 = n17493 ^ n17488 ;
  assign n17495 = n17493 ^ n17436 ;
  assign n17496 = n17495 ^ n17493 ;
  assign n17497 = n17494 & n17496 ;
  assign n17498 = n17497 ^ n17493 ;
  assign n17499 = ~n17472 & n17498 ;
  assign n17517 = n17516 ^ n17499 ;
  assign n17471 = n17437 & ~n17448 ;
  assign n17518 = n17517 ^ n17471 ;
  assign n17519 = n17518 ^ n17470 ;
  assign n17520 = n17519 ^ n14781 ;
  assign n17440 = ~n17378 & n17439 ;
  assign n17521 = n17520 ^ n17440 ;
  assign n17911 = n17521 ^ x109 ;
  assign n18175 = n17910 & n17911 ;
  assign n18089 = n18029 & ~n18088 ;
  assign n18082 = n18081 ^ n18076 ;
  assign n18083 = n18063 & n18082 ;
  assign n18046 = n18045 ^ n18027 ;
  assign n18049 = n18048 ^ n18045 ;
  assign n18055 = n18054 ^ n18049 ;
  assign n18056 = n18055 ^ n18049 ;
  assign n18057 = n18049 ^ n18026 ;
  assign n18058 = n18057 ^ n18049 ;
  assign n18059 = n18056 & n18058 ;
  assign n18060 = n18059 ^ n18049 ;
  assign n18061 = n18046 & ~n18060 ;
  assign n18062 = n18061 ^ n18027 ;
  assign n18084 = n18083 ^ n18062 ;
  assign n18090 = n18089 ^ n18084 ;
  assign n18091 = ~n18044 & ~n18090 ;
  assign n18092 = ~n18042 & n18091 ;
  assign n18099 = n18074 ^ n18027 ;
  assign n18093 = n18076 ^ n17991 ;
  assign n18097 = n18096 ^ n18093 ;
  assign n18098 = n18027 & n18097 ;
  assign n18100 = n18099 ^ n18098 ;
  assign n18101 = n18098 ^ n18026 ;
  assign n18102 = n18101 ^ n18098 ;
  assign n18103 = n18100 & ~n18102 ;
  assign n18104 = n18103 ^ n18098 ;
  assign n18105 = n18092 & ~n18104 ;
  assign n18106 = ~n18038 & n18105 ;
  assign n18107 = ~n18032 & n18106 ;
  assign n18108 = n18107 ^ n15765 ;
  assign n18109 = n18108 ^ x126 ;
  assign n16260 = n16259 ^ n16253 ;
  assign n16261 = n16260 ^ n16244 ;
  assign n16262 = n16261 ^ n15001 ;
  assign n16170 = n16167 & ~n16169 ;
  assign n16163 = ~n15102 & n16162 ;
  assign n16171 = n16170 ^ n16163 ;
  assign n16230 = n16218 ^ n16174 ;
  assign n16222 = n16169 ^ n15725 ;
  assign n16223 = n16222 ^ n16200 ;
  assign n16224 = n16223 ^ n16169 ;
  assign n16225 = n16185 ^ n16169 ;
  assign n16226 = n16225 ^ n16169 ;
  assign n16227 = ~n16224 & ~n16226 ;
  assign n16228 = n16227 ^ n16169 ;
  assign n16229 = ~n16221 & ~n16228 ;
  assign n16231 = n16185 & n16229 ;
  assign n16232 = n16230 & n16231 ;
  assign n16233 = n16232 ^ n16229 ;
  assign n16188 = n16187 ^ n16166 ;
  assign n16195 = n16194 ^ n16188 ;
  assign n16196 = ~n16168 & n16195 ;
  assign n16234 = n16233 ^ n16196 ;
  assign n16186 = n16184 & ~n16185 ;
  assign n16235 = n16234 ^ n16186 ;
  assign n16177 = n16174 ^ n15101 ;
  assign n16178 = n16177 ^ n16174 ;
  assign n16179 = n15495 & n16178 ;
  assign n16180 = n16179 ^ n16174 ;
  assign n16181 = n16161 & n16180 ;
  assign n16236 = n16235 ^ n16181 ;
  assign n16237 = ~n16171 & ~n16236 ;
  assign n16263 = n16262 ^ n16237 ;
  assign n18110 = n16263 ^ x69 ;
  assign n18111 = n18109 & n18110 ;
  assign n18112 = n18111 ^ n18110 ;
  assign n17920 = n17919 ^ n17184 ;
  assign n17921 = n17920 ^ n17188 ;
  assign n17922 = n17075 & n17921 ;
  assign n17923 = n17922 ^ n17215 ;
  assign n17914 = n17913 ^ n17213 ;
  assign n17939 = n17923 ^ n17914 ;
  assign n17209 = n17183 ^ n17075 ;
  assign n17210 = n17209 ^ n17183 ;
  assign n17217 = n17216 ^ n17183 ;
  assign n17936 = n17210 & n17217 ;
  assign n17937 = n17936 ^ n17183 ;
  assign n17938 = n17192 & n17937 ;
  assign n17940 = n17939 ^ n17938 ;
  assign n17191 = n17076 & n17171 ;
  assign n17941 = n17940 ^ n17191 ;
  assign n17925 = n17184 ^ n17181 ;
  assign n17927 = n17926 ^ n17925 ;
  assign n17928 = n17927 ^ n17923 ;
  assign n17924 = n17923 ^ n17918 ;
  assign n17929 = n17928 ^ n17924 ;
  assign n17930 = n17928 ^ n17075 ;
  assign n17931 = n17930 ^ n17928 ;
  assign n17932 = n17929 & n17931 ;
  assign n17933 = n17932 ^ n17928 ;
  assign n17934 = ~n17074 & n17933 ;
  assign n17942 = n17941 ^ n17934 ;
  assign n17193 = n17184 ^ n17174 ;
  assign n17198 = n17197 ^ n17193 ;
  assign n17199 = ~n17075 & n17198 ;
  assign n17200 = n17199 ^ n17184 ;
  assign n17915 = n17914 ^ n17200 ;
  assign n17916 = n17192 & ~n17915 ;
  assign n17943 = n17942 ^ n17916 ;
  assign n17951 = n17943 & ~n17950 ;
  assign n17955 = ~n17163 & ~n17954 ;
  assign n17956 = n17951 & n17955 ;
  assign n17957 = n17956 ^ n16696 ;
  assign n17958 = n17957 ^ x76 ;
  assign n17658 = ~n17536 & n17657 ;
  assign n17659 = n17658 ^ n17656 ;
  assign n17622 = n17595 & ~n17621 ;
  assign n17623 = n17622 ^ n17593 ;
  assign n17624 = n17594 & ~n17623 ;
  assign n17625 = n17624 ^ n17593 ;
  assign n17626 = n17536 & n17625 ;
  assign n17650 = n17649 ^ n17626 ;
  assign n17662 = n17659 ^ n17650 ;
  assign n17663 = n17660 & n17662 ;
  assign n17664 = n17663 ^ n17659 ;
  assign n17959 = n17664 ^ n16701 ;
  assign n17960 = n17959 ^ x86 ;
  assign n17961 = n17958 & ~n17960 ;
  assign n17962 = n17961 ^ n17960 ;
  assign n18114 = n17962 ^ n17958 ;
  assign n18115 = n18114 ^ n17960 ;
  assign n18147 = n18112 & n18115 ;
  assign n18113 = ~n17962 & n18112 ;
  assign n18155 = n18147 ^ n18113 ;
  assign n18153 = n17961 & n18112 ;
  assign n18154 = n18153 ^ n18112 ;
  assign n18156 = n18155 ^ n18154 ;
  assign n18152 = n18111 & n18115 ;
  assign n18157 = n18156 ^ n18152 ;
  assign n18149 = n17961 & n18111 ;
  assign n18150 = n18149 ^ n18147 ;
  assign n18143 = n18110 & n18114 ;
  assign n18151 = n18150 ^ n18143 ;
  assign n18158 = n18157 ^ n18151 ;
  assign n18148 = n18147 ^ n18111 ;
  assign n18159 = n18158 ^ n18148 ;
  assign n19991 = n18159 ^ n18153 ;
  assign n19992 = n18175 & n19991 ;
  assign n20410 = n19992 ^ n16796 ;
  assign n18176 = n18175 ^ n17910 ;
  assign n18116 = n18112 ^ n18109 ;
  assign n18167 = n17961 & ~n18116 ;
  assign n18162 = n18159 ^ n18156 ;
  assign n18163 = n18162 ^ n18149 ;
  assign n18117 = n18115 & ~n18116 ;
  assign n18165 = n18163 ^ n18117 ;
  assign n18140 = n18116 ^ n18110 ;
  assign n18145 = n18114 & n18140 ;
  assign n18144 = n18143 ^ n18114 ;
  assign n18146 = n18145 ^ n18144 ;
  assign n18166 = n18165 ^ n18146 ;
  assign n18168 = n18167 ^ n18166 ;
  assign n18164 = n18163 ^ n18116 ;
  assign n18169 = n18168 ^ n18164 ;
  assign n18172 = n18169 ^ n18145 ;
  assign n18141 = n18115 & n18140 ;
  assign n18173 = n18172 ^ n18141 ;
  assign n18160 = n18159 ^ n18146 ;
  assign n18132 = n18109 ^ n17960 ;
  assign n18138 = n18110 & ~n18132 ;
  assign n18126 = n18109 ^ n17958 ;
  assign n18127 = n18126 ^ n18110 ;
  assign n18128 = n18127 ^ n17960 ;
  assign n18129 = n18128 ^ n18109 ;
  assign n18130 = n18129 ^ n18110 ;
  assign n18131 = n18110 ^ n18109 ;
  assign n18133 = n18132 ^ n18109 ;
  assign n18134 = ~n18131 & n18133 ;
  assign n18135 = n18134 ^ n18109 ;
  assign n18136 = ~n18130 & ~n18135 ;
  assign n18137 = n18136 ^ n18127 ;
  assign n18139 = n18138 ^ n18137 ;
  assign n18142 = n18141 ^ n18139 ;
  assign n18161 = n18160 ^ n18142 ;
  assign n18170 = n18169 ^ n18161 ;
  assign n18171 = n18170 ^ n18140 ;
  assign n18174 = n18173 ^ n18171 ;
  assign n19637 = n18176 ^ n18174 ;
  assign n19638 = n18175 ^ n17911 ;
  assign n18189 = n18167 ^ n18141 ;
  assign n19639 = n19638 ^ n18189 ;
  assign n19640 = n18189 ^ n18176 ;
  assign n19641 = n19640 ^ n18189 ;
  assign n19642 = ~n19639 & ~n19641 ;
  assign n19643 = n19642 ^ n18189 ;
  assign n19644 = ~n19637 & n19643 ;
  assign n19645 = n19644 ^ n18174 ;
  assign n20393 = n18146 ^ n18138 ;
  assign n20392 = n18150 ^ n18141 ;
  assign n20394 = n20393 ^ n20392 ;
  assign n20395 = ~n17911 & n20394 ;
  assign n20396 = n20395 ^ n20392 ;
  assign n18184 = n18161 ^ n18146 ;
  assign n18197 = n18184 ^ n18169 ;
  assign n18198 = n18175 & n18197 ;
  assign n20407 = n20396 ^ n18198 ;
  assign n20398 = n18167 ^ n18147 ;
  assign n18185 = n18184 ^ n18152 ;
  assign n18183 = n18149 ^ n18113 ;
  assign n18186 = n18185 ^ n18183 ;
  assign n20399 = n20398 ^ n18186 ;
  assign n20400 = n20399 ^ n20396 ;
  assign n20397 = n20396 ^ n18137 ;
  assign n20401 = n20400 ^ n20397 ;
  assign n20402 = n20400 ^ n17911 ;
  assign n20403 = n20402 ^ n20400 ;
  assign n20404 = ~n20401 & ~n20403 ;
  assign n20405 = n20404 ^ n20400 ;
  assign n20406 = ~n17910 & ~n20405 ;
  assign n20408 = n20407 ^ n20406 ;
  assign n20409 = n19645 & ~n20408 ;
  assign n20411 = n20410 ^ n20409 ;
  assign n20768 = n20411 ^ x83 ;
  assign n16264 = n16263 ^ x77 ;
  assign n17661 = n17660 ^ n17659 ;
  assign n17665 = n17664 ^ n17661 ;
  assign n17666 = n17665 ^ n17650 ;
  assign n17667 = n17666 ^ n14956 ;
  assign n17668 = n17667 ^ x91 ;
  assign n17671 = ~n16264 & n17668 ;
  assign n17719 = n17671 ^ n16264 ;
  assign n17720 = n17719 ^ n17668 ;
  assign n17227 = n17194 ^ n17166 ;
  assign n17228 = n17227 ^ n17196 ;
  assign n17229 = n17075 & ~n17228 ;
  assign n17230 = n17229 ^ n17196 ;
  assign n17235 = n17234 ^ n17230 ;
  assign n17224 = n17213 ^ n17194 ;
  assign n17226 = n17225 ^ n17224 ;
  assign n17231 = n17230 ^ n17226 ;
  assign n17223 = ~n17075 & ~n17211 ;
  assign n17232 = n17231 ^ n17223 ;
  assign n17233 = ~n17074 & ~n17232 ;
  assign n17236 = n17235 ^ n17233 ;
  assign n17237 = n17236 ^ n17183 ;
  assign n17222 = ~n17075 & n17168 ;
  assign n17238 = n17237 ^ n17222 ;
  assign n17219 = ~n17210 & n17216 ;
  assign n17220 = n17219 ^ n17183 ;
  assign n17221 = n17192 & n17220 ;
  assign n17239 = n17238 ^ n17221 ;
  assign n17240 = n17239 ^ n17181 ;
  assign n17204 = n17181 ^ n17074 ;
  assign n17205 = n17204 ^ n17181 ;
  assign n17206 = n17188 & ~n17205 ;
  assign n17207 = n17206 ^ n17181 ;
  assign n17208 = ~n17075 & n17207 ;
  assign n17241 = n17240 ^ n17208 ;
  assign n17201 = n17192 & n17200 ;
  assign n17242 = n17241 ^ n17201 ;
  assign n17243 = ~n17191 & ~n17242 ;
  assign n17244 = n17190 & n17243 ;
  assign n17245 = n17244 ^ n14729 ;
  assign n17246 = n17245 ^ x78 ;
  assign n17522 = n17521 ^ x67 ;
  assign n17523 = n17246 & ~n17522 ;
  assign n16631 = n16626 ^ n16349 ;
  assign n16632 = ~n16630 & n16631 ;
  assign n16633 = n16632 ^ n16349 ;
  assign n16634 = n16623 ^ n16586 ;
  assign n16635 = n16634 ^ n16623 ;
  assign n16636 = n16635 ^ n16626 ;
  assign n16637 = n16633 & ~n16636 ;
  assign n16638 = n16637 ^ n16634 ;
  assign n16649 = n16648 ^ n16638 ;
  assign n16641 = n16598 ^ n16543 ;
  assign n16620 = n16619 ^ n16585 ;
  assign n16627 = n16626 ^ n16620 ;
  assign n16642 = n16641 ^ n16627 ;
  assign n16643 = n16642 ^ n16640 ;
  assign n16644 = n16349 & ~n16643 ;
  assign n16639 = n16638 ^ n16605 ;
  assign n16645 = n16644 ^ n16639 ;
  assign n16646 = ~n16353 & n16645 ;
  assign n16650 = n16649 ^ n16646 ;
  assign n16651 = n16650 ^ n16597 ;
  assign n16652 = n16651 ^ n14828 ;
  assign n16616 = n16597 ^ n16587 ;
  assign n16628 = n16627 ^ n16616 ;
  assign n16629 = ~n16615 & ~n16628 ;
  assign n16653 = n16652 ^ n16629 ;
  assign n16608 = n16607 ^ n16590 ;
  assign n16588 = n16587 ^ n16544 ;
  assign n16609 = n16608 ^ n16588 ;
  assign n16610 = n16588 ^ n16349 ;
  assign n16611 = n16610 ^ n16588 ;
  assign n16612 = n16609 & ~n16611 ;
  assign n16613 = n16612 ^ n16588 ;
  assign n16614 = n16353 & n16613 ;
  assign n16654 = n16653 ^ n16614 ;
  assign n16655 = n16654 ^ x116 ;
  assign n17052 = n16838 & n17051 ;
  assign n17053 = n17052 ^ n16988 ;
  assign n17054 = n17053 ^ n16838 ;
  assign n17055 = n17054 ^ n17053 ;
  assign n17056 = n17053 ^ n17006 ;
  assign n17057 = n17056 ^ n17053 ;
  assign n17058 = n17055 & n17057 ;
  assign n17059 = n17058 ^ n17053 ;
  assign n17060 = ~n16797 & n17059 ;
  assign n17061 = n17060 ^ n17053 ;
  assign n17045 = n16997 & ~n17002 ;
  assign n17025 = n17009 ^ n16988 ;
  assign n17023 = n17011 ^ n16978 ;
  assign n17024 = n17023 ^ n17022 ;
  assign n17026 = n17025 ^ n17024 ;
  assign n17027 = n17026 ^ n17022 ;
  assign n17028 = ~n16797 & n17027 ;
  assign n17029 = n17028 ^ n17024 ;
  assign n17044 = n17043 ^ n17029 ;
  assign n17046 = n17045 ^ n17044 ;
  assign n17062 = n17061 ^ n17046 ;
  assign n17063 = n17062 ^ n14693 ;
  assign n16996 = n16995 ^ n16994 ;
  assign n17030 = n17029 ^ n16996 ;
  assign n17031 = n17030 ^ n17022 ;
  assign n17013 = n17012 ^ n17011 ;
  assign n17007 = n17006 ^ n16994 ;
  assign n17014 = n17013 ^ n17007 ;
  assign n17015 = ~n16797 & n17014 ;
  assign n17032 = n17031 ^ n17015 ;
  assign n17033 = n17032 ^ n16983 ;
  assign n17034 = ~n16839 & ~n17033 ;
  assign n17064 = n17063 ^ n17034 ;
  assign n17003 = n16983 ^ n16976 ;
  assign n17004 = n17003 ^ n16981 ;
  assign n17005 = ~n17002 & ~n17004 ;
  assign n17065 = n17064 ^ n17005 ;
  assign n16998 = n16997 ^ n16996 ;
  assign n17066 = n17065 ^ n16998 ;
  assign n16990 = n16989 ^ n16988 ;
  assign n16993 = n16992 ^ n16990 ;
  assign n16999 = n16998 ^ n16993 ;
  assign n17000 = ~n16838 & n16999 ;
  assign n17067 = n17066 ^ n17000 ;
  assign n17068 = n17067 ^ n17065 ;
  assign n16985 = ~n16839 & n16976 ;
  assign n17069 = n17068 ^ n16985 ;
  assign n17070 = n16797 & n17069 ;
  assign n17071 = n17070 ^ n17067 ;
  assign n17072 = n17071 ^ x101 ;
  assign n17073 = n16655 & ~n17072 ;
  assign n17526 = n17073 ^ n16655 ;
  assign n17688 = n17523 & n17526 ;
  assign n17527 = n17523 ^ n17246 ;
  assign n17681 = n17073 & n17527 ;
  assign n17709 = n17688 ^ n17681 ;
  assign n17531 = n17073 ^ n17072 ;
  assign n17679 = n17527 & ~n17531 ;
  assign n17710 = n17709 ^ n17679 ;
  assign n17708 = n17073 & n17523 ;
  assign n17711 = n17710 ^ n17708 ;
  assign n17712 = n17711 ^ n17523 ;
  assign n17674 = n17526 ^ n17072 ;
  assign n17677 = n17523 & n17674 ;
  assign n17680 = n17679 ^ n17677 ;
  assign n17682 = n17681 ^ n17680 ;
  assign n17721 = n17712 ^ n17682 ;
  assign n17683 = n17526 & n17527 ;
  assign n17684 = n17683 ^ n17682 ;
  assign n17678 = n17677 ^ n17527 ;
  assign n17685 = n17684 ^ n17678 ;
  assign n17722 = n17721 ^ n17685 ;
  assign n17723 = n17720 & n17722 ;
  assign n20817 = n17723 ^ n16348 ;
  assign n17528 = n17527 ^ n17522 ;
  assign n17673 = n17073 & n17528 ;
  assign n17524 = n17523 ^ n17522 ;
  assign n17532 = ~n17524 & ~n17531 ;
  assign n19936 = n17673 ^ n17532 ;
  assign n17675 = ~n17524 & n17674 ;
  assign n19937 = n19936 ^ n17675 ;
  assign n17529 = n17526 & n17528 ;
  assign n20796 = n19937 ^ n17529 ;
  assign n20797 = n17720 & n20796 ;
  assign n17697 = n17668 ^ n16264 ;
  assign n17525 = n17073 & ~n17524 ;
  assign n19978 = n17685 ^ n17525 ;
  assign n17672 = n17671 ^ n17668 ;
  assign n17689 = n17688 ^ n17683 ;
  assign n17690 = n17689 ^ n17526 ;
  assign n17691 = n17690 ^ n17529 ;
  assign n17686 = n17685 ^ n17677 ;
  assign n17676 = n17675 ^ n17674 ;
  assign n17687 = n17686 ^ n17676 ;
  assign n17692 = n17691 ^ n17687 ;
  assign n17730 = n17672 & n17692 ;
  assign n20790 = n19978 ^ n17730 ;
  assign n17693 = n17692 ^ n17673 ;
  assign n17694 = n17693 ^ n17690 ;
  assign n17695 = n17694 ^ n17528 ;
  assign n19981 = n17695 ^ n17675 ;
  assign n20788 = n19981 ^ n17691 ;
  assign n20789 = ~n17719 & n20788 ;
  assign n20791 = n20790 ^ n20789 ;
  assign n20792 = n20791 ^ n17730 ;
  assign n20779 = n17522 ^ n17246 ;
  assign n20780 = n20779 ^ n16655 ;
  assign n20781 = n20780 ^ n17072 ;
  assign n20782 = n17668 & ~n20781 ;
  assign n17706 = n17522 ^ n16655 ;
  assign n17707 = n17706 ^ n17072 ;
  assign n20784 = n17707 ^ n17706 ;
  assign n20785 = ~n17522 & ~n20784 ;
  assign n20786 = n20785 ^ n17706 ;
  assign n20787 = n20782 & ~n20786 ;
  assign n20793 = n20792 ^ n20787 ;
  assign n20794 = n17697 & n20793 ;
  assign n20795 = n20794 ^ n20791 ;
  assign n20798 = n20797 ^ n20795 ;
  assign n20777 = n17687 ^ n17532 ;
  assign n20778 = n17671 & n20777 ;
  assign n20799 = n20798 ^ n20778 ;
  assign n20800 = n17722 ^ n17688 ;
  assign n20801 = n20800 ^ n17681 ;
  assign n20802 = n20801 ^ n17688 ;
  assign n20803 = n17688 ^ n16264 ;
  assign n20804 = n20803 ^ n17688 ;
  assign n20805 = n20802 & ~n20804 ;
  assign n20806 = n20805 ^ n17688 ;
  assign n20807 = ~n17697 & n20806 ;
  assign n20808 = ~n20799 & ~n20807 ;
  assign n20769 = n17721 ^ n17681 ;
  assign n20772 = n17679 ^ n17668 ;
  assign n20773 = n20772 ^ n17679 ;
  assign n20774 = n20769 & n20773 ;
  assign n20775 = n20774 ^ n17679 ;
  assign n20776 = n16264 & n20775 ;
  assign n20809 = n20808 ^ n20776 ;
  assign n20810 = n19981 ^ n17708 ;
  assign n20811 = n17708 ^ n16264 ;
  assign n20812 = n20811 ^ n17708 ;
  assign n20813 = n20810 & ~n20812 ;
  assign n20814 = n20813 ^ n17708 ;
  assign n20815 = n17697 & n20814 ;
  assign n20816 = n20809 & ~n20815 ;
  assign n20818 = n20817 ^ n20816 ;
  assign n20819 = n20818 ^ x109 ;
  assign n20820 = ~n20768 & ~n20819 ;
  assign n20838 = n20767 & n20820 ;
  assign n20821 = n20820 ^ n20819 ;
  assign n20823 = n20766 ^ n20729 ;
  assign n20825 = n20823 ^ n20765 ;
  assign n20826 = ~n20821 & ~n20825 ;
  assign n20824 = n20820 & n20823 ;
  assign n20827 = n20826 ^ n20824 ;
  assign n20822 = n20767 & ~n20821 ;
  assign n20828 = n20827 ^ n20822 ;
  assign n20853 = n20838 ^ n20828 ;
  assign n20834 = n20821 ^ n20768 ;
  assign n20850 = n20767 & ~n20834 ;
  assign n20851 = n20850 ^ n20827 ;
  assign n20852 = n20851 ^ n20767 ;
  assign n20854 = n20853 ^ n20852 ;
  assign n20835 = n20766 & ~n20834 ;
  assign n20855 = n20854 ^ n20835 ;
  assign n20832 = n20820 ^ n20768 ;
  assign n20849 = n20823 & ~n20832 ;
  assign n20856 = n20855 ^ n20849 ;
  assign n20833 = n20766 & ~n20832 ;
  assign n20836 = n20835 ^ n20833 ;
  assign n20848 = n20836 ^ n20832 ;
  assign n20857 = n20856 ^ n20848 ;
  assign n20847 = n20824 ^ n20822 ;
  assign n20858 = n20857 ^ n20847 ;
  assign n18627 = ~n17402 & n17450 ;
  assign n18624 = n17439 & ~n17453 ;
  assign n18625 = n18624 ^ n18623 ;
  assign n18612 = n17463 ^ n17451 ;
  assign n18613 = n17451 ^ n17402 ;
  assign n18614 = n18613 ^ n17451 ;
  assign n18615 = ~n18612 & ~n18614 ;
  assign n18616 = n18615 ^ n17451 ;
  assign n18617 = n17436 & n18616 ;
  assign n18626 = n18625 ^ n18617 ;
  assign n18628 = n18627 ^ n18626 ;
  assign n18610 = n17446 ^ n17368 ;
  assign n18611 = n18609 & n18610 ;
  assign n18629 = n18628 ^ n18611 ;
  assign n18606 = n17464 ^ n17457 ;
  assign n18607 = n18606 ^ n17363 ;
  assign n18608 = ~n17438 & n18607 ;
  assign n18630 = n18629 ^ n18608 ;
  assign n18598 = n17442 ^ n17375 ;
  assign n18599 = n18598 ^ n17487 ;
  assign n18600 = n18599 ^ n18598 ;
  assign n18601 = n18598 ^ n17436 ;
  assign n18602 = n18601 ^ n18598 ;
  assign n18603 = n18600 & ~n18602 ;
  assign n18604 = n18603 ^ n18598 ;
  assign n18605 = n17402 & n18604 ;
  assign n18631 = n18630 ^ n18605 ;
  assign n18632 = n18631 ^ n17471 ;
  assign n18634 = n18633 ^ n18632 ;
  assign n18635 = n18634 ^ n17470 ;
  assign n18636 = n18635 ^ n15194 ;
  assign n18637 = n18636 ^ x64 ;
  assign n18664 = ~n17077 & n17918 ;
  assign n18661 = n17918 ^ n17213 ;
  assign n18662 = ~n17075 & ~n18661 ;
  assign n18656 = n17194 ^ n17165 ;
  assign n18657 = n18656 ^ n17938 ;
  assign n18652 = n17194 ^ n17186 ;
  assign n18653 = n18652 ^ n17184 ;
  assign n18654 = n18653 ^ n17914 ;
  assign n18655 = n17076 & ~n18654 ;
  assign n18658 = n18657 ^ n18655 ;
  assign n18639 = n17953 ^ n17185 ;
  assign n18640 = n18639 ^ n17183 ;
  assign n18643 = n18640 ^ n17168 ;
  assign n18638 = n17186 ^ n17170 ;
  assign n18641 = n17077 & n18640 ;
  assign n18642 = ~n18638 & n18641 ;
  assign n18644 = n18643 ^ n18642 ;
  assign n18645 = n18644 ^ n17165 ;
  assign n18646 = n17178 ^ n17077 ;
  assign n18649 = ~n18644 & n18646 ;
  assign n18650 = n18649 ^ n17077 ;
  assign n18651 = n18645 & ~n18650 ;
  assign n18659 = n18658 ^ n18651 ;
  assign n18660 = n18659 ^ n18415 ;
  assign n18663 = n18662 ^ n18660 ;
  assign n18665 = n18664 ^ n18663 ;
  assign n18666 = ~n18423 & ~n18665 ;
  assign n18667 = n18666 ^ n17234 ;
  assign n18668 = ~n17189 & n18667 ;
  assign n18669 = n18668 ^ n15450 ;
  assign n18670 = n18669 ^ x73 ;
  assign n18671 = ~n18637 & n18670 ;
  assign n18750 = n18671 ^ n18637 ;
  assign n18704 = n18703 ^ x112 ;
  assign n18707 = n16220 ^ n16206 ;
  assign n18705 = n16211 ^ n16188 ;
  assign n18706 = n18705 ^ n16192 ;
  assign n18708 = n18707 ^ n18706 ;
  assign n18709 = n15987 & n18708 ;
  assign n18710 = n18709 ^ n18706 ;
  assign n18719 = n18710 ^ n16171 ;
  assign n18726 = n18725 ^ n18719 ;
  assign n18729 = n18728 ^ n18726 ;
  assign n18730 = n18729 ^ n18233 ;
  assign n18731 = n18730 ^ n16244 ;
  assign n18732 = n18731 ^ n15408 ;
  assign n18712 = n18710 ^ n16214 ;
  assign n18711 = n18710 ^ n16199 ;
  assign n18713 = n18712 ^ n18711 ;
  assign n18714 = n18711 ^ n16160 ;
  assign n18715 = n18714 ^ n18711 ;
  assign n18716 = ~n18713 & n18715 ;
  assign n18717 = n18716 ^ n18711 ;
  assign n18718 = ~n18224 & ~n18717 ;
  assign n18733 = n18732 ^ n18718 ;
  assign n18734 = n18733 ^ x82 ;
  assign n18735 = n18704 & n18734 ;
  assign n18751 = n18735 ^ n18734 ;
  assign n18752 = ~n18750 & n18751 ;
  assign n18736 = n18671 & n18735 ;
  assign n18756 = n18752 ^ n18736 ;
  assign n18597 = n18596 ^ x105 ;
  assign n18574 = n17045 ^ n15138 ;
  assign n18558 = n18528 ^ n17010 ;
  assign n18552 = n17006 ^ n16997 ;
  assign n18553 = n16997 ^ n16838 ;
  assign n18554 = n18553 ^ n16997 ;
  assign n18555 = n18552 & ~n18554 ;
  assign n18556 = n18555 ^ n16997 ;
  assign n18557 = n16797 & n18556 ;
  assign n18559 = n18558 ^ n18557 ;
  assign n18546 = n17012 ^ n16976 ;
  assign n18545 = n16994 ^ n16980 ;
  assign n18547 = n18546 ^ n18545 ;
  assign n18548 = n18547 ^ n18544 ;
  assign n18549 = n16838 & n18548 ;
  assign n18543 = n17011 ^ n16976 ;
  assign n18550 = n18549 ^ n18543 ;
  assign n18551 = ~n16797 & n18550 ;
  assign n18560 = n18559 ^ n18551 ;
  assign n18536 = n17010 ^ n16797 ;
  assign n18537 = n18536 ^ n17010 ;
  assign n18538 = n17010 ^ n17006 ;
  assign n18539 = n18538 ^ n17010 ;
  assign n18540 = n18537 & n18539 ;
  assign n18541 = n18540 ^ n17010 ;
  assign n18542 = n16838 & n18541 ;
  assign n18561 = n18560 ^ n18542 ;
  assign n18529 = n18528 ^ n16996 ;
  assign n18530 = n18529 ^ n18528 ;
  assign n18531 = n18528 ^ n16838 ;
  assign n18532 = n18531 ^ n18528 ;
  assign n18533 = n18530 & ~n18532 ;
  assign n18534 = n18533 ^ n18528 ;
  assign n18535 = n16839 & n18534 ;
  assign n18562 = n18561 ^ n18535 ;
  assign n18563 = ~n17041 & ~n18562 ;
  assign n18572 = n18571 ^ n18563 ;
  assign n18573 = ~n17061 & n18572 ;
  assign n18575 = n18574 ^ n18573 ;
  assign n18576 = n18575 ^ x123 ;
  assign n19355 = n18597 ^ n18576 ;
  assign n18766 = n18704 ^ n18670 ;
  assign n18737 = n18734 ^ n18637 ;
  assign n18767 = n18766 ^ n18737 ;
  assign n18768 = n18766 ^ n18704 ;
  assign n18759 = ~n18670 & n18704 ;
  assign n18769 = n18768 ^ n18759 ;
  assign n18770 = n18769 ^ n18704 ;
  assign n18771 = n18766 ^ n18637 ;
  assign n18772 = n18771 ^ n18704 ;
  assign n18773 = ~n18770 & ~n18772 ;
  assign n18774 = n18773 ^ n18704 ;
  assign n18775 = n18767 & n18774 ;
  assign n18776 = n18775 ^ n18759 ;
  assign n18762 = n18734 ^ n18704 ;
  assign n18758 = n18734 ^ n18670 ;
  assign n18760 = n18759 ^ n18637 ;
  assign n18761 = n18758 & n18760 ;
  assign n18763 = n18762 ^ n18761 ;
  assign n18738 = n18670 ^ n18637 ;
  assign n18745 = n18704 ^ n18637 ;
  assign n18746 = n18738 & ~n18745 ;
  assign n18747 = n18746 ^ n18704 ;
  assign n18757 = n18747 ^ n18670 ;
  assign n18764 = n18763 ^ n18757 ;
  assign n18744 = n18737 ^ n18704 ;
  assign n18748 = ~n18744 & ~n18747 ;
  assign n18749 = n18748 ^ n18637 ;
  assign n18753 = n18752 ^ n18749 ;
  assign n18765 = n18764 ^ n18753 ;
  assign n18777 = n18776 ^ n18765 ;
  assign n18739 = ~n18737 & n18738 ;
  assign n18740 = n18704 & n18739 ;
  assign n18787 = n18777 ^ n18740 ;
  assign n18783 = n18737 ^ n18671 ;
  assign n18784 = n18744 & ~n18783 ;
  assign n18785 = n18784 ^ n18766 ;
  assign n18788 = n18787 ^ n18785 ;
  assign n18786 = n18748 ^ n18739 ;
  assign n18789 = n18788 ^ n18786 ;
  assign n20484 = n18789 ^ n18749 ;
  assign n20485 = ~n18576 & n20484 ;
  assign n20486 = n20485 ^ n18749 ;
  assign n20487 = n20486 ^ n18785 ;
  assign n20488 = n20487 ^ n18788 ;
  assign n20489 = n20488 ^ n20487 ;
  assign n20490 = n20487 ^ n18597 ;
  assign n20491 = n20490 ^ n20487 ;
  assign n20492 = ~n20489 & ~n20491 ;
  assign n20493 = n20492 ^ n20487 ;
  assign n20494 = n19355 & n20493 ;
  assign n20495 = n20494 ^ n20486 ;
  assign n20496 = ~n18756 & ~n20495 ;
  assign n20497 = n20496 ^ n16937 ;
  assign n20862 = n20497 ^ x126 ;
  assign n20863 = ~n20858 & n20862 ;
  assign n20864 = n20863 ^ n20857 ;
  assign n20859 = n20858 ^ n20825 ;
  assign n20830 = n20766 & n20820 ;
  assign n20831 = n20830 ^ n20766 ;
  assign n20837 = n20836 ^ n20831 ;
  assign n20841 = n20837 ^ n20828 ;
  assign n20840 = n20824 ^ n20821 ;
  assign n20842 = n20841 ^ n20840 ;
  assign n20843 = n20842 ^ n20830 ;
  assign n20839 = n20838 ^ n20837 ;
  assign n20844 = n20843 ^ n20839 ;
  assign n20829 = n20828 ^ n20819 ;
  assign n20845 = n20844 ^ n20829 ;
  assign n20846 = n20845 ^ n20828 ;
  assign n20860 = n20859 ^ n20846 ;
  assign n20861 = n20860 ^ n20855 ;
  assign n20865 = n20864 ^ n20861 ;
  assign n20866 = n20865 ^ n20830 ;
  assign n20867 = n20866 ^ n20855 ;
  assign n20868 = n20867 ^ n20865 ;
  assign n20869 = n20865 ^ n20862 ;
  assign n20870 = n20869 ^ n20865 ;
  assign n20871 = n20868 & n20870 ;
  assign n20872 = n20871 ^ n20865 ;
  assign n20873 = n20686 & ~n20872 ;
  assign n20874 = n20873 ^ n20864 ;
  assign n20888 = n20862 ^ n20686 ;
  assign n20903 = n20850 ^ n20833 ;
  assign n20904 = ~n20888 & n20903 ;
  assign n20898 = n20686 & ~n20862 ;
  assign n20899 = n20898 ^ n20888 ;
  assign n20900 = n20857 ^ n20837 ;
  assign n20901 = n20899 & ~n20900 ;
  assign n20875 = n20856 ^ n20844 ;
  assign n20876 = n20686 & ~n20875 ;
  assign n20877 = n20876 ^ n20856 ;
  assign n20890 = n20877 ^ n20824 ;
  assign n20889 = n20877 ^ n20853 ;
  assign n20891 = n20890 ^ n20889 ;
  assign n20894 = ~n20686 & n20891 ;
  assign n20895 = n20894 ^ n20890 ;
  assign n20896 = ~n20888 & n20895 ;
  assign n20878 = n20823 & ~n20834 ;
  assign n20879 = n20878 ^ n20686 ;
  assign n20880 = n20879 ^ n20878 ;
  assign n20881 = n20845 ^ n20842 ;
  assign n20882 = n20881 ^ n20838 ;
  assign n20883 = n20882 ^ n20878 ;
  assign n20884 = n20880 & ~n20883 ;
  assign n20885 = n20884 ^ n20878 ;
  assign n20886 = n20862 & n20885 ;
  assign n20887 = n20886 ^ n20877 ;
  assign n20897 = n20896 ^ n20887 ;
  assign n20902 = n20901 ^ n20897 ;
  assign n20905 = n20904 ^ n20902 ;
  assign n20906 = n20874 & ~n20905 ;
  assign n20907 = n20878 ^ n20857 ;
  assign n20908 = n20857 ^ n20686 ;
  assign n20909 = n20908 ^ n20857 ;
  assign n20910 = ~n20907 & ~n20909 ;
  assign n20911 = n20910 ^ n20857 ;
  assign n20912 = ~n20862 & ~n20911 ;
  assign n20913 = n20906 & ~n20912 ;
  assign n20914 = n20913 ^ n17245 ;
  assign n20915 = n20914 ^ x83 ;
  assign n18741 = n18740 ^ n18736 ;
  assign n18742 = n18597 & n18741 ;
  assign n18743 = n18742 ^ n18740 ;
  assign n19351 = n18737 ^ n18670 ;
  assign n19352 = n19351 ^ n18764 ;
  assign n19360 = n19352 ^ n18740 ;
  assign n19356 = n18776 ^ n18734 ;
  assign n19357 = n19356 ^ n18704 ;
  assign n19358 = n19357 ^ n18637 ;
  assign n19359 = n19358 ^ n18736 ;
  assign n19361 = n19360 ^ n19359 ;
  assign n19362 = ~n18597 & ~n19361 ;
  assign n19363 = n19362 ^ n19359 ;
  assign n19364 = n19363 ^ n18763 ;
  assign n19365 = n19364 ^ n19363 ;
  assign n19348 = n18734 ^ n18671 ;
  assign n19349 = ~n18704 & ~n19348 ;
  assign n19350 = n19349 ^ n18738 ;
  assign n19366 = n19365 ^ n19350 ;
  assign n19367 = n18597 & n19366 ;
  assign n19368 = n19367 ^ n19364 ;
  assign n19369 = n19368 ^ n18743 ;
  assign n19370 = n19355 & ~n19369 ;
  assign n19371 = n19370 ^ n19350 ;
  assign n19353 = n19352 ^ n19350 ;
  assign n19354 = ~n18597 & n19353 ;
  assign n19372 = n19371 ^ n19354 ;
  assign n19374 = ~n18576 & ~n19372 ;
  assign n19375 = n18743 & n19374 ;
  assign n19373 = n19372 ^ n15494 ;
  assign n19376 = n19375 ^ n19373 ;
  assign n19377 = n19376 ^ x75 ;
  assign n18833 = n18636 ^ x70 ;
  assign n18836 = n17667 ^ x85 ;
  assign n18872 = n18026 & n18045 ;
  assign n18867 = n18095 ^ n18086 ;
  assign n18868 = ~n18030 & ~n18867 ;
  assign n18846 = n18027 ^ n18026 ;
  assign n18847 = n18096 ^ n18079 ;
  assign n18848 = n18847 ^ n18027 ;
  assign n18849 = ~n18846 & ~n18848 ;
  assign n18850 = n18849 ^ n18027 ;
  assign n18853 = n18847 ^ n18076 ;
  assign n18854 = n18850 & ~n18853 ;
  assign n18851 = n18076 ^ n18067 ;
  assign n18855 = n18854 ^ n18851 ;
  assign n18864 = n18855 ^ n18689 ;
  assign n18856 = n18855 ^ n18847 ;
  assign n18857 = n18856 ^ n18036 ;
  assign n18858 = n18857 ^ n18855 ;
  assign n18861 = n18027 & n18858 ;
  assign n18862 = n18861 ^ n18855 ;
  assign n18863 = ~n18846 & ~n18862 ;
  assign n18865 = n18864 ^ n18863 ;
  assign n18845 = n18692 ^ n18029 ;
  assign n18866 = n18865 ^ n18845 ;
  assign n18869 = n18868 ^ n18866 ;
  assign n18838 = n18047 ^ n18029 ;
  assign n18839 = n18043 ^ n18031 ;
  assign n18842 = ~n18047 & ~n18839 ;
  assign n18843 = n18842 ^ n18031 ;
  assign n18844 = n18838 & n18843 ;
  assign n18870 = n18869 ^ n18844 ;
  assign n18837 = n18027 & n18039 ;
  assign n18871 = n18870 ^ n18837 ;
  assign n18873 = n18872 ^ n18871 ;
  assign n18874 = ~n18032 & n18873 ;
  assign n18875 = n18874 ^ n16426 ;
  assign n18876 = n18875 ^ x83 ;
  assign n18877 = n18836 & ~n18876 ;
  assign n18878 = n18877 ^ n18836 ;
  assign n18914 = n18878 ^ n18876 ;
  assign n18908 = n17734 & n17844 ;
  assign n18902 = n18901 ^ n17735 ;
  assign n18894 = n17884 ^ n17864 ;
  assign n18895 = n18329 ^ n17846 ;
  assign n18898 = n17884 & ~n18895 ;
  assign n18899 = n18898 ^ n17846 ;
  assign n18900 = ~n18894 & ~n18899 ;
  assign n18903 = n18902 ^ n18900 ;
  assign n18884 = n18339 ^ n17839 ;
  assign n18885 = n17852 ^ n17778 ;
  assign n18886 = n18885 ^ n18329 ;
  assign n18887 = n18884 & n18886 ;
  assign n18889 = n18888 ^ n18887 ;
  assign n18893 = n18889 ^ n17907 ;
  assign n18904 = n18903 ^ n18893 ;
  assign n18905 = n18904 ^ n16453 ;
  assign n18883 = n17851 ^ n17840 ;
  assign n18890 = n18889 ^ n18883 ;
  assign n18880 = n17840 ^ n17827 ;
  assign n18881 = n18880 ^ n17848 ;
  assign n18882 = ~n17734 & ~n18881 ;
  assign n18891 = n18890 ^ n18882 ;
  assign n18892 = n17824 & ~n18891 ;
  assign n18906 = n18905 ^ n18892 ;
  assign n18879 = ~n17830 & n18350 ;
  assign n18907 = n18906 ^ n18879 ;
  assign n18909 = n18908 ^ n18907 ;
  assign n18910 = n18909 ^ x102 ;
  assign n18911 = n18575 ^ x108 ;
  assign n18912 = ~n18910 & n18911 ;
  assign n18917 = n18912 ^ n18911 ;
  assign n18918 = n18917 ^ n18910 ;
  assign n18921 = n18918 ^ n18911 ;
  assign n18941 = n18914 & ~n18921 ;
  assign n18937 = n18878 & n18918 ;
  assign n18915 = n18914 ^ n18836 ;
  assign n18919 = ~n18915 & n18918 ;
  assign n18938 = n18937 ^ n18919 ;
  assign n18934 = n18912 & ~n18915 ;
  assign n18913 = n18878 & n18912 ;
  assign n18935 = n18934 ^ n18913 ;
  assign n18932 = n18877 & n18912 ;
  assign n18933 = n18932 ^ n18912 ;
  assign n18936 = n18935 ^ n18933 ;
  assign n18939 = n18938 ^ n18936 ;
  assign n18925 = n18910 ^ n18876 ;
  assign n18930 = ~n18911 & n18925 ;
  assign n18923 = n18910 ^ n18836 ;
  assign n18924 = n18911 ^ n18876 ;
  assign n18926 = n18925 ^ n18876 ;
  assign n18927 = ~n18924 & n18926 ;
  assign n18928 = n18927 ^ n18876 ;
  assign n18929 = ~n18923 & n18928 ;
  assign n18931 = n18930 ^ n18929 ;
  assign n18940 = n18939 ^ n18931 ;
  assign n18942 = n18941 ^ n18940 ;
  assign n18943 = n18942 ^ n18919 ;
  assign n18944 = n18943 ^ n18930 ;
  assign n18945 = n18944 ^ n18938 ;
  assign n18946 = n18945 ^ n18918 ;
  assign n18922 = n18877 & ~n18921 ;
  assign n18947 = n18946 ^ n18922 ;
  assign n18948 = n18947 ^ n18942 ;
  assign n18949 = n18948 ^ n18911 ;
  assign n18950 = n18949 ^ n18945 ;
  assign n18951 = n18950 ^ n18934 ;
  assign n18920 = n18919 ^ n18915 ;
  assign n18952 = n18951 ^ n18920 ;
  assign n19012 = n18952 ^ n18934 ;
  assign n19003 = n18936 ^ n18914 ;
  assign n18970 = n18946 ^ n18941 ;
  assign n19004 = n19003 ^ n18970 ;
  assign n19013 = n19012 ^ n19004 ;
  assign n18834 = n17245 ^ x84 ;
  assign n19014 = n19004 ^ n18834 ;
  assign n19015 = n19014 ^ n19004 ;
  assign n19016 = n19013 & n19015 ;
  assign n19017 = n19016 ^ n19004 ;
  assign n19018 = n18833 & n19017 ;
  assign n18956 = n18877 & n18917 ;
  assign n18957 = n18956 ^ n18936 ;
  assign n19378 = n18833 & ~n18834 ;
  assign n19379 = n19378 ^ n18834 ;
  assign n19380 = n18957 & ~n19379 ;
  assign n18835 = n18834 ^ n18833 ;
  assign n19005 = n19004 ^ n18935 ;
  assign n19006 = n18935 ^ n18834 ;
  assign n19007 = n19006 ^ n18935 ;
  assign n19008 = n19005 & n19007 ;
  assign n19009 = n19008 ^ n18935 ;
  assign n19010 = n18835 & n19009 ;
  assign n19381 = n19380 ^ n19010 ;
  assign n19395 = n18937 ^ n18934 ;
  assign n19396 = n19395 ^ n18942 ;
  assign n19397 = n19396 ^ n18947 ;
  assign n19398 = ~n18833 & n19397 ;
  assign n19391 = n18936 ^ n18911 ;
  assign n19392 = ~n18833 & ~n19391 ;
  assign n19393 = n19392 ^ n18948 ;
  assign n19394 = n19393 ^ n18943 ;
  assign n19399 = n19398 ^ n19394 ;
  assign n19400 = ~n18834 & n19399 ;
  assign n19401 = n19400 ^ n19393 ;
  assign n18990 = n18878 & n18917 ;
  assign n19389 = n19378 ^ n18833 ;
  assign n19390 = n18990 & n19389 ;
  assign n19402 = n19401 ^ n19390 ;
  assign n19403 = n19402 ^ n18913 ;
  assign n19384 = n18913 ^ n18833 ;
  assign n19385 = n19384 ^ n18913 ;
  assign n19386 = n18956 & n19385 ;
  assign n19387 = n19386 ^ n18913 ;
  assign n19388 = ~n18834 & n19387 ;
  assign n19404 = n19403 ^ n19388 ;
  assign n19405 = ~n19381 & ~n19404 ;
  assign n19406 = n18833 & n18947 ;
  assign n19407 = n19406 ^ n18946 ;
  assign n19408 = n19407 ^ n18932 ;
  assign n19409 = n19408 ^ n19407 ;
  assign n19412 = ~n18833 & n19409 ;
  assign n19413 = n19412 ^ n19407 ;
  assign n19414 = ~n18835 & n19413 ;
  assign n19415 = n19414 ^ n19407 ;
  assign n19416 = n19405 & ~n19415 ;
  assign n19417 = ~n19018 & n19416 ;
  assign n19418 = n19417 ^ n16541 ;
  assign n19419 = n19418 ^ x124 ;
  assign n19895 = n19377 & n19419 ;
  assign n19897 = n19895 ^ n19377 ;
  assign n19896 = n19895 ^ n19419 ;
  assign n19898 = n19897 ^ n19896 ;
  assign n19607 = n18143 ^ n18117 ;
  assign n19613 = n19607 ^ n18159 ;
  assign n19610 = n18155 ^ n18152 ;
  assign n19611 = n19610 ^ n19607 ;
  assign n19612 = n17911 & n19611 ;
  assign n19614 = n19613 ^ n19612 ;
  assign n19615 = n18161 & ~n19614 ;
  assign n19616 = n17910 & ~n19615 ;
  assign n18177 = n18176 ^ n17911 ;
  assign n19608 = n19607 ^ n18170 ;
  assign n19609 = ~n18177 & n19608 ;
  assign n19617 = n19616 ^ n19609 ;
  assign n19602 = n18167 ^ n17910 ;
  assign n19603 = n19602 ^ n18167 ;
  assign n19604 = n18168 & ~n19603 ;
  assign n19605 = n19604 ^ n18167 ;
  assign n19606 = n17911 & n19605 ;
  assign n19618 = n19617 ^ n19606 ;
  assign n19619 = n18145 ^ n18113 ;
  assign n19620 = n18113 ^ n17911 ;
  assign n19621 = n19620 ^ n18113 ;
  assign n19622 = n19619 & ~n19621 ;
  assign n19623 = n19622 ^ n18113 ;
  assign n19624 = ~n17910 & n19623 ;
  assign n19625 = ~n19618 & ~n19624 ;
  assign n19626 = n17910 & ~n18173 ;
  assign n19627 = n19626 ^ n18141 ;
  assign n19628 = n19627 ^ n18152 ;
  assign n19629 = n19628 ^ n18153 ;
  assign n19630 = n19629 ^ n19627 ;
  assign n19633 = ~n17910 & n19630 ;
  assign n19634 = n19633 ^ n19627 ;
  assign n19635 = ~n17911 & n19634 ;
  assign n19636 = n19635 ^ n19627 ;
  assign n19646 = ~n19636 & n19645 ;
  assign n19647 = n19625 & n19646 ;
  assign n19648 = n19647 ^ n17774 ;
  assign n19649 = n19648 ^ x100 ;
  assign n18491 = ~n18457 & ~n18488 ;
  assign n18492 = n18491 ^ n18449 ;
  assign n18493 = ~n18393 & n18492 ;
  assign n19667 = n18466 ^ n18455 ;
  assign n19668 = n19667 ^ n18464 ;
  assign n19659 = n18456 ^ n18452 ;
  assign n18474 = n18473 ^ n18444 ;
  assign n19660 = n19659 ^ n18474 ;
  assign n19661 = n19660 ^ n18452 ;
  assign n19662 = n18452 ^ n18434 ;
  assign n19663 = n19662 ^ n18452 ;
  assign n19664 = ~n19661 & n19663 ;
  assign n19665 = n19664 ^ n18452 ;
  assign n19666 = ~n18463 & ~n19665 ;
  assign n19669 = n19668 ^ n19666 ;
  assign n19670 = n19669 ^ n18479 ;
  assign n19671 = n19670 ^ n19666 ;
  assign n19672 = n19666 ^ n18434 ;
  assign n19673 = n19672 ^ n19666 ;
  assign n19674 = ~n19671 & ~n19673 ;
  assign n19675 = n19674 ^ n19666 ;
  assign n19676 = ~n18393 & ~n19675 ;
  assign n19677 = n19676 ^ n19666 ;
  assign n19651 = n18458 ^ n18358 ;
  assign n19650 = n18473 ^ n18447 ;
  assign n19652 = n19651 ^ n19650 ;
  assign n19655 = n19654 ^ n19652 ;
  assign n19656 = ~n18393 & n19655 ;
  assign n19657 = n19656 ^ n19651 ;
  assign n19658 = n18434 & ~n19657 ;
  assign n19678 = n19677 ^ n19658 ;
  assign n19679 = ~n18493 & n19678 ;
  assign n18501 = n18500 ^ n18393 ;
  assign n18504 = n18438 & n18501 ;
  assign n18502 = n18466 ^ n18454 ;
  assign n18503 = n18501 & n18502 ;
  assign n18505 = n18504 ^ n18503 ;
  assign n19680 = n19679 ^ n18505 ;
  assign n19687 = n19680 & ~n19686 ;
  assign n19688 = n19687 ^ n17802 ;
  assign n19689 = n19688 ^ x85 ;
  assign n19690 = n19649 & ~n19689 ;
  assign n19691 = n19690 ^ n19649 ;
  assign n19422 = n18316 ^ x75 ;
  assign n19421 = n18108 ^ x93 ;
  assign n19457 = n18392 ^ x68 ;
  assign n19474 = n16992 ^ n16980 ;
  assign n19475 = n19474 ^ n17003 ;
  assign n19468 = n17051 ^ n17009 ;
  assign n19469 = n19468 ^ n18545 ;
  assign n19465 = n17051 ^ n16992 ;
  assign n19466 = n19465 ^ n18544 ;
  assign n19467 = n16838 & n19466 ;
  assign n19470 = n19469 ^ n19467 ;
  assign n19476 = n19475 ^ n19470 ;
  assign n19472 = n17047 ^ n17013 ;
  assign n19473 = n19472 ^ n19470 ;
  assign n19477 = n19476 ^ n19473 ;
  assign n19478 = ~n16797 & ~n19477 ;
  assign n19479 = n19478 ^ n19476 ;
  assign n19480 = n16839 & ~n19479 ;
  assign n19471 = n19470 ^ n18557 ;
  assign n19481 = n19480 ^ n19471 ;
  assign n19482 = n19481 ^ n18557 ;
  assign n19483 = n17010 ^ n16983 ;
  assign n19484 = n19483 ^ n16989 ;
  assign n19485 = ~n19049 & ~n19484 ;
  assign n19486 = ~n19482 & n19485 ;
  assign n19487 = n19486 ^ n19481 ;
  assign n19464 = n17001 & n17047 ;
  assign n19488 = n19487 ^ n19464 ;
  assign n19458 = n17013 ^ n16978 ;
  assign n19459 = n16978 ^ n16838 ;
  assign n19460 = n19459 ^ n16978 ;
  assign n19461 = n19458 & ~n19460 ;
  assign n19462 = n19461 ^ n16978 ;
  assign n19463 = n16797 & n19462 ;
  assign n19489 = n19488 ^ n19463 ;
  assign n19490 = ~n17045 & ~n19489 ;
  assign n19491 = n19490 ^ n15874 ;
  assign n19492 = n19491 ^ x110 ;
  assign n19493 = n19457 & n19492 ;
  assign n19424 = n17909 ^ x125 ;
  assign n19439 = n17507 ^ n17454 ;
  assign n19438 = n17500 ^ n17446 ;
  assign n19440 = n19439 ^ n19438 ;
  assign n19441 = n19438 ^ n17436 ;
  assign n19442 = n19441 ^ n19438 ;
  assign n19443 = ~n19440 & ~n19442 ;
  assign n19444 = n19443 ^ n19438 ;
  assign n19445 = ~n17402 & n19444 ;
  assign n19446 = n19445 ^ n18624 ;
  assign n19436 = n17465 ^ n17365 ;
  assign n19437 = n17437 & ~n19436 ;
  assign n19447 = n19446 ^ n19437 ;
  assign n19435 = ~n17438 & n17461 ;
  assign n19448 = n19447 ^ n19435 ;
  assign n19428 = n17485 ^ n17460 ;
  assign n19425 = n17489 ^ n17275 ;
  assign n19426 = n19425 ^ n17311 ;
  assign n19427 = n19426 ^ n17372 ;
  assign n19429 = n19428 ^ n19427 ;
  assign n19430 = n19427 ^ n17436 ;
  assign n19431 = n19430 ^ n19427 ;
  assign n19432 = n19429 & ~n19431 ;
  assign n19433 = n19432 ^ n19427 ;
  assign n19434 = n17402 & n19433 ;
  assign n19449 = n19448 ^ n19434 ;
  assign n19450 = n19449 ^ n19113 ;
  assign n19451 = ~n17471 & ~n19450 ;
  assign n19452 = n19451 ^ n18633 ;
  assign n19453 = ~n17376 & n19452 ;
  assign n19454 = n19453 ^ n15902 ;
  assign n19455 = n19454 ^ x124 ;
  assign n19456 = ~n19424 & n19455 ;
  assign n19496 = n19456 ^ n19424 ;
  assign n19516 = n19496 ^ n19455 ;
  assign n19572 = n19493 & n19516 ;
  assign n19577 = n19572 ^ n19516 ;
  assign n19520 = n19493 ^ n19457 ;
  assign n19521 = n19516 & n19520 ;
  assign n19519 = n19456 ^ n19455 ;
  assign n19522 = n19521 ^ n19519 ;
  assign n19517 = n19492 & n19516 ;
  assign n19518 = n19517 ^ n19424 ;
  assign n19523 = n19522 ^ n19518 ;
  assign n19578 = n19577 ^ n19523 ;
  assign n19494 = n19493 ^ n19492 ;
  assign n19505 = n19494 ^ n19457 ;
  assign n19509 = n19456 & ~n19505 ;
  assign n19506 = ~n19496 & ~n19505 ;
  assign n19503 = ~n19424 & n19493 ;
  assign n19498 = n19456 & n19493 ;
  assign n19504 = n19503 ^ n19498 ;
  assign n19507 = n19506 ^ n19504 ;
  assign n19510 = n19509 ^ n19507 ;
  assign n19497 = n19494 & ~n19496 ;
  assign n19502 = n19497 ^ n19496 ;
  assign n19508 = n19507 ^ n19502 ;
  assign n19511 = n19510 ^ n19508 ;
  assign n19499 = n19498 ^ n19497 ;
  assign n19495 = n19456 & n19494 ;
  assign n19500 = n19499 ^ n19495 ;
  assign n19501 = n19500 ^ n19424 ;
  assign n19512 = n19511 ^ n19501 ;
  assign n19529 = n19512 ^ n19508 ;
  assign n19528 = n19521 ^ n19520 ;
  assign n19530 = n19529 ^ n19528 ;
  assign n19579 = n19578 ^ n19530 ;
  assign n19580 = ~n19421 & ~n19579 ;
  assign n19583 = n19580 ^ n19530 ;
  assign n19536 = n19494 & n19519 ;
  assign n19586 = n19583 ^ n19536 ;
  assign n19587 = n19586 ^ n19583 ;
  assign n19588 = n19421 & n19587 ;
  assign n19589 = n19588 ^ n19583 ;
  assign n19590 = ~n19422 & ~n19589 ;
  assign n19591 = n19590 ^ n19583 ;
  assign n19524 = n19523 ^ n19509 ;
  assign n19515 = n19506 ^ n19505 ;
  assign n19525 = n19524 ^ n19515 ;
  assign n19559 = ~n19421 & ~n19422 ;
  assign n19560 = n19559 ^ n19422 ;
  assign n19561 = n19560 ^ n19421 ;
  assign n19573 = n19561 ^ n19422 ;
  assign n19576 = ~n19525 & ~n19573 ;
  assign n19592 = n19591 ^ n19576 ;
  assign n19574 = n19572 & ~n19573 ;
  assign n19534 = n19525 ^ n19521 ;
  assign n19535 = n19534 ^ n19530 ;
  assign n19537 = n19536 ^ n19535 ;
  assign n19538 = n19537 ^ n19522 ;
  assign n19566 = n19538 ^ n19523 ;
  assign n19567 = n19523 ^ n19422 ;
  assign n19568 = n19567 ^ n19523 ;
  assign n19569 = n19566 & ~n19568 ;
  assign n19570 = n19569 ^ n19523 ;
  assign n19571 = n19421 & n19570 ;
  assign n19575 = n19574 ^ n19571 ;
  assign n19593 = n19592 ^ n19575 ;
  assign n19533 = n19506 ^ n19497 ;
  assign n19539 = n19538 ^ n19533 ;
  assign n19514 = n19492 ^ n19457 ;
  assign n19526 = n19525 ^ n19514 ;
  assign n19513 = n19512 ^ n19504 ;
  assign n19527 = n19526 ^ n19513 ;
  assign n19531 = n19530 ^ n19527 ;
  assign n19532 = ~n19421 & ~n19531 ;
  assign n19540 = n19539 ^ n19532 ;
  assign n19594 = n19593 ^ n19540 ;
  assign n19563 = n19504 ^ n19495 ;
  assign n19564 = ~n19561 & n19563 ;
  assign n19562 = n19509 & ~n19561 ;
  assign n19565 = n19564 ^ n19562 ;
  assign n19595 = n19594 ^ n19565 ;
  assign n19548 = n19536 ^ n19497 ;
  assign n19549 = ~n19422 & n19548 ;
  assign n19550 = n19549 ^ n19497 ;
  assign n19551 = n19550 ^ n19422 ;
  assign n19552 = n19551 ^ n19550 ;
  assign n19553 = n19550 ^ n19534 ;
  assign n19554 = n19553 ^ n19550 ;
  assign n19555 = ~n19552 & ~n19554 ;
  assign n19556 = n19555 ^ n19550 ;
  assign n19557 = n19421 & n19556 ;
  assign n19558 = n19557 ^ n19550 ;
  assign n19596 = n19595 ^ n19558 ;
  assign n19597 = n19596 ^ n15986 ;
  assign n19423 = n19422 ^ n19421 ;
  assign n19541 = n19540 ^ n19511 ;
  assign n19542 = n19541 ^ n19529 ;
  assign n19543 = n19542 ^ n19536 ;
  assign n19544 = n19543 ^ n19540 ;
  assign n19545 = ~n19421 & n19544 ;
  assign n19546 = n19545 ^ n19541 ;
  assign n19547 = n19423 & ~n19546 ;
  assign n19598 = n19597 ^ n19547 ;
  assign n19599 = n19598 ^ x125 ;
  assign n19833 = n19776 & ~n19832 ;
  assign n19826 = n19825 ^ n19783 ;
  assign n19827 = ~n19696 & ~n19826 ;
  assign n19828 = n19827 ^ n19783 ;
  assign n19804 = ~n19694 & ~n19790 ;
  assign n19778 = n19697 & n19777 ;
  assign n19779 = n19778 ^ n19757 ;
  assign n19792 = n19791 ^ n19779 ;
  assign n19793 = n19792 ^ n19752 ;
  assign n19795 = n19794 ^ n19793 ;
  assign n19796 = n19766 ^ n19696 ;
  assign n19797 = n19793 ^ n19696 ;
  assign n19798 = n19797 ^ n19696 ;
  assign n19799 = ~n19796 & ~n19798 ;
  assign n19800 = n19799 ^ n19696 ;
  assign n19801 = n19795 & n19800 ;
  assign n19802 = n19801 ^ n19794 ;
  assign n19803 = n19802 ^ n19769 ;
  assign n19805 = n19804 ^ n19803 ;
  assign n19829 = n19828 ^ n19805 ;
  assign n19818 = n19758 ^ n19694 ;
  assign n19819 = n19818 ^ n19758 ;
  assign n19820 = n19759 & n19819 ;
  assign n19821 = n19820 ^ n19758 ;
  assign n19822 = ~n19696 & n19821 ;
  assign n19823 = n19822 ^ n19758 ;
  assign n19830 = n19829 ^ n19823 ;
  assign n19806 = n19805 ^ n19802 ;
  assign n19807 = n19806 ^ n19695 ;
  assign n19808 = n19807 ^ n19806 ;
  assign n19814 = n19808 & ~n19811 ;
  assign n19815 = n19814 ^ n19806 ;
  assign n19816 = n19696 & ~n19815 ;
  assign n19831 = n19830 ^ n19816 ;
  assign n19834 = n19833 ^ n19831 ;
  assign n19841 = ~n19834 & ~n19840 ;
  assign n19842 = n19841 ^ n16305 ;
  assign n19843 = n19842 ^ x118 ;
  assign n19844 = ~n19599 & n19843 ;
  assign n19845 = n19844 ^ n19599 ;
  assign n19910 = n19691 & ~n19845 ;
  assign n19860 = n19690 & ~n19845 ;
  assign n19911 = n19910 ^ n19860 ;
  assign n19692 = n19691 ^ n19689 ;
  assign n19882 = n19692 & ~n19845 ;
  assign n19883 = n19882 ^ n19845 ;
  assign n19912 = n19911 ^ n19883 ;
  assign n19846 = n19845 ^ n19843 ;
  assign n19855 = n19690 & n19846 ;
  assign n19927 = n19912 ^ n19855 ;
  assign n19852 = n19690 ^ n19689 ;
  assign n19906 = n19844 & ~n19852 ;
  assign n19907 = n19906 ^ n19882 ;
  assign n19899 = n19691 & n19844 ;
  assign n19926 = n19907 ^ n19899 ;
  assign n19928 = n19927 ^ n19926 ;
  assign n19924 = n19689 ^ n19599 ;
  assign n19875 = n19843 ^ n19599 ;
  assign n19876 = n19843 ^ n19649 ;
  assign n19877 = n19689 ^ n19649 ;
  assign n19878 = n19877 ^ n19649 ;
  assign n19879 = ~n19876 & ~n19878 ;
  assign n19880 = n19879 ^ n19649 ;
  assign n19881 = ~n19875 & n19880 ;
  assign n19925 = n19924 ^ n19881 ;
  assign n19929 = n19928 ^ n19925 ;
  assign n19930 = ~n19419 & n19929 ;
  assign n19931 = n19930 ^ n19925 ;
  assign n19932 = ~n19898 & ~n19931 ;
  assign n19847 = n19846 ^ n19599 ;
  assign n19858 = n19690 & n19847 ;
  assign n19862 = n19858 ^ n19855 ;
  assign n19861 = n19860 ^ n19690 ;
  assign n19863 = n19862 ^ n19861 ;
  assign n19908 = n19907 ^ n19863 ;
  assign n19900 = n19899 ^ n19882 ;
  assign n19905 = n19900 ^ n19844 ;
  assign n19909 = n19908 ^ n19905 ;
  assign n19913 = n19912 ^ n19909 ;
  assign n19884 = n19883 ^ n19881 ;
  assign n19850 = n19692 & n19846 ;
  assign n19885 = n19884 ^ n19850 ;
  assign n19886 = n19885 ^ n19858 ;
  assign n19693 = n19599 & n19692 ;
  assign n19848 = n19847 ^ n19693 ;
  assign n19887 = n19886 ^ n19848 ;
  assign n19888 = n19887 ^ n19855 ;
  assign n19914 = n19913 ^ n19888 ;
  assign n19915 = ~n19419 & n19914 ;
  assign n19901 = n19898 & n19900 ;
  assign n19853 = n19846 & ~n19852 ;
  assign n19889 = n19888 ^ n19853 ;
  assign n19890 = n19853 ^ n19377 ;
  assign n19891 = n19890 ^ n19853 ;
  assign n19892 = ~n19889 & ~n19891 ;
  assign n19893 = n19892 ^ n19853 ;
  assign n19894 = n19419 & n19893 ;
  assign n19902 = n19901 ^ n19894 ;
  assign n19903 = n19902 ^ n18909 ;
  assign n19420 = n19419 ^ n19377 ;
  assign n19851 = n19850 ^ n19693 ;
  assign n19854 = n19853 ^ n19851 ;
  assign n19856 = n19855 ^ n19854 ;
  assign n19849 = n19848 ^ n19599 ;
  assign n19857 = n19856 ^ n19849 ;
  assign n19859 = n19858 ^ n19857 ;
  assign n19864 = n19863 ^ n19859 ;
  assign n19865 = ~n19419 & n19864 ;
  assign n19866 = n19865 ^ n19863 ;
  assign n19867 = n19866 ^ n19860 ;
  assign n19868 = n19867 ^ n19866 ;
  assign n19869 = n19866 ^ n19377 ;
  assign n19870 = n19869 ^ n19866 ;
  assign n19871 = n19868 & n19870 ;
  assign n19872 = n19871 ^ n19866 ;
  assign n19873 = ~n19420 & n19872 ;
  assign n19874 = n19873 ^ n19866 ;
  assign n19904 = n19903 ^ n19874 ;
  assign n19916 = n19915 ^ n19904 ;
  assign n19919 = n19916 ^ n18909 ;
  assign n19920 = n19919 ^ n19874 ;
  assign n19917 = n19884 ^ n19854 ;
  assign n19918 = n19917 ^ n19902 ;
  assign n19921 = n19920 ^ n19918 ;
  assign n19922 = ~n19377 & ~n19921 ;
  assign n19923 = n19922 ^ n19916 ;
  assign n19933 = n19932 ^ n19923 ;
  assign n19934 = n19933 ^ x70 ;
  assign n18178 = ~n18174 & ~n18177 ;
  assign n17912 = n17911 ^ n17910 ;
  assign n18118 = n18117 ^ n18113 ;
  assign n18119 = n18118 ^ n18117 ;
  assign n18120 = n18117 ^ n17910 ;
  assign n18121 = n18120 ^ n18117 ;
  assign n18122 = n18119 & n18121 ;
  assign n18123 = n18122 ^ n18117 ;
  assign n18124 = n17912 & n18123 ;
  assign n18125 = n18124 ^ n18117 ;
  assign n18179 = n18178 ^ n18125 ;
  assign n20000 = n18167 ^ n18159 ;
  assign n20001 = n20000 ^ n18161 ;
  assign n20002 = ~n17910 & ~n20001 ;
  assign n20003 = n20002 ^ n18184 ;
  assign n20004 = ~n17911 & ~n20003 ;
  assign n20005 = n20004 ^ n18151 ;
  assign n19995 = n18151 ^ n17910 ;
  assign n19996 = n19995 ^ n18151 ;
  assign n19997 = n18157 & n19996 ;
  assign n19998 = n19997 ^ n18151 ;
  assign n19999 = ~n17912 & n19998 ;
  assign n20006 = n20005 ^ n19999 ;
  assign n20007 = n18141 ^ n17910 ;
  assign n20008 = n20007 ^ n18141 ;
  assign n20009 = n17911 & n18170 ;
  assign n20010 = n20009 ^ n18141 ;
  assign n20011 = ~n20008 & n20010 ;
  assign n20012 = n20011 ^ n18141 ;
  assign n20013 = ~n20006 & n20012 ;
  assign n20014 = n20013 ^ n20006 ;
  assign n20015 = ~n19624 & ~n20014 ;
  assign n20016 = ~n18179 & n20015 ;
  assign n20017 = ~n19636 & n20016 ;
  assign n19993 = n19992 ^ n18018 ;
  assign n20018 = n20017 ^ n19993 ;
  assign n20019 = n20018 ^ x104 ;
  assign n20053 = n19833 ^ n17988 ;
  assign n20028 = n19748 ^ n19721 ;
  assign n20027 = n20026 ^ n19772 ;
  assign n20029 = n20028 ^ n20027 ;
  assign n20023 = n20022 ^ n19760 ;
  assign n20024 = n20023 ^ n19752 ;
  assign n20025 = n20024 ^ n19773 ;
  assign n20030 = n20029 ^ n20025 ;
  assign n20031 = n19694 & n20030 ;
  assign n20032 = n20031 ^ n20027 ;
  assign n20033 = n20032 ^ n19763 ;
  assign n20020 = n19764 ^ n19749 ;
  assign n20021 = ~n19694 & n20020 ;
  assign n20034 = n20033 ^ n20021 ;
  assign n20035 = ~n19695 & n20034 ;
  assign n20036 = n20035 ^ n20032 ;
  assign n20040 = n19695 & n19779 ;
  assign n20038 = n19696 & n20022 ;
  assign n20037 = n19787 ^ n19757 ;
  assign n20039 = n20038 ^ n20037 ;
  assign n20041 = n20040 ^ n20039 ;
  assign n20042 = n20041 ^ n19695 ;
  assign n20045 = n19765 ^ n19759 ;
  assign n20046 = n20045 ^ n19694 ;
  assign n20047 = ~n20041 & n20046 ;
  assign n20048 = n20047 ^ n19694 ;
  assign n20049 = ~n20042 & ~n20048 ;
  assign n20050 = n20049 ^ n19695 ;
  assign n20051 = n19828 & n20050 ;
  assign n20052 = n20036 & n20051 ;
  assign n20054 = n20053 ^ n20052 ;
  assign n20055 = n20054 ^ x97 ;
  assign n20100 = n19512 ^ n19507 ;
  assign n20101 = n19507 ^ n19421 ;
  assign n20102 = n20101 ^ n19507 ;
  assign n20103 = n20100 & n20102 ;
  assign n20104 = n20103 ^ n19507 ;
  assign n20105 = n19422 & n20104 ;
  assign n20106 = n20105 ^ n16837 ;
  assign n20081 = n19572 ^ n19525 ;
  assign n20082 = n20081 ^ n19495 ;
  assign n20083 = n19495 ^ n19422 ;
  assign n20084 = n20083 ^ n19495 ;
  assign n20085 = ~n20082 & ~n20084 ;
  assign n20086 = n20085 ^ n19495 ;
  assign n20087 = ~n19421 & n20086 ;
  assign n20088 = n20087 ^ n19571 ;
  assign n20068 = n19517 ^ n19500 ;
  assign n20066 = n19538 ^ n19508 ;
  assign n20058 = n19529 ^ n19524 ;
  assign n20059 = n20058 ^ n19572 ;
  assign n20060 = n20059 ^ n19529 ;
  assign n20061 = n19529 ^ n19421 ;
  assign n20062 = n20061 ^ n19529 ;
  assign n20063 = n20060 & n20062 ;
  assign n20064 = n20063 ^ n19529 ;
  assign n20065 = ~n19422 & ~n20064 ;
  assign n20067 = n20066 ^ n20065 ;
  assign n20069 = n20068 ^ n20067 ;
  assign n20070 = n20069 ^ n20065 ;
  assign n20071 = n19421 & ~n20070 ;
  assign n20072 = n20071 ^ n20067 ;
  assign n20089 = n20088 ^ n20072 ;
  assign n20090 = n20089 ^ n19592 ;
  assign n20073 = n20072 ^ n20065 ;
  assign n20076 = n20073 ^ n19578 ;
  assign n20077 = n20076 ^ n20073 ;
  assign n20078 = ~n19421 & n20077 ;
  assign n20079 = n20078 ^ n20073 ;
  assign n20080 = ~n19422 & ~n20079 ;
  assign n20091 = n20090 ^ n20080 ;
  assign n20092 = n19499 ^ n19421 ;
  assign n20093 = n20092 ^ n19499 ;
  assign n20096 = n19500 & n20093 ;
  assign n20097 = n20096 ^ n19499 ;
  assign n20098 = ~n19422 & n20097 ;
  assign n20099 = ~n20091 & ~n20098 ;
  assign n20107 = n20106 ^ n20099 ;
  assign n20108 = n20107 ^ x123 ;
  assign n19001 = n18834 & n18937 ;
  assign n18993 = ~n18834 & n18990 ;
  assign n18985 = n18952 ^ n18950 ;
  assign n18986 = ~n18834 & ~n18985 ;
  assign n18987 = n18986 ^ n18950 ;
  assign n18994 = n18993 ^ n18987 ;
  assign n18995 = ~n18833 & ~n18994 ;
  assign n18996 = n18995 ^ n18987 ;
  assign n18916 = n18915 ^ n18913 ;
  assign n18953 = n18952 ^ n18916 ;
  assign n18954 = n18953 ^ n18910 ;
  assign n18955 = n18954 ^ n18940 ;
  assign n18958 = n18957 ^ n18955 ;
  assign n18959 = n18834 & n18958 ;
  assign n18960 = n18959 ^ n18954 ;
  assign n18997 = n18996 ^ n18960 ;
  assign n18978 = n18970 ^ n18947 ;
  assign n18979 = n18978 ^ n18946 ;
  assign n18980 = n18946 ^ n18834 ;
  assign n18981 = n18980 ^ n18946 ;
  assign n18982 = n18979 & n18981 ;
  assign n18983 = n18982 ^ n18946 ;
  assign n18984 = n18835 & n18983 ;
  assign n18998 = n18997 ^ n18984 ;
  assign n18973 = n18941 ^ n18834 ;
  assign n18974 = n18973 ^ n18941 ;
  assign n18975 = n18970 & n18974 ;
  assign n18976 = n18975 ^ n18941 ;
  assign n18977 = n18833 & n18976 ;
  assign n18999 = n18998 ^ n18977 ;
  assign n18963 = n18960 ^ n18944 ;
  assign n18961 = n18952 ^ n18932 ;
  assign n18962 = n18961 ^ n18960 ;
  assign n18964 = n18963 ^ n18962 ;
  assign n18965 = n18963 ^ n18833 ;
  assign n18966 = n18965 ^ n18963 ;
  assign n18967 = n18964 & ~n18966 ;
  assign n18968 = n18967 ^ n18963 ;
  assign n18969 = n18835 & n18968 ;
  assign n19000 = n18999 ^ n18969 ;
  assign n19002 = n19001 ^ n19000 ;
  assign n19011 = n19002 & ~n19010 ;
  assign n19019 = n19011 & ~n19018 ;
  assign n19020 = n18950 ^ n18944 ;
  assign n19021 = n19020 ^ n18990 ;
  assign n19022 = n18834 & ~n19021 ;
  assign n19023 = n19022 ^ n18990 ;
  assign n19024 = n19023 ^ n19004 ;
  assign n19025 = n19024 ^ n19023 ;
  assign n19026 = n19023 ^ n18833 ;
  assign n19027 = n19026 ^ n19023 ;
  assign n19028 = n19025 & ~n19027 ;
  assign n19029 = n19028 ^ n19023 ;
  assign n19030 = ~n18835 & n19029 ;
  assign n19031 = n19030 ^ n19023 ;
  assign n19032 = n19019 & ~n19031 ;
  assign n19033 = n19032 ^ n17435 ;
  assign n20109 = n19033 ^ x114 ;
  assign n20110 = n20108 & ~n20109 ;
  assign n20121 = n20055 & n20110 ;
  assign n20131 = n20019 & n20121 ;
  assign n20056 = n20019 & ~n20055 ;
  assign n20127 = n20056 ^ n20019 ;
  assign n20132 = n20131 ^ n20127 ;
  assign n20111 = n20110 ^ n20109 ;
  assign n20129 = ~n20111 & n20127 ;
  assign n20112 = n20111 ^ n20108 ;
  assign n20128 = n20112 & n20127 ;
  assign n20130 = n20129 ^ n20128 ;
  assign n20133 = n20132 ^ n20130 ;
  assign n20057 = n20056 ^ n20055 ;
  assign n20116 = n20110 ^ n20108 ;
  assign n20125 = ~n20057 & n20116 ;
  assign n20147 = n20133 ^ n20125 ;
  assign n20113 = ~n20057 & n20112 ;
  assign n20148 = n20147 ^ n20113 ;
  assign n20119 = ~n20057 & n20110 ;
  assign n20134 = n20133 ^ n20119 ;
  assign n20146 = n20134 ^ n20057 ;
  assign n20149 = n20148 ^ n20146 ;
  assign n20117 = n20057 ^ n20019 ;
  assign n20140 = n20109 & n20117 ;
  assign n20118 = n20116 & n20117 ;
  assign n20141 = n20140 ^ n20118 ;
  assign n20150 = n20149 ^ n20141 ;
  assign n20144 = n20140 ^ n20117 ;
  assign n20137 = n20131 ^ n20121 ;
  assign n20145 = n20144 ^ n20137 ;
  assign n20151 = n20150 ^ n20145 ;
  assign n19935 = n17722 ^ n17689 ;
  assign n19945 = n17525 ^ n16264 ;
  assign n19947 = n17683 ^ n17525 ;
  assign n19946 = n17682 ^ n17525 ;
  assign n19948 = n19947 ^ n19946 ;
  assign n19949 = n19947 ^ n17668 ;
  assign n19950 = n19949 ^ n19947 ;
  assign n19951 = n19948 & n19950 ;
  assign n19952 = n19951 ^ n19947 ;
  assign n19953 = n19945 & ~n19952 ;
  assign n19954 = n19953 ^ n16264 ;
  assign n19938 = n19937 ^ n17525 ;
  assign n19939 = n19938 ^ n17711 ;
  assign n19940 = n17711 ^ n17668 ;
  assign n19941 = n19940 ^ n17711 ;
  assign n19942 = n19939 & n19941 ;
  assign n19943 = n19942 ^ n17711 ;
  assign n19944 = ~n16264 & n19943 ;
  assign n19955 = n19954 ^ n19944 ;
  assign n19956 = n19955 ^ n17723 ;
  assign n19960 = ~n17668 & n17693 ;
  assign n19961 = n19960 ^ n17690 ;
  assign n19962 = n17697 & n19961 ;
  assign n19963 = n19962 ^ n17690 ;
  assign n19964 = ~n19956 & n19963 ;
  assign n19965 = n19964 ^ n19956 ;
  assign n19966 = ~n17668 & ~n19965 ;
  assign n19967 = n17532 ^ n16264 ;
  assign n19968 = n19967 ^ n17532 ;
  assign n19971 = n17695 & ~n19968 ;
  assign n19972 = n19971 ^ n17532 ;
  assign n19973 = n19966 & n19972 ;
  assign n19974 = n19973 ^ n19965 ;
  assign n19975 = n17671 & ~n19974 ;
  assign n19976 = n19935 & n19975 ;
  assign n19977 = n19976 ^ n19974 ;
  assign n19979 = n19978 ^ n17532 ;
  assign n19980 = n19979 ^ n17689 ;
  assign n19983 = n19980 ^ n17672 ;
  assign n19984 = ~n19981 & ~n19983 ;
  assign n19985 = n19984 ^ n17672 ;
  assign n19982 = n19981 ^ n19980 ;
  assign n19986 = n19985 ^ n19982 ;
  assign n19987 = ~n19977 & n19986 ;
  assign n19988 = n19987 ^ n16971 ;
  assign n19989 = n19988 ^ x99 ;
  assign n18498 = n18497 ^ n18493 ;
  assign n18481 = n18434 & ~n18480 ;
  assign n18477 = n18448 ^ n18442 ;
  assign n18482 = n18481 ^ n18477 ;
  assign n18499 = n18498 ^ n18482 ;
  assign n18506 = n18505 ^ n18499 ;
  assign n18520 = n18519 ^ n18506 ;
  assign n18483 = n18482 ^ n18458 ;
  assign n18484 = n18483 ^ n18474 ;
  assign n18470 = n18469 ^ n18456 ;
  assign n18465 = n18464 ^ n18444 ;
  assign n18471 = n18470 ^ n18465 ;
  assign n18459 = n18458 ^ n18454 ;
  assign n18472 = n18471 ^ n18459 ;
  assign n18475 = n18474 ^ n18472 ;
  assign n18476 = n18434 & ~n18475 ;
  assign n18485 = n18484 ^ n18476 ;
  assign n18486 = ~n18435 & ~n18485 ;
  assign n18521 = n18520 ^ n18486 ;
  assign n18522 = ~n18358 & ~n18521 ;
  assign n18523 = n18522 ^ n17274 ;
  assign n19990 = n18523 ^ x72 ;
  assign n20183 = n19989 & ~n19990 ;
  assign n20184 = n20183 ^ n19990 ;
  assign n20185 = n20184 ^ n19989 ;
  assign n20188 = n20185 ^ n19990 ;
  assign n20211 = ~n20151 & n20188 ;
  assign n20126 = n20125 ^ n20121 ;
  assign n20135 = n20134 ^ n20126 ;
  assign n20120 = n20119 ^ n20110 ;
  assign n20122 = n20121 ^ n20120 ;
  assign n20123 = n20122 ^ n20118 ;
  assign n20124 = n20123 ^ n20108 ;
  assign n20136 = n20135 ^ n20124 ;
  assign n20198 = n20136 ^ n20131 ;
  assign n20199 = n20198 ^ n20125 ;
  assign n20196 = n20129 & ~n20184 ;
  assign n20169 = n19990 ^ n19989 ;
  assign n20190 = n20137 ^ n20123 ;
  assign n20191 = n20137 ^ n19989 ;
  assign n20192 = n20191 ^ n20137 ;
  assign n20193 = n20190 & ~n20192 ;
  assign n20194 = n20193 ^ n20137 ;
  assign n20195 = n20169 & n20194 ;
  assign n20197 = n20196 ^ n20195 ;
  assign n20200 = n20199 ^ n20197 ;
  assign n20189 = n20122 & n20188 ;
  assign n20201 = n20200 ^ n20189 ;
  assign n20142 = n20141 ^ n20129 ;
  assign n20143 = n20142 ^ n20111 ;
  assign n20152 = n20151 ^ n20143 ;
  assign n20208 = n20201 ^ n20152 ;
  assign n20203 = n20152 ^ n20141 ;
  assign n20204 = n20203 ^ n20128 ;
  assign n20205 = ~n19990 & n20204 ;
  assign n20202 = n20201 ^ n20197 ;
  assign n20206 = n20205 ^ n20202 ;
  assign n20207 = ~n19989 & n20206 ;
  assign n20209 = n20208 ^ n20207 ;
  assign n20186 = n20137 ^ n20133 ;
  assign n20187 = n20185 & n20186 ;
  assign n20210 = n20209 ^ n20187 ;
  assign n20212 = n20211 ^ n20210 ;
  assign n20138 = n20137 ^ n20119 ;
  assign n20139 = n20138 ^ n20136 ;
  assign n20153 = n20152 ^ n20139 ;
  assign n20177 = n20153 ^ n20152 ;
  assign n20178 = n20152 ^ n19990 ;
  assign n20179 = n20178 ^ n20152 ;
  assign n20180 = n20177 & ~n20179 ;
  assign n20181 = n20180 ^ n20152 ;
  assign n20182 = ~n20169 & n20181 ;
  assign n20213 = n20212 ^ n20182 ;
  assign n20214 = n20213 ^ n20113 ;
  assign n20170 = n20129 ^ n19989 ;
  assign n20171 = n20170 ^ n20129 ;
  assign n20174 = n20130 & ~n20171 ;
  assign n20175 = n20174 ^ n20129 ;
  assign n20176 = n20169 & n20175 ;
  assign n20215 = n20214 ^ n20176 ;
  assign n20163 = n20128 ^ n20125 ;
  assign n20164 = n20128 ^ n19989 ;
  assign n20165 = n20164 ^ n20128 ;
  assign n20166 = n20163 & ~n20165 ;
  assign n20167 = n20166 ^ n20128 ;
  assign n20168 = ~n19990 & n20167 ;
  assign n20216 = n20215 ^ n20168 ;
  assign n20217 = n20216 ^ n18875 ;
  assign n20114 = n20113 ^ n19990 ;
  assign n20115 = n20114 ^ n20113 ;
  assign n20154 = n20138 ^ n20122 ;
  assign n20155 = n20154 ^ n20056 ;
  assign n20156 = n20155 ^ n20153 ;
  assign n20157 = n20156 ^ n20145 ;
  assign n20160 = n20115 & n20157 ;
  assign n20161 = n20160 ^ n20113 ;
  assign n20162 = ~n19989 & n20161 ;
  assign n20218 = n20217 ^ n20162 ;
  assign n20219 = n20218 ^ x118 ;
  assign n20387 = n19934 & n20219 ;
  assign n20388 = n20387 ^ n19934 ;
  assign n20389 = n20388 ^ n20219 ;
  assign n20390 = n20389 ^ n19934 ;
  assign n20236 = n18435 & ~n18458 ;
  assign n20229 = n18471 ^ n18455 ;
  assign n20231 = n20230 ^ n20229 ;
  assign n20232 = ~n18434 & n20231 ;
  assign n20227 = n18462 ^ n18442 ;
  assign n20222 = n18474 ^ n18460 ;
  assign n20221 = n19668 ^ n18449 ;
  assign n20223 = n20222 ^ n20221 ;
  assign n20224 = n18434 & n20223 ;
  assign n20225 = n20224 ^ n20222 ;
  assign n20228 = n20227 ^ n20225 ;
  assign n20233 = n20232 ^ n20228 ;
  assign n20234 = ~n18393 & n20233 ;
  assign n20226 = n20225 ^ n18503 ;
  assign n20235 = n20234 ^ n20226 ;
  assign n20237 = n20236 ^ n20235 ;
  assign n20238 = ~n18518 & ~n20237 ;
  assign n20239 = ~n19686 & n20238 ;
  assign n20240 = n20239 ^ n15724 ;
  assign n20241 = n20240 ^ x107 ;
  assign n18180 = ~n17910 & n18139 ;
  assign n18181 = n18180 ^ n18138 ;
  assign n18199 = n18198 ^ n18181 ;
  assign n18190 = n18189 ^ n18169 ;
  assign n18188 = n18163 ^ n18152 ;
  assign n18191 = n18190 ^ n18188 ;
  assign n18192 = n18191 ^ n18181 ;
  assign n18182 = n18181 ^ n18156 ;
  assign n18187 = n18186 ^ n18182 ;
  assign n18193 = n18192 ^ n18187 ;
  assign n18194 = ~n17910 & n18193 ;
  assign n18195 = n18194 ^ n18192 ;
  assign n18196 = ~n17911 & ~n18195 ;
  assign n18200 = n18199 ^ n18196 ;
  assign n18201 = ~n18179 & ~n18200 ;
  assign n18202 = n18201 ^ n17346 ;
  assign n20242 = n18202 ^ x89 ;
  assign n20314 = n18950 ^ n18937 ;
  assign n20315 = n20314 ^ n18952 ;
  assign n20316 = ~n18833 & ~n20315 ;
  assign n20327 = n20316 ^ n18996 ;
  assign n20328 = n20327 ^ n18984 ;
  assign n20329 = n20328 ^ n19381 ;
  assign n20325 = n18940 & ~n19379 ;
  assign n20326 = n20325 ^ n19415 ;
  assign n20330 = n20329 ^ n20326 ;
  assign n20331 = n20330 ^ n17592 ;
  assign n20318 = n18961 ^ n18937 ;
  assign n20319 = n20318 ^ n18990 ;
  assign n20320 = n20319 ^ n20316 ;
  assign n20313 = n18956 ^ n18935 ;
  assign n20317 = n20316 ^ n20313 ;
  assign n20321 = n20320 ^ n20317 ;
  assign n20322 = ~n18833 & n20321 ;
  assign n20323 = n20322 ^ n20320 ;
  assign n20324 = n18834 & n20323 ;
  assign n20332 = n20331 ^ n20324 ;
  assign n20312 = n18939 & n19378 ;
  assign n20333 = n20332 ^ n20312 ;
  assign n20305 = n18944 ^ n18833 ;
  assign n20306 = n20305 ^ n18944 ;
  assign n20309 = n18942 & n20306 ;
  assign n20310 = n20309 ^ n18944 ;
  assign n20311 = n18834 & n20310 ;
  assign n20334 = n20333 ^ n20311 ;
  assign n20335 = n20334 ^ x66 ;
  assign n20262 = n19575 ^ n19565 ;
  assign n20245 = n19525 ^ n19517 ;
  assign n20246 = n20245 ^ n19537 ;
  assign n20247 = n19421 & ~n20246 ;
  assign n20248 = n20247 ^ n19537 ;
  assign n20263 = n20262 ^ n20248 ;
  assign n19581 = n19580 ^ n19578 ;
  assign n20259 = n20248 ^ n19581 ;
  assign n20257 = n19534 ^ n19499 ;
  assign n20258 = ~n19421 & ~n20257 ;
  assign n20260 = n20259 ^ n20258 ;
  assign n20261 = n19422 & n20260 ;
  assign n20264 = n20263 ^ n20261 ;
  assign n20254 = n19506 ^ n19498 ;
  assign n20255 = n20254 ^ n19508 ;
  assign n20256 = ~n19560 & ~n20255 ;
  assign n20265 = n20264 ^ n20256 ;
  assign n20243 = n19536 ^ n19421 ;
  assign n20244 = n20243 ^ n19536 ;
  assign n20250 = n19536 ^ n19507 ;
  assign n20251 = ~n20244 & n20250 ;
  assign n20252 = n20251 ^ n19536 ;
  assign n20253 = ~n19423 & n20252 ;
  assign n20266 = n20265 ^ n20253 ;
  assign n20267 = ~n20098 & ~n20266 ;
  assign n20268 = ~n20105 & n20267 ;
  assign n20269 = n20268 ^ n17620 ;
  assign n20270 = n20269 ^ x122 ;
  assign n20337 = n20335 ^ n20270 ;
  assign n19256 = n19183 ^ n19178 ;
  assign n19257 = ~n19035 & n19256 ;
  assign n19258 = n19257 ^ n19178 ;
  assign n19261 = n19258 ^ n19172 ;
  assign n19262 = n19261 ^ n19258 ;
  assign n19263 = ~n19035 & n19262 ;
  assign n19264 = n19263 ^ n19258 ;
  assign n19265 = ~n19073 & n19264 ;
  assign n19266 = n19265 ^ n19258 ;
  assign n19241 = n19240 ^ n19073 ;
  assign n19255 = ~n19241 & ~n19249 ;
  assign n19267 = n19266 ^ n19255 ;
  assign n19242 = n19212 ^ n19193 ;
  assign n19243 = ~n19241 & ~n19242 ;
  assign n19228 = n19227 ^ n19223 ;
  assign n19230 = n19229 ^ n19228 ;
  assign n19232 = n19231 ^ n19230 ;
  assign n19233 = n19232 ^ n19228 ;
  assign n19234 = n19228 ^ n19073 ;
  assign n19235 = n19234 ^ n19228 ;
  assign n19236 = ~n19233 & ~n19235 ;
  assign n19237 = n19236 ^ n19228 ;
  assign n19238 = n19201 & ~n19237 ;
  assign n19239 = n19238 ^ n19228 ;
  assign n19244 = n19243 ^ n19239 ;
  assign n19214 = n19213 ^ n19196 ;
  assign n19210 = n19209 ^ n19179 ;
  assign n19207 = n19206 ^ n19137 ;
  assign n19211 = n19210 ^ n19207 ;
  assign n19215 = n19214 ^ n19211 ;
  assign n19216 = n19215 ^ n19214 ;
  assign n19217 = n19216 ^ n19214 ;
  assign n19218 = n19214 ^ n19035 ;
  assign n19219 = n19218 ^ n19214 ;
  assign n19220 = ~n19217 & ~n19219 ;
  assign n19221 = n19220 ^ n19214 ;
  assign n19222 = n19073 & ~n19221 ;
  assign n19245 = n19244 ^ n19222 ;
  assign n19202 = n19186 ^ n19176 ;
  assign n19203 = ~n19073 & n19202 ;
  assign n19204 = n19203 ^ n19186 ;
  assign n19205 = n19201 & n19204 ;
  assign n19246 = n19245 ^ n19205 ;
  assign n19254 = n19246 & ~n19253 ;
  assign n19268 = n19267 ^ n19254 ;
  assign n19269 = ~n19200 & n19268 ;
  assign n19276 = n19269 & ~n19275 ;
  assign n19277 = n19276 ^ n17401 ;
  assign n20271 = n19277 ^ x96 ;
  assign n20364 = n20270 & n20271 ;
  assign n20292 = n19766 ^ n19752 ;
  assign n20293 = n20292 ^ n20025 ;
  assign n20294 = n19694 & ~n20293 ;
  assign n20281 = n19824 ^ n19763 ;
  assign n20280 = n19810 ^ n19761 ;
  assign n20282 = n20281 ^ n20280 ;
  assign n20283 = n19694 & n20282 ;
  assign n20284 = n20283 ^ n20281 ;
  assign n20290 = n20284 ^ n19752 ;
  assign n20286 = n19787 ^ n19783 ;
  assign n20289 = n20286 ^ n19773 ;
  assign n20291 = n20290 ^ n20289 ;
  assign n20295 = n20294 ^ n20291 ;
  assign n20296 = ~n19696 & ~n20295 ;
  assign n20285 = n20284 ^ n19823 ;
  assign n20287 = n20286 ^ n20285 ;
  assign n20288 = n20287 ^ n20279 ;
  assign n20297 = n20296 ^ n20288 ;
  assign n20298 = n20297 ^ n19833 ;
  assign n20273 = ~n19695 & n19791 ;
  assign n20299 = n20298 ^ n20273 ;
  assign n20300 = ~n19840 & ~n20299 ;
  assign n20301 = n20300 ^ n16159 ;
  assign n20302 = n20301 ^ x113 ;
  assign n20365 = n20364 ^ n20302 ;
  assign n20366 = ~n20337 & ~n20365 ;
  assign n20343 = n20335 ^ n20271 ;
  assign n20367 = n20366 ^ n20343 ;
  assign n20338 = n20271 & n20337 ;
  assign n20363 = n20338 ^ n20270 ;
  assign n20368 = n20367 ^ n20363 ;
  assign n20369 = n20368 ^ n20343 ;
  assign n20303 = n20302 ^ n20270 ;
  assign n20272 = n20271 ^ n20270 ;
  assign n20304 = n20303 ^ n20272 ;
  assign n20355 = n20302 & n20335 ;
  assign n20356 = n20355 ^ n20302 ;
  assign n20357 = n20337 & n20356 ;
  assign n20358 = n20357 ^ n20270 ;
  assign n20359 = ~n20304 & n20358 ;
  assign n20360 = n20359 ^ n20355 ;
  assign n20361 = n20360 ^ n20270 ;
  assign n20362 = n20361 ^ n20302 ;
  assign n20370 = n20369 ^ n20362 ;
  assign n20371 = n20370 ^ n20369 ;
  assign n20346 = n20302 ^ n20271 ;
  assign n20372 = n20364 ^ n20346 ;
  assign n20373 = n20335 & ~n20372 ;
  assign n20376 = ~n20371 & ~n20373 ;
  assign n20377 = n20376 ^ n20369 ;
  assign n20378 = n20242 & ~n20377 ;
  assign n20379 = n20378 ^ n20369 ;
  assign n20347 = ~n20335 & ~n20346 ;
  assign n20348 = n20347 ^ n20271 ;
  assign n20349 = ~n20270 & n20348 ;
  assign n20344 = n20343 ^ n20302 ;
  assign n20350 = n20349 ^ n20344 ;
  assign n20345 = n20344 ^ n20338 ;
  assign n20351 = n20350 ^ n20345 ;
  assign n20336 = n20335 ^ n20303 ;
  assign n20339 = n20338 ^ n20336 ;
  assign n20340 = n20339 ^ n20272 ;
  assign n20341 = n20304 & ~n20340 ;
  assign n20342 = n20341 ^ n20336 ;
  assign n20352 = n20351 ^ n20342 ;
  assign n20353 = ~n20242 & n20352 ;
  assign n20354 = n20353 ^ n20350 ;
  assign n20380 = n20379 ^ n20354 ;
  assign n20381 = n20241 & ~n20380 ;
  assign n20382 = n20381 ^ n20241 ;
  assign n20383 = n20382 ^ n20379 ;
  assign n20384 = n20383 ^ n17667 ;
  assign n20385 = n20384 ^ x116 ;
  assign n20391 = n20107 ^ x112 ;
  assign n20412 = n20411 ^ x105 ;
  assign n20413 = ~n20391 & n20412 ;
  assign n20414 = n20413 ^ n20412 ;
  assign n20434 = n19215 ^ n19175 ;
  assign n20438 = n20437 ^ n20434 ;
  assign n20439 = n19035 & n20438 ;
  assign n20440 = n20439 ^ n19231 ;
  assign n20441 = ~n19073 & n20440 ;
  assign n20432 = n19035 & ~n20431 ;
  assign n20418 = n19182 ^ n19173 ;
  assign n20419 = n20418 ^ n19229 ;
  assign n20420 = n19229 ^ n19073 ;
  assign n20421 = n19201 & ~n20420 ;
  assign n20422 = n20421 ^ n19073 ;
  assign n20423 = ~n20419 & n20422 ;
  assign n20424 = n20423 ^ n19229 ;
  assign n20425 = n20424 ^ n19195 ;
  assign n20426 = n20425 ^ n19186 ;
  assign n20429 = n20426 ^ n19266 ;
  assign n20415 = n19209 ^ n19206 ;
  assign n20416 = n20415 ^ n19225 ;
  assign n20417 = n19073 & ~n20416 ;
  assign n20427 = n20426 ^ n20417 ;
  assign n20428 = n19201 & n20427 ;
  assign n20430 = n20429 ^ n20428 ;
  assign n20433 = n20432 ^ n20430 ;
  assign n20442 = n20441 ^ n20433 ;
  assign n20443 = ~n19255 & ~n20442 ;
  assign n20455 = n20443 & n20454 ;
  assign n20456 = n20455 ^ n16878 ;
  assign n20457 = n20456 ^ x64 ;
  assign n20498 = n20497 ^ x81 ;
  assign n20543 = ~n20457 & ~n20498 ;
  assign n20462 = n18942 ^ n18932 ;
  assign n20463 = n20462 ^ n18957 ;
  assign n20460 = n18929 ^ n18925 ;
  assign n20461 = n18833 & n20460 ;
  assign n20464 = n20463 ^ n20461 ;
  assign n20476 = n20464 ^ n20326 ;
  assign n20477 = n20476 ^ n18977 ;
  assign n20458 = n18957 ^ n18946 ;
  assign n20459 = n20458 ^ n18951 ;
  assign n20465 = n20464 ^ n20459 ;
  assign n20466 = n20465 ^ n20464 ;
  assign n20467 = n20466 ^ n18945 ;
  assign n20468 = n20467 ^ n20466 ;
  assign n20469 = n20466 ^ n19012 ;
  assign n20470 = n20469 ^ n20466 ;
  assign n20471 = ~n20468 & ~n20470 ;
  assign n20472 = n20471 ^ n20466 ;
  assign n20473 = ~n18833 & n20472 ;
  assign n20474 = n20473 ^ n20465 ;
  assign n20475 = ~n18834 & ~n20474 ;
  assign n20478 = n20477 ^ n20475 ;
  assign n20479 = ~n19031 & ~n20478 ;
  assign n20480 = n20479 ^ n16917 ;
  assign n20481 = n20480 ^ x90 ;
  assign n20482 = ~n20457 & n20481 ;
  assign n20483 = n20482 ^ n20457 ;
  assign n20499 = n19988 ^ x115 ;
  assign n20500 = ~n20498 & n20499 ;
  assign n20501 = n20500 ^ n20498 ;
  assign n20527 = ~n20483 & ~n20501 ;
  assign n20515 = n20482 & n20500 ;
  assign n20528 = n20527 ^ n20515 ;
  assign n20544 = n20543 ^ n20528 ;
  assign n20511 = n20457 & ~n20499 ;
  assign n20512 = n20481 ^ n20457 ;
  assign n20513 = n20511 & ~n20512 ;
  assign n20524 = n20513 ^ n20512 ;
  assign n20525 = ~n20498 & ~n20524 ;
  assign n20526 = n20525 ^ n20500 ;
  assign n20529 = n20528 ^ n20526 ;
  assign n20502 = n20501 ^ n20499 ;
  assign n20504 = n20483 ^ n20481 ;
  assign n20521 = n20502 & n20504 ;
  assign n20505 = n20502 ^ n20498 ;
  assign n20519 = ~n20483 & n20505 ;
  assign n20522 = n20521 ^ n20519 ;
  assign n20506 = n20504 & n20505 ;
  assign n20523 = n20522 ^ n20506 ;
  assign n20530 = n20529 ^ n20523 ;
  assign n20520 = n20519 ^ n20504 ;
  assign n20531 = n20530 ^ n20520 ;
  assign n20534 = n20531 ^ n20515 ;
  assign n20535 = n20534 ^ n20527 ;
  assign n20509 = n20482 ^ n20481 ;
  assign n20510 = n20502 & n20509 ;
  assign n20514 = n20513 ^ n20510 ;
  assign n20516 = n20515 ^ n20514 ;
  assign n20533 = n20516 ^ n20501 ;
  assign n20536 = n20535 ^ n20533 ;
  assign n20545 = n20544 ^ n20536 ;
  assign n20546 = n20545 ^ n20534 ;
  assign n20532 = n20531 ^ n20529 ;
  assign n20542 = n20532 ^ n20500 ;
  assign n20547 = n20546 ^ n20542 ;
  assign n20548 = n20547 ^ n20536 ;
  assign n20508 = n20482 & n20502 ;
  assign n20549 = n20548 ^ n20508 ;
  assign n20540 = n20481 & n20499 ;
  assign n20541 = n20540 ^ n20482 ;
  assign n20550 = n20549 ^ n20541 ;
  assign n20612 = n20550 ^ n20531 ;
  assign n20613 = n20414 & n20612 ;
  assign n20614 = n20613 ^ n18575 ;
  assign n20606 = n20547 ^ n20510 ;
  assign n20607 = n20510 ^ n20412 ;
  assign n20608 = n20607 ^ n20510 ;
  assign n20609 = ~n20606 & n20608 ;
  assign n20610 = n20609 ^ n20510 ;
  assign n20611 = n20391 & n20610 ;
  assign n20615 = n20614 ^ n20611 ;
  assign n20579 = n20413 ^ n20391 ;
  assign n20580 = n20514 & ~n20579 ;
  assign n20551 = n20550 ^ n20522 ;
  assign n20552 = n20551 ^ n20510 ;
  assign n20537 = n20536 ^ n20532 ;
  assign n20538 = n20537 ^ n20525 ;
  assign n20517 = n20516 ^ n20508 ;
  assign n20503 = ~n20483 & n20502 ;
  assign n20507 = n20506 ^ n20503 ;
  assign n20518 = n20517 ^ n20507 ;
  assign n20539 = n20538 ^ n20518 ;
  assign n20553 = n20552 ^ n20539 ;
  assign n20565 = n20553 ^ n20521 ;
  assign n20564 = n20550 ^ n20548 ;
  assign n20566 = n20565 ^ n20564 ;
  assign n20567 = ~n20391 & n20566 ;
  assign n20568 = n20567 ^ n20549 ;
  assign n20556 = n20545 ^ n20510 ;
  assign n20577 = n20568 ^ n20556 ;
  assign n20569 = n20568 ^ n20507 ;
  assign n20570 = n20569 ^ n20550 ;
  assign n20571 = n20570 ^ n20568 ;
  assign n20574 = ~n20391 & n20571 ;
  assign n20575 = n20574 ^ n20568 ;
  assign n20576 = n20412 & n20575 ;
  assign n20578 = n20577 ^ n20576 ;
  assign n20581 = n20580 ^ n20578 ;
  assign n20557 = n20556 ^ n20530 ;
  assign n20558 = n20557 ^ n20556 ;
  assign n20559 = n20556 ^ n20391 ;
  assign n20560 = n20559 ^ n20556 ;
  assign n20561 = n20558 & n20560 ;
  assign n20562 = n20561 ^ n20556 ;
  assign n20563 = ~n20412 & ~n20562 ;
  assign n20582 = n20581 ^ n20563 ;
  assign n20583 = n20412 ^ n20391 ;
  assign n20584 = n20529 ^ n20527 ;
  assign n20585 = n20529 ^ n20412 ;
  assign n20586 = n20585 ^ n20529 ;
  assign n20587 = n20584 & n20586 ;
  assign n20588 = n20587 ^ n20529 ;
  assign n20589 = ~n20583 & n20588 ;
  assign n20590 = n20582 & ~n20589 ;
  assign n20554 = n20553 ^ n20503 ;
  assign n20555 = n20414 & n20554 ;
  assign n20591 = n20590 ^ n20555 ;
  assign n20594 = n20532 & ~n20586 ;
  assign n20595 = n20594 ^ n20529 ;
  assign n20596 = ~n20391 & n20595 ;
  assign n20597 = n20591 & ~n20596 ;
  assign n20598 = n20534 ^ n20412 ;
  assign n20599 = n20598 ^ n20534 ;
  assign n20602 = ~n20546 & ~n20599 ;
  assign n20603 = n20602 ^ n20534 ;
  assign n20604 = ~n20391 & n20603 ;
  assign n20605 = n20597 & ~n20604 ;
  assign n20616 = n20615 ^ n20605 ;
  assign n20617 = n20616 ^ x76 ;
  assign n20618 = ~n20385 & ~n20617 ;
  assign n20619 = n20618 ^ n20385 ;
  assign n20621 = n20619 ^ n20617 ;
  assign n20636 = n20621 ^ n20385 ;
  assign n20644 = n20390 & ~n20636 ;
  assign n20643 = n20387 & n20618 ;
  assign n20645 = n20644 ^ n20643 ;
  assign n20637 = n20388 & ~n20636 ;
  assign n20646 = n20645 ^ n20637 ;
  assign n18203 = n18202 ^ x74 ;
  assign n18793 = n18789 ^ n17357 ;
  assign n18790 = n18789 ^ n18756 ;
  assign n18791 = n18790 ^ n18785 ;
  assign n18792 = n18597 & n18791 ;
  assign n18794 = n18793 ^ n18792 ;
  assign n18795 = n18794 ^ n17357 ;
  assign n18754 = n18753 ^ n18597 ;
  assign n18755 = n18754 ^ n18753 ;
  assign n18778 = n18777 ^ n18756 ;
  assign n18779 = n18778 ^ n18753 ;
  assign n18780 = ~n18755 & ~n18779 ;
  assign n18781 = n18780 ^ n18753 ;
  assign n18782 = ~n18743 & ~n18781 ;
  assign n18796 = n18795 ^ n18782 ;
  assign n18797 = ~n18576 & n18796 ;
  assign n18798 = n18797 ^ n18794 ;
  assign n18799 = n18798 ^ x121 ;
  assign n18800 = n18203 & n18799 ;
  assign n18801 = n18800 ^ n18799 ;
  assign n17725 = n17686 ^ n17674 ;
  assign n17726 = n17720 & n17725 ;
  assign n17713 = n17712 ^ n17707 ;
  assign n17714 = ~n16264 & n17713 ;
  assign n17715 = n17714 ^ n17709 ;
  assign n17716 = n17668 & n17715 ;
  assign n17717 = n17716 ^ n17709 ;
  assign n17699 = n17686 ^ n17673 ;
  assign n17698 = n17689 ^ n17680 ;
  assign n17700 = n17699 ^ n17698 ;
  assign n17701 = n17699 ^ n16264 ;
  assign n17702 = n17701 ^ n17699 ;
  assign n17703 = n17700 & n17702 ;
  assign n17704 = n17703 ^ n17699 ;
  assign n17705 = ~n17697 & n17704 ;
  assign n17718 = n17717 ^ n17705 ;
  assign n17724 = n17723 ^ n17718 ;
  assign n17727 = n17726 ^ n17724 ;
  assign n17696 = n17672 & n17695 ;
  assign n17728 = n17727 ^ n17696 ;
  assign n17530 = n17529 ^ n17525 ;
  assign n17533 = n17532 ^ n17530 ;
  assign n17669 = n17533 & ~n17668 ;
  assign n17535 = n16264 & n17532 ;
  assign n17670 = n17669 ^ n17535 ;
  assign n17729 = n17728 ^ n17670 ;
  assign n17731 = n17730 ^ n17729 ;
  assign n17732 = n17731 ^ n17310 ;
  assign n17733 = n17732 ^ x120 ;
  assign n18524 = n18523 ^ x65 ;
  assign n18803 = ~n17733 & ~n18524 ;
  assign n18804 = n18803 ^ n18524 ;
  assign n18806 = n18804 ^ n17733 ;
  assign n18826 = n18801 & ~n18806 ;
  assign n18807 = n18806 ^ n18524 ;
  assign n18808 = n18800 & ~n18807 ;
  assign n18829 = n18826 ^ n18808 ;
  assign n18817 = n18800 & n18803 ;
  assign n18816 = n18801 & n18803 ;
  assign n18818 = n18817 ^ n18816 ;
  assign n18819 = n18818 ^ n18803 ;
  assign n18810 = n18801 ^ n18203 ;
  assign n18814 = n18810 ^ n18799 ;
  assign n18815 = n18803 & n18814 ;
  assign n18820 = n18819 ^ n18815 ;
  assign n18813 = ~n18806 & ~n18810 ;
  assign n18821 = n18820 ^ n18813 ;
  assign n18811 = ~n18804 & ~n18810 ;
  assign n18812 = n18811 ^ n18810 ;
  assign n18822 = n18821 ^ n18812 ;
  assign n18830 = n18829 ^ n18822 ;
  assign n18805 = n18801 & ~n18804 ;
  assign n18809 = n18808 ^ n18805 ;
  assign n18823 = n18822 ^ n18809 ;
  assign n18824 = n18823 ^ n18821 ;
  assign n18204 = n18203 ^ n17733 ;
  assign n18525 = n18524 ^ n17733 ;
  assign n18526 = ~n18204 & ~n18525 ;
  assign n18527 = n18526 ^ n18524 ;
  assign n18802 = n18801 ^ n18527 ;
  assign n18825 = n18824 ^ n18802 ;
  assign n18827 = n18826 ^ n18825 ;
  assign n18828 = n18827 ^ n18807 ;
  assign n18831 = n18830 ^ n18828 ;
  assign n18832 = n18831 ^ n18825 ;
  assign n19034 = n19033 ^ x98 ;
  assign n19278 = n19277 ^ x88 ;
  assign n19279 = n19034 & ~n19278 ;
  assign n19280 = n18832 & n19279 ;
  assign n19281 = n19278 ^ n19034 ;
  assign n19297 = ~n18806 & n18814 ;
  assign n19298 = ~n19281 & n19297 ;
  assign n19291 = n18813 ^ n18811 ;
  assign n19294 = ~n19278 & n19291 ;
  assign n19295 = n19294 ^ n18811 ;
  assign n19296 = ~n19034 & n19295 ;
  assign n19299 = n19298 ^ n19296 ;
  assign n19317 = ~n18804 & n18814 ;
  assign n19308 = n18831 ^ n18815 ;
  assign n19309 = n19308 ^ n18817 ;
  assign n19301 = n19297 ^ n18816 ;
  assign n19302 = n19301 ^ n18526 ;
  assign n19303 = n19302 ^ n18820 ;
  assign n19306 = n19303 ^ n18831 ;
  assign n19307 = n19306 ^ n18815 ;
  assign n19310 = n19309 ^ n19307 ;
  assign n19305 = n18808 ^ n18800 ;
  assign n19311 = n19310 ^ n19305 ;
  assign n19312 = n19311 ^ n18820 ;
  assign n19325 = n19317 ^ n19312 ;
  assign n19319 = n18817 ^ n18805 ;
  assign n19322 = n19279 ^ n19278 ;
  assign n19323 = n19319 & ~n19322 ;
  assign n19324 = n19323 ^ n18811 ;
  assign n19326 = n19325 ^ n19324 ;
  assign n19318 = n19317 ^ n18826 ;
  assign n19320 = n19319 ^ n19318 ;
  assign n19321 = n19034 & n19320 ;
  assign n19327 = n19326 ^ n19321 ;
  assign n19328 = n19327 ^ n19321 ;
  assign n19329 = n19319 ^ n19311 ;
  assign n19330 = ~n19279 & ~n19329 ;
  assign n19331 = n19328 & n19330 ;
  assign n19332 = n19331 ^ n19327 ;
  assign n19333 = ~n19278 & n19332 ;
  assign n19334 = n19333 ^ n19321 ;
  assign n19300 = n18832 ^ n18809 ;
  assign n19304 = n19303 ^ n19300 ;
  assign n19313 = n19312 ^ n19304 ;
  assign n19314 = n19278 & n19313 ;
  assign n19315 = n19314 ^ n19303 ;
  assign n19316 = ~n19034 & n19315 ;
  assign n19335 = n19334 ^ n19316 ;
  assign n19336 = ~n19299 & ~n19335 ;
  assign n19282 = n19279 ^ n19034 ;
  assign n19285 = n19278 ^ n18816 ;
  assign n19286 = n19285 ^ n19281 ;
  assign n19287 = n19282 & ~n19286 ;
  assign n19288 = n19287 ^ n19281 ;
  assign n19289 = ~n18815 & ~n19288 ;
  assign n19290 = n19289 ^ n19281 ;
  assign n19337 = n19336 ^ n19290 ;
  assign n19338 = ~n19280 & ~n19337 ;
  assign n19339 = n18813 ^ n18808 ;
  assign n19340 = n19339 ^ n18826 ;
  assign n19341 = n19278 & n19340 ;
  assign n19342 = n19341 ^ n18830 ;
  assign n19343 = n19281 & ~n19342 ;
  assign n19344 = n19343 ^ n18822 ;
  assign n19345 = n19338 & n19344 ;
  assign n19346 = n19345 ^ n18636 ;
  assign n19347 = n19346 ^ x101 ;
  assign n20952 = n20645 ^ n19347 ;
  assign n20953 = n20952 ^ n20645 ;
  assign n20956 = n20646 & ~n20953 ;
  assign n20957 = n20956 ^ n20645 ;
  assign n20958 = n20915 & n20957 ;
  assign n20631 = ~n20389 & ~n20619 ;
  assign n20627 = ~n20389 & ~n20621 ;
  assign n20632 = n20631 ^ n20627 ;
  assign n20622 = n20387 & ~n20621 ;
  assign n20620 = n20390 & ~n20619 ;
  assign n20623 = n20622 ^ n20620 ;
  assign n20633 = n20632 ^ n20623 ;
  assign n20629 = n20385 ^ n19934 ;
  assign n20630 = n20617 & n20629 ;
  assign n20634 = n20633 ^ n20630 ;
  assign n20628 = n20627 ^ n20617 ;
  assign n20635 = n20634 ^ n20628 ;
  assign n20638 = n20637 ^ n20635 ;
  assign n20625 = n20388 & n20618 ;
  assign n20626 = n20625 ^ n20388 ;
  assign n20639 = n20638 ^ n20626 ;
  assign n20640 = n20639 ^ n20627 ;
  assign n20624 = n20623 ^ n20617 ;
  assign n20641 = n20640 ^ n20624 ;
  assign n20220 = n20219 ^ n19934 ;
  assign n20386 = n20385 ^ n20220 ;
  assign n20642 = n20641 ^ n20386 ;
  assign n20647 = n20646 ^ n20642 ;
  assign n20654 = n20647 ^ n20644 ;
  assign n20655 = n20654 ^ n20625 ;
  assign n20921 = n20655 ^ n20618 ;
  assign n20922 = n20921 ^ n20645 ;
  assign n20648 = n20647 ^ n20389 ;
  assign n20649 = n20648 ^ n20632 ;
  assign n20923 = n20922 ^ n20649 ;
  assign n20934 = n20923 ^ n20647 ;
  assign n20932 = n20649 ^ n20637 ;
  assign n20931 = n20644 ^ n20636 ;
  assign n20933 = n20932 ^ n20931 ;
  assign n20935 = n20934 ^ n20933 ;
  assign n20929 = n20639 ^ n20622 ;
  assign n20928 = n20635 ^ n20631 ;
  assign n20930 = n20929 ^ n20928 ;
  assign n20936 = n20935 ^ n20930 ;
  assign n20937 = ~n19347 & ~n20936 ;
  assign n20938 = n20937 ^ n20935 ;
  assign n20959 = n20958 ^ n20938 ;
  assign n20939 = n20635 ^ n20623 ;
  assign n20942 = n20939 ^ n20619 ;
  assign n20943 = n20942 ^ n20930 ;
  assign n20944 = n20943 ^ n20627 ;
  assign n20651 = n20622 ^ n20619 ;
  assign n20652 = n20651 ^ n20634 ;
  assign n20941 = n20652 ^ n20622 ;
  assign n20945 = n20944 ^ n20941 ;
  assign n20946 = n20945 ^ n20938 ;
  assign n20940 = n20939 ^ n20625 ;
  assign n20947 = n20946 ^ n20940 ;
  assign n20948 = n20947 ^ n20938 ;
  assign n20949 = n19347 & n20948 ;
  assign n20950 = n20949 ^ n20946 ;
  assign n20951 = n20915 & ~n20950 ;
  assign n20960 = n20959 ^ n20951 ;
  assign n20924 = n19347 & n20915 ;
  assign n20926 = n20924 ^ n19347 ;
  assign n20927 = n20640 & n20926 ;
  assign n20961 = n20960 ^ n20927 ;
  assign n20925 = ~n20923 & n20924 ;
  assign n20962 = n20961 ^ n20925 ;
  assign n20650 = n20649 ^ n20643 ;
  assign n20653 = n20652 ^ n20650 ;
  assign n20656 = n20655 ^ n20653 ;
  assign n20918 = n20656 & ~n20915 ;
  assign n20919 = n20918 ^ n20655 ;
  assign n20920 = ~n19347 & ~n20919 ;
  assign n20963 = n20962 ^ n20920 ;
  assign n20969 = n20620 & n20926 ;
  assign n20964 = n20637 ^ n19347 ;
  assign n20965 = n20964 ^ n20637 ;
  assign n20966 = n20638 & n20965 ;
  assign n20967 = n20966 ^ n20637 ;
  assign n20968 = ~n20915 & n20967 ;
  assign n20970 = n20969 ^ n20968 ;
  assign n20971 = n20963 & ~n20970 ;
  assign n20972 = n20971 ^ n19033 ;
  assign n20973 = n19598 ^ x68 ;
  assign n20974 = n20301 ^ x117 ;
  assign n20975 = ~n20973 & n20974 ;
  assign n20976 = n20975 ^ n20973 ;
  assign n21040 = n19227 ^ n19172 ;
  assign n21039 = n20674 ^ n19204 ;
  assign n21041 = n21040 ^ n21039 ;
  assign n21042 = n21041 ^ n19204 ;
  assign n21043 = n19073 & ~n21042 ;
  assign n21044 = n21043 ^ n21039 ;
  assign n21045 = ~n19201 & n21044 ;
  assign n21034 = n19226 ^ n19204 ;
  assign n21018 = n19212 ^ n19192 ;
  assign n21019 = n21018 ^ n19073 ;
  assign n21020 = n19201 ^ n19073 ;
  assign n21021 = n21019 & ~n21020 ;
  assign n21022 = n21021 ^ n19073 ;
  assign n21023 = n19229 ^ n19213 ;
  assign n21024 = n21023 ^ n19229 ;
  assign n21025 = n21024 ^ n21018 ;
  assign n21026 = ~n21022 & n21025 ;
  assign n21027 = n21026 ^ n21023 ;
  assign n21035 = n21034 ^ n21027 ;
  assign n21029 = n19249 ^ n19187 ;
  assign n21030 = n21029 ^ n19225 ;
  assign n21031 = n19073 & n21030 ;
  assign n21017 = n19199 ^ n19187 ;
  assign n21028 = n21027 ^ n21017 ;
  assign n21032 = n21031 ^ n21028 ;
  assign n21033 = ~n19035 & n21032 ;
  assign n21036 = n21035 ^ n21033 ;
  assign n21016 = n19175 & n19240 ;
  assign n21037 = n21036 ^ n21016 ;
  assign n21009 = n19226 ^ n19210 ;
  assign n21010 = n21009 ^ n19226 ;
  assign n21011 = n19226 ^ n19073 ;
  assign n21012 = n21011 ^ n19226 ;
  assign n21013 = n21010 & n21012 ;
  assign n21014 = n21013 ^ n19226 ;
  assign n21015 = n19201 & n21014 ;
  assign n21038 = n21037 ^ n21015 ;
  assign n21046 = n21045 ^ n21038 ;
  assign n21047 = ~n19255 & n21046 ;
  assign n21048 = ~n19275 & n21047 ;
  assign n21049 = n21048 ^ n14642 ;
  assign n21050 = n21049 ^ x67 ;
  assign n21051 = n20240 ^ x92 ;
  assign n21052 = n21050 & n21051 ;
  assign n21070 = n21052 ^ n21051 ;
  assign n20977 = n19376 ^ x69 ;
  assign n20997 = n17730 ^ n17668 ;
  assign n20989 = n17692 ^ n17680 ;
  assign n20990 = n20989 ^ n17530 ;
  assign n20988 = n20769 ^ n17686 ;
  assign n20991 = n20990 ^ n20988 ;
  assign n20992 = n20990 ^ n17668 ;
  assign n20993 = n20992 ^ n20990 ;
  assign n20994 = ~n20991 & n20993 ;
  assign n20995 = n20994 ^ n20990 ;
  assign n20996 = ~n16264 & ~n20995 ;
  assign n20998 = n20997 ^ n20996 ;
  assign n20986 = n19981 ^ n17720 ;
  assign n20987 = n19985 & n20986 ;
  assign n20999 = n20998 ^ n20987 ;
  assign n20985 = n17668 & n17673 ;
  assign n21000 = n20999 ^ n20985 ;
  assign n20984 = ~n17697 & n20769 ;
  assign n21001 = n21000 ^ n20984 ;
  assign n20978 = n17691 ^ n17683 ;
  assign n20979 = n17683 ^ n16264 ;
  assign n20980 = n20979 ^ n17683 ;
  assign n20981 = n20978 & ~n20980 ;
  assign n20982 = n20981 ^ n17683 ;
  assign n20983 = n17668 & n20982 ;
  assign n21002 = n21001 ^ n20983 ;
  assign n21003 = ~n20815 & n21002 ;
  assign n21004 = n21003 ^ n15099 ;
  assign n21005 = n21004 ^ x86 ;
  assign n21006 = n20977 & ~n21005 ;
  assign n21077 = n21006 ^ n20977 ;
  assign n21080 = n21070 & n21077 ;
  assign n21074 = n21006 & n21070 ;
  assign n21081 = n21080 ^ n21074 ;
  assign n21007 = n21006 ^ n21005 ;
  assign n21071 = ~n21007 & n21070 ;
  assign n21079 = n21071 ^ n21070 ;
  assign n21082 = n21081 ^ n21079 ;
  assign n21083 = n21082 ^ n21080 ;
  assign n21078 = n21052 & n21077 ;
  assign n21084 = n21083 ^ n21078 ;
  assign n21008 = n21007 ^ n20977 ;
  assign n21073 = n21008 & n21052 ;
  assign n21075 = n21074 ^ n21073 ;
  assign n21069 = n21006 & n21052 ;
  assign n21072 = n21071 ^ n21069 ;
  assign n21076 = n21075 ^ n21072 ;
  assign n21085 = n21084 ^ n21076 ;
  assign n21086 = n21085 ^ n21051 ;
  assign n21090 = n21086 ^ n21069 ;
  assign n21053 = n21052 ^ n21050 ;
  assign n21063 = n21006 & n21053 ;
  assign n21089 = n21080 ^ n21063 ;
  assign n21091 = n21090 ^ n21089 ;
  assign n21087 = n21086 ^ n21081 ;
  assign n21088 = n21087 ^ n21006 ;
  assign n21092 = n21091 ^ n21088 ;
  assign n21061 = n21008 & n21053 ;
  assign n21093 = n21092 ^ n21061 ;
  assign n21059 = ~n21007 & n21053 ;
  assign n21094 = n21093 ^ n21059 ;
  assign n21095 = n21094 ^ n21051 ;
  assign n21056 = ~n21007 & ~n21051 ;
  assign n21060 = n21059 ^ n21056 ;
  assign n21062 = n21061 ^ n21060 ;
  assign n21064 = n21063 ^ n21062 ;
  assign n21054 = n21053 ^ n21051 ;
  assign n21057 = n21056 ^ n21054 ;
  assign n21058 = n21057 ^ n21051 ;
  assign n21065 = n21064 ^ n21058 ;
  assign n21055 = n21008 & ~n21054 ;
  assign n21066 = n21065 ^ n21055 ;
  assign n21067 = n21066 ^ n21060 ;
  assign n21068 = n21067 ^ n21063 ;
  assign n21096 = n21095 ^ n21068 ;
  assign n21097 = ~n20976 & ~n21096 ;
  assign n21140 = ~n20976 & n21082 ;
  assign n21105 = n20976 ^ n20974 ;
  assign n21137 = ~n21057 & n21105 ;
  assign n21127 = n20974 ^ n20973 ;
  assign n21132 = n21090 ^ n21075 ;
  assign n21128 = n21089 ^ n20974 ;
  assign n21129 = n21127 & ~n21128 ;
  assign n21130 = n21129 ^ n20974 ;
  assign n21131 = n21091 & n21130 ;
  assign n21133 = n21132 ^ n21131 ;
  assign n21115 = n21070 ^ n21006 ;
  assign n21116 = n21115 ^ n21061 ;
  assign n21117 = n20974 & n21116 ;
  assign n21134 = n21133 ^ n21117 ;
  assign n21135 = ~n21127 & n21134 ;
  assign n21118 = n21071 ^ n21059 ;
  assign n21119 = n21071 ^ n20973 ;
  assign n21120 = n21119 ^ n21071 ;
  assign n21121 = n21118 & ~n21120 ;
  assign n21122 = n21121 ^ n21071 ;
  assign n21123 = ~n20974 & n21122 ;
  assign n21124 = n21123 ^ n21065 ;
  assign n21125 = n21124 ^ n21117 ;
  assign n21108 = n21086 ^ n21078 ;
  assign n21109 = n21108 ^ n21096 ;
  assign n21110 = n21096 ^ n20974 ;
  assign n21111 = n21110 ^ n21096 ;
  assign n21112 = ~n21109 & ~n21111 ;
  assign n21113 = n21112 ^ n21096 ;
  assign n21114 = n20973 & ~n21113 ;
  assign n21126 = n21125 ^ n21114 ;
  assign n21136 = n21135 ^ n21126 ;
  assign n21138 = n21137 ^ n21136 ;
  assign n21106 = n21105 ^ n20973 ;
  assign n21107 = n21067 & n21106 ;
  assign n21139 = n21138 ^ n21107 ;
  assign n21141 = n21140 ^ n21139 ;
  assign n21098 = n21065 ^ n20974 ;
  assign n21099 = n21098 ^ n21065 ;
  assign n21102 = n21074 & ~n21099 ;
  assign n21103 = n21102 ^ n21065 ;
  assign n21104 = n20973 & n21103 ;
  assign n21142 = n21141 ^ n21104 ;
  assign n21143 = ~n21097 & ~n21142 ;
  assign n21144 = n21143 ^ n19169 ;
  assign n21145 = n21144 ^ x82 ;
  assign n21173 = n20129 ^ n20113 ;
  assign n21174 = n20185 & n21173 ;
  assign n21159 = ~n20184 & ~n20186 ;
  assign n21169 = n20056 & ~n20116 ;
  assign n21170 = n21159 & n21169 ;
  assign n21165 = n20156 & n20183 ;
  assign n21166 = n21165 ^ n20176 ;
  assign n21161 = n20198 ^ n20119 ;
  assign n21162 = n21161 ^ n20203 ;
  assign n21163 = n20188 & n21162 ;
  assign n21156 = n20149 ^ n20128 ;
  assign n21157 = n20188 & ~n21156 ;
  assign n21158 = n21157 ^ n20184 ;
  assign n21160 = n21159 ^ n21158 ;
  assign n21164 = n21163 ^ n21160 ;
  assign n21167 = n21166 ^ n21164 ;
  assign n21168 = n21167 ^ n20195 ;
  assign n21171 = n21170 ^ n21168 ;
  assign n21146 = n20131 ^ n20125 ;
  assign n21147 = n21146 ^ n20145 ;
  assign n21148 = n21147 ^ n20131 ;
  assign n21149 = n21148 ^ n20123 ;
  assign n21150 = n21149 ^ n21147 ;
  assign n21151 = n21147 ^ n19990 ;
  assign n21152 = n21151 ^ n21147 ;
  assign n21153 = n21150 & ~n21152 ;
  assign n21154 = n21153 ^ n21147 ;
  assign n21155 = n20169 & n21154 ;
  assign n21172 = n21171 ^ n21155 ;
  assign n21175 = n21174 ^ n21172 ;
  assign n21176 = n20149 ^ n20118 ;
  assign n21177 = n21176 ^ n20140 ;
  assign n21178 = n21177 ^ n20118 ;
  assign n21179 = n20118 ^ n19989 ;
  assign n21180 = n21179 ^ n20118 ;
  assign n21181 = ~n21178 & ~n21180 ;
  assign n21182 = n21181 ^ n20118 ;
  assign n21183 = ~n20169 & n21182 ;
  assign n21184 = n21175 & ~n21183 ;
  assign n21185 = ~n20168 & n21184 ;
  assign n21186 = n21185 ^ n18703 ;
  assign n21187 = n21186 ^ x72 ;
  assign n21188 = ~n21145 & n21187 ;
  assign n21189 = n21188 ^ n21187 ;
  assign n21509 = n21189 ^ n21145 ;
  assign n21190 = n19842 ^ x93 ;
  assign n21191 = n20818 ^ x84 ;
  assign n21286 = n21190 & n21191 ;
  assign n21287 = n21286 ^ n21191 ;
  assign n21223 = n19422 & n19581 ;
  assign n21201 = n19529 ^ n19499 ;
  assign n21200 = n20255 ^ n19509 ;
  assign n21202 = n21201 ^ n21200 ;
  assign n21203 = n21200 ^ n19421 ;
  assign n21205 = n19422 & ~n21203 ;
  assign n21206 = n21205 ^ n19421 ;
  assign n21207 = n21202 & n21206 ;
  assign n21208 = n21207 ^ n21200 ;
  assign n21217 = n21208 ^ n19591 ;
  assign n21209 = n21208 ^ n20254 ;
  assign n21210 = n21209 ^ n19525 ;
  assign n21211 = n21210 ^ n21208 ;
  assign n21212 = n21208 ^ n19421 ;
  assign n21213 = n21212 ^ n21208 ;
  assign n21214 = ~n21211 & n21213 ;
  assign n21215 = n21214 ^ n21208 ;
  assign n21216 = n19422 & ~n21215 ;
  assign n21218 = n21217 ^ n21216 ;
  assign n21199 = n19538 & n19559 ;
  assign n21219 = n21218 ^ n21199 ;
  assign n21192 = n19572 ^ n19421 ;
  assign n21193 = n21192 ^ n19572 ;
  assign n21194 = n19523 ^ n19513 ;
  assign n21195 = n21194 ^ n19572 ;
  assign n21196 = ~n21193 & n21195 ;
  assign n21197 = n21196 ^ n19572 ;
  assign n21198 = n19423 & n21197 ;
  assign n21220 = n21219 ^ n21198 ;
  assign n21221 = ~n19564 & ~n21220 ;
  assign n21222 = n21221 ^ n20087 ;
  assign n21224 = n21223 ^ n21222 ;
  assign n21225 = ~n19558 & n21224 ;
  assign n21226 = n21225 ^ n16390 ;
  assign n21227 = n21226 ^ x91 ;
  assign n21229 = ~n18576 & n19368 ;
  assign n21228 = n19363 ^ n16393 ;
  assign n21230 = n21229 ^ n21228 ;
  assign n21231 = n21230 ^ x70 ;
  assign n21232 = ~n21227 & ~n21231 ;
  assign n21233 = n21232 ^ n21231 ;
  assign n21236 = n20685 ^ x110 ;
  assign n21237 = n19418 ^ x116 ;
  assign n21238 = n21236 & n21237 ;
  assign n21249 = n21238 ^ n21236 ;
  assign n21250 = n21249 ^ n21237 ;
  assign n21265 = ~n21233 & ~n21250 ;
  assign n21234 = n21233 ^ n21227 ;
  assign n21235 = n21234 ^ n21231 ;
  assign n21262 = ~n21235 & ~n21250 ;
  assign n21257 = n21236 ^ n21231 ;
  assign n21258 = n21257 ^ n21237 ;
  assign n21259 = n21249 & ~n21258 ;
  assign n21260 = n21259 ^ n21249 ;
  assign n21256 = n21232 & n21249 ;
  assign n21261 = n21260 ^ n21256 ;
  assign n21263 = n21262 ^ n21261 ;
  assign n21291 = n21265 ^ n21263 ;
  assign n21251 = n21250 ^ n21236 ;
  assign n21252 = ~n21234 & n21251 ;
  assign n21241 = n21231 ^ n21227 ;
  assign n21242 = n21237 ^ n21231 ;
  assign n21243 = n21242 ^ n21237 ;
  assign n21244 = n21237 ^ n21236 ;
  assign n21245 = n21244 ^ n21237 ;
  assign n21246 = ~n21243 & ~n21245 ;
  assign n21247 = n21246 ^ n21237 ;
  assign n21248 = ~n21241 & n21247 ;
  assign n21253 = n21252 ^ n21248 ;
  assign n21254 = n21236 & n21253 ;
  assign n21289 = n21254 ^ n21253 ;
  assign n21290 = n21289 ^ n21261 ;
  assign n21292 = n21291 ^ n21290 ;
  assign n21324 = n21292 ^ n21250 ;
  assign n21325 = n21287 & ~n21324 ;
  assign n21295 = n21291 ^ n21235 ;
  assign n21239 = ~n21235 & n21238 ;
  assign n21240 = n21239 ^ n21238 ;
  assign n21255 = n21254 ^ n21240 ;
  assign n21269 = n21265 ^ n21255 ;
  assign n21270 = n21269 ^ n21252 ;
  assign n21267 = n21227 & ~n21244 ;
  assign n21268 = n21267 ^ n21234 ;
  assign n21271 = n21270 ^ n21268 ;
  assign n21272 = n21271 ^ n21259 ;
  assign n21273 = n21272 ^ n21261 ;
  assign n21266 = n21265 ^ n21239 ;
  assign n21274 = n21273 ^ n21266 ;
  assign n21296 = n21295 ^ n21274 ;
  assign n21323 = n21287 & n21296 ;
  assign n21326 = n21325 ^ n21323 ;
  assign n21317 = n21289 ^ n21191 ;
  assign n21318 = n21317 ^ n21289 ;
  assign n21294 = n21271 ^ n21262 ;
  assign n21297 = n21296 ^ n21294 ;
  assign n21298 = n21297 ^ n21261 ;
  assign n21293 = n21270 ^ n21239 ;
  assign n21299 = n21298 ^ n21293 ;
  assign n21277 = n21274 ^ n21258 ;
  assign n21300 = n21299 ^ n21277 ;
  assign n21301 = n21300 ^ n21292 ;
  assign n21302 = n21301 ^ n21254 ;
  assign n21319 = n21302 ^ n21289 ;
  assign n21320 = n21318 & ~n21319 ;
  assign n21321 = n21320 ^ n21289 ;
  assign n21322 = ~n21190 & n21321 ;
  assign n21327 = n21326 ^ n21322 ;
  assign n21328 = n21327 ^ n18596 ;
  assign n21303 = n21302 ^ n21256 ;
  assign n21288 = n21253 ^ n21232 ;
  assign n21304 = n21303 ^ n21288 ;
  assign n21305 = n21304 ^ n21239 ;
  assign n21306 = n21287 & ~n21305 ;
  assign n21275 = n21274 ^ n21259 ;
  assign n21276 = n21191 & n21275 ;
  assign n21278 = n21277 ^ n21276 ;
  assign n21307 = n21306 ^ n21278 ;
  assign n21279 = n21258 ^ n21248 ;
  assign n21280 = n21279 ^ n21278 ;
  assign n21264 = n21263 ^ n21255 ;
  assign n21281 = n21280 ^ n21264 ;
  assign n21282 = n21281 ^ n21278 ;
  assign n21283 = n21191 & ~n21282 ;
  assign n21284 = n21283 ^ n21280 ;
  assign n21285 = ~n21190 & n21284 ;
  assign n21308 = n21307 ^ n21285 ;
  assign n21309 = n21191 ^ n21190 ;
  assign n21310 = n21304 ^ n21294 ;
  assign n21311 = n21294 ^ n21191 ;
  assign n21312 = n21311 ^ n21294 ;
  assign n21313 = n21310 & ~n21312 ;
  assign n21314 = n21313 ^ n21294 ;
  assign n21315 = ~n21309 & ~n21314 ;
  assign n21316 = n21308 & ~n21315 ;
  assign n21329 = n21328 ^ n21316 ;
  assign n21330 = n21329 ^ x123 ;
  assign n21392 = n20519 ^ n20506 ;
  assign n21393 = n21392 ^ n20548 ;
  assign n21394 = ~n20391 & n21393 ;
  assign n21402 = n21394 ^ n20518 ;
  assign n21401 = n20543 ^ n20540 ;
  assign n21403 = n21402 ^ n21401 ;
  assign n21404 = n21403 ^ n21394 ;
  assign n21405 = n20391 & n21404 ;
  assign n21406 = n21405 ^ n21402 ;
  assign n21407 = ~n20412 & n21406 ;
  assign n21396 = n20510 & ~n20579 ;
  assign n21395 = n20414 & n20508 ;
  assign n21397 = n21396 ^ n21395 ;
  assign n21398 = n21397 ^ n21394 ;
  assign n21388 = n20529 ^ n20510 ;
  assign n21389 = ~n20608 & n21388 ;
  assign n21390 = n21389 ^ n20510 ;
  assign n21391 = n20583 & n21390 ;
  assign n21399 = n21398 ^ n21391 ;
  assign n21400 = n21399 ^ n20604 ;
  assign n21408 = n21407 ^ n21400 ;
  assign n21383 = n20550 ^ n20508 ;
  assign n21384 = n21383 ^ n20506 ;
  assign n21385 = n21384 ^ n20535 ;
  assign n21381 = n20551 ^ n20481 ;
  assign n21382 = n21381 ^ n20517 ;
  assign n21386 = n21385 ^ n21382 ;
  assign n21387 = n20414 & ~n21386 ;
  assign n21409 = n21408 ^ n21387 ;
  assign n21410 = n21409 ^ n20521 ;
  assign n21411 = n21410 ^ n20613 ;
  assign n21412 = n21411 ^ n19072 ;
  assign n21413 = n21412 ^ x114 ;
  assign n21427 = n20357 ^ n20348 ;
  assign n21428 = n21427 ^ n20369 ;
  assign n21429 = n21428 ^ n20344 ;
  assign n21430 = n21429 ^ n20342 ;
  assign n21431 = n20242 & n21430 ;
  assign n21432 = n21431 ^ n21429 ;
  assign n21435 = n21432 ^ n19747 ;
  assign n21421 = n20362 ^ n20272 ;
  assign n21422 = n21421 ^ n20367 ;
  assign n21415 = n20373 ^ n20271 ;
  assign n21416 = n21415 ^ n20360 ;
  assign n21414 = n20373 ^ n20364 ;
  assign n21417 = n21416 ^ n21414 ;
  assign n21418 = n21417 ^ n20360 ;
  assign n21419 = n20303 & n21418 ;
  assign n21420 = n21419 ^ n21416 ;
  assign n21423 = n21422 ^ n21420 ;
  assign n21424 = n21423 ^ n20367 ;
  assign n21425 = n20242 & n21424 ;
  assign n21426 = n21425 ^ n21423 ;
  assign n21433 = n21432 ^ n21426 ;
  assign n21434 = n20241 & n21433 ;
  assign n21436 = n21435 ^ n21434 ;
  assign n21437 = n21436 ^ x105 ;
  assign n21438 = ~n21413 & ~n21437 ;
  assign n21449 = n21330 & n21438 ;
  assign n21510 = n21449 ^ n21438 ;
  assign n21331 = n19860 ^ n19854 ;
  assign n21332 = n21331 ^ n19860 ;
  assign n21333 = n19860 ^ n19377 ;
  assign n21334 = n21333 ^ n19860 ;
  assign n21335 = n21332 & ~n21334 ;
  assign n21336 = n21335 ^ n19860 ;
  assign n21337 = ~n19420 & n21336 ;
  assign n21338 = n21337 ^ n19860 ;
  assign n21361 = n19899 ^ n19859 ;
  assign n21362 = n21361 ^ n19885 ;
  assign n21363 = n21362 ^ n19859 ;
  assign n21364 = n19859 ^ n19377 ;
  assign n21365 = n21364 ^ n19859 ;
  assign n21366 = ~n21363 & n21365 ;
  assign n21367 = n21366 ^ n19859 ;
  assign n21368 = n19420 & n21367 ;
  assign n21369 = n21368 ^ n19859 ;
  assign n21354 = n19926 ^ n19887 ;
  assign n21352 = n19910 ^ n19863 ;
  assign n21353 = n21352 ^ n19900 ;
  assign n21355 = n21354 ^ n21353 ;
  assign n21356 = n21353 ^ n19419 ;
  assign n21357 = n21356 ^ n21353 ;
  assign n21358 = ~n21355 & n21357 ;
  assign n21359 = n21358 ^ n21353 ;
  assign n21360 = ~n19898 & n21359 ;
  assign n21370 = n21369 ^ n21360 ;
  assign n21371 = n21370 ^ n19912 ;
  assign n21346 = n19909 ^ n19906 ;
  assign n21347 = n19906 ^ n19419 ;
  assign n21348 = n21347 ^ n19906 ;
  assign n21349 = n21346 & n21348 ;
  assign n21350 = n21349 ^ n19906 ;
  assign n21351 = n19898 & n21350 ;
  assign n21372 = n21371 ^ n21351 ;
  assign n21339 = n19912 ^ n19896 ;
  assign n21340 = n19897 ^ n19693 ;
  assign n21343 = n19912 & ~n21340 ;
  assign n21344 = n21343 ^ n19897 ;
  assign n21345 = ~n21339 & ~n21344 ;
  assign n21373 = n21372 ^ n21345 ;
  assign n21374 = ~n21338 & n21373 ;
  assign n21375 = ~n19874 & n21374 ;
  assign n21376 = ~n19894 & n21375 ;
  assign n21377 = n21376 ^ n19720 ;
  assign n21378 = n21377 ^ x104 ;
  assign n21379 = ~n21330 & n21378 ;
  assign n21380 = n21379 ^ n21378 ;
  assign n21446 = n21380 ^ n21330 ;
  assign n21448 = ~n21413 & n21446 ;
  assign n21450 = n21449 ^ n21448 ;
  assign n21439 = n21438 ^ n21413 ;
  assign n21447 = ~n21439 & n21446 ;
  assign n21451 = n21450 ^ n21447 ;
  assign n21444 = n21379 & ~n21439 ;
  assign n21452 = n21451 ^ n21444 ;
  assign n21443 = n21380 & ~n21439 ;
  assign n21445 = n21444 ^ n21443 ;
  assign n21453 = n21452 ^ n21445 ;
  assign n21511 = n21510 ^ n21453 ;
  assign n21512 = n21509 & n21511 ;
  assign n21440 = n21439 ^ n21437 ;
  assign n21441 = n21380 & ~n21440 ;
  assign n21442 = n21441 ^ n21380 ;
  assign n21454 = n21453 ^ n21442 ;
  assign n21455 = n21189 & n21454 ;
  assign n21456 = n21379 & ~n21440 ;
  assign n21457 = n21145 & n21456 ;
  assign n21458 = n21187 ^ n21145 ;
  assign n21487 = n21447 ^ n21439 ;
  assign n21488 = n21487 ^ n21445 ;
  assign n21460 = n21379 ^ n21330 ;
  assign n21461 = ~n21440 & ~n21460 ;
  assign n21462 = n21461 ^ n21441 ;
  assign n21463 = n21462 ^ n21440 ;
  assign n21464 = n21463 ^ n21456 ;
  assign n21475 = n21464 ^ n21451 ;
  assign n21470 = n21437 ^ n21413 ;
  assign n21472 = n21413 ^ n21378 ;
  assign n21473 = n21472 ^ n21330 ;
  assign n21474 = ~n21470 & n21473 ;
  assign n21476 = n21475 ^ n21474 ;
  assign n21471 = n21470 ^ n21456 ;
  assign n21477 = n21476 ^ n21471 ;
  assign n21478 = n21477 ^ n21447 ;
  assign n21479 = n21478 ^ n21413 ;
  assign n21480 = n21479 ^ n21452 ;
  assign n21468 = n21437 ^ n21330 ;
  assign n21469 = n21468 ^ n21378 ;
  assign n21481 = n21480 ^ n21469 ;
  assign n21459 = n21448 ^ n21446 ;
  assign n21465 = n21464 ^ n21459 ;
  assign n21466 = n21465 ^ n21462 ;
  assign n21482 = n21481 ^ n21466 ;
  assign n21500 = n21488 ^ n21482 ;
  assign n21501 = n21500 ^ n21449 ;
  assign n21499 = n21447 ^ n21413 ;
  assign n21502 = n21501 ^ n21499 ;
  assign n21503 = ~n21145 & n21502 ;
  assign n21497 = n21461 ^ n21459 ;
  assign n21483 = n21482 ^ n21454 ;
  assign n21484 = n21483 ^ n21464 ;
  assign n21485 = n21484 ^ n21456 ;
  assign n21467 = n21466 ^ n21413 ;
  assign n21486 = n21485 ^ n21467 ;
  assign n21489 = n21488 ^ n21441 ;
  assign n21490 = n21489 ^ n21483 ;
  assign n21491 = n21488 ^ n21187 ;
  assign n21492 = n21458 & n21491 ;
  assign n21493 = n21492 ^ n21187 ;
  assign n21494 = ~n21490 & ~n21493 ;
  assign n21495 = n21494 ^ n21488 ;
  assign n21496 = ~n21486 & n21495 ;
  assign n21498 = n21497 ^ n21496 ;
  assign n21504 = n21503 ^ n21498 ;
  assign n21505 = n21458 & ~n21504 ;
  assign n21506 = n21505 ^ n21496 ;
  assign n21507 = ~n21457 & n21506 ;
  assign n21508 = ~n21455 & n21507 ;
  assign n21513 = n21512 ^ n21508 ;
  assign n21514 = n21458 ^ n21448 ;
  assign n21516 = n21452 ^ n21448 ;
  assign n21515 = n21452 ^ n21187 ;
  assign n21517 = n21516 ^ n21515 ;
  assign n21518 = n21516 ^ n21453 ;
  assign n21519 = n21518 ^ n21516 ;
  assign n21520 = ~n21517 & n21519 ;
  assign n21521 = n21520 ^ n21516 ;
  assign n21522 = ~n21514 & n21521 ;
  assign n21523 = n21522 ^ n21448 ;
  assign n21524 = n21513 & ~n21523 ;
  assign n21525 = n21524 ^ n20301 ;
  assign n21526 = n21525 ^ x93 ;
  assign n21536 = n19989 & n20126 ;
  assign n21544 = n21536 ^ n20157 ;
  assign n21542 = n20123 & ~n20184 ;
  assign n21543 = n21542 ^ n21157 ;
  assign n21545 = n21544 ^ n21543 ;
  assign n21538 = n20141 ^ n20113 ;
  assign n21539 = ~n19989 & n21538 ;
  assign n21534 = n20134 ^ n20113 ;
  assign n21535 = n21534 ^ n20152 ;
  assign n21537 = n21536 ^ n21535 ;
  assign n21540 = n21539 ^ n21537 ;
  assign n21541 = n20169 & n21540 ;
  assign n21546 = n21545 ^ n21541 ;
  assign n21529 = n20157 ^ n19990 ;
  assign n21530 = n21529 ^ n20157 ;
  assign n21531 = n20198 & ~n21530 ;
  assign n21532 = n21531 ^ n20157 ;
  assign n21533 = ~n19989 & n21532 ;
  assign n21547 = n21546 ^ n21533 ;
  assign n21548 = ~n21174 & ~n21547 ;
  assign n21549 = ~n21183 & n21548 ;
  assign n21550 = ~n20197 & n21549 ;
  assign n21551 = ~n20168 & n21550 ;
  assign n21552 = n21551 ^ n18108 ;
  assign n21553 = n21552 ^ x124 ;
  assign n21554 = n21425 ^ n21420 ;
  assign n21555 = n21554 ^ n21432 ;
  assign n21556 = n21432 ^ n20241 ;
  assign n21557 = n21556 ^ n21432 ;
  assign n21558 = n21555 & ~n21557 ;
  assign n21559 = n21558 ^ n21432 ;
  assign n21560 = n21422 & n21559 ;
  assign n21561 = n21560 ^ n18316 ;
  assign n21562 = n21561 ^ x110 ;
  assign n21711 = n21553 & n21562 ;
  assign n21712 = n21711 ^ n21562 ;
  assign n21713 = n21712 ^ n21553 ;
  assign n21584 = n21351 ^ n19857 ;
  assign n21576 = n19910 ^ n19907 ;
  assign n21577 = n21576 ^ n19909 ;
  assign n21581 = n21577 ^ n19886 ;
  assign n21575 = n19887 ^ n19850 ;
  assign n21578 = n21577 ^ n21575 ;
  assign n21571 = n19855 ^ n19690 ;
  assign n21572 = n21571 ^ n19885 ;
  assign n21573 = n21572 ^ n19881 ;
  assign n21574 = n21573 ^ n19856 ;
  assign n21579 = n21578 ^ n21574 ;
  assign n21580 = ~n19419 & n21579 ;
  assign n21582 = n21581 ^ n21580 ;
  assign n21583 = ~n19898 & ~n21582 ;
  assign n21585 = n21584 ^ n21583 ;
  assign n21570 = ~n19419 & n19856 ;
  assign n21586 = n21585 ^ n21570 ;
  assign n21563 = n19896 ^ n19857 ;
  assign n21564 = n19906 ^ n19897 ;
  assign n21565 = n19897 ^ n19857 ;
  assign n21566 = n21565 ^ n19897 ;
  assign n21567 = ~n21564 & ~n21566 ;
  assign n21568 = n21567 ^ n19897 ;
  assign n21569 = n21563 & ~n21568 ;
  assign n21587 = n21586 ^ n21569 ;
  assign n21588 = ~n19902 & ~n21587 ;
  assign n21589 = ~n21338 & n21588 ;
  assign n21590 = n21589 ^ n17909 ;
  assign n21591 = n21590 ^ x93 ;
  assign n21600 = n18827 ^ n18813 ;
  assign n21601 = n21600 ^ n19301 ;
  assign n21602 = n19034 & ~n21601 ;
  assign n21603 = n21602 ^ n19301 ;
  assign n21610 = n21603 ^ n19317 ;
  assign n21611 = n21610 ^ n19290 ;
  assign n21605 = n19311 ^ n18822 ;
  assign n21606 = n21605 ^ n19319 ;
  assign n21607 = n19034 & ~n21606 ;
  assign n21599 = n19319 ^ n18820 ;
  assign n21604 = n21603 ^ n21599 ;
  assign n21608 = n21607 ^ n21604 ;
  assign n21609 = n19281 & n21608 ;
  assign n21612 = n21611 ^ n21609 ;
  assign n21592 = n19317 ^ n19306 ;
  assign n21593 = n19322 ^ n19282 ;
  assign n21594 = n21593 ^ n19279 ;
  assign n21595 = n19306 ^ n19279 ;
  assign n21596 = n21594 & ~n21595 ;
  assign n21597 = n21596 ^ n19279 ;
  assign n21598 = ~n21592 & n21597 ;
  assign n21613 = n21612 ^ n21598 ;
  assign n21614 = n19297 ^ n18817 ;
  assign n21615 = n21614 ^ n19306 ;
  assign n21616 = n19306 ^ n19278 ;
  assign n21617 = n21616 ^ n19306 ;
  assign n21618 = ~n21615 & ~n21617 ;
  assign n21619 = n21618 ^ n19306 ;
  assign n21620 = n19034 & ~n21619 ;
  assign n21621 = n21613 & ~n21620 ;
  assign n21622 = n18827 ^ n18808 ;
  assign n21625 = ~n19278 & ~n21622 ;
  assign n21626 = n21625 ^ n18827 ;
  assign n21627 = ~n19034 & ~n21626 ;
  assign n21628 = n21621 & ~n21627 ;
  assign n21629 = n21628 ^ n19323 ;
  assign n21630 = ~n18826 & n21629 ;
  assign n21631 = n21630 ^ n19454 ;
  assign n21632 = n21631 ^ x92 ;
  assign n21633 = n21591 & ~n21632 ;
  assign n21714 = n21633 ^ n21632 ;
  assign n21715 = n21714 ^ n21591 ;
  assign n21716 = n21715 ^ n21632 ;
  assign n21634 = n21286 ^ n21190 ;
  assign n21653 = n21279 ^ n21267 ;
  assign n21651 = n21261 ^ n21233 ;
  assign n21652 = n21651 ^ n21269 ;
  assign n21654 = n21653 ^ n21652 ;
  assign n21655 = n21634 & n21654 ;
  assign n21647 = n21289 ^ n21255 ;
  assign n21644 = n21254 ^ n21244 ;
  assign n21645 = n21644 ^ n21227 ;
  assign n21646 = n21191 & ~n21645 ;
  assign n21648 = n21647 ^ n21646 ;
  assign n21649 = ~n21309 & n21648 ;
  assign n21650 = n21649 ^ n21647 ;
  assign n21656 = n21655 ^ n21650 ;
  assign n21637 = n21301 ^ n21252 ;
  assign n21638 = n21637 ^ n21277 ;
  assign n21639 = n21277 ^ n21191 ;
  assign n21640 = n21639 ^ n21277 ;
  assign n21641 = n21638 & n21640 ;
  assign n21642 = n21641 ^ n21277 ;
  assign n21643 = ~n21190 & ~n21642 ;
  assign n21657 = n21656 ^ n21643 ;
  assign n21636 = ~n21273 & n21287 ;
  assign n21658 = n21657 ^ n21636 ;
  assign n21659 = n21658 ^ n21325 ;
  assign n21660 = n21659 ^ n21323 ;
  assign n21661 = n21660 ^ n18392 ;
  assign n21635 = ~n21302 & n21634 ;
  assign n21662 = n21661 ^ n21635 ;
  assign n21663 = n21662 ^ x67 ;
  assign n21681 = n20414 & n20506 ;
  assign n21678 = n20522 ^ n20503 ;
  assign n21679 = n20413 & n21678 ;
  assign n21664 = n20412 & ~n20538 ;
  assign n21665 = n21664 ^ n20525 ;
  assign n21674 = n21665 ^ n20596 ;
  assign n21667 = n21665 ^ n20551 ;
  assign n21666 = n21665 ^ n20517 ;
  assign n21668 = n21667 ^ n21666 ;
  assign n21669 = n21667 ^ n20391 ;
  assign n21670 = n21669 ^ n21667 ;
  assign n21671 = n21668 & ~n21670 ;
  assign n21672 = n21671 ^ n21667 ;
  assign n21673 = n20583 & n21672 ;
  assign n21675 = n21674 ^ n21673 ;
  assign n21676 = ~n20611 & ~n21675 ;
  assign n21677 = n21676 ^ n21397 ;
  assign n21680 = n21679 ^ n21677 ;
  assign n21682 = n21681 ^ n21680 ;
  assign n21683 = n21682 ^ n21397 ;
  assign n21686 = n20535 ^ n20391 ;
  assign n21687 = n21686 ^ n20535 ;
  assign n21688 = n21385 & ~n21687 ;
  assign n21689 = n21688 ^ n20535 ;
  assign n21690 = ~n20412 & n21689 ;
  assign n21691 = n21683 & n21690 ;
  assign n21692 = n21691 ^ n21682 ;
  assign n21693 = ~n20555 & n21692 ;
  assign n21694 = ~n21391 & n21693 ;
  assign n21695 = n21694 ^ n19491 ;
  assign n21696 = n21695 ^ x78 ;
  assign n21697 = n21663 & n21696 ;
  assign n21717 = n21697 ^ n21663 ;
  assign n21718 = n21716 & n21717 ;
  assign n21719 = ~n21713 & n21718 ;
  assign n21698 = n21697 ^ n21696 ;
  assign n21699 = n21698 ^ n21663 ;
  assign n21700 = n21633 & ~n21699 ;
  assign n21701 = n21700 ^ n21562 ;
  assign n21702 = n21701 ^ n21700 ;
  assign n21703 = n21696 ^ n21663 ;
  assign n21704 = n21633 & n21703 ;
  assign n21705 = n21704 ^ n21700 ;
  assign n21708 = n21702 & n21705 ;
  assign n21709 = n21708 ^ n21700 ;
  assign n21710 = ~n21553 & n21709 ;
  assign n21720 = n21719 ^ n21710 ;
  assign n21721 = n21713 ^ n21562 ;
  assign n21722 = n21718 & n21721 ;
  assign n21727 = n21698 & n21715 ;
  assign n21726 = n21715 & n21717 ;
  assign n21728 = n21727 ^ n21726 ;
  assign n21724 = n21697 & n21715 ;
  assign n21725 = n21724 ^ n21715 ;
  assign n21729 = n21728 ^ n21725 ;
  assign n21723 = ~n21714 & n21717 ;
  assign n21730 = n21729 ^ n21723 ;
  assign n21731 = n21730 ^ n21727 ;
  assign n21732 = ~n21713 & n21731 ;
  assign n21733 = n21724 ^ n21700 ;
  assign n21734 = n21700 ^ n21553 ;
  assign n21735 = n21734 ^ n21700 ;
  assign n21736 = n21733 & n21735 ;
  assign n21737 = n21736 ^ n21700 ;
  assign n21738 = n21562 & n21737 ;
  assign n21772 = n21705 ^ n21633 ;
  assign n21748 = n21698 & n21716 ;
  assign n21773 = n21772 ^ n21748 ;
  assign n21774 = n21773 ^ n21718 ;
  assign n21775 = n21718 ^ n21562 ;
  assign n21776 = n21775 ^ n21718 ;
  assign n21777 = n21774 & ~n21776 ;
  assign n21778 = n21777 ^ n21718 ;
  assign n21779 = ~n21553 & n21778 ;
  assign n21741 = n21698 & ~n21714 ;
  assign n21763 = n21741 ^ n21712 ;
  assign n21749 = n21697 & n21716 ;
  assign n21764 = n21749 ^ n21721 ;
  assign n21767 = ~n21741 & ~n21764 ;
  assign n21768 = n21767 ^ n21721 ;
  assign n21769 = n21763 & n21768 ;
  assign n21770 = n21769 ^ n21712 ;
  assign n21742 = n21741 ^ n21729 ;
  assign n21743 = n21742 ^ n21714 ;
  assign n21739 = ~n21699 & ~n21714 ;
  assign n21740 = n21739 ^ n21730 ;
  assign n21744 = n21743 ^ n21740 ;
  assign n21745 = n21633 & ~n21696 ;
  assign n21746 = n21745 ^ n21705 ;
  assign n21750 = n21749 ^ n21746 ;
  assign n21755 = n21750 ^ n21739 ;
  assign n21751 = n21750 ^ n21748 ;
  assign n21752 = n21751 ^ n21718 ;
  assign n21747 = n21746 ^ n21716 ;
  assign n21753 = n21752 ^ n21747 ;
  assign n21754 = n21753 ^ n21723 ;
  assign n21756 = n21755 ^ n21754 ;
  assign n21757 = n21754 ^ n21562 ;
  assign n21758 = n21757 ^ n21754 ;
  assign n21759 = n21756 & ~n21758 ;
  assign n21760 = n21759 ^ n21754 ;
  assign n21761 = n21744 & ~n21760 ;
  assign n21762 = n21553 & ~n21761 ;
  assign n21771 = n21770 ^ n21762 ;
  assign n21780 = n21779 ^ n21771 ;
  assign n21781 = n21780 ^ n21562 ;
  assign n21782 = n21781 ^ n21780 ;
  assign n21783 = n21780 ^ n21724 ;
  assign n21784 = n21783 ^ n21780 ;
  assign n21788 = ~n21782 & n21784 ;
  assign n21789 = n21788 ^ n21782 ;
  assign n21790 = n21789 ^ n21781 ;
  assign n21791 = ~n21738 & ~n21790 ;
  assign n21792 = n21773 ^ n21753 ;
  assign n21793 = n21753 ^ n21562 ;
  assign n21794 = n21793 ^ n21753 ;
  assign n21795 = n21792 & n21794 ;
  assign n21796 = n21795 ^ n21753 ;
  assign n21797 = n21553 & n21796 ;
  assign n21798 = n21791 & ~n21797 ;
  assign n21799 = ~n21732 & n21798 ;
  assign n21800 = ~n21722 & n21799 ;
  assign n21801 = ~n21720 & n21800 ;
  assign n21803 = n21739 ^ n21726 ;
  assign n21802 = n21727 ^ n21723 ;
  assign n21804 = n21803 ^ n21802 ;
  assign n21805 = n21803 ^ n21553 ;
  assign n21806 = n21805 ^ n21803 ;
  assign n21807 = n21804 & ~n21806 ;
  assign n21808 = n21807 ^ n21803 ;
  assign n21809 = n21562 & n21808 ;
  assign n21810 = n21801 & ~n21809 ;
  assign n21811 = n21810 ^ n19598 ;
  assign n21812 = n21811 ^ x75 ;
  assign n22633 = n21526 & ~n21812 ;
  assign n22634 = n22633 ^ n21812 ;
  assign n22459 = n20616 ^ x120 ;
  assign n22460 = n21329 ^ x73 ;
  assign n22490 = n21186 ^ x80 ;
  assign n22473 = n21082 ^ n21053 ;
  assign n22474 = n22473 ^ n21060 ;
  assign n22475 = n22474 ^ n21055 ;
  assign n22476 = n20974 & n22475 ;
  assign n22477 = n22476 ^ n21064 ;
  assign n22478 = ~n20973 & n22477 ;
  assign n22479 = n22478 ^ n21097 ;
  assign n22472 = n21072 & n21127 ;
  assign n22480 = n22479 ^ n22472 ;
  assign n22469 = n21083 ^ n21065 ;
  assign n21946 = n21092 ^ n21060 ;
  assign n22470 = n22469 ^ n21946 ;
  assign n22471 = n21106 & n22470 ;
  assign n22481 = n22480 ^ n22471 ;
  assign n22482 = n22481 ^ n21073 ;
  assign n21974 = n21108 ^ n21094 ;
  assign n21975 = n21094 ^ n20974 ;
  assign n21976 = n21975 ^ n21094 ;
  assign n21977 = n21974 & n21976 ;
  assign n21978 = n21977 ^ n21094 ;
  assign n21979 = n20973 & n21978 ;
  assign n22483 = n22482 ^ n21979 ;
  assign n22468 = ~n20976 & n21087 ;
  assign n22484 = n22483 ^ n22468 ;
  assign n22461 = n21073 ^ n21066 ;
  assign n22462 = n22461 ^ n21073 ;
  assign n22463 = n21073 ^ n20974 ;
  assign n22464 = n22463 ^ n21073 ;
  assign n22465 = n22462 & ~n22464 ;
  assign n22466 = n22465 ^ n21073 ;
  assign n22467 = n20973 & n22466 ;
  assign n22485 = n22484 ^ n22467 ;
  assign n21937 = n20975 & n21074 ;
  assign n21942 = n21082 ^ n21063 ;
  assign n21943 = n20974 & n21942 ;
  assign n21944 = n21943 ^ n21082 ;
  assign n21945 = n20973 & n21944 ;
  assign n22486 = ~n21937 & ~n21945 ;
  assign n22487 = ~n22485 & n22486 ;
  assign n22488 = n22487 ^ n18733 ;
  assign n22489 = n22488 ^ x115 ;
  assign n22550 = n22490 ^ n22489 ;
  assign n22493 = n19346 ^ x97 ;
  assign n22553 = n22550 ^ n22493 ;
  assign n22150 = n20878 & n20898 ;
  assign n22494 = ~n20886 & ~n22150 ;
  assign n22502 = n20836 ^ n20822 ;
  assign n22503 = n20857 & ~n20888 ;
  assign n22504 = n20862 & n22503 ;
  assign n22505 = n22502 & n22504 ;
  assign n22506 = n22505 ^ n22503 ;
  assign n22507 = n22506 ^ n20888 ;
  assign n22508 = n22507 ^ n20851 ;
  assign n22496 = n20830 ^ n20826 ;
  assign n22151 = n20845 ^ n20837 ;
  assign n22497 = n22496 ^ n22151 ;
  assign n22495 = n20860 ^ n20854 ;
  assign n22498 = n22497 ^ n22495 ;
  assign n22499 = ~n20862 & n22498 ;
  assign n22500 = n22499 ^ n20851 ;
  assign n22501 = n20686 & n22500 ;
  assign n22509 = n22508 ^ n22501 ;
  assign n22510 = n20849 ^ n20686 ;
  assign n22511 = n22510 ^ n20849 ;
  assign n22514 = ~n20843 & ~n20862 ;
  assign n22515 = n22514 ^ n20849 ;
  assign n22516 = ~n22511 & n22515 ;
  assign n22517 = n22516 ^ n20849 ;
  assign n22518 = n22509 & ~n22517 ;
  assign n22180 = n20855 ^ n20843 ;
  assign n22181 = n22180 ^ n20855 ;
  assign n22182 = n20862 & ~n22181 ;
  assign n22183 = n22182 ^ n20855 ;
  assign n22184 = ~n20686 & n22183 ;
  assign n22519 = n22518 ^ n22184 ;
  assign n22520 = n22494 & n22519 ;
  assign n22521 = n22520 ^ n18669 ;
  assign n22522 = n22521 ^ x106 ;
  assign n22565 = n22493 & ~n22522 ;
  assign n22566 = n22565 ^ n22490 ;
  assign n22567 = n22553 & n22566 ;
  assign n22528 = n22522 ^ n22490 ;
  assign n22568 = n22567 ^ n22528 ;
  assign n22523 = n22522 ^ n22493 ;
  assign n22554 = n22493 ^ n22490 ;
  assign n22557 = n22523 & n22554 ;
  assign n22558 = n22557 ^ n22490 ;
  assign n22559 = ~n22553 & n22558 ;
  assign n22560 = n22559 ^ n22550 ;
  assign n22569 = n22568 ^ n22560 ;
  assign n22491 = ~n22489 & ~n22490 ;
  assign n22492 = n22491 ^ n22489 ;
  assign n22525 = n22493 ^ n22489 ;
  assign n22526 = n22525 ^ n22523 ;
  assign n22527 = n22525 ^ n22522 ;
  assign n22529 = ~n22527 & n22528 ;
  assign n22530 = n22529 ^ n22522 ;
  assign n22531 = ~n22526 & ~n22530 ;
  assign n22532 = n22531 ^ n22523 ;
  assign n22533 = n22491 & n22532 ;
  assign n22524 = n22493 & n22523 ;
  assign n22534 = n22533 ^ n22524 ;
  assign n22535 = n22534 ^ n22493 ;
  assign n22536 = n22535 ^ n22522 ;
  assign n22537 = n22536 ^ n22534 ;
  assign n22538 = n22492 & ~n22537 ;
  assign n22539 = n22538 ^ n22535 ;
  assign n22562 = n22539 ^ n22490 ;
  assign n22570 = n22569 ^ n22562 ;
  assign n22571 = n22570 ^ n22527 ;
  assign n22561 = n22553 ^ n22534 ;
  assign n22572 = n22571 ^ n22561 ;
  assign n22573 = n22572 ^ n22560 ;
  assign n22574 = n22460 & ~n22573 ;
  assign n22575 = n22574 ^ n22571 ;
  assign n22551 = n22550 ^ n22539 ;
  assign n22540 = n22523 ^ n22489 ;
  assign n22541 = n22540 ^ n22539 ;
  assign n22542 = n22541 ^ n22524 ;
  assign n22543 = n22542 ^ n22489 ;
  assign n22544 = n22543 ^ n22541 ;
  assign n22545 = n22541 ^ n22490 ;
  assign n22546 = n22545 ^ n22541 ;
  assign n22547 = ~n22544 & ~n22546 ;
  assign n22548 = n22547 ^ n22541 ;
  assign n22549 = n22460 & n22548 ;
  assign n22552 = n22551 ^ n22549 ;
  assign n22576 = n22575 ^ n22552 ;
  assign n22577 = ~n22459 & ~n22576 ;
  assign n22578 = n22577 ^ n22459 ;
  assign n22579 = n22578 ^ n22552 ;
  assign n22580 = n22579 ^ n19376 ;
  assign n22581 = n22580 ^ x108 ;
  assign n21936 = n20384 ^ x126 ;
  assign n21898 = n20914 ^ x109 ;
  assign n21910 = n18816 ^ n18805 ;
  assign n21911 = n19279 & n21910 ;
  assign n21905 = n19344 ^ n18816 ;
  assign n21906 = n21905 ^ n21620 ;
  assign n21907 = n21906 ^ n21627 ;
  assign n21900 = n18799 ^ n18524 ;
  assign n21901 = n21900 ^ n18203 ;
  assign n21902 = n21901 ^ n17733 ;
  assign n21903 = ~n18527 & ~n19281 ;
  assign n21904 = n21902 & n21903 ;
  assign n21908 = n21907 ^ n21904 ;
  assign n21899 = ~n18825 & ~n19322 ;
  assign n21909 = n21908 ^ n21899 ;
  assign n21912 = n21911 ^ n21909 ;
  assign n21913 = n19317 ^ n18821 ;
  assign n21914 = n21913 ^ n18824 ;
  assign n21915 = n21914 ^ n21913 ;
  assign n21916 = n21913 ^ n19034 ;
  assign n21917 = n21916 ^ n21913 ;
  assign n21918 = ~n21915 & ~n21917 ;
  assign n21919 = n21918 ^ n21913 ;
  assign n21920 = n19281 & n21919 ;
  assign n21921 = n21912 & ~n21920 ;
  assign n21922 = n21921 ^ n17521 ;
  assign n21923 = n21922 ^ x102 ;
  assign n21924 = n21898 & n21923 ;
  assign n21925 = n21924 ^ n21898 ;
  assign n21844 = n20613 ^ n17071 ;
  assign n21845 = n21844 ^ n20611 ;
  assign n21839 = ~n20391 & ~n20545 ;
  assign n21838 = n20412 & n20516 ;
  assign n21840 = n21839 ^ n21838 ;
  assign n21814 = n20527 ^ n20481 ;
  assign n21815 = n21814 ^ n20551 ;
  assign n21816 = ~n20412 & ~n21815 ;
  assign n21817 = n21816 ^ n20536 ;
  assign n21818 = n20583 & ~n21817 ;
  assign n21819 = ~n20528 & ~n20552 ;
  assign n21820 = n20565 ^ n20507 ;
  assign n21821 = n20412 & n21820 ;
  assign n21822 = n21821 ^ n20413 ;
  assign n21823 = n21822 ^ n20391 ;
  assign n21824 = n21823 ^ n21821 ;
  assign n21825 = n21819 & ~n21824 ;
  assign n21826 = n21825 ^ n21822 ;
  assign n21827 = n21826 ^ n20391 ;
  assign n21828 = n21827 ^ n21826 ;
  assign n21829 = n21827 ^ n20506 ;
  assign n21830 = n21829 ^ n21827 ;
  assign n21831 = n21827 ^ n21821 ;
  assign n21832 = n21831 ^ n21827 ;
  assign n21833 = ~n21830 & n21832 ;
  assign n21834 = n21828 & n21833 ;
  assign n21835 = n21834 ^ n21828 ;
  assign n21836 = n21835 ^ n21826 ;
  assign n21837 = ~n21818 & n21836 ;
  assign n21841 = n21840 ^ n21837 ;
  assign n21842 = n21841 ^ n21395 ;
  assign n21843 = ~n20589 & n21842 ;
  assign n21846 = n21845 ^ n21843 ;
  assign n21847 = n21846 ^ x69 ;
  assign n21894 = n21325 ^ n16654 ;
  assign n21876 = n21290 ^ n21272 ;
  assign n21877 = n21876 ^ n21265 ;
  assign n21874 = n21294 ^ n21269 ;
  assign n21875 = n21874 ^ n21637 ;
  assign n21878 = n21877 ^ n21875 ;
  assign n21879 = ~n21190 & ~n21878 ;
  assign n21880 = n21879 ^ n21877 ;
  assign n21881 = ~n21191 & ~n21880 ;
  assign n21853 = n21652 ^ n21255 ;
  assign n21854 = n21853 ^ n21304 ;
  assign n21855 = n21304 ^ n21191 ;
  assign n21856 = n21309 ^ n21191 ;
  assign n21857 = ~n21855 & ~n21856 ;
  assign n21858 = n21857 ^ n21191 ;
  assign n21859 = n21854 & n21858 ;
  assign n21860 = n21859 ^ n21304 ;
  assign n21861 = n21860 ^ n21239 ;
  assign n21862 = n21861 ^ n21296 ;
  assign n21871 = n21862 ^ n21306 ;
  assign n21863 = n21862 ^ n21301 ;
  assign n21864 = n21863 ^ n21265 ;
  assign n21865 = n21864 ^ n21862 ;
  assign n21866 = n21862 ^ n21191 ;
  assign n21867 = n21866 ^ n21862 ;
  assign n21868 = ~n21865 & n21867 ;
  assign n21869 = n21868 ^ n21862 ;
  assign n21870 = ~n21190 & ~n21869 ;
  assign n21872 = n21871 ^ n21870 ;
  assign n21852 = n21286 & ~n21324 ;
  assign n21873 = n21872 ^ n21852 ;
  assign n21882 = n21881 ^ n21873 ;
  assign n21883 = ~n21315 & n21882 ;
  assign n21848 = n21271 ^ n21256 ;
  assign n21849 = ~n21190 & ~n21848 ;
  assign n21850 = n21849 ^ n21256 ;
  assign n21851 = n21191 & n21850 ;
  assign n21884 = n21883 ^ n21851 ;
  assign n21885 = ~n21636 & n21884 ;
  assign n21888 = n21256 ^ n21190 ;
  assign n21889 = n21888 ^ n21256 ;
  assign n21890 = ~n21303 & n21889 ;
  assign n21891 = n21890 ^ n21256 ;
  assign n21892 = ~n21191 & n21891 ;
  assign n21893 = n21885 & ~n21892 ;
  assign n21895 = n21894 ^ n21893 ;
  assign n21896 = n21895 ^ x84 ;
  assign n21897 = ~n21847 & n21896 ;
  assign n21928 = n21897 ^ n21847 ;
  assign n21929 = n21928 ^ n21896 ;
  assign n21932 = n21929 ^ n21847 ;
  assign n22024 = n21925 & n21932 ;
  assign n21991 = n21924 ^ n21923 ;
  assign n22006 = n21932 & n21991 ;
  assign n22034 = n22024 ^ n22006 ;
  assign n22032 = n21897 & n21924 ;
  assign n22008 = n21929 & n21991 ;
  assign n21926 = n21925 ^ n21923 ;
  assign n21933 = ~n21926 & n21932 ;
  assign n21934 = n21933 ^ n21926 ;
  assign n21930 = ~n21926 & n21929 ;
  assign n21927 = n21897 & ~n21926 ;
  assign n21931 = n21930 ^ n21927 ;
  assign n21935 = n21934 ^ n21931 ;
  assign n22031 = n22008 ^ n21935 ;
  assign n22033 = n22032 ^ n22031 ;
  assign n22035 = n22034 ^ n22033 ;
  assign n22036 = n21936 & ~n22035 ;
  assign n22021 = n21924 & ~n21928 ;
  assign n22020 = n21897 & n21925 ;
  assign n22022 = n22021 ^ n22020 ;
  assign n22041 = n22036 ^ n22022 ;
  assign n21939 = ~n20973 & n21080 ;
  assign n21938 = n20974 & n21071 ;
  assign n21940 = n21939 ^ n21938 ;
  assign n21947 = n21082 ^ n21068 ;
  assign n21948 = n21947 ^ n21946 ;
  assign n21949 = ~n20974 & n21948 ;
  assign n21950 = n21949 ^ n21068 ;
  assign n21967 = n21950 ^ n21097 ;
  assign n21968 = n21967 ^ n21114 ;
  assign n21960 = n21074 ^ n21062 ;
  assign n21958 = n21078 ^ n21073 ;
  assign n21959 = n21958 ^ n21069 ;
  assign n21961 = n21960 ^ n21959 ;
  assign n21962 = n21959 ^ n20974 ;
  assign n21963 = n21962 ^ n21959 ;
  assign n21964 = n21961 & n21963 ;
  assign n21965 = n21964 ^ n21959 ;
  assign n21966 = ~n21127 & n21965 ;
  assign n21969 = n21968 ^ n21966 ;
  assign n21953 = n21950 ^ n21080 ;
  assign n21954 = n21953 ^ n21950 ;
  assign n21955 = ~n20974 & n21954 ;
  assign n21956 = n21955 ^ n21950 ;
  assign n21957 = n20973 & n21956 ;
  assign n21970 = n21969 ^ n21957 ;
  assign n21971 = ~n21945 & ~n21970 ;
  assign n21941 = n21063 & n21105 ;
  assign n21972 = n21971 ^ n21941 ;
  assign n21973 = ~n21940 & n21972 ;
  assign n21980 = n21973 & ~n21979 ;
  assign n21981 = ~n21937 & n21980 ;
  assign n21983 = n20975 & n21086 ;
  assign n21984 = n21981 & n21983 ;
  assign n21982 = n21981 ^ n16263 ;
  assign n21985 = n21984 ^ n21982 ;
  assign n21986 = n21985 ^ x108 ;
  assign n22037 = n21924 & n21929 ;
  assign n21992 = ~n21928 & n21991 ;
  assign n22007 = n22006 ^ n21992 ;
  assign n22009 = n22008 ^ n22007 ;
  assign n22010 = n22009 ^ n21991 ;
  assign n22011 = n22010 ^ n21933 ;
  assign n22038 = n22037 ^ n22011 ;
  assign n22039 = n22038 ^ n22036 ;
  assign n22040 = n21986 & n22039 ;
  assign n22042 = n22041 ^ n22040 ;
  assign n21987 = n21936 & ~n21986 ;
  assign n22002 = n21987 ^ n21986 ;
  assign n22003 = n22002 ^ n21936 ;
  assign n22004 = n22003 ^ n21987 ;
  assign n22028 = n21930 & n21986 ;
  assign n22027 = n22022 ^ n21930 ;
  assign n22029 = n22028 ^ n22027 ;
  assign n22030 = ~n22004 & n22029 ;
  assign n22043 = n22042 ^ n22030 ;
  assign n21990 = n21924 & n21932 ;
  assign n22023 = n22022 ^ n21990 ;
  assign n22025 = n22024 ^ n22023 ;
  assign n22026 = ~n22002 & n22025 ;
  assign n22044 = n22043 ^ n22026 ;
  assign n22045 = n22044 ^ n21992 ;
  assign n22018 = n22006 ^ n21930 ;
  assign n22019 = n22003 & n22018 ;
  assign n22046 = n22045 ^ n22019 ;
  assign n22005 = n21925 & ~n21928 ;
  assign n22012 = n22011 ^ n22005 ;
  assign n22013 = n22011 ^ n21986 ;
  assign n22014 = n22013 ^ n22011 ;
  assign n22015 = n22012 & n22014 ;
  assign n22016 = n22015 ^ n22011 ;
  assign n22017 = ~n22004 & n22016 ;
  assign n22047 = n22046 ^ n22017 ;
  assign n21994 = n21925 & n21929 ;
  assign n21993 = n21992 ^ n21990 ;
  assign n21995 = n21994 ^ n21993 ;
  assign n21996 = n21995 ^ n21992 ;
  assign n21997 = n21992 ^ n21986 ;
  assign n21998 = n21997 ^ n21992 ;
  assign n21999 = n21996 & n21998 ;
  assign n22000 = n21999 ^ n21992 ;
  assign n22001 = n21936 & n22000 ;
  assign n22048 = n22047 ^ n22001 ;
  assign n21988 = n21987 ^ n21936 ;
  assign n21989 = ~n21935 & n21988 ;
  assign n22049 = n22048 ^ n21989 ;
  assign n22054 = n21931 & n21986 ;
  assign n22055 = n22054 ^ n21930 ;
  assign n22056 = n21936 & n22055 ;
  assign n22057 = ~n22049 & ~n22056 ;
  assign n22058 = n22057 ^ n21004 ;
  assign n22059 = n22058 ^ x125 ;
  assign n22291 = n21662 ^ x89 ;
  assign n22166 = ~n20686 & n20841 ;
  assign n22156 = n20833 ^ n20686 ;
  assign n22158 = n20839 ^ n20827 ;
  assign n22159 = ~n20862 & n22158 ;
  assign n22157 = n20846 ^ n20833 ;
  assign n22160 = n22159 ^ n22157 ;
  assign n22161 = n22156 & ~n22160 ;
  assign n22162 = n22161 ^ n20686 ;
  assign n22165 = n20849 & ~n22162 ;
  assign n22167 = n22166 ^ n22165 ;
  assign n22168 = n22167 ^ n20860 ;
  assign n22169 = ~n20888 & n22168 ;
  assign n22163 = n22162 ^ n20860 ;
  assign n22152 = n22151 ^ n20878 ;
  assign n22153 = ~n20880 & n22152 ;
  assign n22154 = n22153 ^ n20878 ;
  assign n22155 = n20862 & n22154 ;
  assign n22164 = n22163 ^ n22155 ;
  assign n22170 = n22169 ^ n22164 ;
  assign n22171 = n20850 ^ n20849 ;
  assign n22172 = n20850 ^ n20686 ;
  assign n22173 = n22172 ^ n20850 ;
  assign n22174 = n22171 & ~n22173 ;
  assign n22175 = n22174 ^ n20850 ;
  assign n22176 = n20862 & n22175 ;
  assign n22177 = ~n22170 & ~n22176 ;
  assign n22185 = n22177 & ~n22184 ;
  assign n22186 = ~n22150 & n22185 ;
  assign n22187 = ~n20912 & n22186 ;
  assign n22188 = n22187 ^ n18433 ;
  assign n22292 = n22188 ^ x96 ;
  assign n22439 = n22291 & n22292 ;
  assign n22440 = n22439 ^ n22291 ;
  assign n22441 = n22440 ^ n22292 ;
  assign n22294 = n21561 ^ x65 ;
  assign n22083 = n19862 & n19898 ;
  assign n22064 = n19912 ^ n19857 ;
  assign n22065 = n22064 ^ n19377 ;
  assign n22066 = ~n19420 & ~n22065 ;
  assign n22067 = n22066 ^ n19377 ;
  assign n22070 = n22064 ^ n19911 ;
  assign n22071 = ~n22067 & ~n22070 ;
  assign n22068 = n19911 ^ n19899 ;
  assign n22072 = n22071 ^ n22068 ;
  assign n22073 = n22072 ^ n19909 ;
  assign n22080 = n22073 ^ n18354 ;
  assign n22075 = n19853 ^ n19419 ;
  assign n22076 = n22075 ^ n19885 ;
  assign n22077 = ~n19377 & ~n22076 ;
  assign n22063 = n19908 ^ n19857 ;
  assign n22074 = n22073 ^ n22063 ;
  assign n22078 = n22077 ^ n22074 ;
  assign n22079 = ~n19898 & n22078 ;
  assign n22081 = n22080 ^ n22079 ;
  assign n22061 = n19888 ^ n19885 ;
  assign n22062 = n19895 & n22061 ;
  assign n22082 = n22081 ^ n22062 ;
  assign n22084 = n22083 ^ n22082 ;
  assign n22060 = n19854 & n19896 ;
  assign n22085 = n22084 ^ n22060 ;
  assign n22086 = n22085 ^ n18354 ;
  assign n22087 = n19860 ^ n19693 ;
  assign n22088 = n21334 & n22087 ;
  assign n22089 = n22088 ^ n19860 ;
  assign n22090 = ~n19419 & n22089 ;
  assign n22091 = ~n22086 & n22090 ;
  assign n22092 = n22091 ^ n22085 ;
  assign n22295 = n22092 ^ x99 ;
  assign n22296 = ~n22294 & n22295 ;
  assign n22377 = n22296 ^ n22294 ;
  assign n22380 = n22377 ^ n22295 ;
  assign n22314 = n21080 ^ n21061 ;
  assign n22315 = ~n20976 & n22314 ;
  assign n22308 = n21065 ^ n21059 ;
  assign n22311 = n22308 ^ n21937 ;
  assign n22304 = n21087 ^ n21069 ;
  assign n22305 = n22304 ^ n21093 ;
  assign n22306 = n22305 ^ n21055 ;
  assign n22307 = n20974 & n22306 ;
  assign n22309 = n22308 ^ n22307 ;
  assign n22310 = ~n21127 & n22309 ;
  assign n22312 = n22311 ^ n22310 ;
  assign n22299 = n21084 ^ n20974 ;
  assign n22300 = n22299 ^ n21084 ;
  assign n22301 = n21085 & ~n22300 ;
  assign n22302 = n22301 ^ n21084 ;
  assign n22303 = ~n20973 & n22302 ;
  assign n22313 = n22312 ^ n22303 ;
  assign n22316 = n22315 ^ n22313 ;
  assign n22317 = n21063 ^ n21060 ;
  assign n22318 = n22317 ^ n21096 ;
  assign n22319 = n22318 ^ n21958 ;
  assign n22320 = ~n20974 & ~n22319 ;
  assign n22321 = n22320 ^ n21060 ;
  assign n22322 = n21127 & n22321 ;
  assign n22323 = ~n22316 & ~n22322 ;
  assign n22324 = ~n21123 & n22323 ;
  assign n22325 = n21944 ^ n21092 ;
  assign n22326 = n21092 ^ n20973 ;
  assign n22327 = n22326 ^ n21092 ;
  assign n22328 = n22325 & n22327 ;
  assign n22329 = n22328 ^ n21092 ;
  assign n22330 = n22324 & ~n22329 ;
  assign n22331 = n22330 ^ n18247 ;
  assign n22332 = n22331 ^ x74 ;
  assign n22340 = n20108 ^ n20019 ;
  assign n22341 = n22340 ^ n20109 ;
  assign n22342 = n22341 ^ n20140 ;
  assign n22343 = n19989 & n22342 ;
  assign n22338 = n20152 ^ n20119 ;
  assign n22339 = n22338 ^ n21173 ;
  assign n22344 = n22343 ^ n22339 ;
  assign n22345 = n22344 ^ n20125 ;
  assign n22346 = n22345 ^ n20154 ;
  assign n22347 = n22346 ^ n22344 ;
  assign n22350 = n19989 & n22347 ;
  assign n22351 = n22350 ^ n22344 ;
  assign n22352 = n19990 & n22351 ;
  assign n22353 = n22352 ^ n22344 ;
  assign n22335 = n20136 ^ n20118 ;
  assign n22336 = n22335 ^ n20121 ;
  assign n22337 = n20185 & n22336 ;
  assign n22354 = n22353 ^ n22337 ;
  assign n22355 = n22354 ^ n20113 ;
  assign n22356 = n22355 ^ n21166 ;
  assign n22357 = n22356 ^ n21543 ;
  assign n22358 = n22357 ^ n18294 ;
  assign n22334 = n20142 & n20188 ;
  assign n22359 = n22358 ^ n22334 ;
  assign n22362 = n22359 ^ n20149 ;
  assign n22360 = n22359 ^ n20113 ;
  assign n22333 = ~n19989 & n20147 ;
  assign n22361 = n22360 ^ n22333 ;
  assign n22363 = n22362 ^ n22361 ;
  assign n22364 = n22363 ^ n22338 ;
  assign n22365 = n22364 ^ n20149 ;
  assign n22366 = n22365 ^ n22363 ;
  assign n22369 = n19990 & ~n22366 ;
  assign n22370 = n22369 ^ n22363 ;
  assign n22371 = n20169 & ~n22370 ;
  assign n22372 = n22371 ^ n22361 ;
  assign n22373 = n22372 ^ x113 ;
  assign n22374 = n22332 & n22373 ;
  assign n22388 = n22374 ^ n22332 ;
  assign n22389 = n22388 ^ n22373 ;
  assign n22444 = n22380 & ~n22389 ;
  assign n22375 = n22374 ^ n22373 ;
  assign n22404 = n22380 ^ n22294 ;
  assign n22405 = n22375 & n22404 ;
  assign n22406 = n22405 ^ n22375 ;
  assign n22402 = n22375 & ~n22377 ;
  assign n22376 = n22296 & n22375 ;
  assign n22403 = n22402 ^ n22376 ;
  assign n22407 = n22406 ^ n22403 ;
  assign n22383 = n22374 ^ n22295 ;
  assign n22384 = n22294 & n22383 ;
  assign n22385 = n22384 ^ n22294 ;
  assign n22381 = n22374 & n22380 ;
  assign n22382 = n22381 ^ n22380 ;
  assign n22386 = n22385 ^ n22382 ;
  assign n22408 = n22407 ^ n22386 ;
  assign n22448 = n22444 ^ n22408 ;
  assign n22449 = n22448 ^ n22385 ;
  assign n22390 = n22296 & ~n22389 ;
  assign n22391 = n22390 ^ n22381 ;
  assign n22437 = n22391 ^ n22386 ;
  assign n22395 = n22373 ^ n22332 ;
  assign n22396 = n22295 ^ n22294 ;
  assign n22399 = ~n22373 & n22396 ;
  assign n22400 = n22399 ^ n22294 ;
  assign n22401 = ~n22395 & n22400 ;
  assign n22438 = n22437 ^ n22401 ;
  assign n22450 = n22449 ^ n22438 ;
  assign n22451 = ~n22441 & n22450 ;
  assign n22393 = ~n22377 & ~n22389 ;
  assign n22447 = n22393 & n22439 ;
  assign n22452 = n22451 ^ n22447 ;
  assign n22445 = n22444 ^ n22405 ;
  assign n22446 = n22440 & n22445 ;
  assign n22453 = n22452 ^ n22446 ;
  assign n22424 = n22373 ^ n22295 ;
  assign n22378 = n22374 & ~n22377 ;
  assign n22414 = n22378 ^ n22377 ;
  assign n22422 = n22414 ^ n22376 ;
  assign n22413 = n22402 ^ n22393 ;
  assign n22415 = n22414 ^ n22413 ;
  assign n22416 = n22415 ^ n22381 ;
  assign n22417 = n22416 ^ n22389 ;
  assign n22410 = n22374 ^ n22296 ;
  assign n22379 = n22378 ^ n22376 ;
  assign n22387 = n22386 ^ n22379 ;
  assign n22392 = n22391 ^ n22387 ;
  assign n22411 = n22410 ^ n22392 ;
  assign n22412 = n22411 ^ n22378 ;
  assign n22418 = n22417 ^ n22412 ;
  assign n22419 = n22291 & ~n22418 ;
  assign n22409 = n22408 ^ n22381 ;
  assign n22420 = n22419 ^ n22409 ;
  assign n22421 = n22292 & n22420 ;
  assign n22423 = n22422 ^ n22421 ;
  assign n22425 = n22424 ^ n22423 ;
  assign n22426 = n22425 ^ n22401 ;
  assign n22427 = ~n22292 & ~n22426 ;
  assign n22428 = n22427 ^ n22423 ;
  assign n22454 = n22453 ^ n22428 ;
  assign n22442 = n22441 ^ n22291 ;
  assign n22443 = n22438 & n22442 ;
  assign n22455 = n22454 ^ n22443 ;
  assign n22456 = n22455 ^ n20240 ;
  assign n22293 = n22292 ^ n22291 ;
  assign n22429 = n22428 ^ n22421 ;
  assign n22394 = n22393 ^ n22392 ;
  assign n22430 = n22429 ^ n22394 ;
  assign n22431 = n22430 ^ n22429 ;
  assign n22432 = n22429 ^ n22291 ;
  assign n22433 = n22432 ^ n22429 ;
  assign n22434 = n22431 & ~n22433 ;
  assign n22435 = n22434 ^ n22429 ;
  assign n22436 = ~n22293 & ~n22435 ;
  assign n22457 = n22456 ^ n22436 ;
  assign n22458 = n22457 ^ x68 ;
  assign n22598 = n22059 & ~n22458 ;
  assign n22599 = ~n22581 & n22598 ;
  assign n22648 = n22599 ^ n22598 ;
  assign n22582 = n22458 & ~n22581 ;
  assign n22616 = n22582 ^ n22458 ;
  assign n22210 = n21412 ^ x121 ;
  assign n22093 = n22092 ^ x112 ;
  assign n22237 = n22210 ^ n22093 ;
  assign n22149 = n21144 ^ x98 ;
  assign n22189 = n22188 ^ x107 ;
  assign n22190 = ~n22149 & n22189 ;
  assign n22191 = n22190 ^ n22189 ;
  assign n22192 = n22191 ^ n22149 ;
  assign n22193 = n22192 ^ n22189 ;
  assign n22108 = n18818 & ~n19278 ;
  assign n22105 = n19312 ^ n18827 ;
  assign n22106 = ~n19281 & ~n22105 ;
  assign n22102 = n19299 ^ n19280 ;
  assign n22103 = n22102 ^ n21920 ;
  assign n22104 = n22103 ^ n19136 ;
  assign n22107 = n22106 ^ n22104 ;
  assign n22109 = n22108 ^ n22107 ;
  assign n22101 = n19279 & n19303 ;
  assign n22110 = n22109 ^ n22101 ;
  assign n22096 = n19309 ^ n19034 ;
  assign n22097 = n22096 ^ n19309 ;
  assign n22098 = n19310 & ~n22097 ;
  assign n22099 = n22098 ^ n19309 ;
  assign n22100 = n19278 & ~n22099 ;
  assign n22111 = n22110 ^ n22100 ;
  assign n22112 = n22111 ^ x81 ;
  assign n22113 = n21652 ^ n21304 ;
  assign n22114 = n22113 ^ n21301 ;
  assign n22138 = n22114 ^ n21323 ;
  assign n22126 = n21190 & ~n21299 ;
  assign n22127 = n22126 ^ n21293 ;
  assign n22139 = n22138 ^ n22127 ;
  assign n22140 = n22139 ^ n21322 ;
  assign n22141 = n22140 ^ n21892 ;
  assign n22142 = n22141 ^ n19109 ;
  assign n22128 = n22127 ^ n21291 ;
  assign n22129 = n22128 ^ n21850 ;
  assign n22130 = n22129 ^ n21290 ;
  assign n22131 = n22130 ^ n21291 ;
  assign n22132 = n22131 ^ n22129 ;
  assign n22135 = ~n21190 & n22132 ;
  assign n22136 = n22135 ^ n22129 ;
  assign n22137 = n21191 & n22136 ;
  assign n22143 = n22142 ^ n22137 ;
  assign n22123 = n21293 ^ n21265 ;
  assign n22124 = n22123 ^ n21304 ;
  assign n22125 = n21286 & ~n22124 ;
  assign n22144 = n22143 ^ n22125 ;
  assign n22115 = n22114 ^ n21324 ;
  assign n22116 = n22115 ^ n21272 ;
  assign n22117 = n22116 ^ n22114 ;
  assign n22118 = n22114 ^ n21191 ;
  assign n22119 = n22118 ^ n22114 ;
  assign n22120 = n22117 & ~n22119 ;
  assign n22121 = n22120 ^ n22114 ;
  assign n22122 = ~n21309 & ~n22121 ;
  assign n22145 = n22144 ^ n22122 ;
  assign n22146 = n22145 ^ x88 ;
  assign n22147 = n22112 & n22146 ;
  assign n22148 = n22147 ^ n22112 ;
  assign n22195 = n22148 ^ n22146 ;
  assign n22203 = ~n22193 & ~n22195 ;
  assign n22201 = n22147 & n22192 ;
  assign n22248 = n22203 ^ n22201 ;
  assign n22208 = n22148 & n22191 ;
  assign n22249 = n22248 ^ n22208 ;
  assign n22196 = n22195 ^ n22112 ;
  assign n22238 = n22190 & n22196 ;
  assign n22239 = n22238 ^ n22203 ;
  assign n22240 = n22239 ^ n22196 ;
  assign n22197 = n22192 & n22196 ;
  assign n22205 = n22201 ^ n22197 ;
  assign n22200 = ~n22193 & n22196 ;
  assign n22202 = n22201 ^ n22200 ;
  assign n22204 = n22203 ^ n22202 ;
  assign n22206 = n22205 ^ n22204 ;
  assign n22241 = n22240 ^ n22206 ;
  assign n22194 = n22148 & ~n22193 ;
  assign n22247 = n22241 ^ n22194 ;
  assign n22250 = n22249 ^ n22247 ;
  assign n22251 = n22093 & n22250 ;
  assign n22252 = n22251 ^ n22208 ;
  assign n22253 = n22237 & n22252 ;
  assign n22242 = n22147 & n22190 ;
  assign n22243 = n22242 ^ n22241 ;
  assign n22244 = ~n22237 & n22243 ;
  assign n22254 = n22253 ^ n22244 ;
  assign n22219 = n22192 & ~n22195 ;
  assign n22234 = n22219 ^ n22192 ;
  assign n22235 = n22234 ^ n22205 ;
  assign n22236 = n22235 ^ n22202 ;
  assign n22245 = ~n22093 & ~n22244 ;
  assign n22246 = n22236 & n22245 ;
  assign n22255 = n22254 ^ n22246 ;
  assign n22216 = n22191 & ~n22195 ;
  assign n22217 = n22216 ^ n22203 ;
  assign n22218 = n22217 ^ n22195 ;
  assign n22220 = n22219 ^ n22218 ;
  assign n22256 = n22255 ^ n22220 ;
  assign n22222 = ~n22093 & ~n22210 ;
  assign n22223 = n22222 ^ n22093 ;
  assign n22221 = n22220 ^ n22210 ;
  assign n22224 = n22223 ^ n22221 ;
  assign n22226 = n22203 ^ n22197 ;
  assign n22225 = n22147 & n22191 ;
  assign n22227 = n22226 ^ n22225 ;
  assign n22228 = n22227 ^ n22223 ;
  assign n22229 = n22223 ^ n22220 ;
  assign n22230 = n22229 ^ n22223 ;
  assign n22231 = n22228 & n22230 ;
  assign n22232 = n22231 ^ n22223 ;
  assign n22233 = n22224 & n22232 ;
  assign n22257 = n22256 ^ n22233 ;
  assign n22198 = n22197 ^ n22194 ;
  assign n22199 = n22198 ^ n22193 ;
  assign n22207 = n22206 ^ n22199 ;
  assign n22209 = n22208 ^ n22207 ;
  assign n22213 = ~n22209 & n22210 ;
  assign n22214 = n22213 ^ n22208 ;
  assign n22215 = ~n22093 & n22214 ;
  assign n22258 = n22257 ^ n22215 ;
  assign n22259 = n22219 ^ n22207 ;
  assign n22260 = n22259 ^ n22238 ;
  assign n22261 = n22238 ^ n22210 ;
  assign n22262 = n22261 ^ n22238 ;
  assign n22263 = ~n22260 & n22262 ;
  assign n22264 = n22263 ^ n22238 ;
  assign n22265 = n22093 & n22264 ;
  assign n22266 = n22258 & ~n22265 ;
  assign n22274 = n22093 & ~n22210 ;
  assign n22275 = n22242 & n22274 ;
  assign n22267 = n22203 ^ n22093 ;
  assign n22268 = n22267 ^ n22203 ;
  assign n22271 = n22217 & n22268 ;
  assign n22272 = n22271 ^ n22203 ;
  assign n22273 = ~n22210 & n22272 ;
  assign n22276 = n22275 ^ n22273 ;
  assign n22283 = n22093 & n22238 ;
  assign n22277 = n22148 & n22190 ;
  assign n22278 = n22277 ^ n22216 ;
  assign n22279 = n22278 ^ n22235 ;
  assign n22280 = ~n22093 & n22279 ;
  assign n22281 = n22280 ^ n22235 ;
  assign n22282 = n22281 ^ n22238 ;
  assign n22284 = n22283 ^ n22282 ;
  assign n22285 = ~n22237 & n22284 ;
  assign n22286 = n22285 ^ n22281 ;
  assign n22287 = ~n22276 & ~n22286 ;
  assign n22288 = n22266 & n22287 ;
  assign n22289 = n22288 ^ n21049 ;
  assign n22290 = n22289 ^ x110 ;
  assign n22587 = n22290 & n22581 ;
  assign n22588 = n22458 & n22587 ;
  assign n22617 = n22616 ^ n22588 ;
  assign n22615 = n22587 ^ n22581 ;
  assign n22618 = n22617 ^ n22615 ;
  assign n22626 = n22618 ^ n22458 ;
  assign n22603 = n22290 & n22599 ;
  assign n22604 = n22603 ^ n22599 ;
  assign n22601 = n22598 ^ n22458 ;
  assign n22602 = n22587 & ~n22601 ;
  assign n22605 = n22604 ^ n22602 ;
  assign n22606 = n22605 ^ n22603 ;
  assign n22597 = n22582 ^ n22581 ;
  assign n22600 = n22599 ^ n22597 ;
  assign n22607 = n22606 ^ n22600 ;
  assign n22627 = n22626 ^ n22607 ;
  assign n22649 = n22648 ^ n22627 ;
  assign n22650 = n22649 ^ n22604 ;
  assign n22651 = n22650 ^ n22627 ;
  assign n22644 = n22290 ^ n22059 ;
  assign n22645 = n22644 ^ n22581 ;
  assign n22646 = ~n22458 & ~n22645 ;
  assign n22647 = n22646 ^ n22626 ;
  assign n22652 = n22651 ^ n22647 ;
  assign n22689 = ~n22634 & ~n22652 ;
  assign n22583 = n22290 & n22582 ;
  assign n22584 = n22583 ^ n22582 ;
  assign n22585 = ~n22059 & n22584 ;
  assign n22586 = n22585 ^ n22584 ;
  assign n22635 = n22634 ^ n21526 ;
  assign n22688 = n22586 & n22635 ;
  assign n22690 = n22689 ^ n22688 ;
  assign n22621 = n22059 & n22583 ;
  assign n22676 = n22627 ^ n22621 ;
  assign n22677 = n22627 ^ n21812 ;
  assign n22678 = n22677 ^ n22627 ;
  assign n22679 = n22676 & ~n22678 ;
  assign n22680 = n22679 ^ n22627 ;
  assign n22681 = n21526 & n22680 ;
  assign n22622 = n22621 ^ n22583 ;
  assign n22589 = ~n22059 & n22588 ;
  assign n22623 = n22622 ^ n22589 ;
  assign n22624 = n22623 ^ n22585 ;
  assign n22620 = n22601 ^ n22059 ;
  assign n22625 = n22624 ^ n22620 ;
  assign n22639 = n22625 ^ n22617 ;
  assign n22663 = n22639 ^ n22621 ;
  assign n22660 = n22649 ^ n22618 ;
  assign n22661 = n22660 ^ n22604 ;
  assign n21813 = n21812 ^ n21526 ;
  assign n22653 = n22652 ^ n22600 ;
  assign n22643 = n22625 ^ n22585 ;
  assign n22654 = n22653 ^ n22643 ;
  assign n22655 = n22643 ^ n21526 ;
  assign n22656 = n22655 ^ n22643 ;
  assign n22657 = n22654 & n22656 ;
  assign n22658 = n22657 ^ n22643 ;
  assign n22659 = ~n21813 & n22658 ;
  assign n22662 = n22661 ^ n22659 ;
  assign n22664 = n22663 ^ n22662 ;
  assign n22665 = n22664 ^ n22659 ;
  assign n22666 = ~n21526 & n22665 ;
  assign n22667 = n22666 ^ n22662 ;
  assign n22682 = n22681 ^ n22667 ;
  assign n22668 = n22667 ^ n22659 ;
  assign n22637 = n22589 ^ n22588 ;
  assign n22669 = n22668 ^ n22637 ;
  assign n22670 = n22669 ^ n22668 ;
  assign n22671 = n22668 ^ n21812 ;
  assign n22672 = n22671 ^ n22668 ;
  assign n22673 = n22670 & ~n22672 ;
  assign n22674 = n22673 ^ n22668 ;
  assign n22675 = n21813 & n22674 ;
  assign n22683 = n22682 ^ n22675 ;
  assign n22636 = n22635 ^ n21812 ;
  assign n22640 = n22639 ^ n22586 ;
  assign n22638 = n22637 ^ n22622 ;
  assign n22641 = n22640 ^ n22638 ;
  assign n22642 = n22636 & n22641 ;
  assign n22684 = n22683 ^ n22642 ;
  assign n22628 = n22627 ^ n22625 ;
  assign n22614 = n22603 ^ n22589 ;
  assign n22619 = n22618 ^ n22614 ;
  assign n22629 = n22628 ^ n22619 ;
  assign n22630 = ~n21526 & n22629 ;
  assign n22631 = n22630 ^ n22628 ;
  assign n22632 = n21813 & n22631 ;
  assign n22685 = n22684 ^ n22632 ;
  assign n22686 = n22685 ^ n22600 ;
  assign n22609 = n22600 ^ n21526 ;
  assign n22610 = n22609 ^ n22600 ;
  assign n22611 = n22606 & ~n22610 ;
  assign n22612 = n22611 ^ n22600 ;
  assign n22613 = ~n21813 & ~n22612 ;
  assign n22687 = n22686 ^ n22613 ;
  assign n22691 = n22690 ^ n22687 ;
  assign n22590 = n22589 ^ n22586 ;
  assign n22591 = n22590 ^ n22585 ;
  assign n22592 = n22585 ^ n21526 ;
  assign n22593 = n22592 ^ n22585 ;
  assign n22594 = n22591 & n22593 ;
  assign n22595 = n22594 ^ n22585 ;
  assign n22596 = n21813 & n22595 ;
  assign n22692 = n22691 ^ n22596 ;
  assign n22693 = n22692 ^ n21144 ;
  assign n22985 = n20972 ^ x74 ;
  assign n22941 = n22449 ^ n22402 ;
  assign n22942 = n22440 & n22941 ;
  assign n22938 = n22442 & n22448 ;
  assign n22935 = ~n22405 & n22441 ;
  assign n22936 = n22384 & ~n22935 ;
  assign n22929 = n22412 ^ n22390 ;
  assign n22930 = n22929 ^ n22393 ;
  assign n22931 = n22440 & n22930 ;
  assign n22927 = n22411 & n22442 ;
  assign n22928 = n22927 ^ n22447 ;
  assign n22932 = n22931 ^ n22928 ;
  assign n22922 = n22415 ^ n22292 ;
  assign n22923 = n22922 ^ n22415 ;
  assign n22924 = ~n22416 & ~n22923 ;
  assign n22925 = n22924 ^ n22415 ;
  assign n22926 = n22293 & ~n22925 ;
  assign n22933 = n22932 ^ n22926 ;
  assign n22934 = n22933 ^ n18523 ;
  assign n22937 = n22936 ^ n22934 ;
  assign n22939 = n22938 ^ n22937 ;
  assign n22912 = n22438 ^ n22408 ;
  assign n22914 = n22912 ^ n22411 ;
  assign n22901 = n22403 ^ n22393 ;
  assign n22915 = n22914 ^ n22901 ;
  assign n22916 = n22915 ^ n22424 ;
  assign n22917 = n22916 ^ n22394 ;
  assign n22913 = n22912 ^ n22415 ;
  assign n22918 = n22917 ^ n22913 ;
  assign n22919 = n22439 & ~n22918 ;
  assign n22940 = n22939 ^ n22919 ;
  assign n22943 = n22942 ^ n22940 ;
  assign n22911 = n22379 & n22442 ;
  assign n22944 = n22943 ^ n22911 ;
  assign n22902 = n22414 ^ n22383 ;
  assign n22903 = n22902 ^ n22385 ;
  assign n22904 = n22903 ^ n22901 ;
  assign n22905 = n22904 ^ n22903 ;
  assign n22906 = n22903 ^ n22291 ;
  assign n22907 = n22906 ^ n22903 ;
  assign n22908 = n22905 & ~n22907 ;
  assign n22909 = n22908 ^ n22903 ;
  assign n22910 = ~n22293 & n22909 ;
  assign n22945 = n22944 ^ n22910 ;
  assign n22946 = n22945 ^ x106 ;
  assign n22954 = n22550 ^ n22522 ;
  assign n22955 = n22490 & ~n22954 ;
  assign n22956 = n22955 ^ n22550 ;
  assign n22957 = n22523 & n22956 ;
  assign n22958 = n22957 ^ n22550 ;
  assign n22960 = ~n22459 & ~n22958 ;
  assign n22959 = n22958 ^ n22459 ;
  assign n22961 = n22960 ^ n22959 ;
  assign n22962 = n22961 ^ n22532 ;
  assign n22970 = n22962 ^ n18798 ;
  assign n22947 = n22534 ^ n22532 ;
  assign n22948 = n22947 ^ n22570 ;
  assign n22951 = n22948 ^ n22568 ;
  assign n22963 = n22962 ^ n22951 ;
  assign n22950 = n22560 ^ n22532 ;
  assign n22964 = n22963 ^ n22950 ;
  assign n22967 = ~n22459 & ~n22964 ;
  assign n22968 = n22967 ^ n22963 ;
  assign n22969 = n22460 & ~n22968 ;
  assign n22971 = n22970 ^ n22969 ;
  assign n22949 = ~n22459 & n22948 ;
  assign n22972 = n22971 ^ n22949 ;
  assign n22973 = n22972 ^ x97 ;
  assign n22974 = n22946 & ~n22973 ;
  assign n22995 = n22974 ^ n22946 ;
  assign n22996 = n22995 ^ n22973 ;
  assign n22745 = n20881 ^ n20835 ;
  assign n22746 = n22745 ^ n20903 ;
  assign n22747 = n20862 & ~n22746 ;
  assign n22748 = n22747 ^ n20855 ;
  assign n22749 = ~n20686 & n22748 ;
  assign n22750 = n22749 ^ n20855 ;
  assign n22741 = n22495 ^ n20849 ;
  assign n22742 = ~n20862 & n22741 ;
  assign n22743 = n22742 ^ n20849 ;
  assign n22744 = ~n20888 & n22743 ;
  assign n22751 = n22750 ^ n22744 ;
  assign n22752 = n22751 ^ n20841 ;
  assign n22732 = n22496 ^ n20839 ;
  assign n22731 = n22496 ^ n20881 ;
  assign n22733 = n22732 ^ n22731 ;
  assign n22734 = n22731 ^ n20862 ;
  assign n22735 = n22734 ^ n22731 ;
  assign n22736 = ~n22733 & ~n22735 ;
  assign n22737 = n22736 ^ n22731 ;
  assign n22738 = ~n20888 & ~n22737 ;
  assign n22739 = n22738 ^ n20841 ;
  assign n22740 = ~n20898 & n22739 ;
  assign n22753 = n22752 ^ n22740 ;
  assign n22754 = ~n22176 & ~n22753 ;
  assign n22755 = n22754 ^ n22150 ;
  assign n22756 = ~n20912 & n22755 ;
  assign n22757 = n22756 ^ n17957 ;
  assign n22730 = ~n20686 & ~n20864 ;
  assign n22760 = n22757 ^ n22730 ;
  assign n22761 = n22760 ^ x75 ;
  assign n22762 = n21985 ^ x100 ;
  assign n22763 = n22761 & n22762 ;
  assign n22764 = n22763 ^ n22761 ;
  assign n22765 = n21552 ^ x94 ;
  assign n22767 = n20381 ^ n20354 ;
  assign n22768 = n22767 ^ n17959 ;
  assign n22769 = n22768 ^ x117 ;
  assign n22770 = n22765 & n22769 ;
  assign n22783 = n22770 ^ n22765 ;
  assign n22784 = n22783 ^ n22769 ;
  assign n22791 = n22764 & ~n22784 ;
  assign n22792 = n22791 ^ n22764 ;
  assign n22814 = n22792 ^ n22783 ;
  assign n22804 = n22769 ^ n22761 ;
  assign n22797 = n22765 ^ n22761 ;
  assign n22805 = ~n22761 & ~n22797 ;
  assign n22806 = n22805 ^ n22763 ;
  assign n22807 = ~n22804 & ~n22806 ;
  assign n22815 = n22814 ^ n22807 ;
  assign n22773 = n22764 ^ n22762 ;
  assign n22774 = n22773 ^ n22761 ;
  assign n22776 = n22770 ^ n22769 ;
  assign n22777 = n22774 & n22776 ;
  assign n22851 = n22815 ^ n22777 ;
  assign n22780 = n21922 ^ x77 ;
  assign n22729 = n21590 ^ x68 ;
  assign n22785 = n22784 ^ n22770 ;
  assign n22803 = n22785 ^ n22762 ;
  assign n22808 = n22807 ^ n22803 ;
  assign n22801 = n22763 & n22770 ;
  assign n22778 = n22777 ^ n22774 ;
  assign n22775 = n22765 & n22774 ;
  assign n22779 = n22778 ^ n22775 ;
  assign n22802 = n22801 ^ n22779 ;
  assign n22809 = n22808 ^ n22802 ;
  assign n22799 = ~n22773 & ~n22784 ;
  assign n22798 = n22797 ^ n22762 ;
  assign n22800 = n22799 ^ n22798 ;
  assign n22810 = n22809 ^ n22800 ;
  assign n22771 = n22764 & n22770 ;
  assign n22766 = n22764 & n22765 ;
  assign n22772 = n22771 ^ n22766 ;
  assign n22813 = n22810 ^ n22772 ;
  assign n22816 = n22815 ^ n22813 ;
  assign n22795 = n22770 & n22774 ;
  assign n22796 = n22795 ^ n22775 ;
  assign n22811 = n22810 ^ n22796 ;
  assign n22812 = n22811 ^ n22783 ;
  assign n22817 = n22816 ^ n22812 ;
  assign n22794 = ~n22773 & n22776 ;
  assign n22818 = n22817 ^ n22794 ;
  assign n22793 = n22792 ^ n22766 ;
  assign n22819 = n22818 ^ n22793 ;
  assign n22781 = ~n22729 & n22780 ;
  assign n22782 = n22781 ^ n22780 ;
  assign n22786 = n22762 & ~n22785 ;
  assign n22787 = ~n22782 & n22786 ;
  assign n22788 = ~n22779 & n22787 ;
  assign n22789 = n22788 ^ n22786 ;
  assign n22790 = n22789 ^ n22772 ;
  assign n22820 = n22819 ^ n22790 ;
  assign n22821 = n22820 ^ n22789 ;
  assign n22822 = n22789 ^ n22780 ;
  assign n22823 = n22822 ^ n22789 ;
  assign n22824 = n22821 & ~n22823 ;
  assign n22825 = n22824 ^ n22789 ;
  assign n22826 = ~n22729 & n22825 ;
  assign n22827 = n22826 ^ n22789 ;
  assign n22831 = n22799 ^ n22771 ;
  assign n22829 = n22801 ^ n22791 ;
  assign n22828 = n22796 ^ n22793 ;
  assign n22830 = n22829 ^ n22828 ;
  assign n22832 = n22831 ^ n22830 ;
  assign n22833 = ~n22780 & n22832 ;
  assign n22834 = n22833 ^ n22793 ;
  assign n22835 = n22834 ^ n22808 ;
  assign n22836 = n22835 ^ n22809 ;
  assign n22837 = n22836 ^ n22835 ;
  assign n22840 = ~n22780 & ~n22837 ;
  assign n22841 = n22840 ^ n22835 ;
  assign n22842 = ~n22729 & ~n22841 ;
  assign n22843 = n22842 ^ n22834 ;
  assign n22844 = ~n22827 & ~n22843 ;
  assign n22852 = ~n22780 & n22844 ;
  assign n22853 = n22851 & n22852 ;
  assign n22847 = n22799 ^ n22772 ;
  assign n22848 = n22782 & n22847 ;
  assign n22846 = n22782 & n22794 ;
  assign n22849 = n22848 ^ n22846 ;
  assign n22845 = n22844 ^ n18202 ;
  assign n22850 = n22849 ^ n22845 ;
  assign n22854 = n22853 ^ n22850 ;
  assign n22855 = n22854 ^ x115 ;
  assign n22893 = n22021 ^ n21994 ;
  assign n22894 = n21987 & n22893 ;
  assign n22892 = ~n22002 & n22037 ;
  assign n22895 = n22894 ^ n22892 ;
  assign n22856 = ~n22002 & n22005 ;
  assign n22857 = n22856 ^ n22019 ;
  assign n22885 = n22031 ^ n22011 ;
  assign n22886 = n22885 ^ n22022 ;
  assign n22887 = ~n22002 & ~n22886 ;
  assign n22875 = n22037 ^ n21994 ;
  assign n22873 = n21897 & ~n21898 ;
  assign n22874 = n22873 ^ n22032 ;
  assign n22876 = n22875 ^ n22874 ;
  assign n22877 = n22876 ^ n21987 ;
  assign n22878 = n22003 & ~n22877 ;
  assign n22879 = n22878 ^ n21987 ;
  assign n22864 = n22008 ^ n21933 ;
  assign n22865 = ~n21987 & ~n22864 ;
  assign n22866 = n22865 ^ n22006 ;
  assign n22867 = n21936 & ~n22866 ;
  assign n22881 = n22867 ^ n22003 ;
  assign n22880 = n22867 ^ n22024 ;
  assign n22882 = n22881 ^ n22880 ;
  assign n22883 = n22879 & n22882 ;
  assign n22884 = n22883 ^ n22881 ;
  assign n22888 = n22887 ^ n22884 ;
  assign n22860 = n21992 ^ n21927 ;
  assign n22861 = n22860 ^ n21990 ;
  assign n22862 = n22861 ^ n22031 ;
  assign n22863 = n22862 ^ n21990 ;
  assign n22870 = n22863 & n22867 ;
  assign n22871 = n22870 ^ n21990 ;
  assign n22872 = n21987 & n22871 ;
  assign n22889 = n22888 ^ n22872 ;
  assign n22858 = n22023 ^ n21994 ;
  assign n22859 = n21988 & n22858 ;
  assign n22890 = n22889 ^ n22859 ;
  assign n22891 = ~n22857 & ~n22890 ;
  assign n22896 = n22895 ^ n22891 ;
  assign n22897 = n22896 ^ n21989 ;
  assign n22898 = n22897 ^ n17732 ;
  assign n22899 = n22898 ^ x96 ;
  assign n22900 = n22855 & n22899 ;
  assign n22978 = n22900 ^ n22899 ;
  assign n23000 = n22978 ^ n22855 ;
  assign n23001 = n22996 & ~n23000 ;
  assign n23059 = n22985 & n23001 ;
  assign n23024 = n22974 & ~n23000 ;
  assign n23023 = n22900 & n22974 ;
  assign n23025 = n23024 ^ n23023 ;
  assign n23021 = n22974 & n22978 ;
  assign n23022 = n23021 ^ n22974 ;
  assign n23026 = n23025 ^ n23022 ;
  assign n22722 = n22222 & n22225 ;
  assign n22695 = n22241 ^ n22220 ;
  assign n22719 = n22222 & ~n22695 ;
  assign n22710 = n22277 ^ n22238 ;
  assign n22711 = n22710 ^ n22219 ;
  assign n22712 = n22219 ^ n22093 ;
  assign n22713 = n22712 ^ n22219 ;
  assign n22714 = n22711 & n22713 ;
  assign n22715 = n22714 ^ n22219 ;
  assign n22716 = n22237 & n22715 ;
  assign n22717 = n22716 ^ n22283 ;
  assign n22705 = n22242 ^ n22202 ;
  assign n22706 = n22705 ^ n22247 ;
  assign n22707 = ~n22093 & n22706 ;
  assign n22718 = n22717 ^ n22707 ;
  assign n22720 = n22719 ^ n22718 ;
  assign n22721 = n22720 ^ n22276 ;
  assign n22723 = n22722 ^ n22721 ;
  assign n22704 = n22259 ^ n22235 ;
  assign n22708 = n22707 ^ n22704 ;
  assign n22709 = ~n22237 & ~n22708 ;
  assign n22724 = n22723 ^ n22709 ;
  assign n22696 = n22695 ^ n22200 ;
  assign n22697 = n22696 ^ n22208 ;
  assign n22694 = n22227 ^ n22207 ;
  assign n22698 = n22697 ^ n22694 ;
  assign n22699 = n22694 ^ n22210 ;
  assign n22700 = n22699 ^ n22694 ;
  assign n22701 = n22698 & n22700 ;
  assign n22702 = n22701 ^ n22694 ;
  assign n22703 = n22093 & ~n22702 ;
  assign n22725 = n22724 ^ n22703 ;
  assign n22726 = ~n22286 & ~n22725 ;
  assign n22727 = n22726 ^ n19277 ;
  assign n22728 = n22727 ^ x64 ;
  assign n22991 = n22985 ^ n22728 ;
  assign n22992 = ~n22985 & n22991 ;
  assign n23055 = n23026 ^ n22992 ;
  assign n22980 = n22900 ^ n22855 ;
  assign n23008 = n22980 & n22995 ;
  assign n22993 = n22992 ^ n22728 ;
  assign n22994 = n22993 ^ n22985 ;
  assign n23056 = n23008 ^ n22994 ;
  assign n23057 = n23055 & n23056 ;
  assign n23007 = n22978 & n22995 ;
  assign n23009 = n23008 ^ n23007 ;
  assign n23037 = n22992 ^ n22985 ;
  assign n23051 = n23009 & ~n23037 ;
  assign n23047 = n22993 & n23007 ;
  assign n23010 = n22995 & ~n23000 ;
  assign n23011 = n23010 ^ n22995 ;
  assign n23012 = n23011 ^ n23009 ;
  assign n23045 = n23021 ^ n23012 ;
  assign n23046 = n22992 & n23045 ;
  assign n23048 = n23047 ^ n23046 ;
  assign n22999 = n22978 & n22996 ;
  assign n23002 = n23001 ^ n22999 ;
  assign n22997 = n22900 & n22996 ;
  assign n22998 = n22997 ^ n22996 ;
  assign n23003 = n23002 ^ n22998 ;
  assign n23042 = n22992 & n23003 ;
  assign n23041 = n22991 & n22999 ;
  assign n23043 = n23042 ^ n23041 ;
  assign n22975 = n22974 ^ n22973 ;
  assign n22981 = ~n22975 & n22980 ;
  assign n22979 = ~n22975 & n22978 ;
  assign n22982 = n22981 ^ n22979 ;
  assign n22976 = n22900 & ~n22975 ;
  assign n22977 = n22976 ^ n22975 ;
  assign n22983 = n22982 ^ n22977 ;
  assign n22984 = n22983 ^ n22979 ;
  assign n23038 = ~n22984 & ~n23037 ;
  assign n23027 = n23026 ^ n23010 ;
  assign n23028 = n23027 ^ n23025 ;
  assign n23031 = n23028 ^ n22728 ;
  assign n23032 = n23031 ^ n23028 ;
  assign n23033 = n23024 & n23032 ;
  assign n23034 = n23033 ^ n23028 ;
  assign n23035 = ~n22991 & n23034 ;
  assign n23036 = n23035 ^ n23025 ;
  assign n23039 = n23038 ^ n23036 ;
  assign n23006 = n22997 ^ n22976 ;
  assign n23040 = n23039 ^ n23006 ;
  assign n23044 = n23043 ^ n23040 ;
  assign n23049 = n23048 ^ n23044 ;
  assign n23013 = n23012 ^ n22981 ;
  assign n23016 = n23006 ^ n22728 ;
  assign n23017 = n23016 ^ n23006 ;
  assign n23018 = n23013 & ~n23017 ;
  assign n23019 = n23018 ^ n23006 ;
  assign n23020 = n22991 & n23019 ;
  assign n23050 = n23049 ^ n23020 ;
  assign n23052 = n23051 ^ n23050 ;
  assign n23004 = n22994 & n23003 ;
  assign n22988 = ~n22984 & ~n22985 ;
  assign n22989 = n22988 ^ n22979 ;
  assign n22990 = n22728 & n22989 ;
  assign n23005 = n23004 ^ n22990 ;
  assign n23053 = n23052 ^ n23005 ;
  assign n23054 = n23053 ^ n19346 ;
  assign n23058 = n23057 ^ n23054 ;
  assign n23060 = n23059 ^ n23058 ;
  assign n23079 = n21459 ^ n21456 ;
  assign n23080 = n23079 ^ n21500 ;
  assign n23081 = n21188 & ~n23080 ;
  assign n23076 = ~n21458 & ~n21480 ;
  assign n23069 = n21440 ^ n21413 ;
  assign n23070 = n23069 ^ n21454 ;
  assign n23071 = n23070 ^ n21456 ;
  assign n23072 = ~n21145 & ~n23071 ;
  assign n23073 = n23072 ^ n21485 ;
  assign n23074 = ~n21187 & ~n23073 ;
  assign n23066 = n21188 & n21486 ;
  assign n23065 = n21478 & n21509 ;
  assign n23067 = n23066 ^ n23065 ;
  assign n23064 = n21455 ^ n19842 ;
  assign n23068 = n23067 ^ n23064 ;
  assign n23075 = n23074 ^ n23068 ;
  assign n23077 = n23076 ^ n23075 ;
  assign n23062 = n21486 ^ n21462 ;
  assign n23063 = n21189 & n23062 ;
  assign n23078 = n23077 ^ n23063 ;
  assign n23082 = n23081 ^ n23078 ;
  assign n23061 = n21452 & n21458 ;
  assign n23083 = n23082 ^ n23061 ;
  assign n23112 = n23003 & ~n23037 ;
  assign n23110 = n23024 ^ n23008 ;
  assign n23111 = n22993 & n23110 ;
  assign n23113 = n23112 ^ n23111 ;
  assign n23114 = n23113 ^ n23043 ;
  assign n23109 = n22994 & n23045 ;
  assign n23115 = n23114 ^ n23109 ;
  assign n23116 = n23115 ^ n23027 ;
  assign n23107 = n23046 ^ n23004 ;
  assign n23097 = n22728 & n23002 ;
  assign n23098 = n23097 ^ n23001 ;
  assign n23099 = n23098 ^ n22979 ;
  assign n23100 = n23099 ^ n23098 ;
  assign n23101 = n23098 ^ n22728 ;
  assign n23102 = n23101 ^ n23098 ;
  assign n23103 = n23100 & n23102 ;
  assign n23104 = n23103 ^ n23098 ;
  assign n23105 = n22991 & n23104 ;
  assign n23106 = n23105 ^ n23098 ;
  assign n23108 = n23107 ^ n23106 ;
  assign n23117 = n23116 ^ n23108 ;
  assign n23090 = n23021 ^ n23001 ;
  assign n23091 = n23090 ^ n22981 ;
  assign n23094 = n22985 & n23091 ;
  assign n23095 = n23094 ^ n22981 ;
  assign n23096 = n22728 & n23095 ;
  assign n23118 = n23117 ^ n23096 ;
  assign n23086 = n23025 ^ n22976 ;
  assign n23087 = ~n22728 & n23086 ;
  assign n23085 = n23027 ^ n22983 ;
  assign n23088 = n23087 ^ n23085 ;
  assign n23089 = ~n22991 & ~n23088 ;
  assign n23119 = n23118 ^ n23089 ;
  assign n23120 = n23119 ^ n23051 ;
  assign n23121 = n23120 ^ n21922 ;
  assign n23084 = n22985 & n23006 ;
  assign n23122 = n23121 ^ n23084 ;
  assign n23133 = n22781 ^ n22729 ;
  assign n23134 = n23133 ^ n22780 ;
  assign n23156 = n22817 & n23134 ;
  assign n23125 = n22779 ^ n22766 ;
  assign n23126 = n23125 ^ n22810 ;
  assign n23127 = n23126 ^ n22818 ;
  assign n23128 = ~n22729 & ~n23127 ;
  assign n23124 = n22815 ^ n22771 ;
  assign n23129 = n23128 ^ n23124 ;
  assign n23130 = n22780 & n23129 ;
  assign n23157 = n23156 ^ n23130 ;
  assign n23138 = n22763 & ~n22784 ;
  assign n23135 = n22794 ^ n22771 ;
  assign n23136 = n23135 ^ n22779 ;
  assign n23137 = n23134 & n23136 ;
  assign n23139 = n23138 ^ n23137 ;
  assign n23158 = n23157 ^ n23139 ;
  assign n23148 = n22810 ^ n22795 ;
  assign n23149 = n23148 ^ n22775 ;
  assign n23150 = n23149 ^ n22795 ;
  assign n23151 = n22795 ^ n22780 ;
  assign n23152 = n23151 ^ n22795 ;
  assign n23153 = ~n23150 & n23152 ;
  assign n23154 = n23153 ^ n22795 ;
  assign n23155 = n22729 & n23154 ;
  assign n23159 = n23158 ^ n23155 ;
  assign n23160 = n23159 ^ n22849 ;
  assign n23161 = n23160 ^ n20411 ;
  assign n23141 = n23138 ^ n22780 ;
  assign n23142 = n23141 ^ n23138 ;
  assign n23143 = n23138 ^ n22808 ;
  assign n23144 = n23143 ^ n23138 ;
  assign n23145 = ~n23142 & ~n23144 ;
  assign n23146 = n23145 ^ n23138 ;
  assign n23147 = ~n22729 & n23146 ;
  assign n23162 = n23161 ^ n23147 ;
  assign n23123 = n22780 ^ n22729 ;
  assign n23132 = n22829 & n23123 ;
  assign n23163 = n23162 ^ n23132 ;
  assign n23164 = n23083 ^ x69 ;
  assign n23187 = n21986 & n22032 ;
  assign n23184 = n22858 ^ n21935 ;
  assign n23185 = n22003 & ~n23184 ;
  assign n23166 = n22865 ^ n21992 ;
  assign n23169 = n22011 ^ n21935 ;
  assign n23170 = ~n21988 & n23169 ;
  assign n23171 = ~n23166 & n23170 ;
  assign n23165 = n22020 ^ n21990 ;
  assign n23167 = n23166 ^ n23165 ;
  assign n23172 = n23171 ^ n23167 ;
  assign n23175 = n23172 ^ n22860 ;
  assign n23176 = n23175 ^ n22034 ;
  assign n23177 = n23176 ^ n23172 ;
  assign n23178 = n23172 ^ n21986 ;
  assign n23179 = n23178 ^ n23172 ;
  assign n23180 = n23177 & ~n23179 ;
  assign n23181 = n23180 ^ n23172 ;
  assign n23182 = ~n21936 & ~n23181 ;
  assign n23173 = n22857 ^ n22017 ;
  assign n23174 = n23173 ^ n23172 ;
  assign n23183 = n23182 ^ n23174 ;
  assign n23186 = n23185 ^ n23183 ;
  assign n23188 = n23187 ^ n23186 ;
  assign n23189 = ~n22892 & n23188 ;
  assign n23190 = ~n22894 & n23189 ;
  assign n23191 = ~n22056 & n23190 ;
  assign n23192 = n23191 ^ n20818 ;
  assign n23193 = n23192 ^ x91 ;
  assign n23194 = n23164 & ~n23193 ;
  assign n23195 = n23194 ^ n23193 ;
  assign n23196 = n23195 ^ n23164 ;
  assign n23238 = n21749 ^ n21700 ;
  assign n23239 = ~n21553 & n23238 ;
  assign n23240 = n23239 ^ n21700 ;
  assign n23243 = n23240 ^ n21803 ;
  assign n23244 = n23243 ^ n23240 ;
  assign n23245 = ~n21553 & n23244 ;
  assign n23246 = n23245 ^ n23240 ;
  assign n23247 = n21562 & n23246 ;
  assign n23248 = n23247 ^ n23240 ;
  assign n23255 = n21744 ^ n21729 ;
  assign n23256 = n23255 ^ n21773 ;
  assign n23257 = n21553 & ~n23256 ;
  assign n23258 = n23257 ^ n21773 ;
  assign n23253 = n21748 ^ n21722 ;
  assign n23252 = n21749 ^ n21704 ;
  assign n23254 = n23253 ^ n23252 ;
  assign n23259 = n23258 ^ n23254 ;
  assign n23260 = n23259 ^ n23258 ;
  assign n23261 = n21750 ^ n21718 ;
  assign n23262 = ~n21711 & ~n23261 ;
  assign n23263 = n23260 & n23262 ;
  assign n23264 = n23263 ^ n23259 ;
  assign n23265 = n23264 ^ n23258 ;
  assign n23249 = n21753 ^ n21744 ;
  assign n23250 = n23249 ^ n21724 ;
  assign n23251 = ~n21562 & ~n23250 ;
  assign n23266 = n23265 ^ n23251 ;
  assign n23267 = ~n21553 & n23266 ;
  assign n23268 = n23267 ^ n23264 ;
  assign n23269 = n23268 ^ n23258 ;
  assign n23270 = n21742 ^ n21553 ;
  assign n23271 = n23270 ^ n21742 ;
  assign n23274 = n21802 & n23271 ;
  assign n23275 = n23274 ^ n21742 ;
  assign n23276 = ~n23269 & n23275 ;
  assign n23277 = n23276 ^ n23258 ;
  assign n23278 = ~n21562 & n23277 ;
  assign n23279 = n23278 ^ n23268 ;
  assign n23280 = ~n23248 & ~n23279 ;
  assign n23281 = ~n21720 & n23280 ;
  assign n23282 = ~n21809 & n23281 ;
  assign n23283 = n23282 ^ n21226 ;
  assign n23284 = n23283 ^ x67 ;
  assign n23290 = n20933 ^ n20625 ;
  assign n23302 = n23290 ^ n20637 ;
  assign n23303 = n23302 ^ n20922 ;
  assign n23296 = n20385 ^ n20219 ;
  assign n23297 = n20617 & ~n23296 ;
  assign n23295 = n20935 ^ n20641 ;
  assign n23298 = n23297 ^ n23295 ;
  assign n23299 = ~n20915 & ~n23298 ;
  assign n23300 = n23299 ^ n23297 ;
  assign n23301 = n23300 ^ n20652 ;
  assign n23304 = n23303 ^ n23301 ;
  assign n23305 = n23304 ^ n23300 ;
  assign n23308 = ~n20915 & ~n23305 ;
  assign n23309 = n23308 ^ n23300 ;
  assign n23310 = n19347 & n23309 ;
  assign n23311 = n23310 ^ n23300 ;
  assign n23288 = n20635 ^ n20389 ;
  assign n23289 = n23288 ^ n20922 ;
  assign n23291 = n23290 ^ n23289 ;
  assign n23292 = n19347 & ~n23291 ;
  assign n23293 = n23292 ^ n20934 ;
  assign n23294 = n20915 & n23293 ;
  assign n23312 = n23311 ^ n23294 ;
  assign n23313 = ~n20958 & ~n23312 ;
  assign n23286 = n20926 & ~n20944 ;
  assign n23285 = n20637 & n20924 ;
  assign n23287 = n23286 ^ n23285 ;
  assign n23314 = n23313 ^ n23287 ;
  assign n23315 = ~n20969 & n23314 ;
  assign n23316 = n23315 ^ n19418 ;
  assign n23317 = n23316 ^ x92 ;
  assign n23318 = ~n23284 & n23317 ;
  assign n23321 = n23318 ^ n23317 ;
  assign n23325 = n23321 ^ n23284 ;
  assign n23230 = n22722 ^ n20685 ;
  assign n23217 = n22198 & ~n22237 ;
  assign n23200 = n22277 ^ n22203 ;
  assign n23198 = n22242 ^ n22208 ;
  assign n23197 = n22696 ^ n22225 ;
  assign n23199 = n23198 ^ n23197 ;
  assign n23201 = n23200 ^ n23199 ;
  assign n23202 = n22210 & ~n23201 ;
  assign n23203 = n23202 ^ n23198 ;
  assign n23212 = n23203 ^ n22265 ;
  assign n23213 = n23212 ^ n22273 ;
  assign n23214 = n23213 ^ n22717 ;
  assign n23215 = n23214 ^ n22719 ;
  assign n23205 = n23203 ^ n22216 ;
  assign n23204 = n23203 ^ n22236 ;
  assign n23206 = n23205 ^ n23204 ;
  assign n23209 = ~n22210 & n23206 ;
  assign n23210 = n23209 ^ n23205 ;
  assign n23211 = n22093 & n23210 ;
  assign n23216 = n23215 ^ n23211 ;
  assign n23218 = n23217 ^ n23216 ;
  assign n23219 = n22093 & ~n22704 ;
  assign n23220 = n23219 ^ n22235 ;
  assign n23223 = n23220 ^ n23198 ;
  assign n23224 = n23223 ^ n23220 ;
  assign n23225 = n22093 & n23224 ;
  assign n23226 = n23225 ^ n23220 ;
  assign n23227 = ~n22237 & n23226 ;
  assign n23228 = n23227 ^ n23220 ;
  assign n23229 = ~n23218 & ~n23228 ;
  assign n23231 = n23230 ^ n23229 ;
  assign n23232 = n23231 ^ x86 ;
  assign n23233 = n22577 ^ n22575 ;
  assign n23234 = n23233 ^ n21230 ;
  assign n23235 = n23234 ^ x109 ;
  assign n23236 = ~n23232 & n23235 ;
  assign n23237 = n23236 ^ n23235 ;
  assign n23329 = n23237 ^ n23232 ;
  assign n23334 = n23325 & n23329 ;
  assign n23319 = n23318 ^ n23284 ;
  assign n23330 = ~n23319 & n23329 ;
  assign n23326 = n23236 & n23325 ;
  assign n23324 = n23236 & n23318 ;
  assign n23327 = n23326 ^ n23324 ;
  assign n23322 = n23236 & n23321 ;
  assign n23323 = n23322 ^ n23236 ;
  assign n23328 = n23327 ^ n23323 ;
  assign n23331 = n23330 ^ n23328 ;
  assign n23332 = n23331 ^ n23319 ;
  assign n23320 = n23237 & ~n23319 ;
  assign n23333 = n23332 ^ n23320 ;
  assign n23335 = n23334 ^ n23333 ;
  assign n23336 = n23335 ^ n23328 ;
  assign n23337 = n23196 & ~n23336 ;
  assign n23338 = n23194 ^ n23164 ;
  assign n23339 = n23326 ^ n23325 ;
  assign n23340 = n23339 ^ n23334 ;
  assign n23341 = n23338 & n23340 ;
  assign n23348 = n23321 & n23329 ;
  assign n23360 = n23348 ^ n23324 ;
  assign n23353 = n23329 ^ n23235 ;
  assign n23354 = n23318 & ~n23353 ;
  assign n23361 = n23360 ^ n23354 ;
  assign n23350 = n23334 ^ n23330 ;
  assign n23349 = n23348 ^ n23329 ;
  assign n23351 = n23350 ^ n23349 ;
  assign n23362 = n23361 ^ n23351 ;
  assign n23359 = n23348 ^ n23318 ;
  assign n23363 = n23362 ^ n23359 ;
  assign n23364 = n23363 ^ n23360 ;
  assign n23365 = n23364 ^ n23322 ;
  assign n23357 = n23321 & ~n23353 ;
  assign n23358 = n23357 ^ n23351 ;
  assign n23366 = n23365 ^ n23358 ;
  assign n23356 = n23354 ^ n23317 ;
  assign n23367 = n23366 ^ n23356 ;
  assign n23389 = n23367 ^ n23331 ;
  assign n23388 = n23354 ^ n23338 ;
  assign n23390 = n23389 ^ n23388 ;
  assign n23368 = n23363 ^ n23357 ;
  assign n23391 = n23368 ^ n23195 ;
  assign n23392 = n23389 ^ n23368 ;
  assign n23393 = n23392 ^ n23354 ;
  assign n23394 = n23393 ^ n23368 ;
  assign n23395 = n23391 & n23394 ;
  assign n23396 = n23395 ^ n23368 ;
  assign n23397 = n23390 & ~n23396 ;
  assign n23398 = n23397 ^ n23193 ;
  assign n23344 = n23237 & n23325 ;
  assign n23381 = n23344 ^ n23339 ;
  assign n23380 = n23358 ^ n23344 ;
  assign n23382 = n23381 ^ n23380 ;
  assign n23383 = n23381 ^ n23193 ;
  assign n23384 = n23383 ^ n23381 ;
  assign n23385 = ~n23382 & n23384 ;
  assign n23386 = n23385 ^ n23381 ;
  assign n23387 = ~n23164 & n23386 ;
  assign n23399 = n23398 ^ n23387 ;
  assign n23372 = n23348 ^ n23322 ;
  assign n23400 = n23399 ^ n23372 ;
  assign n23369 = n23368 ^ n23367 ;
  assign n23345 = n23344 ^ n23334 ;
  assign n23346 = n23345 ^ n23328 ;
  assign n23342 = n23317 ^ n23284 ;
  assign n23343 = n23342 ^ n23232 ;
  assign n23347 = n23346 ^ n23343 ;
  assign n23352 = n23351 ^ n23347 ;
  assign n23355 = n23354 ^ n23352 ;
  assign n23370 = n23369 ^ n23355 ;
  assign n23371 = n23370 ^ n23343 ;
  assign n23373 = n23372 ^ n23371 ;
  assign n23374 = n23373 ^ n23372 ;
  assign n23375 = n23372 ^ n23193 ;
  assign n23376 = n23375 ^ n23372 ;
  assign n23377 = ~n23374 & ~n23376 ;
  assign n23378 = n23377 ^ n23372 ;
  assign n23379 = n23164 & n23378 ;
  assign n23401 = n23400 ^ n23379 ;
  assign n23402 = ~n23341 & ~n23401 ;
  assign n23403 = ~n23337 & n23402 ;
  assign n23404 = n23403 ^ n21662 ;
  assign n23430 = n23135 ^ n22805 ;
  assign n23406 = n22816 ^ n22795 ;
  assign n23431 = n23430 ^ n23406 ;
  assign n23432 = ~n23133 & n23431 ;
  assign n23417 = n22781 ^ n22777 ;
  assign n23418 = n23134 ^ n22779 ;
  assign n23421 = ~n22781 & ~n23418 ;
  assign n23422 = n23421 ^ n22779 ;
  assign n23423 = n23417 & n23422 ;
  assign n23424 = n23423 ^ n22777 ;
  assign n23425 = n23424 ^ n23137 ;
  assign n23426 = n23425 ^ n23406 ;
  assign n23427 = n23426 ^ n20018 ;
  assign n23408 = n22785 ^ n22761 ;
  assign n23409 = n23408 ^ n22762 ;
  assign n23407 = n23406 ^ n22766 ;
  assign n23410 = n23409 ^ n23407 ;
  assign n23411 = n23410 ^ n23406 ;
  assign n23412 = n23406 ^ n22780 ;
  assign n23413 = n23412 ^ n23406 ;
  assign n23414 = ~n23411 & n23413 ;
  assign n23415 = n23414 ^ n23406 ;
  assign n23416 = ~n23123 & ~n23415 ;
  assign n23428 = n23427 ^ n23416 ;
  assign n23405 = n22781 & n22831 ;
  assign n23429 = n23428 ^ n23405 ;
  assign n23433 = n23432 ^ n23429 ;
  assign n23435 = n23196 & n23320 ;
  assign n23448 = n23345 ^ n23339 ;
  assign n23449 = ~n23193 & n23448 ;
  assign n23453 = n23449 ^ n23193 ;
  assign n23447 = n23344 ^ n23335 ;
  assign n23450 = n23449 ^ n23447 ;
  assign n23445 = n23334 ^ n23327 ;
  assign n23446 = n23193 & ~n23445 ;
  assign n23451 = n23450 ^ n23446 ;
  assign n23452 = ~n23164 & ~n23451 ;
  assign n23454 = n23453 ^ n23452 ;
  assign n23439 = n23346 ^ n23195 ;
  assign n23442 = n23354 & n23439 ;
  assign n23443 = n23442 ^ n23346 ;
  assign n23444 = n23388 & ~n23443 ;
  assign n23455 = n23454 ^ n23444 ;
  assign n23456 = n23455 ^ n23358 ;
  assign n23438 = n23194 & n23320 ;
  assign n23457 = n23456 ^ n23438 ;
  assign n23436 = n23193 ^ n23164 ;
  assign n23437 = n23366 & ~n23436 ;
  assign n23458 = n23457 ^ n23437 ;
  assign n23459 = ~n23435 & ~n23458 ;
  assign n23434 = n23194 & n23389 ;
  assign n23460 = n23459 ^ n23434 ;
  assign n23461 = n23367 ^ n23326 ;
  assign n23462 = n23326 ^ n23193 ;
  assign n23463 = n23462 ^ n23326 ;
  assign n23464 = n23461 & n23463 ;
  assign n23465 = n23464 ^ n23326 ;
  assign n23466 = n23436 & n23465 ;
  assign n23467 = n23460 & ~n23466 ;
  assign n23468 = n23467 ^ n22145 ;
  assign n23502 = n21803 ^ n21727 ;
  assign n23503 = n21711 & n23502 ;
  assign n23485 = n21745 ^ n21743 ;
  assign n23486 = n23485 ^ n21749 ;
  assign n23487 = n23486 ^ n21753 ;
  assign n23488 = n21553 & ~n23487 ;
  assign n23489 = n23488 ^ n21743 ;
  assign n23499 = n23489 ^ n20269 ;
  assign n23500 = n23499 ^ n21738 ;
  assign n23483 = n21562 ^ n21553 ;
  assign n23490 = n21772 ^ n21718 ;
  assign n23491 = n23490 ^ n21704 ;
  assign n23492 = n23491 ^ n23489 ;
  assign n23484 = n21752 ^ n21743 ;
  assign n23493 = n23492 ^ n23484 ;
  assign n23494 = n23492 ^ n21553 ;
  assign n23495 = n23494 ^ n23492 ;
  assign n23496 = n23493 & ~n23495 ;
  assign n23497 = n23496 ^ n23492 ;
  assign n23498 = ~n23483 & ~n23497 ;
  assign n23501 = n23500 ^ n23498 ;
  assign n23504 = n23503 ^ n23501 ;
  assign n23475 = n21744 ^ n21742 ;
  assign n23476 = n23475 ^ n21726 ;
  assign n23477 = n23476 ^ n21744 ;
  assign n23478 = n21744 ^ n21553 ;
  assign n23479 = n23478 ^ n21744 ;
  assign n23480 = n23477 & n23479 ;
  assign n23481 = n23480 ^ n21744 ;
  assign n23482 = ~n21562 & ~n23481 ;
  assign n23505 = n23504 ^ n23482 ;
  assign n23469 = n21751 ^ n21740 ;
  assign n23470 = n21740 ^ n21562 ;
  assign n23471 = n23470 ^ n21740 ;
  assign n23472 = n23469 & n23471 ;
  assign n23473 = n23472 ^ n21740 ;
  assign n23474 = ~n21553 & n23473 ;
  assign n23506 = n23505 ^ n23474 ;
  assign n23524 = n23192 ^ x85 ;
  assign n23544 = n22917 ^ n22407 ;
  assign n23539 = n22403 ^ n22386 ;
  assign n23538 = n22415 ^ n22390 ;
  assign n23540 = n23539 ^ n23538 ;
  assign n23541 = ~n22292 & ~n23540 ;
  assign n23525 = n22917 ^ n22903 ;
  assign n23534 = n23525 ^ n22402 ;
  assign n23526 = n22412 ^ n22403 ;
  assign n23527 = n23526 ^ n23525 ;
  assign n23528 = n23527 ^ n23526 ;
  assign n23529 = n23526 ^ n22292 ;
  assign n23530 = n23529 ^ n23526 ;
  assign n23531 = n23528 & n23530 ;
  assign n23532 = n23531 ^ n23526 ;
  assign n23533 = ~n22291 & n23532 ;
  assign n23535 = n22292 & n23533 ;
  assign n23536 = ~n23534 & n23535 ;
  assign n23537 = n23536 ^ n23533 ;
  assign n23542 = n23541 ^ n23537 ;
  assign n23543 = n23542 ^ n23536 ;
  assign n23545 = n23544 ^ n23543 ;
  assign n23546 = n23545 ^ n23533 ;
  assign n23547 = ~n22293 & n23546 ;
  assign n23548 = n23547 ^ n23542 ;
  assign n23557 = n23548 ^ n22453 ;
  assign n23549 = n22292 & ~n23548 ;
  assign n23550 = n22445 ^ n22386 ;
  assign n23551 = n23550 ^ n22392 ;
  assign n23552 = n22392 ^ n22291 ;
  assign n23553 = n23552 ^ n22392 ;
  assign n23554 = n23551 & ~n23553 ;
  assign n23555 = n23554 ^ n22392 ;
  assign n23556 = n23549 & n23555 ;
  assign n23558 = n23557 ^ n23556 ;
  assign n23559 = ~n22443 & ~n23558 ;
  assign n23560 = ~n22926 & n23559 ;
  assign n23561 = n23560 ^ n20764 ;
  assign n23562 = n23561 ^ x70 ;
  assign n23563 = n23524 & ~n23562 ;
  assign n23564 = n23563 ^ n23524 ;
  assign n23566 = n23163 ^ x126 ;
  assign n23580 = n21509 ^ n21187 ;
  assign n23581 = n21456 ^ n21454 ;
  assign n23582 = ~n23580 & n23581 ;
  assign n23583 = n23582 ^ n21457 ;
  assign n23573 = n23062 ^ n21478 ;
  assign n23574 = n21145 & n23573 ;
  assign n23575 = n23574 ^ n21478 ;
  assign n23584 = n23583 ^ n23575 ;
  assign n23579 = n21188 & n21452 ;
  assign n23585 = n23584 ^ n23579 ;
  assign n23576 = n23575 ^ n21466 ;
  assign n23570 = n21488 ^ n21462 ;
  assign n23571 = n23570 ^ n21459 ;
  assign n23572 = ~n21145 & ~n23571 ;
  assign n23577 = n23576 ^ n23572 ;
  assign n23578 = ~n21458 & ~n23577 ;
  assign n23586 = n23585 ^ n23578 ;
  assign n23568 = n21459 ^ n21440 ;
  assign n23569 = n21188 & ~n23568 ;
  assign n23587 = n23586 ^ n23569 ;
  assign n23567 = n21189 & ~n21501 ;
  assign n23588 = n23587 ^ n23567 ;
  assign n23589 = n21454 ^ n21443 ;
  assign n23590 = n23589 ^ n21516 ;
  assign n23591 = n21516 ^ n21145 ;
  assign n23592 = n23591 ^ n21516 ;
  assign n23593 = n23590 & n23592 ;
  assign n23594 = n23593 ^ n21516 ;
  assign n23595 = ~n21187 & n23594 ;
  assign n23596 = ~n23588 & ~n23595 ;
  assign n23597 = ~n23065 & n23596 ;
  assign n23598 = n23597 ^ n20728 ;
  assign n23599 = n23598 ^ x84 ;
  assign n23600 = ~n23566 & n23599 ;
  assign n23606 = n23564 & n23600 ;
  assign n23601 = n23600 ^ n23566 ;
  assign n23604 = n23601 ^ n23599 ;
  assign n23669 = n23606 ^ n23604 ;
  assign n23507 = n22960 ^ n22532 ;
  assign n23509 = n23507 ^ n22568 ;
  assign n23508 = n23507 ^ n22560 ;
  assign n23510 = n23509 ^ n23508 ;
  assign n23513 = n22459 & ~n23510 ;
  assign n23514 = n23513 ^ n23509 ;
  assign n23515 = n22460 & ~n23514 ;
  assign n23516 = n23515 ^ n23507 ;
  assign n23517 = ~n22948 & ~n23516 ;
  assign n23518 = n23517 ^ n20497 ;
  assign n23519 = n23518 ^ x102 ;
  assign n23520 = n23231 ^ x116 ;
  assign n23521 = n23519 & ~n23520 ;
  assign n23674 = ~n23521 & n23562 ;
  assign n23522 = n23521 ^ n23520 ;
  assign n23523 = n23522 ^ n23519 ;
  assign n23675 = n23674 ^ n23523 ;
  assign n23676 = n23524 & n23675 ;
  assign n23677 = n23669 & ~n23676 ;
  assign n23641 = n23523 ^ n23520 ;
  assign n23609 = n23563 ^ n23562 ;
  assign n23610 = n23600 & ~n23609 ;
  assign n23605 = n23564 & n23604 ;
  assign n23607 = n23606 ^ n23605 ;
  assign n23602 = n23564 & ~n23601 ;
  assign n23603 = n23602 ^ n23564 ;
  assign n23608 = n23607 ^ n23603 ;
  assign n23611 = n23610 ^ n23608 ;
  assign n23657 = n23611 ^ n23606 ;
  assign n23624 = n23563 & n23604 ;
  assign n23619 = n23563 & n23600 ;
  assign n23625 = n23624 ^ n23619 ;
  assign n23658 = n23657 ^ n23625 ;
  assign n23565 = n23564 ^ n23562 ;
  assign n23616 = n23565 & n23599 ;
  assign n23659 = n23658 ^ n23616 ;
  assign n23655 = n23624 ^ n23600 ;
  assign n23656 = n23655 ^ n23608 ;
  assign n23660 = n23659 ^ n23656 ;
  assign n23661 = n23660 ^ n23565 ;
  assign n23614 = n23565 & n23604 ;
  assign n23615 = n23614 ^ n23565 ;
  assign n23617 = n23616 ^ n23615 ;
  assign n23662 = n23661 ^ n23617 ;
  assign n23663 = n23641 & n23662 ;
  assign n23621 = n23604 ^ n23566 ;
  assign n23622 = n23563 & n23621 ;
  assign n23623 = n23622 ^ n23563 ;
  assign n23626 = n23625 ^ n23623 ;
  assign n23652 = ~n23522 & n23626 ;
  assign n23651 = n23622 & n23641 ;
  assign n23653 = n23652 ^ n23651 ;
  assign n23646 = n23604 & ~n23609 ;
  assign n23645 = ~n23601 & ~n23609 ;
  assign n23647 = n23646 ^ n23645 ;
  assign n23642 = n23610 ^ n23609 ;
  assign n23643 = n23642 ^ n23616 ;
  assign n23644 = ~n23641 & ~n23643 ;
  assign n23648 = n23647 ^ n23644 ;
  assign n23633 = n23625 ^ n23519 ;
  assign n23634 = n23633 ^ n23625 ;
  assign n23635 = n23625 ^ n23602 ;
  assign n23636 = n23635 ^ n23625 ;
  assign n23637 = ~n23634 & n23636 ;
  assign n23638 = n23637 ^ n23625 ;
  assign n23639 = n23520 & n23638 ;
  assign n23640 = n23639 ^ n23625 ;
  assign n23649 = n23648 ^ n23640 ;
  assign n23620 = n23619 ^ n23608 ;
  assign n23627 = n23626 ^ n23620 ;
  assign n23628 = n23626 ^ n23520 ;
  assign n23629 = n23628 ^ n23626 ;
  assign n23630 = n23627 & n23629 ;
  assign n23631 = n23630 ^ n23626 ;
  assign n23632 = n23519 & n23631 ;
  assign n23650 = n23649 ^ n23632 ;
  assign n23654 = n23653 ^ n23650 ;
  assign n23664 = n23663 ^ n23654 ;
  assign n23665 = n23664 ^ n22521 ;
  assign n23666 = n23665 ^ n23604 ;
  assign n23618 = ~n23520 & n23617 ;
  assign n23667 = n23666 ^ n23618 ;
  assign n23612 = n23611 ^ n23565 ;
  assign n23613 = n23523 & n23612 ;
  assign n23668 = n23667 ^ n23613 ;
  assign n23678 = n23677 ^ n23668 ;
  assign n23706 = n22928 ^ n22443 ;
  assign n23692 = ~n22407 & n22935 ;
  assign n23693 = n23692 ^ n22449 ;
  assign n23694 = ~n22442 & ~n23693 ;
  assign n23695 = n23544 ^ n22376 ;
  assign n23696 = n23695 ^ n22381 ;
  assign n23697 = n23694 & ~n23696 ;
  assign n23698 = n23697 ^ n23693 ;
  assign n23707 = n23706 ^ n23698 ;
  assign n23699 = n23698 ^ n22915 ;
  assign n23700 = n23699 ^ n22381 ;
  assign n23701 = n23700 ^ n23550 ;
  assign n23702 = n23701 ^ n23698 ;
  assign n23703 = n22292 & n23702 ;
  assign n23704 = n23703 ^ n23699 ;
  assign n23705 = n22291 & ~n23704 ;
  assign n23708 = n23707 ^ n23705 ;
  assign n23691 = ~n22293 & ~n23538 ;
  assign n23709 = n23708 ^ n23691 ;
  assign n23686 = n22402 ^ n22291 ;
  assign n23687 = n23686 ^ n22402 ;
  assign n23688 = n22413 & ~n23687 ;
  assign n23689 = n23688 ^ n22402 ;
  assign n23690 = n22292 & n23689 ;
  assign n23710 = n23709 ^ n23690 ;
  assign n23679 = n22903 ^ n22292 ;
  assign n23680 = n23679 ^ n22903 ;
  assign n23681 = n22903 ^ n22378 ;
  assign n23682 = n23681 ^ n22903 ;
  assign n23683 = ~n23680 & n23682 ;
  assign n23684 = n23683 ^ n22903 ;
  assign n23685 = ~n22291 & n23684 ;
  assign n23711 = n23710 ^ n23685 ;
  assign n23712 = ~n22926 & n23711 ;
  assign n23713 = n23712 ^ n19688 ;
  assign n23714 = n23163 ^ x81 ;
  assign n23742 = n21732 ^ n20107 ;
  assign n23743 = n23742 ^ n21797 ;
  assign n23738 = n23248 ^ n21770 ;
  assign n23725 = n21745 ^ n21730 ;
  assign n23723 = n21741 ^ n21704 ;
  assign n23715 = n21728 ^ n21724 ;
  assign n23716 = n23715 ^ n23490 ;
  assign n23717 = n23716 ^ n21728 ;
  assign n23718 = n21728 ^ n21562 ;
  assign n23719 = n23718 ^ n21728 ;
  assign n23720 = n23717 & ~n23719 ;
  assign n23721 = n23720 ^ n21728 ;
  assign n23722 = n21553 & n23721 ;
  assign n23724 = n23723 ^ n23722 ;
  assign n23726 = n23725 ^ n23724 ;
  assign n23727 = n23726 ^ n23722 ;
  assign n23728 = n21553 & n23727 ;
  assign n23729 = n23728 ^ n23724 ;
  assign n23739 = n23738 ^ n23729 ;
  assign n23730 = n23729 ^ n23722 ;
  assign n23731 = n23730 ^ n23249 ;
  assign n23732 = n23731 ^ n23730 ;
  assign n23733 = n23730 ^ n21553 ;
  assign n23734 = n23733 ^ n23730 ;
  assign n23735 = ~n23732 & ~n23734 ;
  assign n23736 = n23735 ^ n23730 ;
  assign n23737 = n23483 & n23736 ;
  assign n23740 = n23739 ^ n23737 ;
  assign n23741 = ~n21710 & ~n23740 ;
  assign n23744 = n23743 ^ n23741 ;
  assign n23745 = n23744 ^ x88 ;
  assign n23878 = ~n23714 & n23745 ;
  assign n23747 = n23518 ^ x122 ;
  assign n23764 = n22032 ^ n22005 ;
  assign n23760 = n22005 ^ n21935 ;
  assign n23761 = n23760 ^ n22024 ;
  assign n23762 = n23761 ^ n22021 ;
  assign n23763 = n21986 & ~n23762 ;
  assign n23765 = n23764 ^ n23763 ;
  assign n23766 = n22004 & n23765 ;
  assign n23755 = ~n21847 & ~n21898 ;
  assign n23756 = ~n21986 & n23755 ;
  assign n23750 = n22873 ^ n22037 ;
  assign n23751 = n23750 ^ n23165 ;
  assign n23752 = n21986 & n23751 ;
  assign n23753 = n23752 ^ n22873 ;
  assign n23754 = n23753 ^ n22011 ;
  assign n23757 = n23756 ^ n23754 ;
  assign n23758 = ~n21936 & n23757 ;
  assign n23759 = n23758 ^ n23753 ;
  assign n23767 = n23766 ^ n23759 ;
  assign n23768 = n23767 ^ n21989 ;
  assign n23769 = n23768 ^ n22894 ;
  assign n23748 = n23165 ^ n21994 ;
  assign n23749 = ~n22002 & n23748 ;
  assign n23770 = n23769 ^ n23749 ;
  assign n23771 = ~n22028 & ~n23770 ;
  assign n23772 = n22008 ^ n21986 ;
  assign n23773 = n23772 ^ n21936 ;
  assign n23774 = n23773 ^ n22008 ;
  assign n23775 = n22009 ^ n22008 ;
  assign n23776 = n21936 & n23775 ;
  assign n23777 = n23776 ^ n22008 ;
  assign n23778 = ~n23774 & n23777 ;
  assign n23779 = n23778 ^ n22008 ;
  assign n23780 = n23771 & n23779 ;
  assign n23781 = n23780 ^ n23771 ;
  assign n23782 = ~n22892 & n23781 ;
  assign n23783 = ~n22056 & n23782 ;
  assign n23784 = n23783 ^ n19988 ;
  assign n23785 = n23784 ^ x120 ;
  assign n23786 = n23747 & ~n23785 ;
  assign n23787 = n23786 ^ n23747 ;
  assign n23797 = n23200 ^ n22206 ;
  assign n23798 = n23797 ^ n22239 ;
  assign n23799 = n22239 ^ n22210 ;
  assign n23800 = n23799 ^ n22239 ;
  assign n23801 = n23798 & ~n23800 ;
  assign n23802 = n23801 ^ n22239 ;
  assign n23803 = ~n22093 & n23802 ;
  assign n23795 = n23228 ^ n22247 ;
  assign n23796 = n23795 ^ n22215 ;
  assign n23804 = n23803 ^ n23796 ;
  assign n23805 = n23804 ^ n22722 ;
  assign n23806 = n23805 ^ n22286 ;
  assign n23807 = n23806 ^ n20456 ;
  assign n23793 = n22219 ^ n22204 ;
  assign n23794 = ~n22237 & n23793 ;
  assign n23808 = n23807 ^ n23794 ;
  assign n23788 = n22238 ^ n22198 ;
  assign n23789 = n23788 ^ n23198 ;
  assign n23790 = n22093 & n23789 ;
  assign n23791 = n23790 ^ n22247 ;
  assign n23792 = ~n22210 & n23791 ;
  assign n23809 = n23808 ^ n23792 ;
  assign n23810 = n23809 ^ x105 ;
  assign n23838 = n20970 ^ n20480 ;
  assign n23832 = n20941 ^ n20647 ;
  assign n23833 = n23832 ^ n20643 ;
  assign n23834 = n20926 & n23833 ;
  assign n23811 = n20915 ^ n19347 ;
  assign n23824 = n20923 ^ n20644 ;
  assign n23821 = n20654 ^ n20620 ;
  assign n23822 = n23821 ^ n20650 ;
  assign n23823 = n23822 ^ n20944 ;
  assign n23825 = n23824 ^ n23823 ;
  assign n23826 = n23823 ^ n20915 ;
  assign n23827 = n23826 ^ n23823 ;
  assign n23828 = ~n23825 & ~n23827 ;
  assign n23829 = n23828 ^ n23823 ;
  assign n23830 = ~n23811 & n23829 ;
  assign n23813 = n20932 ^ n20630 ;
  assign n23814 = n23813 ^ n20634 ;
  assign n23815 = n23814 ^ n20630 ;
  assign n23816 = n20915 ^ n20630 ;
  assign n23817 = n23816 ^ n20630 ;
  assign n23818 = n23815 & n23817 ;
  assign n23819 = n23818 ^ n20630 ;
  assign n23820 = ~n19347 & n23819 ;
  assign n23831 = n23830 ^ n23820 ;
  assign n23835 = n23834 ^ n23831 ;
  assign n23812 = ~n23290 & n23811 ;
  assign n23836 = n23835 ^ n23812 ;
  assign n23837 = ~n23285 & ~n23836 ;
  assign n23839 = n23838 ^ n23837 ;
  assign n23840 = n23839 ^ x66 ;
  assign n23841 = ~n23810 & n23840 ;
  assign n23843 = n23841 ^ n23840 ;
  assign n23854 = n23843 ^ n23810 ;
  assign n23855 = n23854 ^ n23840 ;
  assign n23887 = n23787 & ~n23855 ;
  assign n23927 = n23878 & n23887 ;
  assign n23846 = n23787 ^ n23785 ;
  assign n23867 = n23846 ^ n23747 ;
  assign n23871 = n23854 & ~n23867 ;
  assign n23844 = n23786 & n23843 ;
  assign n23842 = n23787 & n23841 ;
  assign n23845 = n23844 ^ n23842 ;
  assign n23919 = n23871 ^ n23845 ;
  assign n23920 = n23745 & n23919 ;
  assign n23879 = n23878 ^ n23714 ;
  assign n23881 = n23844 ^ n23843 ;
  assign n23868 = n23843 & ~n23867 ;
  assign n23866 = n23787 & n23843 ;
  assign n23869 = n23868 ^ n23866 ;
  assign n23882 = n23881 ^ n23869 ;
  assign n23847 = n23841 & n23846 ;
  assign n23883 = n23882 ^ n23847 ;
  assign n23862 = ~n23747 & n23854 ;
  assign n23872 = n23871 ^ n23862 ;
  assign n23880 = n23872 ^ n23846 ;
  assign n23884 = n23883 ^ n23880 ;
  assign n23885 = n23884 ^ n23868 ;
  assign n23886 = n23885 ^ n23872 ;
  assign n23891 = n23878 & n23885 ;
  assign n23892 = n23891 ^ n23882 ;
  assign n23893 = n23892 ^ n23862 ;
  assign n23896 = ~n23886 & n23893 ;
  assign n23897 = n23879 & n23896 ;
  assign n23898 = n23897 ^ n23893 ;
  assign n23889 = n23884 ^ n23855 ;
  assign n23856 = n23786 & ~n23855 ;
  assign n23888 = n23887 ^ n23856 ;
  assign n23890 = n23889 ^ n23888 ;
  assign n23899 = n23898 ^ n23890 ;
  assign n23921 = n23920 ^ n23899 ;
  assign n23924 = n23921 ^ n23882 ;
  assign n23925 = n23714 & ~n23924 ;
  assign n23905 = n23841 & ~n23867 ;
  assign n23857 = n23786 & n23854 ;
  assign n23858 = n23857 ^ n23842 ;
  assign n23913 = n23905 ^ n23858 ;
  assign n23914 = n23878 & n23913 ;
  assign n23908 = n23888 ^ n23745 ;
  assign n23909 = n23908 ^ n23888 ;
  assign n23910 = n23905 & n23909 ;
  assign n23911 = n23910 ^ n23888 ;
  assign n23912 = n23714 & n23911 ;
  assign n23915 = n23914 ^ n23912 ;
  assign n23873 = n23872 ^ n23847 ;
  assign n23863 = n23857 ^ n23854 ;
  assign n23864 = n23863 ^ n23862 ;
  assign n23859 = n23858 ^ n23856 ;
  assign n23860 = n23859 ^ n23786 ;
  assign n23861 = n23860 ^ n23845 ;
  assign n23865 = n23864 ^ n23861 ;
  assign n23870 = n23869 ^ n23865 ;
  assign n23874 = n23873 ^ n23870 ;
  assign n23875 = n23874 ^ n23861 ;
  assign n23876 = n23714 & n23875 ;
  assign n23877 = n23876 ^ n23865 ;
  assign n23901 = n23899 ^ n23745 ;
  assign n23900 = n23899 ^ n23861 ;
  assign n23902 = n23901 ^ n23900 ;
  assign n23903 = ~n23877 & ~n23902 ;
  assign n23904 = n23903 ^ n23901 ;
  assign n23916 = n23915 ^ n23904 ;
  assign n23746 = n23745 ^ n23714 ;
  assign n23848 = n23847 ^ n23845 ;
  assign n23849 = n23847 ^ n23714 ;
  assign n23850 = n23849 ^ n23847 ;
  assign n23851 = n23848 & ~n23850 ;
  assign n23852 = n23851 ^ n23847 ;
  assign n23853 = ~n23746 & n23852 ;
  assign n23917 = n23916 ^ n23853 ;
  assign n23918 = n23917 ^ n21846 ;
  assign n23926 = n23925 ^ n23918 ;
  assign n23928 = n23927 ^ n23926 ;
  assign n23945 = n23882 ^ n23714 ;
  assign n23946 = n23945 ^ n23882 ;
  assign n23949 = n23883 & ~n23946 ;
  assign n23950 = n23949 ^ n23882 ;
  assign n23951 = n23746 & n23950 ;
  assign n23938 = n23884 ^ n23871 ;
  assign n23939 = n23938 ^ n23873 ;
  assign n23940 = ~n23714 & n23939 ;
  assign n23941 = n23940 ^ n23873 ;
  assign n23952 = n23951 ^ n23941 ;
  assign n23937 = n23913 ^ n23885 ;
  assign n23942 = n23941 ^ n23937 ;
  assign n23933 = n23885 ^ n23786 ;
  assign n23934 = n23933 ^ n23890 ;
  assign n23935 = n23934 ^ n23913 ;
  assign n23936 = ~n23714 & ~n23935 ;
  assign n23943 = n23942 ^ n23936 ;
  assign n23944 = ~n23745 & n23943 ;
  assign n23953 = n23952 ^ n23944 ;
  assign n23954 = n23868 ^ n23714 ;
  assign n23955 = n23954 ^ n23868 ;
  assign n23958 = n23869 & ~n23955 ;
  assign n23959 = n23958 ^ n23868 ;
  assign n23960 = ~n23746 & n23959 ;
  assign n23961 = ~n23953 & ~n23960 ;
  assign n23962 = n23873 ^ n23714 ;
  assign n23963 = n23962 ^ n23873 ;
  assign n23964 = n23866 ^ n23861 ;
  assign n23965 = n23964 ^ n23873 ;
  assign n23966 = n23963 & n23965 ;
  assign n23967 = n23966 ^ n23873 ;
  assign n23968 = ~n23746 & n23967 ;
  assign n23969 = n23961 & ~n23968 ;
  assign n23930 = n23864 ^ n23844 ;
  assign n23931 = n23878 & n23930 ;
  assign n23929 = n23915 ^ n21695 ;
  assign n23932 = n23931 ^ n23929 ;
  assign n23970 = n23969 ^ n23932 ;
  assign n23971 = ~n21455 & ~n23582 ;
  assign n24004 = n21189 & n21456 ;
  assign n24001 = ~n21187 & ~n21488 ;
  assign n23983 = n21465 ^ n21187 ;
  assign n23986 = n21145 & ~n21462 ;
  assign n23987 = n23986 ^ n21482 ;
  assign n23990 = n23983 ^ n21465 ;
  assign n23991 = ~n23987 & ~n23990 ;
  assign n23992 = n23991 ^ n21145 ;
  assign n23993 = n23983 & n23992 ;
  assign n23994 = n23993 ^ n21187 ;
  assign n23982 = n21447 & ~n23580 ;
  assign n23995 = n23994 ^ n23982 ;
  assign n23998 = n23995 ^ n23067 ;
  assign n23981 = n21477 ^ n21443 ;
  assign n23996 = ~n21458 & n23995 ;
  assign n23997 = n23981 & n23996 ;
  assign n23999 = n23998 ^ n23997 ;
  assign n23979 = n21461 ^ n21448 ;
  assign n23980 = n21189 & n23979 ;
  assign n24000 = n23999 ^ n23980 ;
  assign n24002 = n24001 ^ n24000 ;
  assign n23974 = n21451 ^ n21187 ;
  assign n23975 = n23974 ^ n21451 ;
  assign n23976 = ~n21476 & n23975 ;
  assign n23977 = n23976 ^ n21451 ;
  assign n23978 = n21458 & n23977 ;
  assign n24003 = n24002 ^ n23978 ;
  assign n24005 = n24004 ^ n24003 ;
  assign n24006 = ~n23579 & n24005 ;
  assign n24007 = n23971 & n24006 ;
  assign n24008 = n24007 ^ n20054 ;
  assign n24030 = n23010 ^ n22976 ;
  assign n24031 = n24030 ^ n23013 ;
  assign n24032 = n22728 & n24031 ;
  assign n24020 = n23023 ^ n23021 ;
  assign n24019 = n22997 ^ n22982 ;
  assign n24021 = n24020 ^ n24019 ;
  assign n24011 = n23026 ^ n23007 ;
  assign n24012 = n24011 ^ n23023 ;
  assign n24018 = n24012 ^ n23012 ;
  assign n24022 = n24021 ^ n24018 ;
  assign n24023 = ~n22728 & n24022 ;
  assign n24024 = n24023 ^ n24018 ;
  assign n24033 = n24032 ^ n24024 ;
  assign n24034 = n22985 & n24033 ;
  assign n24009 = n22992 ^ n22983 ;
  assign n24010 = n24009 ^ n23090 ;
  assign n24013 = n24012 ^ n24010 ;
  assign n24014 = ~n22997 & n24013 ;
  assign n24015 = n24014 ^ n22992 ;
  assign n24017 = n23111 ^ n22994 ;
  assign n24025 = n24024 ^ n24017 ;
  assign n24016 = n23111 ^ n22997 ;
  assign n24026 = n24025 ^ n24016 ;
  assign n24027 = n24026 ^ n24024 ;
  assign n24028 = n24015 & n24027 ;
  assign n24029 = n24028 ^ n24025 ;
  assign n24035 = n24034 ^ n24029 ;
  assign n24036 = n24035 ^ n23042 ;
  assign n24037 = n24036 ^ n23106 ;
  assign n24038 = ~n23051 & ~n24037 ;
  assign n24039 = ~n23005 & n24038 ;
  assign n24040 = n24039 ^ n22111 ;
  assign n24060 = n20641 & n20924 ;
  assign n24053 = n20650 ^ n20620 ;
  assign n24054 = ~n19347 & n24053 ;
  assign n24050 = n20929 ^ n20654 ;
  assign n24044 = n20923 ^ n20643 ;
  assign n24042 = n20941 ^ n20632 ;
  assign n24043 = n24042 ^ n23303 ;
  assign n24045 = n24044 ^ n24043 ;
  assign n24046 = ~n20915 & n24045 ;
  assign n24047 = n24046 ^ n24044 ;
  assign n24051 = n24050 ^ n24047 ;
  assign n24048 = n24047 ^ n23287 ;
  assign n24052 = n24051 ^ n24048 ;
  assign n24055 = n24054 ^ n24052 ;
  assign n24056 = ~n20625 & n24055 ;
  assign n24057 = n24056 ^ n24048 ;
  assign n24058 = n23811 & n24057 ;
  assign n24041 = n20969 ^ n20334 ;
  assign n24049 = n24048 ^ n24041 ;
  assign n24059 = n24058 ^ n24049 ;
  assign n24061 = n24060 ^ n24059 ;
  assign n24088 = n22637 ^ n22585 ;
  assign n24089 = n22633 & n24088 ;
  assign n24073 = n22689 ^ n22635 ;
  assign n24074 = n22652 ^ n22603 ;
  assign n24075 = n24074 ^ n22650 ;
  assign n24076 = n24073 & ~n24075 ;
  assign n24071 = n22652 ^ n22605 ;
  assign n24072 = n22636 & ~n24071 ;
  assign n24077 = n24076 ^ n24072 ;
  assign n24069 = n22660 ^ n22627 ;
  assign n24068 = n22621 ^ n22617 ;
  assign n24070 = n24069 ^ n24068 ;
  assign n24078 = n24077 ^ n24070 ;
  assign n24079 = n24078 ^ n24077 ;
  assign n24080 = n24079 ^ n22646 ;
  assign n24081 = n24080 ^ n24079 ;
  assign n24084 = n21526 & n24081 ;
  assign n24085 = n24084 ^ n24079 ;
  assign n24086 = n21813 & n24085 ;
  assign n24087 = n24086 ^ n24078 ;
  assign n24090 = n24089 ^ n24087 ;
  assign n24062 = n22625 ^ n22589 ;
  assign n24063 = n22589 ^ n21812 ;
  assign n24064 = n24063 ^ n22589 ;
  assign n24065 = n24062 & n24064 ;
  assign n24066 = n24065 ^ n22589 ;
  assign n24067 = ~n21526 & n24066 ;
  assign n24091 = n24090 ^ n24067 ;
  assign n24094 = n22640 ^ n21812 ;
  assign n24095 = n24094 ^ n22640 ;
  assign n24096 = n22641 & n24095 ;
  assign n24097 = n24096 ^ n22640 ;
  assign n24098 = ~n21526 & n24097 ;
  assign n24099 = ~n24091 & ~n24098 ;
  assign n24100 = ~n22596 & n24099 ;
  assign n24101 = n24100 ^ n22488 ;
  assign n24132 = n23409 ^ n22775 ;
  assign n24133 = ~n23133 & ~n24132 ;
  assign n24128 = n22848 ^ n22780 ;
  assign n24118 = n22791 ^ n22772 ;
  assign n24119 = n24118 ^ n22819 ;
  assign n24120 = n22819 ^ n22780 ;
  assign n24121 = ~n23123 & ~n24120 ;
  assign n24122 = n24121 ^ n22780 ;
  assign n24123 = n24119 & ~n24122 ;
  assign n24124 = n24123 ^ n22819 ;
  assign n24125 = n24124 ^ n22771 ;
  assign n24129 = n24128 ^ n24125 ;
  assign n24130 = n24129 ^ n23156 ;
  assign n24110 = n22770 ^ n22761 ;
  assign n24111 = n24110 ^ n22762 ;
  assign n24112 = n24111 ^ n22770 ;
  assign n24115 = ~n22785 & n24112 ;
  assign n24116 = n24115 ^ n22770 ;
  assign n24117 = n22729 & ~n24116 ;
  assign n24126 = n24125 ^ n24117 ;
  assign n24127 = ~n23123 & ~n24126 ;
  assign n24131 = n24130 ^ n24127 ;
  assign n24134 = n24133 ^ n24131 ;
  assign n24109 = n22781 & n22815 ;
  assign n24135 = n24134 ^ n24109 ;
  assign n24102 = n23134 ^ n22796 ;
  assign n24103 = n22793 ^ n22781 ;
  assign n24106 = n23134 & ~n24103 ;
  assign n24107 = n24106 ^ n22781 ;
  assign n24108 = n24102 & n24107 ;
  assign n24136 = n24135 ^ n24108 ;
  assign n24137 = ~n23424 & n24136 ;
  assign n24138 = ~n23155 & n24137 ;
  assign n24139 = n24138 ^ n19648 ;
  assign n24149 = n23369 ^ n23324 ;
  assign n24141 = n23284 ^ n23235 ;
  assign n24142 = n24141 ^ n23232 ;
  assign n24143 = n24142 ^ n23235 ;
  assign n24146 = ~n23342 & n24143 ;
  assign n24147 = n24146 ^ n23235 ;
  assign n24148 = ~n23164 & n24147 ;
  assign n24150 = n24149 ^ n24148 ;
  assign n24151 = ~n23193 & n24150 ;
  assign n24163 = n23362 ^ n23335 ;
  assign n24164 = n23362 ^ n23164 ;
  assign n24165 = n24164 ^ n23362 ;
  assign n24166 = ~n24163 & n24165 ;
  assign n24167 = n24166 ^ n23362 ;
  assign n24168 = ~n23193 & n24167 ;
  assign n24161 = n23338 & n23350 ;
  assign n24152 = n23351 ^ n23193 ;
  assign n24154 = n23354 ^ n23322 ;
  assign n24157 = n24154 ^ n23351 ;
  assign n24153 = n23363 ^ n23327 ;
  assign n24155 = n24154 ^ n24153 ;
  assign n24156 = n23164 & n24155 ;
  assign n24158 = n24157 ^ n24156 ;
  assign n24159 = n24152 & ~n24158 ;
  assign n24160 = n24159 ^ n23193 ;
  assign n24162 = n24161 ^ n24160 ;
  assign n24169 = n24168 ^ n24162 ;
  assign n24170 = ~n23438 & ~n24169 ;
  assign n24171 = ~n23466 & n24170 ;
  assign n24172 = ~n24151 & n24171 ;
  assign n24173 = ~n23435 & n24172 ;
  assign n24174 = ~n23341 & n24173 ;
  assign n24177 = n24174 ^ n21895 ;
  assign n24140 = n23448 ^ n23335 ;
  assign n24175 = n23196 & n24174 ;
  assign n24176 = ~n24140 & n24175 ;
  assign n24178 = n24177 ^ n24176 ;
  assign n24187 = n24019 ^ n23001 ;
  assign n24188 = n24187 ^ n22994 ;
  assign n24190 = ~n23008 & ~n24188 ;
  assign n24191 = n24190 ^ n22994 ;
  assign n24193 = n23087 ^ n22992 ;
  assign n24192 = n23087 ^ n23008 ;
  assign n24194 = n24193 ^ n24192 ;
  assign n24195 = n24191 & n24194 ;
  assign n24196 = n24195 ^ n24193 ;
  assign n24197 = n24196 ^ n23038 ;
  assign n24183 = n23087 ^ n22981 ;
  assign n24180 = n23023 ^ n22997 ;
  assign n24184 = n24183 ^ n24180 ;
  assign n24179 = n24012 ^ n22999 ;
  assign n24181 = n24180 ^ n24179 ;
  assign n24182 = ~n22728 & n24181 ;
  assign n24185 = n24184 ^ n24182 ;
  assign n24186 = ~n22991 & n24185 ;
  assign n24198 = n24197 ^ n24186 ;
  assign n24199 = n24198 ^ n23109 ;
  assign n24200 = n24199 ^ n23048 ;
  assign n24201 = n24200 ^ n23113 ;
  assign n24202 = n24201 ^ n23005 ;
  assign n24203 = n22983 & ~n24202 ;
  assign n24204 = n24203 ^ n21631 ;
  assign n24205 = n23626 & n23641 ;
  assign n24220 = n23647 ^ n23610 ;
  assign n24229 = n24220 ^ n23609 ;
  assign n24230 = n24229 ^ n23602 ;
  assign n24231 = n24230 ^ n23610 ;
  assign n24227 = n24220 ^ n23614 ;
  assign n24214 = n23660 ^ n23645 ;
  assign n24215 = n24214 ^ n23617 ;
  assign n24221 = n24220 ^ n24215 ;
  assign n24223 = n24215 ^ n23519 ;
  assign n24224 = ~n23520 & ~n24223 ;
  assign n24225 = n24224 ^ n23519 ;
  assign n24226 = n24221 & n24225 ;
  assign n24228 = n24227 ^ n24226 ;
  assign n24232 = n24231 ^ n24228 ;
  assign n24233 = n24232 ^ n23608 ;
  assign n24234 = n24233 ^ n24228 ;
  assign n24235 = n24228 ^ n23519 ;
  assign n24236 = n24235 ^ n24228 ;
  assign n24237 = ~n24234 & n24236 ;
  assign n24238 = n24237 ^ n24228 ;
  assign n24239 = ~n23520 & n24238 ;
  assign n24240 = n24239 ^ n24228 ;
  assign n24206 = n23520 ^ n23519 ;
  assign n24219 = n23606 & ~n24206 ;
  assign n24241 = n24240 ^ n24219 ;
  assign n24216 = n24215 ^ n23610 ;
  assign n24217 = ~n23522 & n24216 ;
  assign n24213 = n23621 & n23676 ;
  assign n24218 = n24217 ^ n24213 ;
  assign n24242 = n24241 ^ n24218 ;
  assign n24243 = n24242 ^ n23651 ;
  assign n24244 = n24243 ^ n23640 ;
  assign n24207 = n23662 ^ n23607 ;
  assign n24208 = n23607 ^ n23520 ;
  assign n24209 = n24208 ^ n23607 ;
  assign n24210 = n24207 & ~n24209 ;
  assign n24211 = n24210 ^ n23607 ;
  assign n24212 = n24206 & n24211 ;
  assign n24245 = n24244 ^ n24212 ;
  assign n24246 = ~n24205 & ~n24245 ;
  assign n24247 = n24246 ^ n22188 ;
  assign n24248 = n22945 ^ x113 ;
  assign n24249 = n23784 ^ x104 ;
  assign n24250 = n24248 & ~n24249 ;
  assign n24251 = n24250 ^ n24248 ;
  assign n24252 = n24251 ^ n24249 ;
  assign n24253 = n24252 ^ n24248 ;
  assign n24254 = n23433 ^ x80 ;
  assign n24255 = n20972 ^ x90 ;
  assign n24256 = ~n24254 & ~n24255 ;
  assign n24257 = n24256 ^ n24255 ;
  assign n24263 = n24257 ^ n24254 ;
  assign n24264 = n24263 ^ n24255 ;
  assign n24258 = n23744 ^ x99 ;
  assign n24259 = n24008 ^ x73 ;
  assign n24260 = ~n24258 & ~n24259 ;
  assign n24267 = n24260 ^ n24259 ;
  assign n24278 = ~n24264 & ~n24267 ;
  assign n24268 = n24267 ^ n24258 ;
  assign n24269 = ~n24257 & ~n24268 ;
  assign n24282 = n24278 ^ n24269 ;
  assign n24281 = n24256 & ~n24268 ;
  assign n24283 = n24282 ^ n24281 ;
  assign n24280 = ~n24264 & ~n24268 ;
  assign n24284 = n24283 ^ n24280 ;
  assign n24279 = n24278 ^ n24268 ;
  assign n24285 = n24284 ^ n24279 ;
  assign n24286 = n24285 ^ n24263 ;
  assign n24276 = ~n24263 & ~n24267 ;
  assign n24275 = n24260 & ~n24263 ;
  assign n24277 = n24276 ^ n24275 ;
  assign n24287 = n24286 ^ n24277 ;
  assign n24272 = n24254 & ~n24258 ;
  assign n24265 = n24260 & ~n24264 ;
  assign n24261 = n24260 ^ n24258 ;
  assign n24262 = ~n24257 & ~n24261 ;
  assign n24266 = n24265 ^ n24262 ;
  assign n24273 = n24272 ^ n24266 ;
  assign n24274 = n24273 ^ n24260 ;
  assign n24288 = n24287 ^ n24274 ;
  assign n24289 = n24288 ^ n24275 ;
  assign n24271 = n24265 ^ n24260 ;
  assign n24290 = n24289 ^ n24271 ;
  assign n24291 = n24290 ^ n24265 ;
  assign n24292 = n24291 ^ n24257 ;
  assign n24270 = n24269 ^ n24266 ;
  assign n24293 = n24292 ^ n24270 ;
  assign n24294 = n24293 ^ n24280 ;
  assign n24295 = ~n24253 & ~n24294 ;
  assign n24347 = n24290 ^ n24287 ;
  assign n24354 = n24347 ^ n24288 ;
  assign n24355 = n24252 & n24354 ;
  assign n24332 = n24249 ^ n24248 ;
  assign n24302 = n24293 ^ n24278 ;
  assign n24348 = n24347 ^ n24302 ;
  assign n24349 = n24347 ^ n24249 ;
  assign n24350 = n24349 ^ n24347 ;
  assign n24351 = ~n24348 & n24350 ;
  assign n24352 = n24351 ^ n24347 ;
  assign n24353 = n24332 & n24352 ;
  assign n24356 = n24355 ^ n24353 ;
  assign n24301 = n24276 ^ n24267 ;
  assign n24303 = n24302 ^ n24301 ;
  assign n24304 = n24303 ^ n24285 ;
  assign n24305 = n24304 ^ n24270 ;
  assign n24298 = n24288 ^ n24262 ;
  assign n24297 = ~n24261 & ~n24264 ;
  assign n24299 = n24298 ^ n24297 ;
  assign n24300 = n24299 ^ n24285 ;
  assign n24306 = n24305 ^ n24300 ;
  assign n24296 = n24284 ^ n24254 ;
  assign n24307 = n24306 ^ n24296 ;
  assign n24308 = n24251 & ~n24307 ;
  assign n24318 = ~n24253 & n24298 ;
  assign n24316 = n24275 ^ n24269 ;
  assign n24317 = n24316 ^ n24265 ;
  assign n24319 = n24318 ^ n24317 ;
  assign n24320 = n24319 ^ n24251 ;
  assign n24321 = n24294 ^ n24288 ;
  assign n24322 = n24321 ^ n24253 ;
  assign n24325 = ~n24319 & ~n24322 ;
  assign n24326 = n24325 ^ n24253 ;
  assign n24327 = n24320 & ~n24326 ;
  assign n24328 = n24327 ^ n24251 ;
  assign n24314 = n24297 ^ n24281 ;
  assign n24315 = n24252 & n24314 ;
  assign n24329 = n24328 ^ n24315 ;
  assign n24310 = n24276 ^ n24269 ;
  assign n24311 = n24310 ^ n24280 ;
  assign n24309 = n24307 ^ n24303 ;
  assign n24312 = n24311 ^ n24309 ;
  assign n24313 = n24250 & ~n24312 ;
  assign n24330 = n24329 ^ n24313 ;
  assign n24331 = ~n24308 & ~n24330 ;
  assign n24333 = n24278 ^ n24276 ;
  assign n24334 = n24278 ^ n24249 ;
  assign n24335 = n24334 ^ n24278 ;
  assign n24336 = n24333 & n24335 ;
  assign n24337 = n24336 ^ n24278 ;
  assign n24338 = ~n24332 & n24337 ;
  assign n24339 = n24331 & ~n24338 ;
  assign n24340 = n24297 ^ n24285 ;
  assign n24341 = n24285 ^ n24249 ;
  assign n24342 = n24341 ^ n24285 ;
  assign n24343 = ~n24340 & ~n24342 ;
  assign n24344 = n24343 ^ n24285 ;
  assign n24345 = n24332 & ~n24344 ;
  assign n24346 = n24339 & ~n24345 ;
  assign n24357 = n24356 ^ n24346 ;
  assign n24358 = ~n24295 & n24357 ;
  assign n24359 = n24358 ^ n21186 ;
  assign n24381 = n23522 & ~n23621 ;
  assign n24382 = n24215 & n24381 ;
  assign n24378 = n23646 ^ n23605 ;
  assign n24379 = n24378 ^ n24215 ;
  assign n24369 = n24231 ^ n23646 ;
  assign n24370 = n24369 ^ n23656 ;
  assign n24371 = n23520 & ~n24370 ;
  assign n24372 = n24371 ^ n23658 ;
  assign n24377 = n24372 ^ n23602 ;
  assign n24380 = n24379 ^ n24377 ;
  assign n24383 = n24382 ^ n24380 ;
  assign n24375 = n23622 ^ n23602 ;
  assign n24376 = ~n23520 & n24375 ;
  assign n24384 = n24383 ^ n24376 ;
  assign n24385 = ~n24206 & n24384 ;
  assign n24368 = n23653 ^ n23605 ;
  assign n24373 = n24372 ^ n24368 ;
  assign n24364 = n23625 ^ n23607 ;
  assign n24365 = n24209 & n24364 ;
  assign n24366 = n24365 ^ n23607 ;
  assign n24367 = ~n23519 & n24366 ;
  assign n24374 = n24373 ^ n24367 ;
  assign n24386 = n24385 ^ n24374 ;
  assign n24387 = n24386 ^ n24205 ;
  assign n24388 = n24387 ^ n23663 ;
  assign n24389 = n24388 ^ n20914 ;
  assign n24360 = n24229 ^ n24214 ;
  assign n24361 = n23520 & ~n24360 ;
  assign n24362 = n24361 ^ n24214 ;
  assign n24363 = n23519 & n24362 ;
  assign n24390 = n24389 ^ n24363 ;
  assign n24392 = n23316 ^ x100 ;
  assign n24391 = n22580 ^ x118 ;
  assign n24394 = n23713 ^ x124 ;
  assign n24395 = n24139 ^ x76 ;
  assign n24396 = ~n24394 & n24395 ;
  assign n24397 = n23083 ^ x94 ;
  assign n24398 = n21811 ^ x101 ;
  assign n24399 = n24397 & ~n24398 ;
  assign n24400 = n24399 ^ n24397 ;
  assign n24401 = n24400 ^ n24398 ;
  assign n24413 = n24401 ^ n24397 ;
  assign n24429 = n24396 & ~n24413 ;
  assign n24403 = n24396 ^ n24395 ;
  assign n24414 = n24403 & ~n24413 ;
  assign n24470 = n24429 ^ n24414 ;
  assign n24404 = n24403 ^ n24394 ;
  assign n24426 = n24404 & ~n24413 ;
  assign n24469 = n24426 ^ n24413 ;
  assign n24471 = n24470 ^ n24469 ;
  assign n24450 = n24399 & n24404 ;
  assign n24487 = n24471 ^ n24450 ;
  assign n24488 = n24487 ^ n24429 ;
  assign n24489 = n24488 ^ n24396 ;
  assign n24460 = n24396 & n24400 ;
  assign n24416 = n24394 & n24398 ;
  assign n24465 = n24460 ^ n24416 ;
  assign n24423 = n24401 & n24403 ;
  assign n24461 = n24460 ^ n24423 ;
  assign n24418 = n24396 ^ n24394 ;
  assign n24419 = n24401 & ~n24418 ;
  assign n24405 = n24400 & n24404 ;
  assign n24420 = n24419 ^ n24405 ;
  assign n24402 = n24396 & n24401 ;
  assign n24421 = n24420 ^ n24402 ;
  assign n24417 = n24416 ^ n24401 ;
  assign n24422 = n24421 ^ n24417 ;
  assign n24462 = n24461 ^ n24422 ;
  assign n24463 = n24462 ^ n24405 ;
  assign n24466 = n24465 ^ n24463 ;
  assign n24467 = n24466 ^ n24422 ;
  assign n24485 = n24467 ^ n24460 ;
  assign n24486 = n24485 ^ n24471 ;
  assign n24490 = n24489 ^ n24486 ;
  assign n24491 = n24391 & n24490 ;
  assign n24492 = n24491 ^ n24461 ;
  assign n24493 = ~n24392 & n24492 ;
  assign n24445 = ~n24391 & ~n24392 ;
  assign n24446 = n24445 ^ n24391 ;
  assign n24482 = n24460 ^ n24419 ;
  assign n24483 = ~n24446 & n24482 ;
  assign n24393 = n24392 ^ n24391 ;
  assign n24459 = n24423 ^ n24400 ;
  assign n24464 = n24463 ^ n24459 ;
  assign n24472 = n24471 ^ n24464 ;
  assign n24468 = n24467 ^ n24464 ;
  assign n24473 = n24472 ^ n24468 ;
  assign n24474 = n24472 ^ n24391 ;
  assign n24475 = n24474 ^ n24472 ;
  assign n24476 = ~n24473 & ~n24475 ;
  assign n24477 = n24476 ^ n24472 ;
  assign n24478 = n24393 & ~n24477 ;
  assign n24479 = n24478 ^ n24464 ;
  assign n24480 = n24479 ^ n21590 ;
  assign n24424 = n24423 ^ n24422 ;
  assign n24415 = n24414 ^ n24403 ;
  assign n24425 = n24424 ^ n24415 ;
  assign n24427 = n24426 ^ n24425 ;
  assign n24430 = n24429 ^ n24425 ;
  assign n24428 = n24399 & ~n24418 ;
  assign n24431 = n24430 ^ n24428 ;
  assign n24432 = n24392 & ~n24431 ;
  assign n24433 = n24432 ^ n24431 ;
  assign n24434 = n24433 ^ n24391 ;
  assign n24435 = n24434 ^ n24433 ;
  assign n24438 = n24433 ^ n24414 ;
  assign n24439 = n24438 ^ n24433 ;
  assign n24440 = n24432 & ~n24439 ;
  assign n24441 = n24435 & n24440 ;
  assign n24442 = n24441 ^ n24435 ;
  assign n24443 = n24442 ^ n24434 ;
  assign n24444 = ~n24427 & ~n24443 ;
  assign n24447 = n24446 ^ n24392 ;
  assign n24448 = n24430 & ~n24446 ;
  assign n24449 = n24448 ^ n24414 ;
  assign n24451 = n24450 ^ n24449 ;
  assign n24452 = n24447 & ~n24451 ;
  assign n24453 = n24452 ^ n24391 ;
  assign n24454 = n24452 ^ n24392 ;
  assign n24455 = n24454 ^ n24452 ;
  assign n24456 = n24453 & ~n24455 ;
  assign n24457 = n24456 ^ n24452 ;
  assign n24458 = ~n24444 & ~n24457 ;
  assign n24481 = n24480 ^ n24458 ;
  assign n24484 = n24483 ^ n24481 ;
  assign n24494 = n24493 ^ n24484 ;
  assign n24406 = n24405 ^ n24402 ;
  assign n24407 = n24406 ^ n24405 ;
  assign n24408 = n24405 ^ n24391 ;
  assign n24409 = n24408 ^ n24405 ;
  assign n24410 = n24407 & n24409 ;
  assign n24411 = n24410 ^ n24405 ;
  assign n24412 = ~n24393 & n24411 ;
  assign n24495 = n24494 ^ n24412 ;
  assign n24523 = ~n24447 & n24460 ;
  assign n24524 = n24523 ^ n24419 ;
  assign n24525 = n24524 ^ n24479 ;
  assign n24515 = n24471 ^ n24405 ;
  assign n24516 = n24515 ^ n24486 ;
  assign n24517 = n24516 ^ n24515 ;
  assign n24518 = n24515 ^ n24392 ;
  assign n24519 = n24518 ^ n24515 ;
  assign n24520 = ~n24517 & ~n24519 ;
  assign n24521 = n24520 ^ n24515 ;
  assign n24522 = n24393 & ~n24521 ;
  assign n24526 = n24525 ^ n24522 ;
  assign n24512 = n24448 ^ n24393 ;
  assign n24527 = n24526 ^ n24512 ;
  assign n24509 = n24396 & n24399 ;
  assign n24510 = n24509 ^ n24426 ;
  assign n24508 = n24449 ^ n24405 ;
  assign n24511 = n24510 ^ n24508 ;
  assign n24513 = ~n24445 & ~n24512 ;
  assign n24514 = ~n24511 & n24513 ;
  assign n24528 = n24527 ^ n24514 ;
  assign n24529 = n24528 ^ n24526 ;
  assign n24530 = n24452 ^ n24428 ;
  assign n24531 = ~n24426 & n24530 ;
  assign n24532 = ~n24529 & n24531 ;
  assign n24533 = n24532 ^ n24528 ;
  assign n24507 = n24424 & n24445 ;
  assign n24534 = n24533 ^ n24507 ;
  assign n24499 = n24464 ^ n24402 ;
  assign n24497 = n24431 ^ n24419 ;
  assign n24498 = n24497 ^ n24431 ;
  assign n24500 = n24499 ^ n24498 ;
  assign n24501 = n24500 ^ n24497 ;
  assign n24502 = n24497 ^ n24392 ;
  assign n24503 = n24502 ^ n24497 ;
  assign n24504 = n24501 & n24503 ;
  assign n24505 = n24504 ^ n24497 ;
  assign n24506 = n24393 & n24505 ;
  assign n24535 = n24534 ^ n24506 ;
  assign n24496 = n24423 & ~n24447 ;
  assign n24536 = n24535 ^ n24496 ;
  assign n24537 = n24536 ^ n22092 ;
  assign n24548 = n23368 ^ n23326 ;
  assign n24546 = n23360 ^ n23334 ;
  assign n24549 = n24548 ^ n24546 ;
  assign n24550 = n23193 & n24549 ;
  assign n24539 = n23368 ^ n23366 ;
  assign n24540 = n24539 ^ n23343 ;
  assign n24541 = n23193 & n24540 ;
  assign n24542 = n24541 ^ n23371 ;
  assign n24545 = n24542 ^ n23354 ;
  assign n24547 = n24546 ^ n24545 ;
  assign n24551 = n24550 ^ n24547 ;
  assign n24552 = n23436 & ~n24551 ;
  assign n24538 = n23434 ^ n23337 ;
  assign n24543 = n24542 ^ n24538 ;
  assign n24544 = n24543 ^ n23341 ;
  assign n24553 = n24552 ^ n24544 ;
  assign n24554 = ~n23466 & n24553 ;
  assign n24555 = n24554 ^ n21329 ;
  assign n24596 = n22457 ^ x112 ;
  assign n24556 = n22854 ^ x65 ;
  assign n24560 = n22727 ^ x72 ;
  assign n24558 = n21525 ^ x89 ;
  assign n24598 = n24560 ^ n24558 ;
  assign n24557 = n23506 ^ x98 ;
  assign n24565 = ~n24557 & ~n24560 ;
  assign n24572 = n24565 ^ n24557 ;
  assign n24570 = n24061 ^ x107 ;
  assign n24574 = n24570 ^ n24560 ;
  assign n24575 = n24572 & n24574 ;
  assign n24587 = ~n24558 & n24575 ;
  assign n24609 = n24587 ^ n24558 ;
  assign n24563 = n24557 & ~n24558 ;
  assign n24564 = n24560 & ~n24563 ;
  assign n24566 = n24565 ^ n24564 ;
  assign n24567 = n24566 ^ n24563 ;
  assign n24561 = n24560 ^ n24557 ;
  assign n24562 = n24558 & n24561 ;
  assign n24568 = n24567 ^ n24562 ;
  assign n24583 = n24572 ^ n24568 ;
  assign n24584 = ~n24570 & n24583 ;
  assign n24608 = n24584 ^ n24563 ;
  assign n24610 = n24609 ^ n24608 ;
  assign n24601 = ~n24570 & n24598 ;
  assign n24602 = n24601 ^ n24558 ;
  assign n24603 = n24557 & n24602 ;
  assign n24600 = n24574 ^ n24558 ;
  assign n24604 = n24603 ^ n24600 ;
  assign n24599 = n24570 ^ n24561 ;
  assign n24605 = n24604 ^ n24599 ;
  assign n24606 = n24605 ^ n24561 ;
  assign n24607 = n24606 ^ n24604 ;
  assign n24611 = n24610 ^ n24607 ;
  assign n24612 = n24598 & n24611 ;
  assign n24613 = n24612 ^ n24605 ;
  assign n24614 = ~n24556 & n24613 ;
  assign n24615 = n24614 ^ n24604 ;
  assign n24579 = n24567 ^ n24558 ;
  assign n24588 = n24587 ^ n24579 ;
  assign n24585 = n24584 ^ n24568 ;
  assign n24576 = n24575 ^ n24574 ;
  assign n24586 = n24585 ^ n24576 ;
  assign n24589 = n24588 ^ n24586 ;
  assign n24571 = n24560 & n24570 ;
  assign n24573 = n24572 ^ n24571 ;
  assign n24577 = n24576 ^ n24573 ;
  assign n24578 = n24577 ^ n24575 ;
  assign n24580 = n24579 ^ n24578 ;
  assign n24590 = n24589 ^ n24580 ;
  assign n24591 = n24590 ^ n24579 ;
  assign n24592 = n24591 ^ n24561 ;
  assign n24569 = n24568 ^ n24564 ;
  assign n24581 = n24580 ^ n24569 ;
  assign n24559 = n24558 ^ n24557 ;
  assign n24582 = n24581 ^ n24559 ;
  assign n24593 = n24592 ^ n24582 ;
  assign n24594 = n24556 & n24593 ;
  assign n24595 = n24594 ^ n24592 ;
  assign n24616 = n24615 ^ n24595 ;
  assign n24617 = n24596 & ~n24616 ;
  assign n24618 = n24617 ^ n24615 ;
  assign n24597 = n24596 ^ n24595 ;
  assign n24619 = n24618 ^ n24597 ;
  assign n24620 = n24619 ^ n24615 ;
  assign n24621 = n24620 ^ n20384 ;
  assign n24647 = n24287 ^ n24269 ;
  assign n24648 = n24647 ^ n24288 ;
  assign n24649 = n24648 ^ n24307 ;
  assign n24650 = ~n24248 & ~n24649 ;
  assign n24651 = n24650 ^ n24277 ;
  assign n24652 = n24249 & n24651 ;
  assign n24634 = n24297 ^ n24251 ;
  assign n24635 = n24288 ^ n24253 ;
  assign n24638 = ~n24297 & n24635 ;
  assign n24639 = n24638 ^ n24253 ;
  assign n24640 = n24634 & ~n24639 ;
  assign n24641 = n24640 ^ n24251 ;
  assign n24623 = n24304 ^ n24262 ;
  assign n24642 = n24641 ^ n24623 ;
  assign n24643 = n24642 ^ n24353 ;
  assign n24632 = n24250 & ~n24294 ;
  assign n24633 = n24632 ^ n24308 ;
  assign n24644 = n24643 ^ n24633 ;
  assign n24624 = n24623 ^ n24265 ;
  assign n24625 = n24624 ^ n24283 ;
  assign n24626 = n24625 ^ n24623 ;
  assign n24627 = n24623 ^ n24249 ;
  assign n24628 = n24627 ^ n24623 ;
  assign n24629 = n24626 & ~n24628 ;
  assign n24630 = n24629 ^ n24623 ;
  assign n24631 = n24332 & ~n24630 ;
  assign n24645 = n24644 ^ n24631 ;
  assign n24622 = ~n24253 & n24291 ;
  assign n24646 = n24645 ^ n24622 ;
  assign n24653 = n24652 ^ n24646 ;
  assign n24654 = n24653 ^ n24295 ;
  assign n24655 = n24654 ^ n21552 ;
  assign n24684 = n24074 ^ n22627 ;
  assign n24685 = n22636 & ~n24684 ;
  assign n24666 = n22605 ^ n22585 ;
  assign n24667 = n24666 ^ n22627 ;
  assign n24665 = n22660 ^ n22606 ;
  assign n24668 = n24667 ^ n24665 ;
  assign n24669 = ~n21526 & n24668 ;
  assign n24670 = n24669 ^ n24667 ;
  assign n24678 = n24670 ^ n22690 ;
  assign n24679 = n24678 ^ n22659 ;
  assign n24680 = n24679 ^ n22596 ;
  assign n24681 = n24680 ^ n22331 ;
  assign n24671 = n24670 ^ n22651 ;
  assign n24672 = n24671 ^ n22617 ;
  assign n24673 = n24672 ^ n22623 ;
  assign n24674 = n24673 ^ n24670 ;
  assign n24675 = n21526 & n24674 ;
  assign n24676 = n24675 ^ n24671 ;
  assign n24677 = ~n21813 & n24676 ;
  assign n24682 = n24681 ^ n24677 ;
  assign n24664 = n22635 & n22637 ;
  assign n24683 = n24682 ^ n24664 ;
  assign n24686 = n24685 ^ n24683 ;
  assign n24663 = n21813 & n22621 ;
  assign n24687 = n24686 ^ n24663 ;
  assign n24656 = n22622 ^ n22586 ;
  assign n24657 = n24656 ^ n22639 ;
  assign n24658 = n22639 ^ n21526 ;
  assign n24659 = n24658 ^ n22639 ;
  assign n24660 = n24657 & ~n24659 ;
  assign n24661 = n24660 ^ n22639 ;
  assign n24662 = ~n21812 & n24661 ;
  assign n24688 = n24687 ^ n24662 ;
  assign n24689 = n24471 ^ n24461 ;
  assign n24690 = ~n24392 & ~n24689 ;
  assign n24691 = n24690 ^ n24471 ;
  assign n24692 = n24691 ^ n24392 ;
  assign n24693 = n24692 ^ n24691 ;
  assign n24694 = n24691 ^ n24428 ;
  assign n24695 = n24694 ^ n24691 ;
  assign n24696 = n24693 & n24695 ;
  assign n24697 = n24696 ^ n24691 ;
  assign n24698 = ~n24391 & ~n24697 ;
  assign n24699 = n24698 ^ n24691 ;
  assign n24716 = n24509 ^ n24422 ;
  assign n24714 = n24466 ^ n24420 ;
  assign n24715 = n24445 & n24714 ;
  assign n24717 = n24716 ^ n24715 ;
  assign n24718 = n24717 ^ n24428 ;
  assign n24713 = ~n24447 & n24499 ;
  assign n24719 = n24718 ^ n24713 ;
  assign n24723 = n24719 ^ n24496 ;
  assign n24702 = n24429 ^ n24392 ;
  assign n24703 = n24702 ^ n24429 ;
  assign n24704 = n24470 & n24703 ;
  assign n24705 = n24704 ^ n24429 ;
  assign n24706 = ~n24393 & n24705 ;
  assign n24724 = n24723 ^ n24706 ;
  assign n24712 = n24487 ^ n24427 ;
  assign n24720 = n24719 ^ n24712 ;
  assign n24708 = n24487 ^ n24460 ;
  assign n24709 = n24708 ^ n24421 ;
  assign n24710 = n24709 ^ n24427 ;
  assign n24711 = n24392 & ~n24710 ;
  assign n24721 = n24720 ^ n24711 ;
  assign n24722 = n24393 & ~n24721 ;
  assign n24725 = n24724 ^ n24722 ;
  assign n24707 = ~n24391 & n24426 ;
  assign n24726 = n24725 ^ n24707 ;
  assign n24727 = n24726 ^ n24706 ;
  assign n24728 = n24447 ^ n24391 ;
  assign n24729 = n24420 & ~n24728 ;
  assign n24730 = ~n24727 & n24729 ;
  assign n24731 = n24730 ^ n24726 ;
  assign n24732 = ~n24448 & ~n24731 ;
  assign n24733 = n24699 & n24732 ;
  assign n24734 = n24733 ^ n21377 ;
  assign n24738 = n24463 ^ n24430 ;
  assign n24739 = n24738 ^ n24510 ;
  assign n24740 = ~n24392 & n24739 ;
  assign n24741 = n24740 ^ n24463 ;
  assign n24749 = n24741 ^ n24496 ;
  assign n24745 = n24509 ^ n24414 ;
  assign n24746 = ~n24392 & n24745 ;
  assign n24743 = n24420 & n24445 ;
  assign n24737 = n24523 ^ n24499 ;
  assign n24742 = n24741 ^ n24737 ;
  assign n24744 = n24743 ^ n24742 ;
  assign n24747 = n24746 ^ n24744 ;
  assign n24748 = ~n24393 & n24747 ;
  assign n24750 = n24749 ^ n24748 ;
  assign n24736 = ~n24446 & ~n24488 ;
  assign n24751 = n24750 ^ n24736 ;
  assign n24752 = n24391 & ~n24751 ;
  assign n24753 = n24466 ^ n24392 ;
  assign n24754 = n24753 ^ n24466 ;
  assign n24755 = n24466 ^ n24464 ;
  assign n24756 = n24755 ^ n24466 ;
  assign n24757 = ~n24754 & n24756 ;
  assign n24758 = n24757 ^ n24466 ;
  assign n24759 = n24752 & n24758 ;
  assign n24760 = n24759 ^ n24751 ;
  assign n24761 = n24699 & ~n24760 ;
  assign n24762 = n24761 ^ n19933 ;
  assign n24735 = ~n24393 & n24427 ;
  assign n24765 = n24762 ^ n24735 ;
  assign n24766 = n23624 ^ n23617 ;
  assign n24783 = n24766 ^ n23632 ;
  assign n24784 = n24783 ^ n24362 ;
  assign n24785 = n24784 ^ n24212 ;
  assign n24786 = n24785 ^ n24367 ;
  assign n24776 = n24362 ^ n24216 ;
  assign n24775 = n24369 ^ n24362 ;
  assign n24777 = n24776 ^ n24775 ;
  assign n24780 = ~n23520 & ~n24777 ;
  assign n24781 = n24780 ^ n24776 ;
  assign n24782 = ~n23519 & n24781 ;
  assign n24787 = n24786 ^ n24782 ;
  assign n24767 = n24766 ^ n23620 ;
  assign n24768 = n24767 ^ n23622 ;
  assign n24769 = n24768 ^ n24766 ;
  assign n24770 = n24766 ^ n23520 ;
  assign n24771 = n24770 ^ n24766 ;
  assign n24772 = n24769 & ~n24771 ;
  assign n24773 = n24772 ^ n24766 ;
  assign n24774 = n24206 & n24773 ;
  assign n24788 = n24787 ^ n24774 ;
  assign n24789 = n24788 ^ n24205 ;
  assign n24790 = n24789 ^ n23663 ;
  assign n24791 = n24790 ^ n22760 ;
  assign n24805 = n24355 ^ n24281 ;
  assign n24806 = n24805 ^ n24355 ;
  assign n24807 = n24806 ^ n24265 ;
  assign n24808 = n24807 ^ n24806 ;
  assign n24809 = n24806 ^ n24249 ;
  assign n24810 = n24809 ^ n24806 ;
  assign n24811 = n24808 & n24810 ;
  assign n24812 = n24811 ^ n24806 ;
  assign n24813 = n24332 & n24812 ;
  assign n24814 = n24813 ^ n24805 ;
  assign n24815 = n24814 ^ n24633 ;
  assign n24802 = n24287 ^ n24266 ;
  assign n24803 = n24802 ^ n24303 ;
  assign n24804 = n24251 & n24803 ;
  assign n24816 = n24815 ^ n24804 ;
  assign n24801 = ~n24293 & ~n24332 ;
  assign n24817 = n24816 ^ n24801 ;
  assign n24796 = n24300 ^ n24248 ;
  assign n24797 = n24796 ^ n24300 ;
  assign n24798 = n24306 & n24797 ;
  assign n24799 = n24798 ^ n24300 ;
  assign n24800 = ~n24249 & ~n24799 ;
  assign n24818 = n24817 ^ n24800 ;
  assign n24793 = n24252 & n24311 ;
  assign n24819 = n24818 ^ n24793 ;
  assign n24820 = ~n24338 & ~n24819 ;
  assign n24821 = ~n24345 & n24820 ;
  assign n24822 = n24821 ^ n22372 ;
  assign n24792 = ~n24253 & n24276 ;
  assign n24825 = n24822 ^ n24792 ;
  assign n24835 = n24563 & n24571 ;
  assign n24833 = n24577 ^ n24566 ;
  assign n24832 = n24602 ^ n24586 ;
  assign n24834 = n24833 ^ n24832 ;
  assign n24836 = n24835 ^ n24834 ;
  assign n24826 = n24563 ^ n24558 ;
  assign n24829 = n24574 & n24826 ;
  assign n24830 = n24829 ^ n24563 ;
  assign n24831 = n24585 & ~n24830 ;
  assign n24837 = n24836 ^ n24831 ;
  assign n24838 = ~n24556 & ~n24837 ;
  assign n24839 = n24838 ^ n24836 ;
  assign n24848 = n24839 ^ n21436 ;
  assign n24841 = n24839 ^ n24589 ;
  assign n24840 = n24839 ^ n24580 ;
  assign n24842 = n24841 ^ n24840 ;
  assign n24845 = ~n24556 & ~n24842 ;
  assign n24846 = n24845 ^ n24841 ;
  assign n24847 = n24596 & n24846 ;
  assign n24849 = n24848 ^ n24847 ;
  assign n24859 = n24303 ^ n24249 ;
  assign n24860 = n24332 & n24859 ;
  assign n24861 = n24860 ^ n24249 ;
  assign n24864 = n24303 ^ n24283 ;
  assign n24865 = ~n24861 & n24864 ;
  assign n24862 = n24283 ^ n24276 ;
  assign n24866 = n24865 ^ n24862 ;
  assign n24877 = n24866 ^ n24641 ;
  assign n24871 = n24259 ^ n24254 ;
  assign n24872 = n24255 & n24871 ;
  assign n24869 = n24866 ^ n24284 ;
  assign n24867 = n24259 ^ n24258 ;
  assign n24868 = n24867 ^ n24866 ;
  assign n24870 = n24869 ^ n24868 ;
  assign n24873 = n24872 ^ n24870 ;
  assign n24874 = ~n24249 & ~n24873 ;
  assign n24875 = n24874 ^ n24869 ;
  assign n24876 = n24332 & n24875 ;
  assign n24878 = n24877 ^ n24876 ;
  assign n24857 = n24307 ^ n24289 ;
  assign n24858 = ~n24253 & ~n24857 ;
  assign n24879 = n24878 ^ n24858 ;
  assign n24852 = n24266 ^ n24248 ;
  assign n24853 = n24852 ^ n24266 ;
  assign n24854 = n24273 & ~n24853 ;
  assign n24855 = n24854 ^ n24266 ;
  assign n24856 = n24249 & n24855 ;
  assign n24880 = n24879 ^ n24856 ;
  assign n24881 = ~n24295 & ~n24880 ;
  assign n24882 = n24881 ^ n20218 ;
  assign n24883 = n24618 ^ n22768 ;
  assign n24885 = n24589 ^ n24561 ;
  assign n24886 = n24885 ^ n24613 ;
  assign n24888 = ~n24556 & ~n24596 ;
  assign n24889 = n24886 & n24888 ;
  assign n24884 = n24586 ^ n24580 ;
  assign n24887 = n24886 ^ n24884 ;
  assign n24890 = n24889 ^ n24887 ;
  assign n24891 = n24831 ^ n24588 ;
  assign n24892 = ~n24556 & ~n24891 ;
  assign n24893 = n24892 ^ n24588 ;
  assign n24894 = n24893 ^ n24596 ;
  assign n24895 = n24894 ^ n24556 ;
  assign n24896 = n24895 ^ n24893 ;
  assign n24897 = n24556 & n24836 ;
  assign n24898 = n24897 ^ n24893 ;
  assign n24899 = ~n24896 & n24898 ;
  assign n24900 = n24899 ^ n24893 ;
  assign n24901 = n24890 & n24900 ;
  assign n24902 = n24901 ^ n24890 ;
  assign n24903 = n24586 & n24902 ;
  assign n24904 = n24903 ^ n21561 ;
  assign n24945 = ~n23745 & n23872 ;
  assign n24938 = n23905 ^ n23842 ;
  assign n24939 = n24938 ^ n23938 ;
  assign n24933 = n23857 ^ n23844 ;
  assign n24934 = n24933 ^ n23890 ;
  assign n24935 = n24934 ^ n23887 ;
  assign n24940 = n24939 ^ n24935 ;
  assign n24941 = ~n23745 & ~n24940 ;
  assign n24922 = n23887 ^ n23847 ;
  assign n24923 = n24922 ^ n23864 ;
  assign n24924 = n24923 ^ n23882 ;
  assign n24921 = n23856 ^ n23845 ;
  assign n24925 = n24924 ^ n24921 ;
  assign n24926 = ~n23745 & n24925 ;
  assign n24927 = n24926 ^ n24924 ;
  assign n24936 = n24935 ^ n24927 ;
  assign n24942 = n24941 ^ n24936 ;
  assign n24943 = ~n23714 & ~n24942 ;
  assign n24928 = n24927 ^ n23951 ;
  assign n24917 = n23890 ^ n23882 ;
  assign n24918 = n23946 & ~n24917 ;
  assign n24919 = n24918 ^ n23882 ;
  assign n24920 = n23746 & n24919 ;
  assign n24929 = n24928 ^ n24920 ;
  assign n24930 = n24929 ^ n23960 ;
  assign n24911 = n23905 ^ n23857 ;
  assign n24912 = n23857 ^ n23714 ;
  assign n24913 = n24912 ^ n23857 ;
  assign n24914 = n24911 & ~n24913 ;
  assign n24915 = n24914 ^ n23857 ;
  assign n24916 = n23746 & n24915 ;
  assign n24931 = n24930 ^ n24916 ;
  assign n24905 = n23938 ^ n23856 ;
  assign n24906 = n23856 ^ n23714 ;
  assign n24907 = n24906 ^ n23856 ;
  assign n24908 = n24905 & n24907 ;
  assign n24909 = n24908 ^ n23856 ;
  assign n24910 = ~n23746 & n24909 ;
  assign n24932 = n24931 ^ n24910 ;
  assign n24944 = n24943 ^ n24932 ;
  assign n24946 = n24945 ^ n24944 ;
  assign n24947 = ~n23861 & ~n24946 ;
  assign n24948 = n24947 ^ n21412 ;
  assign n24975 = ~n23861 & n23968 ;
  assign n24970 = n23882 ^ n23859 ;
  assign n24971 = n24970 ^ n23905 ;
  assign n24972 = n24971 ^ n24923 ;
  assign n24973 = ~n23745 & n24972 ;
  assign n24967 = n24923 ^ n23858 ;
  assign n24968 = n23878 & n24967 ;
  assign n24958 = n24920 ^ n23887 ;
  assign n24957 = n24910 ^ n23853 ;
  assign n24959 = n24958 ^ n24957 ;
  assign n24956 = n24923 ^ n23859 ;
  assign n24960 = n24959 ^ n24956 ;
  assign n24954 = n23861 ^ n23856 ;
  assign n24955 = n24954 ^ n24916 ;
  assign n24961 = n24960 ^ n24955 ;
  assign n24962 = n24961 ^ n23931 ;
  assign n24963 = n24962 ^ n23891 ;
  assign n24964 = n24963 ^ n20616 ;
  assign n24951 = n23864 ^ n23847 ;
  assign n24952 = n24951 ^ n23861 ;
  assign n24953 = ~n23714 & n24952 ;
  assign n24965 = n24964 ^ n24953 ;
  assign n24949 = n24923 ^ n23856 ;
  assign n24950 = ~n23887 & n24949 ;
  assign n24966 = n24965 ^ n24950 ;
  assign n24969 = n24968 ^ n24966 ;
  assign n24974 = n24973 ^ n24969 ;
  assign n24976 = n24975 ^ n24974 ;
  assign n24992 = n24074 ^ n22618 ;
  assign n24989 = n22625 ^ n22606 ;
  assign n24990 = n21526 & n24989 ;
  assign n24991 = n24990 ^ n22646 ;
  assign n24993 = n24992 ^ n24991 ;
  assign n24985 = n22643 ^ n22618 ;
  assign n24986 = n24985 ^ n22638 ;
  assign n24987 = n24986 ^ n24074 ;
  assign n24988 = n21526 & ~n24987 ;
  assign n24994 = n24993 ^ n24988 ;
  assign n24995 = ~n21813 & ~n24994 ;
  assign n24996 = n24995 ^ n24991 ;
  assign n24984 = n22624 & n22633 ;
  assign n24997 = n24996 ^ n24984 ;
  assign n24983 = ~n22634 & n24088 ;
  assign n24998 = n24997 ^ n24983 ;
  assign n24977 = n22640 ^ n22606 ;
  assign n24978 = n22606 ^ n21526 ;
  assign n24979 = n24978 ^ n22606 ;
  assign n24980 = n24977 & ~n24979 ;
  assign n24981 = n24980 ^ n22606 ;
  assign n24982 = n21812 & n24981 ;
  assign n24999 = n24998 ^ n24982 ;
  assign n25000 = ~n24098 & ~n24999 ;
  assign n25001 = ~n22681 & n25000 ;
  assign n25002 = n25001 ^ n21985 ;
  assign y0 = ~n20972 ;
  assign y1 = ~n22693 ;
  assign y2 = ~n21525 ;
  assign y3 = ~n23060 ;
  assign y4 = ~n23083 ;
  assign y5 = ~n23122 ;
  assign y6 = ~n23163 ;
  assign y7 = ~n23404 ;
  assign y8 = ~n23433 ;
  assign y9 = ~n23468 ;
  assign y10 = ~n23506 ;
  assign y11 = ~n23678 ;
  assign y12 = ~n23713 ;
  assign y13 = ~n23928 ;
  assign y14 = ~n23561 ;
  assign y15 = ~n23970 ;
  assign y16 = ~n24008 ;
  assign y17 = n24040 ;
  assign y18 = n24061 ;
  assign y19 = n24101 ;
  assign y20 = n24139 ;
  assign y21 = ~n24178 ;
  assign y22 = n23598 ;
  assign y23 = ~n24204 ;
  assign y24 = n23744 ;
  assign y25 = ~n24247 ;
  assign y26 = n22727 ;
  assign y27 = n24359 ;
  assign y28 = n21811 ;
  assign y29 = n24390 ;
  assign y30 = n23192 ;
  assign y31 = ~n24495 ;
  assign y32 = n23784 ;
  assign y33 = ~n24537 ;
  assign y34 = n22854 ;
  assign y35 = n24555 ;
  assign y36 = ~n22580 ;
  assign y37 = ~n24621 ;
  assign y38 = n23231 ;
  assign y39 = n24655 ;
  assign y40 = n23839 ;
  assign y41 = ~n24688 ;
  assign y42 = ~n22898 ;
  assign y43 = ~n24734 ;
  assign y44 = n22058 ;
  assign y45 = n24765 ;
  assign y46 = ~n23283 ;
  assign y47 = n24791 ;
  assign y48 = ~n23809 ;
  assign y49 = n24825 ;
  assign y50 = n22972 ;
  assign y51 = n24849 ;
  assign y52 = n22289 ;
  assign y53 = n24882 ;
  assign y54 = ~n23234 ;
  assign y55 = ~n24883 ;
  assign y56 = n23518 ;
  assign y57 = n24904 ;
  assign y58 = n22945 ;
  assign y59 = ~n24948 ;
  assign y60 = n22457 ;
  assign y61 = n24976 ;
  assign y62 = ~n23316 ;
  assign y63 = ~n25002 ;
endmodule
