module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n226 , n227 , n228 , n229 , n230 , n231 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n271 , n272 , n273 , n274 , n275 ;
  assign n65 = x59 ^ x27 ;
  assign n69 = ~x27 & x59 ;
  assign n67 = ~x25 & ~x57 ;
  assign n66 = x58 ^ x57 ;
  assign n68 = n67 ^ n66 ;
  assign n70 = n69 ^ n68 ;
  assign n73 = x59 ^ x26 ;
  assign n71 = x59 ^ x57 ;
  assign n72 = n71 ^ n67 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~n70 & ~n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = ~n65 & n76 ;
  assign n78 = n77 ^ x27 ;
  assign n79 = ~x28 & x60 ;
  assign n80 = ~x31 & x63 ;
  assign n81 = ~n79 & n80 ;
  assign n82 = n81 ^ x29 ;
  assign n83 = n81 ^ n79 ;
  assign n84 = x61 & ~n83 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = ~x30 & x62 ;
  assign n88 = ~n86 & n87 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = ~n78 & ~n89 ;
  assign n133 = n67 ^ x25 ;
  assign n134 = ~n69 & n133 ;
  assign n135 = ~x26 & x58 ;
  assign n136 = n134 & n135 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = x24 & n137 ;
  assign n91 = x55 ^ x23 ;
  assign n93 = ~x22 & x54 ;
  assign n92 = x54 ^ x22 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = n94 ^ x55 ;
  assign n96 = ~n91 & n95 ;
  assign n97 = n96 ^ x23 ;
  assign n98 = x53 ^ x21 ;
  assign n100 = ~x20 & x52 ;
  assign n99 = x52 ^ x20 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ x53 ;
  assign n103 = ~n98 & n102 ;
  assign n104 = n103 ^ x21 ;
  assign n105 = ~x23 & x55 ;
  assign n106 = ~n93 & n105 ;
  assign n107 = n106 ^ n93 ;
  assign n108 = n104 & ~n107 ;
  assign n109 = x51 ^ x19 ;
  assign n111 = x50 ^ x18 ;
  assign n115 = x50 ^ x49 ;
  assign n116 = n115 ^ x17 ;
  assign n113 = ~x16 & x48 ;
  assign n112 = x48 ^ x16 ;
  assign n114 = n113 ^ n112 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = x49 ^ x17 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = n120 ^ n115 ;
  assign n122 = ~n111 & n121 ;
  assign n110 = x51 ^ x50 ;
  assign n123 = n122 ^ n110 ;
  assign n124 = ~n109 & ~n123 ;
  assign n125 = n124 ^ x19 ;
  assign n126 = ~n100 & ~n107 ;
  assign n127 = ~x21 & x53 ;
  assign n128 = n126 & n127 ;
  assign n129 = n128 ^ n126 ;
  assign n130 = n125 & n129 ;
  assign n131 = ~n108 & ~n130 ;
  assign n132 = ~n97 & n131 ;
  assign n139 = n138 ^ n132 ;
  assign n140 = ~x56 & n137 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = ~n139 & n141 ;
  assign n143 = n142 ^ n138 ;
  assign n144 = n90 & ~n143 ;
  assign n145 = n144 ^ n89 ;
  assign n146 = x63 ^ x31 ;
  assign n148 = x60 ^ x28 ;
  assign n149 = n148 ^ n79 ;
  assign n150 = n149 ^ x62 ;
  assign n147 = x62 ^ x29 ;
  assign n151 = n150 ^ n147 ;
  assign n152 = x62 ^ x61 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = n151 & ~n153 ;
  assign n155 = n154 ^ n150 ;
  assign n157 = x63 ^ x30 ;
  assign n156 = x63 ^ x62 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n155 & ~n158 ;
  assign n160 = n159 ^ n157 ;
  assign n161 = ~n146 & n160 ;
  assign n162 = n161 ^ x31 ;
  assign n163 = ~n109 & ~n111 ;
  assign n164 = ~x15 & x47 ;
  assign n165 = x47 ^ x15 ;
  assign n168 = ~x13 & ~x45 ;
  assign n166 = x46 ^ x45 ;
  assign n167 = n166 ^ n164 ;
  assign n169 = n168 ^ n167 ;
  assign n172 = x47 ^ x14 ;
  assign n170 = x47 ^ x46 ;
  assign n171 = n170 ^ n164 ;
  assign n173 = n172 ^ n171 ;
  assign n174 = ~n169 & ~n173 ;
  assign n175 = n174 ^ n172 ;
  assign n176 = ~n165 & n175 ;
  assign n177 = n176 ^ x15 ;
  assign n178 = ~n164 & ~n177 ;
  assign n179 = n168 ^ x13 ;
  assign n180 = x42 ^ x10 ;
  assign n181 = x43 ^ x11 ;
  assign n182 = ~n180 & ~n181 ;
  assign n184 = x9 & ~x41 ;
  assign n183 = x41 ^ x9 ;
  assign n185 = n184 ^ n183 ;
  assign n188 = x8 & ~n185 ;
  assign n189 = n182 & n188 ;
  assign n186 = ~x40 & ~n185 ;
  assign n187 = n182 & n186 ;
  assign n190 = n189 ^ n187 ;
  assign n192 = x39 ^ x38 ;
  assign n191 = x39 ^ x6 ;
  assign n193 = n192 ^ n191 ;
  assign n216 = x39 ^ x5 ;
  assign n220 = n216 ^ n191 ;
  assign n195 = x34 ^ x2 ;
  assign n196 = x33 ^ x1 ;
  assign n197 = n196 ^ n195 ;
  assign n200 = ~x0 & x32 ;
  assign n201 = n200 ^ x1 ;
  assign n202 = ~n197 & ~n201 ;
  assign n198 = x34 ^ x1 ;
  assign n203 = n202 ^ n198 ;
  assign n204 = ~n195 & ~n203 ;
  assign n194 = x35 ^ x34 ;
  assign n205 = n204 ^ n194 ;
  assign n207 = x36 ^ x3 ;
  assign n206 = x36 ^ x35 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = ~n205 & ~n208 ;
  assign n210 = n209 ^ n207 ;
  assign n212 = x37 ^ x4 ;
  assign n211 = x37 ^ x36 ;
  assign n213 = n212 ^ n211 ;
  assign n214 = n210 & ~n213 ;
  assign n215 = n214 ^ n212 ;
  assign n218 = x37 ^ x5 ;
  assign n219 = n215 & ~n218 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = ~n193 & ~n221 ;
  assign n223 = n222 ^ n192 ;
  assign n226 = x39 ^ x7 ;
  assign n227 = ~n223 & ~n226 ;
  assign n224 = n189 ^ x7 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n190 & n228 ;
  assign n230 = n229 ^ n189 ;
  assign n234 = n184 ^ x43 ;
  assign n231 = x43 ^ x42 ;
  assign n235 = n234 ^ n231 ;
  assign n236 = ~n180 & ~n235 ;
  assign n237 = n236 ^ n231 ;
  assign n238 = ~n181 & n237 ;
  assign n239 = n238 ^ x43 ;
  assign n240 = ~n230 & n239 ;
  assign n241 = n240 ^ x44 ;
  assign n242 = x44 ^ x12 ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = n243 ^ x12 ;
  assign n245 = n179 & n244 ;
  assign n246 = n178 & n245 ;
  assign n254 = x46 & n246 ;
  assign n255 = ~x14 & n254 ;
  assign n256 = n255 ^ x14 ;
  assign n247 = n246 ^ n177 ;
  assign n248 = n247 ^ x14 ;
  assign n257 = n256 ^ n248 ;
  assign n258 = ~n113 & n257 ;
  assign n259 = n163 & n258 ;
  assign n260 = ~n119 & n259 ;
  assign n261 = n129 & n260 ;
  assign n262 = ~n89 & n261 ;
  assign n263 = ~n162 & n262 ;
  assign n271 = ~n140 & n263 ;
  assign n272 = ~n138 & n271 ;
  assign n273 = n272 ^ n138 ;
  assign n264 = n263 ^ n162 ;
  assign n265 = n264 ^ n138 ;
  assign n274 = n273 ^ n265 ;
  assign n275 = n145 & ~n274 ;
  assign y0 = n275 ;
endmodule
