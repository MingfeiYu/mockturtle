module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1481 , n1482 , n1483 , n1484 , n1485 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1584 , n1585 , n1586 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1614 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1641 , n1642 , n1643 , n1644 , n1645 , n1647 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1663 , n1664 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1674 , n1675 , n1676 , n1677 , n1678 , n1681 , n1682 , n1689 , n1690 , n1691 , n1695 , n1696 , n1698 , n1699 , n1701 , n1702 , n1704 , n1706 , n1708 , n1713 , n1717 , n1718 , n1719 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1730 , n1731 , n1732 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1819 , n1822 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1892 , n1893 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2059 , n2060 , n2061 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2090 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2171 , n2172 , n2175 , n2176 , n2177 , n2178 , n2182 , n2183 , n2184 , n2185 , n2186 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2250 , n2251 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2293 , n2294 , n2295 , n2296 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2306 , n2309 , n2310 , n2311 , n2312 , n2313 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2346 , n2347 , n2348 , n2349 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2396 , n2397 , n2398 , n2399 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2439 , n2440 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2455 , n2456 , n2457 , n2458 , n2460 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2766 , n2768 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2852 , n2853 , n2854 , n2855 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2881 , n2882 , n2883 , n2884 , n2885 , n2887 , n2888 , n2889 , n2894 , n2895 , n2896 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2916 , n2917 , n2918 , n2920 , n2921 , n2922 , n2924 , n2925 , n2926 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3058 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3102 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3203 , n3204 , n3205 , n3206 , n3207 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3325 , n3335 , n3346 , n3348 , n3357 , n3358 , n3359 , n3360 , n3362 , n3363 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3375 , n3376 , n3378 , n3379 , n3380 , n3381 , n3382 , n3384 , n3385 , n3386 , n3388 , n3389 , n3390 , n3391 , n3392 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3406 , n3407 , n3408 , n3409 , n3410 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3518 , n3519 , n3520 , n3521 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3534 , n3537 , n3538 , n3539 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3558 , n3559 , n3560 , n3561 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3616 , n3617 , n3618 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3635 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3648 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3809 , n3810 , n3811 , n3812 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3829 , n3830 , n3831 , n3832 , n3833 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4021 , n4022 , n4023 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4042 , n4043 , n4044 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4079 , n4080 , n4081 , n4082 , n4083 , n4085 , n4095 , n4106 , n4108 , n4117 , n4118 , n4119 , n4120 , n4122 , n4123 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4135 , n4136 , n4138 , n4139 , n4140 , n4141 , n4142 , n4144 , n4145 , n4146 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4180 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4198 , n4209 , n4211 , n4220 , n4221 , n4222 , n4223 , n4225 , n4226 , n4227 , n4228 , n4231 , n4232 , n4233 , n4234 , n4238 , n4239 , n4241 , n4242 , n4243 , n4244 , n4245 , n4247 , n4248 , n4249 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4268 , n4269 , n4270 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4388 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4422 , n4423 , n4424 , n4425 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4517 , n4518 , n4519 , n4520 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4553 , n4554 , n4555 , n4556 , n4557 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4659 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4671 , n4673 , n4683 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4701 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4726 , n4727 , n4728 , n4734 , n4735 , n4736 , n4742 , n4743 , n4744 , n4745 , n4748 , n4749 , n4750 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4762 , n4763 , n4764 , n4771 , n4772 , n4773 , n4774 , n4776 , n4777 , n4778 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4828 , n4829 , n4830 , n4831 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4857 , n4858 , n4859 , n4864 , n4865 , n4866 , n4867 , n4868 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4980 , n4981 , n4982 , n4983 , n4985 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5042 , n5043 , n5044 , n5045 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5065 , n5066 , n5074 , n5075 , n5076 , n5077 , n5081 , n5082 , n5087 , n5090 , n5100 , n5102 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5114 , n5115 , n5116 , n5117 , n5119 , n5120 , n5128 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5170 , n5171 , n5172 , n5173 , n5174 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5211 , n5212 , n5213 , n5214 , n5215 , n5218 , n5219 , n5220 , n5221 , n5222 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5271 , n5272 , n5273 , n5274 , n5275 , n5282 , n5283 , n5284 , n5287 , n5288 , n5289 , n5290 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5319 , n5320 , n5321 , n5322 , n5323 , n5325 , n5326 , n5327 , n5328 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5341 , n5342 , n5343 , n5344 , n5345 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5361 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5445 , n5446 , n5447 , n5448 , n5452 , n5453 , n5454 , n5455 , n5456 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5482 , n5485 , n5486 , n5487 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5513 , n5514 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5599 , n5600 , n5601 , n5602 , n5603 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5644 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5660 , n5661 , n5662 , n5663 , n5666 , n5667 , n5668 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5885 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5894 , n5897 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5906 , n5907 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5942 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5951 , n5954 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5963 , n5966 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5975 , n5976 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5989 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5998 , n5999 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6070 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6359 , n6360 , n6361 , n6362 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6559 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6569 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6696 , n6697 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6835 , n6836 , n6837 , n6838 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6882 , n6883 , n6884 , n6885 , n6886 , n6891 , n6892 , n6893 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6922 , n6923 , n6924 , n6925 , n6926 , n6929 , n6930 , n6931 , n6932 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6998 , n6999 , n7000 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7029 , n7030 , n7031 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7045 , n7046 , n7047 , n7048 , n7049 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7061 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7101 , n7102 , n7103 , n7104 , n7106 , n7107 , n7110 , n7113 , n7114 , n7115 , n7116 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7128 , n7131 , n7132 , n7133 , n7134 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7147 , n7148 , n7149 , n7150 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7203 , n7206 , n7207 , n7208 , n7209 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7221 , n7224 , n7225 , n7226 , n7227 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7248 , n7251 , n7252 , n7253 , n7254 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7652 , n7653 , n7654 , n7659 , n7660 , n7661 , n7662 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8657 , n8658 , n8659 , n8660 , n8663 , n8664 , n8665 , n8666 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8803 , n8804 , n8805 , n8806 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8830 , n8831 , n8832 , n8838 , n8842 , n8848 , n8852 , n8853 , n8854 , n8855 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8880 , n8881 , n8883 , n8887 , n8888 , n8889 , n8890 , n8892 , n8893 , n8894 , n8895 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8925 , n8926 , n8927 , n8928 , n8929 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8953 , n8954 , n8955 , n8956 , n8959 , n8960 , n8961 , n8962 , n8965 , n8966 , n8967 , n8968 , n8971 , n8972 , n8973 , n8974 , n8977 , n8978 , n8979 , n8980 , n8983 , n8984 , n8985 , n8986 , n8989 , n8990 , n8991 , n8992 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9008 , n9011 , n9024 , n9025 , n9026 , n9027 , n9029 , n9030 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9042 , n9043 , n9044 , n9046 , n9051 , n9058 , n9059 , n9060 , n9063 , n9064 , n9065 , n9066 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9087 , n9088 , n9089 , n9090 , n9093 , n9094 , n9095 , n9096 , n9099 , n9100 , n9101 , n9102 , n9105 , n9106 , n9107 , n9108 , n9111 , n9112 , n9113 , n9114 , n9117 , n9118 , n9119 , n9120 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9138 , n9139 , n9140 , n9141 , n9144 , n9145 , n9146 , n9147 , n9150 , n9151 , n9152 , n9153 , n9156 , n9157 , n9158 , n9159 , n9162 , n9163 , n9164 , n9165 , n9168 , n9169 , n9170 , n9171 , n9174 , n9175 , n9176 , n9177 , n9180 , n9181 , n9182 , n9183 , n9186 , n9187 , n9188 , n9189 , n9192 , n9193 , n9194 , n9195 , n9198 , n9199 , n9200 , n9201 , n9204 , n9205 , n9206 , n9207 , n9210 , n9211 , n9212 , n9213 , n9216 , n9217 , n9218 , n9219 , n9222 , n9223 , n9224 , n9225 , n9228 , n9229 , n9230 , n9231 , n9234 , n9235 , n9236 , n9237 , n9240 , n9241 , n9242 , n9243 , n9246 , n9247 , n9248 , n9249 , n9252 , n9253 , n9254 , n9255 , n9258 , n9259 , n9260 , n9261 , n9264 , n9265 , n9266 , n9267 , n9270 , n9271 , n9272 , n9273 , n9276 , n9277 , n9278 , n9279 , n9282 , n9283 , n9284 , n9285 , n9288 , n9289 , n9290 , n9291 , n9294 , n9295 , n9296 , n9297 , n9300 , n9301 , n9302 , n9303 , n9306 , n9307 , n9308 , n9309 , n9312 , n9313 , n9314 , n9315 , n9318 , n9319 , n9320 , n9321 , n9324 , n9325 , n9326 , n9327 , n9330 , n9331 , n9332 , n9333 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9352 , n9353 , n9354 , n9355 , n9358 , n9359 , n9360 , n9361 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9378 , n9381 , n9382 , n9383 , n9393 , n9396 , n9400 , n9401 , n9406 , n9408 , n9410 , n9416 , n9417 , n9418 , n9419 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9437 , n9438 , n9448 , n9449 , n9450 , n9454 , n9455 , n9456 , n9457 , n9458 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9500 , n9501 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9514 , n9517 , n9518 , n9519 , n9529 , n9532 , n9536 , n9537 , n9542 , n9544 , n9546 , n9552 , n9553 , n9554 , n9555 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9573 , n9574 , n9584 , n9585 , n9586 , n9590 , n9591 , n9592 , n9593 , n9594 , n9596 , n9597 , n9598 , n9599 , n9600 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9624 , n9625 , n9628 , n9629 , n9630 , n9631 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9644 , n9647 , n9648 , n9649 , n9659 , n9662 , n9666 , n9667 , n9672 , n9674 , n9676 , n9682 , n9683 , n9684 , n9685 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9703 , n9704 , n9714 , n9715 , n9716 , n9720 , n9721 , n9722 , n9723 , n9724 , n9726 , n9727 , n9728 , n9729 , n9730 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9762 , n9765 , n9766 , n9767 , n9777 , n9780 , n9784 , n9785 , n9790 , n9792 , n9794 , n9800 , n9801 , n9802 , n9803 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9821 , n9822 , n9832 , n9833 , n9834 , n9838 , n9839 , n9841 , n9843 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9886 , n9889 , n9890 , n9891 , n9901 , n9904 , n9908 , n9909 , n9914 , n9916 , n9918 , n9924 , n9925 , n9926 , n9927 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9945 , n9946 , n9956 , n9957 , n9958 , n9962 , n9963 , n9965 , n9967 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10028 , n10029 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10078 , n10081 , n10082 , n10083 , n10093 , n10096 , n10100 , n10101 , n10106 , n10108 , n10110 , n10116 , n10117 , n10118 , n10119 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10137 , n10138 , n10148 , n10149 , n10150 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10192 , n10195 , n10196 , n10197 , n10207 , n10210 , n10214 , n10215 , n10220 , n10222 , n10224 , n10230 , n10231 , n10232 , n10233 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10251 , n10252 , n10262 , n10263 , n10264 , n10268 , n10269 , n10271 , n10273 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10322 , n10325 , n10326 , n10327 , n10337 , n10340 , n10344 , n10345 , n10350 , n10352 , n10354 , n10360 , n10361 , n10362 , n10363 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10381 , n10382 , n10392 , n10393 , n10394 , n10398 , n10399 , n10400 , n10401 , n10402 , n10404 , n10405 , n10406 , n10407 , n10408 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10440 , n10443 , n10444 , n10445 , n10455 , n10458 , n10462 , n10463 , n10468 , n10470 , n10472 , n10478 , n10479 , n10480 , n10481 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10499 , n10500 , n10510 , n10511 , n10512 , n10516 , n10517 , n10519 , n10520 , n10521 , n10522 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10570 , n10573 , n10574 , n10575 , n10585 , n10588 , n10592 , n10593 , n10598 , n10600 , n10602 , n10608 , n10609 , n10610 , n10611 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10629 , n10630 , n10640 , n10641 , n10642 , n10646 , n10647 , n10648 , n10649 , n10650 , n10652 , n10653 , n10654 , n10655 , n10656 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10688 , n10691 , n10692 , n10693 , n10703 , n10706 , n10710 , n10711 , n10716 , n10718 , n10720 , n10726 , n10727 , n10728 , n10729 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10747 , n10748 , n10758 , n10759 , n10760 , n10764 , n10765 , n10767 , n10769 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10828 , n10831 , n10832 , n10833 , n10843 , n10846 , n10850 , n10851 , n10856 , n10858 , n10860 , n10866 , n10867 , n10868 , n10869 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10887 , n10888 , n10898 , n10899 , n10900 , n10904 , n10905 , n10907 , n10908 , n10909 , n10910 , n10913 , n10914 , n10915 , n10916 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10936 , n10937 , n10938 , n10939 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10984 , n10987 , n10988 , n10989 , n10999 , n11002 , n11006 , n11007 , n11012 , n11014 , n11016 , n11022 , n11023 , n11024 , n11025 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11043 , n11044 , n11054 , n11055 , n11056 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11102 , n11103 , n11104 , n11105 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11117 , n11120 , n11121 , n11122 , n11132 , n11135 , n11139 , n11140 , n11145 , n11147 , n11149 , n11155 , n11156 , n11157 , n11158 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11176 , n11177 , n11187 , n11188 , n11189 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11220 , n11221 , n11222 , n11223 , n11224 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11236 , n11239 , n11240 , n11241 , n11251 , n11254 , n11258 , n11259 , n11264 , n11266 , n11268 , n11274 , n11275 , n11276 , n11277 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11295 , n11296 , n11306 , n11307 , n11308 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11351 , n11352 , n11353 , n11354 , n11357 , n11358 , n11359 , n11360 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11373 , n11376 , n11377 , n11378 , n11388 , n11391 , n11395 , n11396 , n11401 , n11403 , n11405 , n11411 , n11412 , n11413 , n11414 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11432 , n11433 , n11443 , n11444 , n11445 , n11449 , n11450 , n11452 , n11453 , n11454 , n11455 , n11458 , n11459 , n11460 , n11461 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11489 , n11490 , n11491 , n11492 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11504 , n11507 , n11508 , n11509 , n11519 , n11522 , n11526 , n11527 , n11532 , n11534 , n11536 , n11542 , n11543 , n11544 , n11545 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11563 , n11564 , n11574 , n11575 , n11576 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11618 , n11619 , n11620 , n11621 , n11624 , n11625 , n11626 , n11627 , n11630 , n11631 , n11632 , n11633 , n11636 , n11637 , n11638 , n11639 , n11642 , n11643 , n11644 , n11645 , n11648 , n11649 , n11650 , n11651 , n11654 , n11655 , n11656 , n11657 , n11660 , n11661 , n11662 , n11663 , n11666 , n11667 , n11668 , n11669 , n11672 , n11673 , n11674 , n11675 , n11678 , n11679 , n11680 , n11681 , n11684 , n11685 , n11686 , n11687 , n11690 , n11691 , n11692 , n11693 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11705 , n11708 , n11709 , n11710 , n11720 , n11723 , n11727 , n11728 , n11733 , n11735 , n11737 , n11743 , n11744 , n11745 , n11746 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11764 , n11765 , n11775 , n11776 , n11777 , n11781 , n11782 , n11783 , n11784 , n11785 , n11787 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11832 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11846 , n11849 , n11850 , n11851 , n11861 , n11864 , n11868 , n11869 , n11874 , n11876 , n11878 , n11884 , n11885 , n11886 , n11887 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11905 , n11906 , n11916 , n11917 , n11918 , n11922 , n11923 , n11925 , n11926 , n11927 , n11928 , n11929 , n11931 , n11932 , n11933 , n11934 , n11935 , n11938 , n11939 , n11940 , n11941 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11953 , n11956 , n11957 , n11958 , n11968 , n11971 , n11975 , n11976 , n11981 , n11983 , n11985 , n11991 , n11992 , n11993 , n11994 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12012 , n12013 , n12023 , n12024 , n12025 , n12029 , n12030 , n12031 , n12032 , n12033 , n12035 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12070 , n12073 , n12074 , n12075 , n12085 , n12088 , n12092 , n12093 , n12098 , n12100 , n12102 , n12108 , n12109 , n12110 , n12111 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12129 , n12130 , n12140 , n12141 , n12142 , n12146 , n12147 , n12148 , n12149 , n12150 , n12152 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12187 , n12190 , n12191 , n12192 , n12202 , n12205 , n12209 , n12210 , n12215 , n12217 , n12219 , n12225 , n12226 , n12227 , n12228 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12246 , n12247 , n12257 , n12258 , n12259 , n12263 , n12264 , n12265 , n12266 , n12267 , n12269 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12305 , n12308 , n12309 , n12310 , n12320 , n12323 , n12327 , n12328 , n12333 , n12335 , n12337 , n12343 , n12344 , n12345 , n12346 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12364 , n12365 , n12375 , n12376 , n12377 , n12381 , n12382 , n12384 , n12385 , n12386 , n12387 , n12390 , n12391 , n12392 , n12393 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12422 , n12423 , n12424 , n12426 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12448 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12478 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12496 , n12499 , n12500 , n12501 , n12511 , n12514 , n12518 , n12519 , n12524 , n12526 , n12528 , n12534 , n12535 , n12536 , n12537 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12555 , n12556 , n12566 , n12567 , n12568 , n12572 , n12573 , n12575 , n12576 , n12577 , n12578 , n12581 , n12582 , n12583 , n12584 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12623 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12649 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12667 , n12670 , n12671 , n12672 , n12682 , n12685 , n12689 , n12690 , n12695 , n12697 , n12699 , n12705 , n12706 , n12707 , n12708 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12726 , n12727 , n12737 , n12738 , n12739 , n12743 , n12744 , n12746 , n12747 , n12748 , n12749 , n12752 , n12753 , n12754 , n12755 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12787 , n12790 , n12791 , n12792 , n12802 , n12805 , n12809 , n12810 , n12815 , n12817 , n12819 , n12825 , n12826 , n12827 , n12828 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12846 , n12847 , n12857 , n12858 , n12859 , n12863 , n12864 , n12866 , n12867 , n12868 , n12869 , n12872 , n12873 , n12874 , n12875 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12934 , n12937 , n12938 , n12939 , n12949 , n12952 , n12956 , n12957 , n12962 , n12964 , n12966 , n12972 , n12973 , n12974 , n12975 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12993 , n12994 , n13004 , n13005 , n13006 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13049 , n13050 , n13051 , n13052 , n13055 , n13056 , n13057 , n13058 , n13061 , n13062 , n13063 , n13064 , n13067 , n13068 , n13069 , n13070 , n13073 , n13074 , n13075 , n13076 , n13079 , n13080 , n13081 , n13082 , n13085 , n13086 , n13087 , n13088 , n13091 , n13092 , n13093 , n13094 , n13099 , n13100 , n13101 , n13102 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13124 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13138 , n13141 , n13142 , n13143 , n13153 , n13156 , n13160 , n13161 , n13166 , n13168 , n13170 , n13176 , n13177 , n13178 , n13179 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13197 , n13198 , n13208 , n13209 , n13210 , n13214 , n13215 , n13217 , n13218 , n13219 , n13220 , n13221 , n13223 , n13224 , n13225 , n13226 , n13227 , n13230 , n13231 , n13232 , n13233 , n13236 , n13237 , n13238 , n13239 , n13242 , n13243 , n13244 , n13245 , n13248 , n13249 , n13250 , n13251 , n13254 , n13255 , n13256 , n13257 , n13260 , n13261 , n13262 , n13263 , n13266 , n13267 , n13268 , n13269 , n13272 , n13273 , n13274 , n13275 , n13278 , n13279 , n13280 , n13281 , n13284 , n13285 , n13286 , n13287 , n13290 , n13291 , n13292 , n13293 , n13296 , n13297 , n13298 , n13303 , n13304 , n13305 , n13306 , n13309 , n13310 , n13311 , n13312 , n13315 , n13316 , n13317 , n13318 , n13321 , n13322 , n13323 , n13324 , n13327 , n13328 , n13329 , n13330 , n13333 , n13334 , n13335 , n13336 , n13339 , n13340 , n13341 , n13342 , n13345 , n13346 , n13347 , n13348 , n13351 , n13352 , n13353 , n13354 , n13357 , n13358 , n13359 , n13360 , n13363 , n13364 , n13365 , n13366 , n13369 , n13370 , n13371 , n13372 , n13375 , n13376 , n13377 , n13378 , n13381 , n13382 , n13383 , n13384 , n13387 , n13388 , n13389 , n13390 , n13393 , n13394 , n13395 , n13396 , n13399 , n13400 , n13401 , n13402 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13423 , n13424 , n13425 , n13426 , n13429 , n13430 , n13431 , n13432 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13461 , n13462 , n13463 , n13468 , n13469 , n13470 , n13471 , n13474 , n13475 , n13476 , n13477 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 ;
  assign n1205 = ~x56 & ~x62 ;
  assign n1206 = ~x55 & n1205 ;
  assign n1207 = x57 & ~x59 ;
  assign n1208 = n1207 ^ x59 ;
  assign n1209 = n1206 & ~n1208 ;
  assign n1210 = ~x75 & x100 ;
  assign n1211 = n1210 ^ x75 ;
  assign n1212 = ~x87 & ~n1211 ;
  assign n1213 = ~x38 & ~x54 ;
  assign n1214 = ~x74 & ~x92 ;
  assign n1215 = n1213 & n1214 ;
  assign n1216 = n1212 & n1215 ;
  assign n1217 = x39 & n1216 ;
  assign n1218 = n1217 ^ n1216 ;
  assign n1219 = n1209 & ~n1218 ;
  assign n1220 = n1219 ^ n1209 ;
  assign n1221 = ~x69 & ~x83 ;
  assign n1222 = ~x103 & n1221 ;
  assign n1223 = x82 & ~x111 ;
  assign n1224 = n1223 ^ x111 ;
  assign n1225 = ~x36 & ~n1224 ;
  assign n1226 = ~x66 & n1225 ;
  assign n1227 = n1222 & n1226 ;
  assign n1228 = ~x85 & ~x106 ;
  assign n1229 = ~x76 & n1228 ;
  assign n1230 = ~x48 & ~x61 ;
  assign n1231 = n1229 & n1230 ;
  assign n1233 = x104 & ~n1231 ;
  assign n1232 = n1231 ^ x104 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1235 = n1234 ^ x89 ;
  assign n1236 = ~x49 & ~n1233 ;
  assign n1237 = n1236 ^ x89 ;
  assign n1238 = ~n1235 & ~n1237 ;
  assign n1239 = n1238 ^ x89 ;
  assign n1240 = ~x45 & ~n1239 ;
  assign n1241 = ~x89 & n1234 ;
  assign n1242 = ~x49 & n1241 ;
  assign n1244 = ~n1240 & ~n1242 ;
  assign n1243 = n1242 ^ n1240 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1246 = n1227 & ~n1245 ;
  assign n1247 = ~x73 & n1246 ;
  assign n1248 = ~x88 & ~x98 ;
  assign n1249 = ~x102 & ~x107 ;
  assign n1250 = n1248 & n1249 ;
  assign n1251 = ~x64 & ~x65 ;
  assign n1252 = ~x63 & n1251 ;
  assign n1253 = n1250 & n1252 ;
  assign n1254 = ~x81 & n1253 ;
  assign n1255 = n1247 & n1254 ;
  assign n1256 = ~x67 & ~x68 ;
  assign n1257 = ~x71 & ~x84 ;
  assign n1258 = n1256 & n1257 ;
  assign n1259 = n1255 & n1258 ;
  assign n1260 = ~x91 & ~x109 ;
  assign n1261 = ~x46 & ~x47 ;
  assign n1262 = n1260 & n1261 ;
  assign n1263 = ~x77 & ~x86 ;
  assign n1264 = ~x50 & ~x110 ;
  assign n1265 = n1263 & n1264 ;
  assign n1266 = n1262 & n1265 ;
  assign n1267 = ~x53 & x60 ;
  assign n1268 = n1267 ^ x53 ;
  assign n1269 = ~x58 & ~n1268 ;
  assign n1270 = ~x97 & ~x108 ;
  assign n1271 = ~x94 & n1270 ;
  assign n1272 = n1269 & n1271 ;
  assign n1273 = n1266 & n1272 ;
  assign n1274 = n1259 & n1273 ;
  assign n1275 = x35 & ~x93 ;
  assign n1276 = n1275 ^ x93 ;
  assign n1277 = ~x90 & ~n1276 ;
  assign n1296 = ~x72 & ~x96 ;
  assign n1297 = ~x51 & ~x70 ;
  assign n1298 = n1296 & n1297 ;
  assign n1299 = n1277 & n1298 ;
  assign n1300 = n1274 & n1299 ;
  assign n1511 = ~x40 & x95 ;
  assign n1509 = x40 ^ x32 ;
  assign n1301 = ~x90 & n1274 ;
  assign n1302 = x93 ^ x35 ;
  assign n1303 = n1301 & n1302 ;
  assign n1304 = ~x50 & ~n1268 ;
  assign n1305 = ~x77 & n1304 ;
  assign n1306 = n1270 & n1305 ;
  assign n1308 = x86 & x94 ;
  assign n1307 = x94 ^ x86 ;
  assign n1309 = n1308 ^ n1307 ;
  assign n1310 = n1306 & ~n1309 ;
  assign n1311 = n1259 & n1310 ;
  assign n1312 = x46 & ~x109 ;
  assign n1313 = n1312 ^ x109 ;
  assign n1314 = x53 ^ x50 ;
  assign n1315 = n1314 ^ n1267 ;
  assign n1316 = n1268 ^ x60 ;
  assign n1317 = n1316 ^ n1267 ;
  assign n1318 = n1317 ^ n1268 ;
  assign n1321 = ~x77 & ~n1318 ;
  assign n1322 = n1321 ^ n1268 ;
  assign n1323 = n1315 & n1322 ;
  assign n1324 = n1323 ^ x50 ;
  assign n1325 = ~n1313 & ~n1324 ;
  assign n1326 = n1311 & n1325 ;
  assign n1327 = ~x58 & ~x90 ;
  assign n1328 = ~x47 & ~x110 ;
  assign n1329 = n1327 & n1328 ;
  assign n1330 = ~x91 & ~x93 ;
  assign n1331 = n1329 & n1330 ;
  assign n1332 = ~n1326 & ~n1331 ;
  assign n1333 = x110 ^ x90 ;
  assign n1334 = x90 ^ x58 ;
  assign n1335 = n1333 & ~n1334 ;
  assign n1336 = n1335 ^ x110 ;
  assign n1337 = x91 ^ x47 ;
  assign n1338 = n1327 ^ x91 ;
  assign n1339 = n1337 & ~n1338 ;
  assign n1340 = n1339 ^ x91 ;
  assign n1341 = ~n1276 & ~n1340 ;
  assign n1342 = n1339 ^ n1336 ;
  assign n1343 = n1342 ^ n1341 ;
  assign n1344 = n1339 ^ n1335 ;
  assign n1345 = n1344 ^ n1341 ;
  assign n1346 = n1335 ^ x47 ;
  assign n1347 = n1346 ^ n1336 ;
  assign n1348 = ~n1345 & n1347 ;
  assign n1349 = n1343 & n1348 ;
  assign n1350 = n1349 ^ n1335 ;
  assign n1351 = n1350 ^ n1336 ;
  assign n1352 = n1341 & ~n1351 ;
  assign n1353 = ~n1336 & n1352 ;
  assign n1354 = ~n1332 & n1353 ;
  assign n1496 = ~x46 & ~n1260 ;
  assign n1355 = n1247 & n1258 ;
  assign n1358 = x98 ^ x88 ;
  assign n1359 = n1358 ^ x102 ;
  assign n1360 = n1359 ^ x107 ;
  assign n1361 = x102 ^ x98 ;
  assign n1363 = ~n1358 & n1361 ;
  assign n1364 = n1363 ^ x102 ;
  assign n1365 = n1360 & ~n1364 ;
  assign n1366 = n1365 ^ n1250 ;
  assign n1367 = ~x81 & n1366 ;
  assign n1368 = n1367 ^ n1250 ;
  assign n1375 = n1368 ^ x63 ;
  assign n1371 = ~x102 & n1258 ;
  assign n1372 = ~x81 & n1248 ;
  assign n1373 = n1371 & n1372 ;
  assign n1376 = n1375 ^ n1373 ;
  assign n1356 = x65 ^ x64 ;
  assign n1357 = x65 ^ x63 ;
  assign n1369 = n1368 ^ n1357 ;
  assign n1370 = ~n1356 & n1369 ;
  assign n1374 = n1373 ^ n1370 ;
  assign n1377 = n1376 ^ n1374 ;
  assign n1382 = n1368 & n1374 ;
  assign n1383 = n1382 ^ n1373 ;
  assign n1384 = ~n1377 & n1383 ;
  assign n1385 = n1355 & n1384 ;
  assign n1460 = ~x71 & ~x81 ;
  assign n1461 = n1253 & n1460 ;
  assign n1397 = x68 ^ x66 ;
  assign n1398 = n1397 ^ x73 ;
  assign n1399 = n1398 ^ x84 ;
  assign n1400 = x73 ^ x68 ;
  assign n1401 = x84 ^ x73 ;
  assign n1402 = n1400 & ~n1401 ;
  assign n1403 = n1402 ^ x68 ;
  assign n1404 = ~x66 & ~n1403 ;
  assign n1405 = ~n1399 & n1404 ;
  assign n1406 = ~n1245 & n1405 ;
  assign n1417 = ~x36 & ~x67 ;
  assign n1418 = ~n1224 & n1417 ;
  assign n1455 = n1406 & n1418 ;
  assign n1468 = n1255 & n1455 ;
  assign n1407 = n1222 & n1406 ;
  assign n1408 = x82 ^ x36 ;
  assign n1410 = x82 ^ x67 ;
  assign n1409 = x111 ^ x82 ;
  assign n1411 = n1410 ^ n1409 ;
  assign n1412 = n1411 ^ x82 ;
  assign n1413 = ~n1408 & n1412 ;
  assign n1414 = n1413 ^ n1411 ;
  assign n1415 = n1407 & ~n1414 ;
  assign n1424 = x111 & ~n1413 ;
  assign n1416 = n1415 ^ n1222 ;
  assign n1419 = n1418 ^ n1416 ;
  assign n1425 = n1424 ^ n1419 ;
  assign n1426 = n1415 & n1425 ;
  assign n1427 = n1426 ^ n1419 ;
  assign n1428 = n1427 ^ n1222 ;
  assign n1429 = ~n1416 & ~n1426 ;
  assign n1430 = ~n1428 & n1429 ;
  assign n1431 = n1430 ^ n1427 ;
  assign n1434 = x83 ^ x69 ;
  assign n1435 = x103 ^ x83 ;
  assign n1436 = n1434 & ~n1435 ;
  assign n1437 = n1436 ^ x69 ;
  assign n1456 = n1455 ^ n1437 ;
  assign n1439 = ~n1244 & n1405 ;
  assign n1432 = n1399 & ~n1403 ;
  assign n1433 = ~n1245 & n1432 ;
  assign n1440 = x106 ^ x85 ;
  assign n1441 = x85 ^ x76 ;
  assign n1442 = n1440 & n1441 ;
  assign n1443 = n1442 ^ x85 ;
  assign n1444 = n1230 & ~n1443 ;
  assign n1445 = n1444 ^ x48 ;
  assign n1446 = n1445 ^ x61 ;
  assign n1447 = n1446 ^ n1444 ;
  assign n1450 = n1229 & n1447 ;
  assign n1451 = n1450 ^ n1444 ;
  assign n1452 = ~n1433 & n1451 ;
  assign n1453 = n1439 & n1452 ;
  assign n1438 = n1437 ^ n1433 ;
  assign n1454 = n1453 ^ n1438 ;
  assign n1457 = n1456 ^ n1454 ;
  assign n1458 = n1457 ^ n1455 ;
  assign n1459 = ~n1431 & n1458 ;
  assign n1462 = n1461 ^ n1459 ;
  assign n1469 = n1468 ^ n1462 ;
  assign n1470 = ~n1461 & ~n1469 ;
  assign n1471 = n1470 ^ n1462 ;
  assign n1472 = n1471 ^ n1437 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1474 = n1459 ^ n1455 ;
  assign n1475 = n1470 ^ n1459 ;
  assign n1476 = n1474 & ~n1475 ;
  assign n1477 = n1473 & n1476 ;
  assign n1478 = n1477 ^ n1471 ;
  assign n1481 = ~n1385 & n1478 ;
  assign n1386 = x108 ^ x97 ;
  assign n1387 = n1386 ^ n1305 ;
  assign n1388 = n1387 ^ n1309 ;
  assign n1389 = n1305 ^ x108 ;
  assign n1390 = n1309 ^ x108 ;
  assign n1391 = ~n1389 & n1390 ;
  assign n1392 = n1391 ^ x108 ;
  assign n1393 = ~n1388 & ~n1392 ;
  assign n1394 = n1393 ^ n1259 ;
  assign n1482 = n1481 ^ n1394 ;
  assign n1483 = n1310 & n1482 ;
  assign n1484 = n1483 ^ n1394 ;
  assign n1485 = n1484 ^ n1259 ;
  assign n1487 = n1484 ^ n1310 ;
  assign n1488 = ~n1483 & ~n1487 ;
  assign n1489 = ~n1485 & n1488 ;
  assign n1490 = n1489 ^ n1485 ;
  assign n1491 = n1490 ^ n1259 ;
  assign n1492 = n1325 & ~n1491 ;
  assign n1493 = ~n1308 & n1492 ;
  assign n1497 = n1496 ^ n1493 ;
  assign n1498 = n1311 & n1497 ;
  assign n1499 = n1498 ^ n1493 ;
  assign n1500 = n1329 & n1499 ;
  assign n1501 = n1500 ^ n1329 ;
  assign n1502 = n1354 & ~n1501 ;
  assign n1278 = n1274 & n1277 ;
  assign n1279 = ~x32 & ~x95 ;
  assign n1280 = ~x40 & n1279 ;
  assign n1281 = x96 ^ x51 ;
  assign n1282 = x72 ^ x70 ;
  assign n1283 = n1282 ^ x96 ;
  assign n1284 = ~n1281 & n1283 ;
  assign n1285 = n1284 ^ n1282 ;
  assign n1286 = n1280 & ~n1285 ;
  assign n1287 = n1278 & n1286 ;
  assign n1288 = x72 & ~n1284 ;
  assign n1289 = n1287 & n1288 ;
  assign n1290 = n1289 ^ n1287 ;
  assign n1503 = n1280 & n1298 ;
  assign n1504 = ~n1290 & n1503 ;
  assign n1505 = ~n1502 & n1504 ;
  assign n1506 = ~n1303 & n1505 ;
  assign n1507 = n1506 ^ n1504 ;
  assign n1508 = n1507 ^ n1290 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1512 = n1511 ^ n1510 ;
  assign n1513 = n1512 ^ n1508 ;
  assign n1514 = n1512 ^ x95 ;
  assign n1515 = n1514 ^ n1511 ;
  assign n1516 = n1515 ^ n1512 ;
  assign n1517 = n1513 & n1516 ;
  assign n1518 = n1517 ^ n1512 ;
  assign n1519 = n1300 & n1518 ;
  assign n1520 = n1519 ^ n1508 ;
  assign n1521 = ~x228 & n1520 ;
  assign n1294 = ~x105 & x228 ;
  assign n1295 = n1294 ^ x228 ;
  assign n1522 = n1521 ^ n1295 ;
  assign n1535 = ~x215 & x299 ;
  assign n1525 = x216 & ~x221 ;
  assign n1536 = n1525 ^ x221 ;
  assign n1537 = n1535 & n1536 ;
  assign n1538 = n1537 ^ n1535 ;
  assign n1539 = n1522 & n1538 ;
  assign n1529 = ~x223 & ~x299 ;
  assign n1532 = x224 & n1529 ;
  assign n1530 = x222 & n1529 ;
  assign n1531 = ~x224 & n1530 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1534 = n1533 ^ n1529 ;
  assign n1540 = n1539 ^ n1534 ;
  assign n1291 = x96 & n1290 ;
  assign n1292 = x95 & ~x479 ;
  assign n1293 = ~n1291 & ~n1292 ;
  assign n1543 = ~n1503 & ~n1520 ;
  assign n1594 = ~x95 & n1301 ;
  assign n1595 = n1301 ^ x93 ;
  assign n1596 = ~x40 & ~x51 ;
  assign n1597 = n1296 & n1596 ;
  assign n1598 = n1597 ^ x225 ;
  assign n1601 = ~x35 & n1598 ;
  assign n1602 = n1601 ^ x225 ;
  assign n1603 = n1595 & n1602 ;
  assign n1604 = n1603 ^ x35 ;
  assign n1605 = n1594 & ~n1604 ;
  assign n1606 = n1605 ^ x95 ;
  assign n1607 = ~n1502 & ~n1606 ;
  assign n1544 = ~x97 & ~x137 ;
  assign n1545 = ~x35 & n1544 ;
  assign n1546 = ~n1268 & n1545 ;
  assign n1547 = n1546 ^ n1544 ;
  assign n1548 = n1547 ^ x137 ;
  assign n1549 = x210 ^ x198 ;
  assign n1550 = x299 & n1549 ;
  assign n1551 = n1550 ^ x198 ;
  assign n1552 = x146 ^ x142 ;
  assign n1553 = x299 & n1552 ;
  assign n1554 = n1553 ^ x142 ;
  assign n1557 = ~x152 & ~x166 ;
  assign n1558 = ~x161 & n1557 ;
  assign n1555 = ~x174 & ~x189 ;
  assign n1556 = ~x144 & n1555 ;
  assign n1559 = n1558 ^ n1556 ;
  assign n1560 = ~x299 & n1559 ;
  assign n1561 = n1560 ^ n1558 ;
  assign n1562 = ~n1554 & ~n1561 ;
  assign n1563 = ~n1551 & ~n1562 ;
  assign n1564 = x950 & x1092 ;
  assign n1565 = x829 & n1564 ;
  assign n1566 = x1091 & x1093 ;
  assign n1568 = ~x833 & x957 ;
  assign n1569 = n1566 & n1568 ;
  assign n1567 = n1566 ^ x1093 ;
  assign n1570 = n1569 ^ n1567 ;
  assign n1571 = n1565 & ~n1570 ;
  assign n1572 = ~x841 & n1571 ;
  assign n1588 = n1291 & n1572 ;
  assign n1573 = ~x46 & ~x94 ;
  assign n1574 = x97 ^ x36 ;
  assign n1575 = n1573 & n1574 ;
  assign n1576 = ~x1093 & n1565 ;
  assign n1577 = n1576 ^ n1571 ;
  assign n1578 = n1575 & n1577 ;
  assign n1579 = x97 & n1331 ;
  assign n1580 = n1492 & n1579 ;
  assign n1581 = n1331 & n1503 ;
  assign n1582 = ~x35 & n1581 ;
  assign n1584 = n1580 & n1582 ;
  assign n1585 = n1584 ^ n1291 ;
  assign n1586 = ~n1578 & n1585 ;
  assign n1589 = n1588 ^ n1586 ;
  assign n1590 = n1589 ^ n1585 ;
  assign n1591 = n1563 & n1590 ;
  assign n1592 = ~n1548 & n1591 ;
  assign n1593 = n1592 ^ n1548 ;
  assign n1608 = n1326 & n1328 ;
  assign n1609 = n1311 & ~n1608 ;
  assign n1610 = n1327 & n1609 ;
  assign n1614 = ~x109 & ~x110 ;
  assign n1619 = n1610 & ~n1614 ;
  assign n1620 = ~n1261 & n1619 ;
  assign n1621 = n1620 ^ n1261 ;
  assign n1611 = n1610 ^ n1327 ;
  assign n1612 = n1611 ^ n1261 ;
  assign n1622 = n1621 ^ n1612 ;
  assign n1623 = n1354 & ~n1622 ;
  assign n1624 = n1593 & ~n1623 ;
  assign n1625 = n1607 & n1624 ;
  assign n1626 = n1625 ^ n1593 ;
  assign n1627 = ~n1543 & n1626 ;
  assign n1541 = n1540 ^ x234 ;
  assign n1526 = ~x215 & n1525 ;
  assign n1523 = ~x215 & x221 ;
  assign n1524 = n1523 ^ x215 ;
  assign n1527 = n1526 ^ n1524 ;
  assign n1528 = n1522 & ~n1527 ;
  assign n1542 = n1541 ^ n1528 ;
  assign n1628 = n1627 ^ n1542 ;
  assign n1629 = n1628 ^ n1540 ;
  assign n1630 = n1629 ^ n1528 ;
  assign n1631 = n1293 & n1630 ;
  assign n1632 = n1631 ^ n1542 ;
  assign n1681 = n1632 ^ n1540 ;
  assign n1641 = x153 & ~n1295 ;
  assign n1674 = ~x332 & n1538 ;
  assign n1675 = n1641 & n1674 ;
  assign n1676 = n1675 ^ n1538 ;
  assign n1642 = ~x216 & x833 ;
  assign n1643 = ~x215 & ~x929 ;
  assign n1644 = n1642 & n1643 ;
  assign n1645 = n1644 ^ x215 ;
  assign n1653 = ~x221 & ~n1645 ;
  assign n1654 = x265 & n1653 ;
  assign n1655 = n1654 ^ x265 ;
  assign n1647 = n1644 ^ x265 ;
  assign n1656 = n1655 ^ n1647 ;
  assign n1657 = ~x332 & ~n1656 ;
  assign n1663 = n1523 & n1642 ;
  assign n1664 = n1663 ^ n1524 ;
  assign n1667 = n1657 & n1664 ;
  assign n1668 = ~x1144 & n1667 ;
  assign n1669 = n1668 ^ x1144 ;
  assign n1658 = n1657 ^ x332 ;
  assign n1659 = n1658 ^ x1144 ;
  assign n1670 = n1669 ^ n1659 ;
  assign n1671 = n1527 & n1670 ;
  assign n1672 = x299 & ~n1671 ;
  assign n1677 = n1676 ^ n1672 ;
  assign n1678 = n1677 ^ n1528 ;
  assign n1682 = n1681 ^ n1678 ;
  assign n1633 = ~x40 & n1300 ;
  assign n1634 = n1279 ^ x95 ;
  assign n1635 = n1633 & ~n1634 ;
  assign n1636 = ~x841 & n1551 ;
  assign n1637 = n1636 ^ x841 ;
  assign n1638 = x225 & n1637 ;
  assign n1639 = n1635 & n1638 ;
  assign n1689 = n1682 ^ n1639 ;
  assign n1690 = n1689 ^ n1632 ;
  assign n1698 = n1690 ^ n1677 ;
  assign n1699 = n1698 ^ n1689 ;
  assign n1691 = n1690 ^ n1682 ;
  assign n1717 = n1699 ^ n1691 ;
  assign n1701 = n1699 ^ n1528 ;
  assign n1718 = n1717 ^ n1701 ;
  assign n1719 = n1540 & n1718 ;
  assign n1708 = ~n1677 & ~n1678 ;
  assign n1721 = n1719 ^ n1708 ;
  assign n1695 = n1690 ^ n1639 ;
  assign n1696 = n1695 ^ n1677 ;
  assign n1704 = n1696 ^ n1691 ;
  assign n1722 = n1721 ^ n1704 ;
  assign n1702 = n1701 ^ n1689 ;
  assign n1723 = n1722 ^ n1702 ;
  assign n1724 = n1723 ^ n1691 ;
  assign n1725 = n1724 ^ n1701 ;
  assign n1713 = n1632 ^ n1528 ;
  assign n1735 = n1725 ^ n1713 ;
  assign n1736 = n1735 ^ n1690 ;
  assign n1726 = n1698 ^ n1678 ;
  assign n1730 = n1726 ^ n1681 ;
  assign n1731 = n1730 ^ n1701 ;
  assign n1732 = n1731 ^ n1677 ;
  assign n1737 = n1736 ^ n1732 ;
  assign n1738 = n1737 ^ n1713 ;
  assign n1739 = n1738 ^ n1528 ;
  assign n1706 = n1701 ^ n1698 ;
  assign n1740 = n1739 ^ n1706 ;
  assign n1741 = n1220 & ~n1740 ;
  assign n1742 = ~n1209 & ~n1671 ;
  assign n1743 = n1280 & n1300 ;
  assign n1744 = n1218 & n1743 ;
  assign n1745 = n1205 & n1744 ;
  assign n1746 = n1207 & n1745 ;
  assign n1747 = ~x55 & n1746 ;
  assign n1754 = ~x39 & ~x87 ;
  assign n1755 = ~x38 & n1754 ;
  assign n1756 = ~x92 & ~n1211 ;
  assign n1757 = n1755 & n1756 ;
  assign n1758 = ~x74 & n1757 ;
  assign n1759 = ~x57 & n1205 ;
  assign n1761 = ~x54 & ~x59 ;
  assign n1760 = x59 ^ x54 ;
  assign n1762 = n1761 ^ n1760 ;
  assign n1763 = n1759 & n1762 ;
  assign n1764 = n1761 ^ x55 ;
  assign n1765 = n1763 & ~n1764 ;
  assign n1766 = n1758 & n1765 ;
  assign n1767 = n1743 & n1766 ;
  assign n1748 = n1209 & n1743 ;
  assign n1749 = ~x54 & n1214 ;
  assign n1750 = n1212 & n1749 ;
  assign n1751 = x38 & ~x39 ;
  assign n1752 = n1750 & n1751 ;
  assign n1753 = n1748 & n1752 ;
  assign n1768 = n1767 ^ n1753 ;
  assign n1769 = ~n1747 & ~n1768 ;
  assign n1770 = n1748 & n1755 ;
  assign n1771 = x74 ^ x54 ;
  assign n1772 = n1771 ^ x75 ;
  assign n1773 = n1772 ^ x92 ;
  assign n1774 = x75 ^ x74 ;
  assign n1775 = x92 ^ x74 ;
  assign n1776 = n1774 & n1775 ;
  assign n1777 = n1776 ^ x74 ;
  assign n1778 = n1773 & ~n1777 ;
  assign n1779 = n1770 & n1778 ;
  assign n1780 = ~x100 & n1779 ;
  assign n1781 = n1769 & ~n1780 ;
  assign n1786 = ~x74 & ~x75 ;
  assign n1787 = n1213 & n1786 ;
  assign n1788 = x87 ^ x39 ;
  assign n1789 = n1788 ^ x92 ;
  assign n1790 = n1789 ^ x100 ;
  assign n1791 = x92 ^ x87 ;
  assign n1792 = x100 ^ x87 ;
  assign n1793 = n1791 & n1792 ;
  assign n1794 = n1793 ^ x87 ;
  assign n1795 = n1790 & ~n1794 ;
  assign n1796 = n1787 & n1795 ;
  assign n1797 = n1748 & n1796 ;
  assign n1782 = ~n1208 & n1744 ;
  assign n1783 = x62 ^ x56 ;
  assign n1784 = ~x55 & n1783 ;
  assign n1785 = n1782 & n1784 ;
  assign n1798 = n1797 ^ n1785 ;
  assign n1799 = n1781 & ~n1798 ;
  assign n1800 = ~x137 & ~n1294 ;
  assign n1801 = ~n1527 & n1800 ;
  assign n1802 = n1801 ^ n1527 ;
  assign n1803 = n1641 & ~n1802 ;
  assign n1811 = ~n1208 & n1803 ;
  assign n1812 = ~x228 & n1811 ;
  assign n1813 = n1812 ^ x228 ;
  assign n1804 = n1803 ^ n1802 ;
  assign n1805 = n1804 ^ x228 ;
  assign n1814 = n1813 ^ n1805 ;
  assign n1815 = ~n1799 & ~n1814 ;
  assign n1816 = n1742 & ~n1815 ;
  assign n1819 = n1782 & ~n1799 ;
  assign n1822 = x234 & n1292 ;
  assign n1825 = ~n1819 & ~n1822 ;
  assign n1826 = n1295 & n1825 ;
  assign n1827 = n1826 ^ n1295 ;
  assign n1817 = n1785 ^ n1295 ;
  assign n1828 = n1827 ^ n1817 ;
  assign n1829 = ~n1527 & ~n1828 ;
  assign n1830 = ~x228 & n1819 ;
  assign n1831 = n1641 & ~n1830 ;
  assign n1832 = n1829 & n1831 ;
  assign n1833 = n1832 ^ n1829 ;
  assign n1834 = n1816 & ~n1833 ;
  assign n1838 = ~x332 & ~n1802 ;
  assign n1839 = n1294 & n1838 ;
  assign n1840 = x153 & n1839 ;
  assign n1841 = n1840 ^ n1838 ;
  assign n1842 = n1841 ^ x332 ;
  assign n1843 = n1672 & ~n1842 ;
  assign n1835 = ~x137 & ~x332 ;
  assign n1836 = n1534 & n1835 ;
  assign n1844 = n1843 ^ n1836 ;
  assign n1845 = ~x39 & ~n1216 ;
  assign n1854 = ~n1677 & n1750 ;
  assign n1846 = ~x74 & ~n1211 ;
  assign n1847 = ~n1213 & n1846 ;
  assign n1848 = n1847 ^ n1846 ;
  assign n1849 = n1791 & n1848 ;
  assign n1855 = n1854 ^ n1849 ;
  assign n1856 = n1845 & n1855 ;
  assign n1857 = n1856 ^ n1216 ;
  assign n1858 = ~n1844 & n1857 ;
  assign n1859 = n1743 & n1858 ;
  assign n1860 = n1219 & ~n1859 ;
  assign n1861 = x100 ^ x75 ;
  assign n1862 = n1749 & n1861 ;
  assign n1863 = ~x198 & n1836 ;
  assign n1864 = ~n1556 & n1863 ;
  assign n1865 = ~x142 & n1864 ;
  assign n1866 = n1865 ^ n1863 ;
  assign n1867 = n1866 ^ n1836 ;
  assign n1868 = n1862 & ~n1867 ;
  assign n1869 = x137 & ~n1211 ;
  assign n1870 = n1778 & n1869 ;
  assign n1871 = ~n1868 & ~n1870 ;
  assign n1872 = n1672 & n1835 ;
  assign n1873 = ~x146 & ~n1558 ;
  assign n1874 = ~x210 & ~n1873 ;
  assign n1875 = n1872 & n1874 ;
  assign n1876 = n1875 ^ n1872 ;
  assign n1877 = ~n1871 & ~n1876 ;
  assign n1878 = n1743 & n1877 ;
  assign n1879 = n1755 & n1878 ;
  assign n1880 = n1879 ^ n1677 ;
  assign n1881 = ~x39 & x252 ;
  assign n1882 = ~n1849 & n1881 ;
  assign n1883 = ~n1873 & n1882 ;
  assign n1884 = ~x228 & n1796 ;
  assign n1885 = ~n1883 & n1884 ;
  assign n1886 = n1743 & n1885 ;
  assign n1887 = ~n1527 & n1886 ;
  assign n1888 = ~n1879 & n1887 ;
  assign n1889 = n1888 ^ n1879 ;
  assign n1892 = n1295 & n1538 ;
  assign n1893 = n1892 ^ n1534 ;
  assign n1898 = ~n1822 & n1893 ;
  assign n1899 = ~x332 & n1898 ;
  assign n1900 = n1899 ^ x332 ;
  assign n1890 = n1888 ^ x332 ;
  assign n1901 = n1900 ^ n1890 ;
  assign n1902 = ~n1889 & n1901 ;
  assign n1903 = n1902 ^ n1887 ;
  assign n1904 = ~n1880 & ~n1903 ;
  assign n1905 = n1904 ^ n1879 ;
  assign n1906 = n1860 & ~n1905 ;
  assign n1907 = ~x224 & x833 ;
  assign n1908 = x222 & ~x223 ;
  assign n1909 = ~n1907 & n1908 ;
  assign n1910 = n1909 ^ x223 ;
  assign n1911 = ~x299 & n1209 ;
  assign n1912 = x1144 & n1911 ;
  assign n1913 = n1910 & n1912 ;
  assign n1914 = n1913 ^ n1911 ;
  assign n1915 = x224 ^ x222 ;
  assign n1918 = x833 & x929 ;
  assign n1919 = n1918 ^ x265 ;
  assign n1920 = ~x224 & n1919 ;
  assign n1921 = n1920 ^ x265 ;
  assign n1922 = n1915 & n1921 ;
  assign n1923 = n1922 ^ x222 ;
  assign n1924 = ~x223 & ~n1923 ;
  assign n1925 = n1914 & n1924 ;
  assign n1926 = n1925 ^ n1914 ;
  assign n1927 = ~n1906 & ~n1926 ;
  assign n1928 = ~n1834 & n1927 ;
  assign n1929 = ~n1741 & n1928 ;
  assign n1930 = ~x332 & ~n1929 ;
  assign n1935 = n1531 ^ n1530 ;
  assign n1936 = n1935 ^ n1532 ;
  assign n1937 = x276 & n1936 ;
  assign n1933 = ~x299 & n1910 ;
  assign n1934 = x1146 & n1933 ;
  assign n1938 = n1937 ^ n1934 ;
  assign n1931 = n1530 & n1907 ;
  assign n1932 = x939 & n1931 ;
  assign n1939 = n1938 ^ n1932 ;
  assign n1940 = n1209 & ~n1939 ;
  assign n1953 = n1940 ^ n1209 ;
  assign n1941 = ~n1293 & n1521 ;
  assign n1942 = n1218 & ~n1527 ;
  assign n1943 = x299 & n1942 ;
  assign n1944 = n1218 & n1291 ;
  assign n1946 = n1944 ^ n1292 ;
  assign n1947 = n1893 & n1946 ;
  assign n1948 = n1943 & ~n1947 ;
  assign n1949 = n1941 & n1948 ;
  assign n1950 = n1949 ^ n1947 ;
  assign n1951 = x239 & n1950 ;
  assign n1952 = n1940 & n1951 ;
  assign n1954 = n1953 ^ n1952 ;
  assign n1956 = ~n1295 & ~n1527 ;
  assign n1962 = n1956 ^ n1527 ;
  assign n1963 = ~n1292 & ~n1962 ;
  assign n1964 = n1963 ^ n1962 ;
  assign n1965 = x239 & ~n1964 ;
  assign n1961 = x939 & n1663 ;
  assign n1966 = n1965 ^ n1961 ;
  assign n1958 = x1146 & n1664 ;
  assign n1957 = ~x154 & n1956 ;
  assign n1959 = n1958 ^ n1957 ;
  assign n1955 = x276 & n1526 ;
  assign n1960 = n1959 ^ n1955 ;
  assign n1967 = n1966 ^ n1960 ;
  assign n1968 = ~n1527 & ~n1911 ;
  assign n1969 = n1209 & n1886 ;
  assign n1970 = n1968 & ~n1969 ;
  assign n1971 = n1220 & n1520 ;
  assign n1972 = ~n1819 & ~n1971 ;
  assign n1978 = ~x228 & ~n1972 ;
  assign n1973 = n1968 ^ n1911 ;
  assign n1979 = n1978 ^ n1973 ;
  assign n1980 = n1970 & n1979 ;
  assign n1981 = n1980 ^ n1973 ;
  assign n1982 = n1967 & ~n1981 ;
  assign n1983 = ~n1954 & n1982 ;
  assign n1984 = n1983 ^ n1954 ;
  assign n1987 = ~x274 & n1936 ;
  assign n1986 = x1145 & n1933 ;
  assign n1988 = n1987 ^ n1986 ;
  assign n1985 = x927 & n1931 ;
  assign n1989 = n1988 ^ n1985 ;
  assign n1990 = n1209 & ~n1989 ;
  assign n1992 = x235 & n1950 ;
  assign n1993 = n1990 & n1992 ;
  assign n1991 = n1990 ^ n1209 ;
  assign n1994 = n1993 ^ n1991 ;
  assign n2001 = x927 & n1663 ;
  assign n2000 = x235 & ~n1964 ;
  assign n2002 = n2001 ^ n2000 ;
  assign n1998 = ~x274 & n1526 ;
  assign n1996 = x1145 & n1664 ;
  assign n1995 = ~x151 & n1956 ;
  assign n1997 = n1996 ^ n1995 ;
  assign n1999 = n1998 ^ n1997 ;
  assign n2003 = n2002 ^ n1999 ;
  assign n2004 = ~n1994 & n2003 ;
  assign n2005 = ~n1981 & n2004 ;
  assign n2006 = n2005 ^ n1994 ;
  assign n2018 = ~n1294 & ~n1527 ;
  assign n2019 = x284 & ~n1292 ;
  assign n2020 = n2018 & n2019 ;
  assign n2021 = n2020 ^ n2018 ;
  assign n2012 = x1143 & n1664 ;
  assign n2011 = x146 & n1956 ;
  assign n2013 = n2012 ^ n2011 ;
  assign n2010 = ~x284 & n1963 ;
  assign n2014 = n2013 ^ n2010 ;
  assign n2008 = x944 & n1663 ;
  assign n2007 = ~x264 & n1526 ;
  assign n2009 = n2008 ^ n2007 ;
  assign n2015 = n2014 ^ n2009 ;
  assign n2059 = n2021 ^ n2015 ;
  assign n2067 = x238 & n2021 ;
  assign n2068 = x228 & n2067 ;
  assign n2069 = n2068 ^ x228 ;
  assign n2060 = ~n1527 & n1830 ;
  assign n2061 = n2060 ^ x228 ;
  assign n2070 = n2069 ^ n2061 ;
  assign n2071 = n2059 & n2070 ;
  assign n2072 = n2071 ^ n2015 ;
  assign n2073 = ~n1209 & n2072 ;
  assign n2016 = x299 & ~n1887 ;
  assign n2017 = n2015 & n2016 ;
  assign n2022 = n2021 ^ n2017 ;
  assign n2023 = n1886 ^ n1295 ;
  assign n2024 = n2017 ^ x299 ;
  assign n2025 = ~n1943 & n2024 ;
  assign n2026 = n2023 & n2025 ;
  assign n2027 = n2022 & n2026 ;
  assign n2028 = n2027 ^ n2025 ;
  assign n2029 = n2028 ^ n1943 ;
  assign n2030 = x284 & n1534 ;
  assign n2031 = ~x944 & n1209 ;
  assign n2032 = n1931 & n2031 ;
  assign n2033 = n2032 ^ n1936 ;
  assign n2034 = n2032 ^ n1209 ;
  assign n2035 = x264 & n2034 ;
  assign n2036 = n2033 & n2035 ;
  assign n2037 = n2036 ^ n2034 ;
  assign n2038 = ~x1143 & n1933 ;
  assign n2039 = n2037 & n2038 ;
  assign n2040 = n2039 ^ n2037 ;
  assign n2041 = ~n1946 & n2040 ;
  assign n2042 = n2030 & n2041 ;
  assign n2043 = n2042 ^ n2040 ;
  assign n2044 = n1950 & n2043 ;
  assign n2045 = ~x238 & n2044 ;
  assign n2046 = n2045 ^ n2043 ;
  assign n2047 = n2029 & n2046 ;
  assign n2050 = x284 & n1293 ;
  assign n2051 = n2050 ^ x146 ;
  assign n2052 = n1522 & ~n2051 ;
  assign n2053 = n2052 ^ x146 ;
  assign n2054 = n1942 & n2053 ;
  assign n2055 = n2054 ^ n2045 ;
  assign n2056 = n2047 & ~n2055 ;
  assign n2057 = n2056 ^ n2046 ;
  assign n2074 = n2073 ^ n2057 ;
  assign n2147 = ~x249 & n1534 ;
  assign n2148 = ~n1293 & n2147 ;
  assign n2082 = x216 & ~x277 ;
  assign n2075 = x1142 ^ x932 ;
  assign n2076 = ~n1642 & n2075 ;
  assign n2077 = n2076 ^ x932 ;
  assign n2083 = n2082 ^ n2077 ;
  assign n2084 = ~x221 & n2083 ;
  assign n2085 = n2084 ^ n2077 ;
  assign n2146 = n1535 & ~n2085 ;
  assign n2149 = n2148 ^ n2146 ;
  assign n2150 = n1220 & n2149 ;
  assign n2152 = x249 ^ x172 ;
  assign n2151 = x262 ^ x172 ;
  assign n2153 = n2152 ^ n2151 ;
  assign n2156 = n1293 & ~n2153 ;
  assign n2157 = n2156 ^ n2152 ;
  assign n2158 = n1522 & ~n2157 ;
  assign n2159 = n2158 ^ x172 ;
  assign n2160 = n1538 & ~n2159 ;
  assign n2090 = n1830 ^ n1295 ;
  assign n2095 = ~x172 & ~n1830 ;
  assign n2096 = n2095 ^ n1292 ;
  assign n2097 = ~n1295 & n2096 ;
  assign n2098 = n2097 ^ n1292 ;
  assign n2099 = ~x262 & ~n2098 ;
  assign n2100 = ~n2090 & n2099 ;
  assign n2101 = ~n1969 & n2100 ;
  assign n2102 = n2101 ^ n2099 ;
  assign n2103 = n2102 ^ n2098 ;
  assign n2104 = ~n1527 & n2103 ;
  assign n2086 = n2085 ^ x1142 ;
  assign n2087 = ~x215 & n2086 ;
  assign n2088 = n2087 ^ x1142 ;
  assign n2105 = n2104 ^ n2088 ;
  assign n2106 = n2105 ^ n1887 ;
  assign n2107 = n2106 ^ n1209 ;
  assign n2108 = n1887 ^ x299 ;
  assign n2109 = n2108 ^ n1209 ;
  assign n2110 = x299 ^ x262 ;
  assign n2111 = n2110 ^ n2105 ;
  assign n2112 = n2109 & n2111 ;
  assign n2113 = n2107 & n2112 ;
  assign n2114 = n2113 ^ x299 ;
  assign n2115 = n2114 ^ n2105 ;
  assign n2116 = n1209 & n2115 ;
  assign n2117 = n2105 & n2116 ;
  assign n2118 = n2117 ^ n2105 ;
  assign n2124 = ~x249 & n1292 ;
  assign n2137 = ~n1962 & n2124 ;
  assign n2129 = n2118 ^ n1209 ;
  assign n2121 = ~x277 & n1936 ;
  assign n2120 = x1142 & n1933 ;
  assign n2122 = n2121 ^ n2120 ;
  assign n2119 = x932 & n1931 ;
  assign n2123 = n2122 ^ n2119 ;
  assign n2130 = n2129 ^ n2123 ;
  assign n2125 = n1534 & ~n2124 ;
  assign n2131 = n2130 ^ n2125 ;
  assign n2127 = x262 & ~n1946 ;
  assign n2128 = n2125 & n2127 ;
  assign n2132 = n2131 ^ n2128 ;
  assign n2138 = n2137 ^ n2132 ;
  assign n2139 = n2118 & n2138 ;
  assign n2140 = n2139 ^ n2132 ;
  assign n2141 = n2140 ^ n1209 ;
  assign n2142 = n2140 ^ n2118 ;
  assign n2143 = ~n2139 & ~n2142 ;
  assign n2144 = ~n2141 & n2143 ;
  assign n2145 = n2144 ^ n2140 ;
  assign n2161 = n2160 ^ n2145 ;
  assign n2162 = n2150 & ~n2161 ;
  assign n2163 = n2162 ^ n2145 ;
  assign n2193 = x270 & n1936 ;
  assign n2192 = ~x1141 & n1933 ;
  assign n2194 = n2193 ^ n2192 ;
  assign n2191 = ~x935 & n1931 ;
  assign n2195 = n2194 ^ n2191 ;
  assign n2171 = x861 & ~n1292 ;
  assign n2172 = n2171 ^ x171 ;
  assign n2175 = n1295 & ~n2172 ;
  assign n2176 = n2175 ^ x171 ;
  assign n2177 = ~n1527 & n2176 ;
  assign n2167 = ~x1141 & n1664 ;
  assign n2166 = x270 & n1526 ;
  assign n2168 = n2167 ^ n2166 ;
  assign n2165 = ~x935 & n1663 ;
  assign n2169 = n2168 ^ n2165 ;
  assign n2178 = n2177 ^ n2169 ;
  assign n2196 = x299 & n1218 ;
  assign n2197 = ~n1528 & n2196 ;
  assign n2198 = n2178 & n2197 ;
  assign n2199 = n2198 ^ n2196 ;
  assign n2200 = n2199 ^ x299 ;
  assign n2201 = n1540 & ~n2200 ;
  assign n2202 = n2171 & n2201 ;
  assign n2203 = ~n1291 & n2202 ;
  assign n2204 = n2203 ^ n2201 ;
  assign n2205 = n2204 ^ n2200 ;
  assign n2209 = n2171 ^ x861 ;
  assign n2208 = n2178 ^ n2171 ;
  assign n2210 = n2209 ^ n2208 ;
  assign n2213 = ~n1887 & ~n2210 ;
  assign n2214 = n2213 ^ n2209 ;
  assign n2215 = x299 & n2214 ;
  assign n2216 = n2215 ^ n2171 ;
  assign n2217 = ~n1218 & n2216 ;
  assign n2218 = n2205 & n2217 ;
  assign n2206 = n2195 ^ n1209 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2219 = n2218 ^ n2207 ;
  assign n2220 = ~n2195 & n2219 ;
  assign n2188 = x241 & n1950 ;
  assign n2189 = n1209 & n2188 ;
  assign n2182 = ~n2060 & ~n2210 ;
  assign n2183 = n2182 ^ x861 ;
  assign n2184 = ~n1209 & ~n2183 ;
  assign n2186 = n2184 ^ n1209 ;
  assign n2190 = n2189 ^ n2186 ;
  assign n2221 = n2190 ^ n2184 ;
  assign n2222 = n2220 & n2221 ;
  assign n2223 = n2222 ^ n2190 ;
  assign n2164 = x241 & ~n1964 ;
  assign n2185 = n2164 & n2184 ;
  assign n2224 = n2223 ^ n2185 ;
  assign n2238 = n1209 & ~n1950 ;
  assign n2244 = ~n1292 & n1534 ;
  assign n2245 = x869 & n2244 ;
  assign n2243 = x1140 & n1933 ;
  assign n2246 = n2245 ^ n2243 ;
  assign n2241 = ~x282 & n1936 ;
  assign n2240 = x921 & n1931 ;
  assign n2242 = n2241 ^ n2240 ;
  assign n2247 = n2246 ^ n2242 ;
  assign n2229 = ~x1140 & n1664 ;
  assign n2228 = x282 & n1526 ;
  assign n2230 = n2229 ^ n2228 ;
  assign n2227 = ~x921 & n1663 ;
  assign n2231 = n2230 ^ n2227 ;
  assign n2239 = x299 & ~n2231 ;
  assign n2260 = n2247 ^ n2239 ;
  assign n2257 = x248 & ~n1209 ;
  assign n2258 = n1964 & n2257 ;
  assign n2259 = n2258 ^ x248 ;
  assign n2261 = n2260 ^ n2259 ;
  assign n2250 = x869 ^ x170 ;
  assign n2251 = n1218 & n1521 ;
  assign n2253 = n2251 ^ n2023 ;
  assign n2254 = ~n2250 & n2253 ;
  assign n2255 = n2254 ^ x170 ;
  assign n2256 = n1538 & n2255 ;
  assign n2262 = n2261 ^ n2256 ;
  assign n2263 = n2238 & n2262 ;
  assign n2264 = n2263 ^ n2259 ;
  assign n2225 = n2060 ^ n1963 ;
  assign n2232 = n1527 ^ x869 ;
  assign n2233 = n2232 ^ n2231 ;
  assign n2226 = ~x170 & n1956 ;
  assign n2234 = n2233 ^ n2226 ;
  assign n2235 = ~n2225 & n2234 ;
  assign n2236 = n2235 ^ x869 ;
  assign n2237 = ~n1209 & n2236 ;
  assign n2266 = n2264 ^ n2237 ;
  assign n2278 = x281 & n1526 ;
  assign n2277 = ~x1139 & n1664 ;
  assign n2279 = n2278 ^ n2277 ;
  assign n2275 = ~x920 & n1663 ;
  assign n2274 = x148 & n1956 ;
  assign n2276 = n2275 ^ n2274 ;
  assign n2280 = n2279 ^ n2276 ;
  assign n2284 = n2280 ^ x862 ;
  assign n2285 = n2284 ^ x247 ;
  assign n2286 = ~n1292 & n2285 ;
  assign n2287 = n2286 ^ x247 ;
  assign n2288 = ~n1962 & ~n2287 ;
  assign n2289 = n2288 ^ n2284 ;
  assign n2329 = ~n2060 & ~n2289 ;
  assign n2330 = n2329 ^ x862 ;
  assign n2331 = ~n1209 & n2330 ;
  assign n2306 = x862 ^ x247 ;
  assign n2309 = ~n1946 & n2306 ;
  assign n2310 = n2309 ^ x247 ;
  assign n7674 = n1209 & n1534 ;
  assign n2311 = ~n2310 & n7674 ;
  assign n2267 = ~x920 & n1209 ;
  assign n2268 = n1931 & n2267 ;
  assign n2269 = n2268 ^ n1936 ;
  assign n2270 = n2268 ^ n1209 ;
  assign n2271 = x281 & n2270 ;
  assign n2272 = n2269 & n2271 ;
  assign n2273 = n2272 ^ n2270 ;
  assign n2299 = ~x1139 & n1910 ;
  assign n2290 = n2289 ^ x862 ;
  assign n2293 = ~n1942 & n2290 ;
  assign n2294 = n2293 ^ x862 ;
  assign n2295 = ~n1887 & ~n2294 ;
  assign n2296 = n2295 ^ x862 ;
  assign n2300 = n2299 ^ n2296 ;
  assign n2301 = ~x299 & ~n2300 ;
  assign n2302 = n2301 ^ n2296 ;
  assign n2303 = n2273 & ~n2302 ;
  assign n2304 = n2303 ^ n2273 ;
  assign n2312 = n2311 ^ n2304 ;
  assign n2318 = n1293 & n2306 ;
  assign n2313 = x247 ^ x148 ;
  assign n2319 = n2318 ^ n2313 ;
  assign n2320 = n1522 & ~n2319 ;
  assign n2321 = n2320 ^ x148 ;
  assign n2322 = n1943 & n2321 ;
  assign n2323 = n2312 & n2322 ;
  assign n2324 = n2323 ^ n2312 ;
  assign n2332 = n2331 ^ n2324 ;
  assign n2335 = x269 & n1526 ;
  assign n2334 = ~x1138 & n1664 ;
  assign n2336 = n2335 ^ n2334 ;
  assign n2333 = ~x940 & n1663 ;
  assign n2337 = n2336 ^ n2333 ;
  assign n2338 = x299 & ~n2337 ;
  assign n2339 = x877 & ~n1292 ;
  assign n2340 = n2339 ^ x169 ;
  assign n2355 = n2023 & ~n2340 ;
  assign n2342 = x246 ^ x169 ;
  assign n2341 = x877 ^ x169 ;
  assign n2343 = n2342 ^ n2341 ;
  assign n2346 = n1293 & n2343 ;
  assign n2347 = n2346 ^ n2342 ;
  assign n2348 = n1522 & ~n2347 ;
  assign n2356 = n2355 ^ n2348 ;
  assign n2357 = ~n1218 & n2356 ;
  assign n2349 = n2348 ^ x169 ;
  assign n2358 = n2357 ^ n2349 ;
  assign n2359 = ~n1527 & n2358 ;
  assign n2360 = n2338 & ~n2359 ;
  assign n2364 = x940 & n1931 ;
  assign n2363 = ~x269 & n1936 ;
  assign n2365 = n2364 ^ n2363 ;
  assign n2366 = n2365 ^ x246 ;
  assign n2362 = x877 & n1534 ;
  assign n2367 = n2366 ^ n2362 ;
  assign n2361 = x1138 & n1933 ;
  assign n2368 = n2367 ^ n2361 ;
  assign n2369 = ~n1947 & n2368 ;
  assign n2370 = n2369 ^ x246 ;
  assign n2371 = n1209 & ~n2370 ;
  assign n2372 = ~n2360 & n2371 ;
  assign n2378 = n2090 & ~n2340 ;
  assign n2379 = n2378 ^ x169 ;
  assign n2380 = ~n1527 & n2379 ;
  assign n2381 = n2380 ^ n2337 ;
  assign n2382 = ~n1209 & n2381 ;
  assign n2383 = x246 & ~n1964 ;
  assign n2384 = n2382 & n2383 ;
  assign n2385 = n2384 ^ n2382 ;
  assign n2386 = ~n2372 & ~n2385 ;
  assign n2387 = x240 & n1534 ;
  assign n2389 = x933 & n1663 ;
  assign n2388 = x1137 & n1664 ;
  assign n2390 = n2389 ^ n2388 ;
  assign n2391 = x299 & ~n2390 ;
  assign n2399 = ~x280 & n1526 ;
  assign n2392 = x878 & ~n1292 ;
  assign n2393 = n2392 ^ x168 ;
  assign n2396 = n1295 & ~n2393 ;
  assign n2397 = n2396 ^ x168 ;
  assign n2398 = ~n1527 & ~n2397 ;
  assign n2401 = n2399 ^ n2398 ;
  assign n2402 = n2401 ^ x878 ;
  assign n2403 = ~n1887 & n2402 ;
  assign n2404 = n2403 ^ x878 ;
  assign n2405 = n2391 & ~n2404 ;
  assign n2407 = ~n1218 & ~n1947 ;
  assign n2406 = n1947 ^ n1218 ;
  assign n2408 = n2407 ^ n2406 ;
  assign n2409 = ~n2405 & n2408 ;
  assign n2410 = ~n1943 & n2409 ;
  assign n2411 = n1538 & ~n2407 ;
  assign n2413 = x240 ^ x168 ;
  assign n2412 = x878 ^ x168 ;
  assign n2414 = n2413 ^ n2412 ;
  assign n2417 = n1293 & n2414 ;
  assign n2418 = n2417 ^ n2413 ;
  assign n2419 = n1522 & ~n2418 ;
  assign n2420 = n2419 ^ x168 ;
  assign n2421 = n2411 & ~n2420 ;
  assign n2422 = ~n2410 & ~n2421 ;
  assign n2427 = ~x933 & n1931 ;
  assign n2426 = n1534 & ~n2392 ;
  assign n2428 = n2427 ^ n2426 ;
  assign n2424 = x280 & n1936 ;
  assign n2423 = ~x1137 & n1933 ;
  assign n2425 = n2424 ^ n2423 ;
  assign n2429 = n2428 ^ n2425 ;
  assign n2430 = ~n2422 & ~n2429 ;
  assign n2439 = n1946 & ~n2430 ;
  assign n2440 = n2387 & n2439 ;
  assign n2432 = n2390 ^ x878 ;
  assign n2433 = n2432 ^ n2401 ;
  assign n2431 = x240 & ~n1964 ;
  assign n2434 = n2433 ^ n2431 ;
  assign n2435 = ~n2060 & n2434 ;
  assign n2436 = n2435 ^ x878 ;
  assign n2437 = n2436 ^ n2430 ;
  assign n2442 = n2440 ^ n2437 ;
  assign n2443 = n1209 & n2442 ;
  assign n2444 = n2443 ^ n2436 ;
  assign n2447 = x266 & n1526 ;
  assign n2446 = x1136 & n1664 ;
  assign n2448 = n2447 ^ n2446 ;
  assign n2445 = x928 & n1663 ;
  assign n2449 = n2448 ^ n2445 ;
  assign n2450 = ~n1911 & ~n2449 ;
  assign n2451 = ~x875 & ~n1292 ;
  assign n2452 = n2451 ^ x166 ;
  assign n2455 = n2090 & ~n2452 ;
  assign n2456 = n2455 ^ x166 ;
  assign n2457 = ~n1220 & ~n2456 ;
  assign n2458 = n2457 ^ n1522 ;
  assign n2494 = x875 ^ x245 ;
  assign n2462 = n1293 & n2494 ;
  assign n2460 = n1209 ^ x245 ;
  assign n2463 = n2462 ^ n2460 ;
  assign n2464 = n2463 ^ n1209 ;
  assign n2465 = n1292 ^ x166 ;
  assign n2466 = n2465 ^ n2451 ;
  assign n2467 = n2023 & ~n2466 ;
  assign n2468 = n2467 ^ x166 ;
  assign n2471 = n2463 ^ n1219 ;
  assign n2472 = n2468 & ~n2471 ;
  assign n2473 = ~n2464 & n2472 ;
  assign n2474 = n2473 ^ n2464 ;
  assign n2475 = n2474 ^ n1209 ;
  assign n2476 = ~n2457 & ~n2475 ;
  assign n2477 = n2476 ^ n1209 ;
  assign n2478 = n2458 & ~n2477 ;
  assign n2479 = n2478 ^ n1522 ;
  assign n2480 = n1209 & ~n2468 ;
  assign n2481 = ~n1522 & n2480 ;
  assign n2482 = n2481 ^ n1527 ;
  assign n2483 = ~n1527 & ~n2482 ;
  assign n2484 = ~n2479 & n2483 ;
  assign n2485 = n2450 & ~n2484 ;
  assign n2495 = ~n1946 & n2494 ;
  assign n2496 = n2495 ^ x245 ;
  assign n2497 = ~n2496 & n7674 ;
  assign n2488 = ~x266 & n1936 ;
  assign n2487 = ~x1136 & n1933 ;
  assign n2489 = n2488 ^ n2487 ;
  assign n2486 = ~x928 & n1931 ;
  assign n2490 = n2489 ^ n2486 ;
  assign n2491 = n1209 & ~n2490 ;
  assign n2492 = n2491 ^ n1209 ;
  assign n2498 = n2497 ^ n2492 ;
  assign n2499 = ~n2485 & ~n2498 ;
  assign n2501 = x244 ^ x161 ;
  assign n2500 = x879 ^ x161 ;
  assign n2502 = n2501 ^ n2500 ;
  assign n2505 = ~n1292 & n2502 ;
  assign n2506 = n2505 ^ n2501 ;
  assign n2507 = n2090 & n2506 ;
  assign n2508 = n2507 ^ x161 ;
  assign n2509 = ~n1209 & ~n1527 ;
  assign n2510 = n2508 & n2509 ;
  assign n2511 = n2510 ^ n1209 ;
  assign n2514 = x279 & n1526 ;
  assign n2513 = x1135 & n1664 ;
  assign n2515 = n2514 ^ n2513 ;
  assign n2512 = x938 & n1663 ;
  assign n2516 = n2515 ^ n2512 ;
  assign n2517 = n2511 & ~n2516 ;
  assign n2519 = x938 & n1209 ;
  assign n2520 = n1931 & n2519 ;
  assign n2521 = n2520 ^ n1936 ;
  assign n2522 = n2520 ^ n1209 ;
  assign n2523 = x279 & n2522 ;
  assign n2524 = n2521 & n2523 ;
  assign n2525 = n2524 ^ n2522 ;
  assign n2518 = x879 & ~n1946 ;
  assign n2526 = n2525 ^ n2518 ;
  assign n2527 = x1135 & n1933 ;
  assign n2528 = n2525 & n2527 ;
  assign n2529 = n2528 ^ n2525 ;
  assign n2534 = n1538 & n2023 ;
  assign n2535 = n2534 ^ n1534 ;
  assign n2536 = n2529 & n2535 ;
  assign n2537 = ~n2526 & n2536 ;
  assign n2538 = n2537 ^ n2529 ;
  assign n2539 = x244 & n1950 ;
  assign n2540 = n2538 & n2539 ;
  assign n2541 = n2540 ^ n2538 ;
  assign n2542 = ~n1527 & n2541 ;
  assign n2543 = n2518 ^ x161 ;
  assign n2546 = ~n2253 & n2543 ;
  assign n2547 = n2546 ^ n2518 ;
  assign n2548 = n2542 & n2547 ;
  assign n2549 = n2548 ^ n2541 ;
  assign n2550 = n2517 & ~n2549 ;
  assign n2551 = n2550 ^ n2516 ;
  assign n2552 = ~x299 & n2541 ;
  assign n2553 = n2551 & n2552 ;
  assign n2554 = n2553 ^ n2551 ;
  assign n2570 = x846 ^ x242 ;
  assign n2560 = ~n1292 & n2570 ;
  assign n2555 = x242 ^ x152 ;
  assign n2561 = n2560 ^ n2555 ;
  assign n2562 = n2090 & n2561 ;
  assign n2563 = n2562 ^ x152 ;
  assign n2564 = n2509 & ~n2563 ;
  assign n2565 = n2564 ^ n1209 ;
  assign n2567 = ~x930 & n1663 ;
  assign n2566 = ~x278 & n1526 ;
  assign n2568 = n2567 ^ n2566 ;
  assign n2569 = n2565 & ~n2568 ;
  assign n2571 = ~n1946 & n2570 ;
  assign n2572 = n2571 ^ x242 ;
  assign n2573 = n1534 & ~n2572 ;
  assign n2575 = ~x278 & n1936 ;
  assign n2574 = ~x930 & n1931 ;
  assign n2576 = n2575 ^ n2574 ;
  assign n2577 = n1209 & ~n2576 ;
  assign n2578 = ~n2573 & n2577 ;
  assign n2579 = ~n1527 & n2578 ;
  assign n2580 = n2572 ^ x152 ;
  assign n2583 = ~n2253 & n2580 ;
  assign n2584 = n2583 ^ n2572 ;
  assign n2585 = n2579 & ~n2584 ;
  assign n2586 = n2585 ^ n2578 ;
  assign n2587 = n2569 & ~n2586 ;
  assign n2588 = n2587 ^ n2568 ;
  assign n2598 = ~x299 & n2578 ;
  assign n2592 = n2588 ^ x1134 ;
  assign n2589 = n1933 ^ n1664 ;
  assign n2590 = n1911 & n2589 ;
  assign n2591 = n2590 ^ n1664 ;
  assign n2593 = n2592 ^ n2591 ;
  assign n2599 = n2598 ^ n2593 ;
  assign n2600 = n2588 & ~n2599 ;
  assign n2601 = n2600 ^ n2593 ;
  assign n2602 = n2601 ^ x1134 ;
  assign n2603 = n2601 ^ n2591 ;
  assign n2604 = ~n2600 & n2603 ;
  assign n2605 = ~n2602 & n2604 ;
  assign n2606 = n2605 ^ n2601 ;
  assign n2607 = n1259 & n1271 ;
  assign n2608 = n1354 & ~n2607 ;
  assign n2609 = n1493 & n2608 ;
  assign n2610 = x93 & x841 ;
  assign n2611 = n1303 & n1597 ;
  assign n2612 = ~n2610 & n2611 ;
  assign n2613 = n2612 ^ n1597 ;
  assign n2614 = ~n1623 & n2613 ;
  assign n2615 = ~n2609 & n2614 ;
  assign n2616 = ~n1543 & ~n2615 ;
  assign n2617 = ~n1633 & ~n2616 ;
  assign n2618 = ~x70 & ~x95 ;
  assign n2619 = ~n1268 & n2618 ;
  assign n2620 = x32 & n1633 ;
  assign n2621 = n1637 & n2620 ;
  assign n2622 = n2621 ^ x32 ;
  assign n2623 = n2619 & ~n2622 ;
  assign n2624 = x32 & ~n2623 ;
  assign n2625 = n1220 & ~n1743 ;
  assign n2626 = ~n2624 & n2625 ;
  assign n2627 = ~n2617 & n2626 ;
  assign n2628 = n1785 ^ n1747 ;
  assign n2629 = ~n1799 & ~n2628 ;
  assign n2630 = ~x979 & ~x984 ;
  assign n2631 = ~x287 & n2630 ;
  assign n2632 = ~x252 & ~x1001 ;
  assign n2633 = x835 & ~n2632 ;
  assign n2634 = n2631 & n2633 ;
  assign n2635 = ~x332 & ~x468 ;
  assign n2636 = ~x299 & n2635 ;
  assign n2637 = n2636 ^ n2635 ;
  assign n2642 = x829 & x1092 ;
  assign n2643 = ~n1567 & n2642 ;
  assign n2638 = x824 & n1564 ;
  assign n2644 = ~n1569 & n2638 ;
  assign n2639 = ~x1093 & n2638 ;
  assign n2645 = n2644 ^ n2639 ;
  assign n2646 = ~n2643 & n2645 ;
  assign n2640 = ~n1576 & ~n2639 ;
  assign n2641 = n2640 ^ n1577 ;
  assign n2647 = n2646 ^ n2641 ;
  assign n2648 = ~n2637 & ~n2647 ;
  assign n2656 = ~x969 & ~x971 ;
  assign n2657 = ~x974 & ~x977 ;
  assign n2658 = n2656 & n2657 ;
  assign n2659 = ~x587 & ~x602 ;
  assign n2660 = ~x961 & ~x967 ;
  assign n2661 = n2659 & n2660 ;
  assign n2662 = n2658 & n2661 ;
  assign n2649 = ~x614 & ~x616 ;
  assign n2650 = ~x642 & n2649 ;
  assign n2651 = x603 & n2650 ;
  assign n2652 = ~x661 & ~x662 ;
  assign n2653 = ~x681 & n2652 ;
  assign n2654 = x680 & n2653 ;
  assign n2655 = ~n2651 & ~n2654 ;
  assign n2663 = n2662 ^ n2655 ;
  assign n2664 = ~n2635 & n2663 ;
  assign n2665 = n2664 ^ n2662 ;
  assign n2666 = n2648 & n2665 ;
  assign n2667 = n2666 ^ n2647 ;
  assign n2668 = n2634 & ~n2667 ;
  assign n2669 = n1535 ^ n1529 ;
  assign n2670 = n2668 & ~n2669 ;
  assign n2671 = ~x970 & ~x972 ;
  assign n2672 = ~x975 & ~x978 ;
  assign n2673 = n2671 & n2672 ;
  assign n2674 = ~x907 & ~x947 ;
  assign n2675 = ~x960 & ~x963 ;
  assign n2676 = n2674 & n2675 ;
  assign n2677 = n2673 & n2676 ;
  assign n2678 = n2637 & n2677 ;
  assign n2679 = n2670 & ~n2678 ;
  assign n2680 = ~x250 & n1562 ;
  assign n2681 = ~n2640 & n2680 ;
  assign n2682 = ~x41 & ~x101 ;
  assign n2683 = ~x99 & n2682 ;
  assign n2684 = ~x113 & n2683 ;
  assign n2685 = ~x43 & ~x44 ;
  assign n2686 = ~x42 & ~x114 ;
  assign n2687 = n2685 & n2686 ;
  assign n2688 = ~x115 & ~x116 ;
  assign n2689 = n2687 & n2688 ;
  assign n2690 = n2684 & n2689 ;
  assign n2691 = ~x52 & n2690 ;
  assign n2692 = x683 & ~n2691 ;
  assign n2700 = ~x129 & n2692 ;
  assign n2701 = x250 & n2700 ;
  assign n2702 = n2701 ^ x250 ;
  assign n2693 = n2692 ^ x252 ;
  assign n2694 = n2693 ^ x250 ;
  assign n2703 = n2702 ^ n2694 ;
  assign n2704 = n1562 & n2703 ;
  assign n2705 = n2704 ^ x252 ;
  assign n2706 = n2681 & n2705 ;
  assign n2707 = n2706 ^ n2705 ;
  assign n2708 = n2707 ^ n1755 ;
  assign n2713 = ~x87 & x100 ;
  assign n2714 = n2708 & n2713 ;
  assign n2715 = n2714 ^ n2708 ;
  assign n2716 = n2715 ^ n2707 ;
  assign n2717 = ~x74 & n2716 ;
  assign n2718 = x39 & ~n2717 ;
  assign n2719 = n1577 & n2634 ;
  assign n2721 = n2677 ^ n2655 ;
  assign n2722 = n2635 & n2721 ;
  assign n2723 = n2722 ^ n2655 ;
  assign n2724 = x299 & n1523 ;
  assign n2725 = ~x216 & n2724 ;
  assign n2726 = n2725 ^ n2724 ;
  assign n2727 = ~n2723 & n2726 ;
  assign n2720 = n1935 & ~n2665 ;
  assign n2728 = n2727 ^ n2720 ;
  assign n2729 = n2719 & n2728 ;
  assign n2730 = n2718 & ~n2729 ;
  assign n2731 = ~n2679 & n2730 ;
  assign n2732 = n2731 ^ n2718 ;
  assign n2733 = n2732 ^ n2717 ;
  assign n2734 = n2629 & ~n2733 ;
  assign n2735 = n2734 ^ n2628 ;
  assign n2736 = ~n2627 & ~n2735 ;
  assign n2737 = n1220 & n1508 ;
  assign n2746 = n1279 & n1298 ;
  assign n2747 = x90 & n1334 ;
  assign n2748 = x841 & n2747 ;
  assign n2749 = n2748 ^ n1334 ;
  assign n2750 = n2746 & n2749 ;
  assign n2745 = n1635 & ~n1637 ;
  assign n2751 = n2750 ^ n2745 ;
  assign n2738 = n1251 & n1373 ;
  assign n2739 = n1273 & n2738 ;
  assign n2740 = n1246 & n2739 ;
  assign n2741 = ~x73 & n1299 ;
  assign n2742 = n2740 & n2741 ;
  assign n2743 = ~x32 & n1292 ;
  assign n2744 = n2742 & n2743 ;
  assign n2752 = n2751 ^ n2744 ;
  assign n2753 = ~n1280 & ~n2752 ;
  assign n2754 = n1220 & n1298 ;
  assign n2755 = n1354 & n2754 ;
  assign n2756 = ~n2753 & n2755 ;
  assign n2757 = ~n2737 & ~n2756 ;
  assign n2768 = n1434 ^ n1221 ;
  assign n2771 = ~x67 & n2768 ;
  assign n2772 = n2771 ^ n1221 ;
  assign n2773 = n1225 & n2772 ;
  assign n2774 = n1406 & n2773 ;
  assign n2775 = ~x85 & n1460 ;
  assign n2776 = ~n1433 & n2775 ;
  assign n2777 = ~n2774 & n2776 ;
  assign n2778 = ~x82 & n2777 ;
  assign n2779 = ~n2607 & n2778 ;
  assign n2780 = ~x58 & n1328 ;
  assign n2781 = ~n2779 & n2780 ;
  assign n2761 = x103 & ~x109 ;
  assign n2762 = ~x314 & n2761 ;
  assign n2763 = n2762 ^ x109 ;
  assign n4836 = n1971 & n2763 ;
  assign n2758 = n1220 & n1503 ;
  assign n2759 = n1623 & n2758 ;
  assign n2760 = ~n1971 & ~n2759 ;
  assign n2785 = ~n4836 ^ n2760 ;
  assign n2786 = n2781 & n2785 ;
  assign n2787 = n2613 & n2786 ;
  assign n2788 = n2787 ^ n2613 ;
  assign n2766 = ~n4836 ^ n2613 ;
  assign n2789 = n2788 ^ n2766 ;
  assign n2790 = ~x72 & n2789 ;
  assign n2791 = ~n2757 & ~n2790 ;
  assign n2837 = x109 & x145 ;
  assign n2838 = x180 & x181 ;
  assign n2839 = n2837 & n2838 ;
  assign n2840 = x182 & x232 ;
  assign n2841 = n2839 & n2840 ;
  assign n2824 = x158 & x159 ;
  assign n2825 = x197 & n2824 ;
  assign n2826 = x160 & x232 ;
  assign n2827 = n2825 & n2826 ;
  assign n2842 = n2841 ^ n2827 ;
  assign n2843 = x299 & n2842 ;
  assign n2844 = n2843 ^ n2841 ;
  assign n2845 = n2635 & n2844 ;
  assign n2846 = ~x109 & n2843 ;
  assign n2847 = n2845 & n2846 ;
  assign n2848 = n2847 ^ n2845 ;
  assign n2849 = n2791 & ~n2848 ;
  assign n2850 = ~x228 & n2849 ;
  assign n2798 = ~x228 & n1743 ;
  assign n2799 = n2726 ^ n1935 ;
  assign n2800 = n2719 & n2799 ;
  assign n2801 = n2634 & n2646 ;
  assign n2802 = n2724 ^ n1530 ;
  assign n2803 = n1217 & n2802 ;
  assign n2804 = n2801 & n2803 ;
  assign n2805 = n2804 ^ n1217 ;
  assign n2806 = n2800 & n2805 ;
  assign n2808 = n2806 ^ n2804 ;
  assign n2809 = n2798 & n2808 ;
  assign n2810 = n2809 ^ x228 ;
  assign n2793 = ~x30 & x228 ;
  assign n2794 = ~n1209 & ~n2793 ;
  assign n2811 = n2794 ^ n2793 ;
  assign n2812 = ~n2810 & ~n2811 ;
  assign n2813 = n1749 & n1770 ;
  assign n2814 = n1210 & n2707 ;
  assign n2816 = n2813 & n2814 ;
  assign n2817 = n2816 ^ n1781 ;
  assign n2818 = n2812 & n2817 ;
  assign n2819 = n2818 ^ n2811 ;
  assign n2852 = n2850 ^ n2819 ;
  assign n2853 = ~n2636 & ~n2852 ;
  assign n2854 = n2853 ^ n2852 ;
  assign n2855 = x602 & ~n2854 ;
  assign n2792 = ~x228 & n2791 ;
  assign n2795 = ~x228 & n1781 ;
  assign n2796 = n2794 & n2795 ;
  assign n2797 = n2796 ^ n2794 ;
  assign n2820 = n2819 ^ n2797 ;
  assign n2821 = ~n2792 & n2820 ;
  assign n2834 = ~n2635 & n2654 ;
  assign n2822 = ~x299 & ~n2794 ;
  assign n2823 = x109 & ~x228 ;
  assign n2828 = n2635 & n2827 ;
  assign n2829 = n2823 & n2828 ;
  assign n2830 = n2829 ^ n2635 ;
  assign n2831 = n2822 & n2830 ;
  assign n2832 = n2831 ^ n2830 ;
  assign n2833 = x907 & n2832 ;
  assign n2835 = n2834 ^ n2833 ;
  assign n2836 = ~n2821 & n2835 ;
  assign n2857 = n2855 ^ n2836 ;
  assign n2858 = n2651 ^ x947 ;
  assign n2859 = ~n2635 & n2858 ;
  assign n2860 = n2859 ^ x947 ;
  assign n2868 = ~n2797 & ~n2853 ;
  assign n2861 = n2860 ^ x587 ;
  assign n2862 = n2861 ^ n2853 ;
  assign n2863 = n2862 ^ n2852 ;
  assign n2869 = n2868 ^ n2863 ;
  assign n2870 = n2860 & ~n2869 ;
  assign n2871 = n2870 ^ n2863 ;
  assign n2872 = n2871 ^ x587 ;
  assign n2873 = n2871 ^ n2860 ;
  assign n2874 = ~n2870 & n2873 ;
  assign n2875 = n2872 & n2874 ;
  assign n2876 = n2875 ^ n2871 ;
  assign n2879 = x967 & ~n2854 ;
  assign n2877 = ~n2821 & n2832 ;
  assign n2878 = x970 & n2877 ;
  assign n2881 = n2879 ^ n2878 ;
  assign n2883 = x299 & x972 ;
  assign n2887 = n2883 ^ n2827 ;
  assign n2882 = ~x299 & x961 ;
  assign n2888 = n2887 ^ n2882 ;
  assign n2889 = n2888 ^ x109 ;
  assign n2894 = n2887 ^ n2842 ;
  assign n2895 = ~n2889 & n2894 ;
  assign n2896 = n2895 ^ n2883 ;
  assign n2898 = n2882 & n2894 ;
  assign n2899 = n2898 ^ n2888 ;
  assign n2900 = n2883 & ~n2899 ;
  assign n2901 = n2896 & n2900 ;
  assign n2902 = n2901 ^ n2898 ;
  assign n2903 = n2902 ^ n2827 ;
  assign n2904 = n2903 ^ n2888 ;
  assign n2905 = n2792 & n2904 ;
  assign n2884 = n2883 ^ n2882 ;
  assign n2885 = ~n2819 & n2884 ;
  assign n2906 = n2905 ^ n2885 ;
  assign n2907 = n2635 & ~n2906 ;
  assign n2911 = n2907 ^ n2635 ;
  assign n2908 = n2797 & n2907 ;
  assign n2909 = n2885 ^ x972 ;
  assign n2910 = n2908 & n2909 ;
  assign n2912 = n2911 ^ n2910 ;
  assign n2914 = x960 & n2877 ;
  assign n2913 = x977 & ~n2854 ;
  assign n2916 = n2914 ^ n2913 ;
  assign n2918 = x963 & n2877 ;
  assign n2917 = x969 & ~n2854 ;
  assign n2920 = n2918 ^ n2917 ;
  assign n2922 = x971 & ~n2854 ;
  assign n2921 = x975 & n2877 ;
  assign n2924 = n2922 ^ n2921 ;
  assign n2926 = x974 & ~n2854 ;
  assign n2925 = x978 & n2877 ;
  assign n2928 = n2926 ^ n2925 ;
  assign n2929 = ~x96 & n1280 ;
  assign n2930 = ~x70 & n1277 ;
  assign n2931 = n2929 & n2930 ;
  assign n2932 = n1273 & n2931 ;
  assign n2933 = n1255 & n2932 ;
  assign n2934 = ~x92 & n1848 ;
  assign n2935 = n1209 & n2934 ;
  assign n2936 = n2933 & n2935 ;
  assign n2937 = ~x39 & ~x72 ;
  assign n2938 = n2937 ^ x72 ;
  assign n2939 = n2936 & ~n2938 ;
  assign n2940 = x51 & ~x87 ;
  assign n2941 = n2940 ^ x87 ;
  assign n2942 = n1258 & ~n2941 ;
  assign n2943 = n2939 & n2942 ;
  assign n2951 = n1209 & n1530 ;
  assign n2952 = ~n2665 & n2951 ;
  assign n2949 = n1523 & ~n1911 ;
  assign n2950 = ~n2723 & n2949 ;
  assign n2953 = n2952 ^ n2950 ;
  assign n2954 = n2801 & n2953 ;
  assign n2957 = ~n2729 & ~n2954 ;
  assign n2958 = n2943 & n2957 ;
  assign n2959 = n2958 ^ n2943 ;
  assign n2960 = n2959 ^ n2817 ;
  assign n2961 = ~n2849 & n2960 ;
  assign n2962 = n2961 ^ x24 ;
  assign n2963 = ~x954 & n2962 ;
  assign n2964 = n2963 ^ x24 ;
  assign n2966 = n1797 & n1882 ;
  assign n2967 = ~n1562 & n2966 ;
  assign n2968 = n2967 ^ n1797 ;
  assign n2969 = n2968 ^ n1972 ;
  assign n2970 = n2969 ^ x105 ;
  assign n2971 = ~x228 & ~n2970 ;
  assign n2972 = n2971 ^ x105 ;
  assign n2976 = x119 & ~x468 ;
  assign n2977 = ~x1056 & n2976 ;
  assign n2973 = ~x119 & ~x228 ;
  assign n2974 = x252 & ~x468 ;
  assign n2975 = n2973 & n2974 ;
  assign n2978 = n2977 ^ n2975 ;
  assign n2979 = ~x1077 & n2976 ;
  assign n2980 = n2979 ^ n2975 ;
  assign n2981 = ~x1073 & n2976 ;
  assign n2982 = n2981 ^ n2975 ;
  assign n2983 = ~x1041 & n2976 ;
  assign n2984 = n2983 ^ n2975 ;
  assign n2985 = x1092 & x1093 ;
  assign n2986 = ~x98 & x567 ;
  assign n2987 = n2985 & ~n2986 ;
  assign n2989 = x1161 & x1162 ;
  assign n2988 = x1162 ^ x1161 ;
  assign n2990 = n2989 ^ n2988 ;
  assign n2991 = ~x1163 & ~n2990 ;
  assign n2992 = ~n2987 & n2991 ;
  assign n2993 = n1209 & n2992 ;
  assign n2994 = x591 & ~x592 ;
  assign n3000 = x394 ^ x329 ;
  assign n3001 = n3000 ^ x328 ;
  assign n2998 = x399 ^ x398 ;
  assign n2996 = x408 ^ x400 ;
  assign n2995 = x396 ^ x395 ;
  assign n2997 = n2996 ^ n2995 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n3002 = n3001 ^ n2999 ;
  assign n3016 = x1198 & n3002 ;
  assign n3008 = x335 ^ x334 ;
  assign n3009 = n3008 ^ x333 ;
  assign n3006 = x463 ^ x413 ;
  assign n3004 = x407 ^ x393 ;
  assign n3003 = x392 ^ x391 ;
  assign n3005 = n3004 ^ n3003 ;
  assign n3007 = n3006 ^ n3005 ;
  assign n3010 = n3009 ^ n3007 ;
  assign n3017 = x1197 & n3010 ;
  assign n3018 = ~n3016 & n3017 ;
  assign n3019 = n3018 ^ n3016 ;
  assign n3020 = n2994 & n3019 ;
  assign n3021 = n3020 ^ x591 ;
  assign n3022 = ~x590 & ~x592 ;
  assign n3023 = x588 & n3022 ;
  assign n3038 = x428 ^ x427 ;
  assign n3039 = n3038 ^ x426 ;
  assign n3036 = x451 ^ x449 ;
  assign n3034 = x433 ^ x430 ;
  assign n3033 = x448 ^ x445 ;
  assign n3035 = n3034 ^ n3033 ;
  assign n3037 = n3036 ^ n3035 ;
  assign n3040 = n3039 ^ n3037 ;
  assign n3046 = x421 ^ x420 ;
  assign n3047 = n3046 ^ x419 ;
  assign n3044 = x459 ^ x454 ;
  assign n3042 = x432 ^ x425 ;
  assign n3041 = x424 ^ x423 ;
  assign n3043 = n3042 ^ n3041 ;
  assign n3045 = n3044 ^ n3043 ;
  assign n3048 = n3047 ^ n3045 ;
  assign n3061 = x1198 & n3048 ;
  assign n3062 = x1199 & ~n3061 ;
  assign n3063 = n3040 & n3062 ;
  assign n3054 = x417 ^ x416 ;
  assign n3055 = n3054 ^ x415 ;
  assign n3052 = x464 ^ x453 ;
  assign n3050 = x431 ^ x418 ;
  assign n3049 = x438 ^ x437 ;
  assign n3051 = n3050 ^ n3049 ;
  assign n3053 = n3052 ^ n3051 ;
  assign n3056 = n3055 ^ n3053 ;
  assign n3058 = n3056 ^ x1197 ;
  assign n3064 = n3063 ^ n3058 ;
  assign n3065 = n3063 ^ n3061 ;
  assign n3066 = n3056 & ~n3065 ;
  assign n3067 = ~n3064 & n3066 ;
  assign n3068 = n3067 ^ n3065 ;
  assign n3029 = x429 ^ x422 ;
  assign n3030 = n3029 ^ x414 ;
  assign n3027 = x443 ^ x436 ;
  assign n3025 = x446 ^ x444 ;
  assign n3024 = x435 ^ x434 ;
  assign n3026 = n3025 ^ n3024 ;
  assign n3028 = n3027 ^ n3026 ;
  assign n3031 = n3030 ^ n3028 ;
  assign n3032 = n3031 ^ x588 ;
  assign n3069 = n3068 ^ n3032 ;
  assign n3070 = n3068 ^ n3022 ;
  assign n3071 = x1196 & n3070 ;
  assign n3072 = ~n3069 & n3071 ;
  assign n3073 = n3072 ^ n3070 ;
  assign n3074 = n3023 & ~n3073 ;
  assign n3075 = n3074 ^ x588 ;
  assign n3076 = ~x591 & n3022 ;
  assign n3121 = x343 ^ x327 ;
  assign n3122 = n3121 ^ x323 ;
  assign n3119 = x450 ^ x362 ;
  assign n3117 = x358 ^ x346 ;
  assign n3116 = x345 ^ x344 ;
  assign n3118 = n3117 ^ n3116 ;
  assign n3120 = n3119 ^ n3118 ;
  assign n3123 = n3122 ^ n3120 ;
  assign n3082 = x321 ^ x316 ;
  assign n3083 = n3082 ^ x315 ;
  assign n3080 = x349 ^ x348 ;
  assign n3078 = x359 ^ x350 ;
  assign n3077 = x347 ^ x322 ;
  assign n3079 = n3078 ^ n3077 ;
  assign n3081 = n3080 ^ n3079 ;
  assign n3084 = n3083 ^ n3081 ;
  assign n3090 = x353 ^ x352 ;
  assign n3091 = n3090 ^ x351 ;
  assign n3088 = x462 ^ x461 ;
  assign n3086 = x360 ^ x357 ;
  assign n3085 = x356 ^ x354 ;
  assign n3087 = n3086 ^ n3085 ;
  assign n3089 = n3088 ^ n3087 ;
  assign n3092 = n3091 ^ n3089 ;
  assign n3105 = x1199 & n3092 ;
  assign n3106 = x1198 & ~n3105 ;
  assign n3107 = n3084 & n3106 ;
  assign n3098 = x355 ^ x342 ;
  assign n3099 = n3098 ^ x320 ;
  assign n3096 = x455 ^ x452 ;
  assign n3094 = x460 ^ x458 ;
  assign n3093 = x441 ^ x361 ;
  assign n3095 = n3094 ^ n3093 ;
  assign n3097 = n3096 ^ n3095 ;
  assign n3100 = n3099 ^ n3097 ;
  assign n3102 = n3100 ^ x1196 ;
  assign n3108 = n3107 ^ n3102 ;
  assign n3109 = ~x591 & ~x592 ;
  assign n3110 = n3107 ^ n3105 ;
  assign n3111 = n3109 & ~n3110 ;
  assign n3112 = n3100 & n3111 ;
  assign n3113 = ~n3108 & n3112 ;
  assign n3114 = n3113 ^ n3111 ;
  assign n3126 = x1197 & n3114 ;
  assign n3127 = n3123 & n3126 ;
  assign n3115 = n3114 ^ n3109 ;
  assign n3128 = n3127 ^ n3115 ;
  assign n3134 = x365 ^ x364 ;
  assign n3135 = n3134 ^ x336 ;
  assign n3132 = x447 ^ x389 ;
  assign n3130 = x383 ^ x368 ;
  assign n3129 = x367 ^ x366 ;
  assign n3131 = n3130 ^ n3129 ;
  assign n3133 = n3132 ^ n3131 ;
  assign n3136 = n3135 ^ n3133 ;
  assign n3151 = x371 ^ x370 ;
  assign n3152 = n3151 ^ x369 ;
  assign n3149 = x442 ^ x440 ;
  assign n3147 = x384 ^ x375 ;
  assign n3146 = x374 ^ x373 ;
  assign n3148 = n3147 ^ n3146 ;
  assign n3150 = n3149 ^ n3148 ;
  assign n3153 = n3152 ^ n3150 ;
  assign n3157 = x1198 & n3153 ;
  assign n3158 = x1197 & ~n3157 ;
  assign n3159 = n3136 & n3158 ;
  assign n3175 = n3159 ^ x1196 ;
  assign n3142 = x339 ^ x338 ;
  assign n3143 = n3142 ^ x337 ;
  assign n3140 = x388 ^ x387 ;
  assign n3138 = x372 ^ x363 ;
  assign n3137 = x386 ^ x380 ;
  assign n3139 = n3138 ^ n3137 ;
  assign n3141 = n3140 ^ n3139 ;
  assign n3144 = n3143 ^ n3141 ;
  assign n3160 = n3159 ^ n3157 ;
  assign n3166 = x377 ^ x376 ;
  assign n3167 = n3166 ^ x317 ;
  assign n3164 = x382 ^ x381 ;
  assign n3162 = x439 ^ x385 ;
  assign n3161 = x379 ^ x378 ;
  assign n3163 = n3162 ^ n3161 ;
  assign n3165 = n3164 ^ n3163 ;
  assign n3168 = n3167 ^ n3165 ;
  assign n3169 = ~x591 & x1199 ;
  assign n3170 = n3168 & n3169 ;
  assign n3171 = n3170 ^ x591 ;
  assign n3172 = ~n3160 & ~n3171 ;
  assign n3173 = ~x590 & n3172 ;
  assign n3176 = n3144 & n3173 ;
  assign n3177 = n3175 & n3176 ;
  assign n3174 = n3173 ^ x590 ;
  assign n3178 = n3177 ^ n3174 ;
  assign n3179 = ~n3128 & n3178 ;
  assign n3180 = ~n3076 & n3179 ;
  assign n3181 = n3180 ^ n3076 ;
  assign n3182 = ~n3075 & n3181 ;
  assign n3183 = n3182 ^ x588 ;
  assign n3184 = ~x217 & ~n3183 ;
  assign n3185 = ~x285 & ~x288 ;
  assign n3186 = ~x286 & ~x289 ;
  assign n3187 = n3185 & n3186 ;
  assign n3188 = n1278 & n1297 ;
  assign n3189 = ~x122 & x829 ;
  assign n3190 = ~x841 & n3189 ;
  assign n3191 = n1280 & n3190 ;
  assign n3192 = n3188 & n3191 ;
  assign n3193 = ~n2929 & ~n3192 ;
  assign n3196 = ~x35 & ~x70 ;
  assign n3197 = x90 ^ x51 ;
  assign n3198 = n3197 ^ x93 ;
  assign n3199 = x93 ^ x90 ;
  assign n3200 = x841 ^ x93 ;
  assign n3203 = n3199 & ~n3200 ;
  assign n3204 = n3203 ^ x90 ;
  assign n3205 = n3198 & ~n3204 ;
  assign n3206 = n3196 & n3205 ;
  assign n3207 = n1274 & n3206 ;
  assign n3194 = n1297 & n1502 ;
  assign n3195 = x98 & n3194 ;
  assign n3209 = n3207 ^ n3195 ;
  assign n3210 = ~x96 & ~n3209 ;
  assign n3211 = ~n2647 & ~n3210 ;
  assign n3212 = ~x122 & n1577 ;
  assign n3213 = ~x72 & n1297 ;
  assign n3214 = n1277 & n3213 ;
  assign n3215 = n3212 & n3214 ;
  assign n3216 = x91 & n1608 ;
  assign n3217 = ~x24 & ~x58 ;
  assign n3218 = n3216 & n3217 ;
  assign n3219 = n3218 ^ n1580 ;
  assign n3220 = n3215 & n3219 ;
  assign n3221 = ~x72 & n2640 ;
  assign n3229 = ~x98 & n3221 ;
  assign n3230 = x1091 & n3229 ;
  assign n3231 = n3230 ^ x1091 ;
  assign n3222 = n3221 ^ x72 ;
  assign n3223 = n3222 ^ x1091 ;
  assign n3232 = n3231 ^ n3223 ;
  assign n3233 = ~n3220 & ~n3232 ;
  assign n3234 = n3211 & n3233 ;
  assign n3235 = n3234 ^ n3220 ;
  assign n3236 = ~n3193 & n3235 ;
  assign n3237 = n2929 & n2937 ;
  assign n3238 = ~x87 & n3209 ;
  assign n3239 = n3237 & n3238 ;
  assign n3240 = n3239 ^ x87 ;
  assign n3241 = ~n2647 & n3240 ;
  assign n3242 = x100 ^ x39 ;
  assign n3243 = ~x75 & ~n3242 ;
  assign n3244 = ~n3241 & n3243 ;
  assign n3245 = ~n3236 & n3244 ;
  assign n3246 = ~x24 & ~x100 ;
  assign n3247 = ~x87 & n3246 ;
  assign n3248 = n3212 & n3247 ;
  assign n3249 = x232 & n2635 ;
  assign n3250 = ~n2691 & n3249 ;
  assign n3251 = n1561 & n3250 ;
  assign n3252 = n3251 ^ n2691 ;
  assign n3253 = x252 & n3252 ;
  assign n3254 = n3253 ^ x252 ;
  assign n3255 = n3248 & n3254 ;
  assign n3256 = n1743 & n3255 ;
  assign n3257 = x75 & ~n3256 ;
  assign n3258 = ~x39 & ~x100 ;
  assign n3259 = n1215 & n3258 ;
  assign n3260 = n1743 & n3259 ;
  assign n3261 = ~n3257 & n3260 ;
  assign n3262 = n2725 ^ n1531 ;
  assign n3264 = n1537 & ~n2723 ;
  assign n3263 = n1533 & ~n2665 ;
  assign n3266 = n3264 ^ n3263 ;
  assign n3267 = n3262 & n3266 ;
  assign n3268 = n2719 & n3267 ;
  assign n3269 = x39 & ~n3268 ;
  assign n3270 = ~x87 & ~x92 ;
  assign n3271 = n1787 & n3270 ;
  assign n3272 = n3212 & ~n3252 ;
  assign n3273 = x100 & x228 ;
  assign n3274 = n3272 & n3273 ;
  assign n3275 = n3274 ^ x100 ;
  assign n3276 = n3271 & ~n3275 ;
  assign n3277 = ~n3269 & n3276 ;
  assign n3278 = n1743 & n3277 ;
  assign n3279 = ~n1218 & ~n3278 ;
  assign n3280 = ~n3261 & n3279 ;
  assign n3281 = ~n3245 & ~n3280 ;
  assign n3282 = n1567 & n3281 ;
  assign n3288 = x326 ^ x325 ;
  assign n3289 = n3288 ^ x318 ;
  assign n3286 = x405 ^ x403 ;
  assign n3284 = x409 ^ x406 ;
  assign n3283 = x402 ^ x401 ;
  assign n3285 = n3284 ^ n3283 ;
  assign n3287 = n3286 ^ n3285 ;
  assign n3290 = n3289 ^ n3287 ;
  assign n3304 = x1199 & n3290 ;
  assign n3296 = x390 ^ x324 ;
  assign n3297 = n3296 ^ x319 ;
  assign n3294 = x456 ^ x412 ;
  assign n3292 = x404 ^ x397 ;
  assign n3291 = x411 ^ x410 ;
  assign n3293 = n3292 ^ n3291 ;
  assign n3295 = n3294 ^ n3293 ;
  assign n3298 = n3297 ^ n3295 ;
  assign n3305 = x1196 & n3298 ;
  assign n3306 = ~n3304 & n3305 ;
  assign n3307 = n3306 ^ n3304 ;
  assign n3308 = n3022 & n3307 ;
  assign n3309 = n3021 & n3184 ;
  assign n3310 = x567 & n3309 ;
  assign n3311 = n3308 & n3310 ;
  assign n3312 = n3311 ^ n3309 ;
  assign n3313 = n3312 ^ n3184 ;
  assign n3314 = n3282 & n3313 ;
  assign n3315 = n3314 ^ n3281 ;
  assign n3316 = ~n3187 & ~n3315 ;
  assign n3317 = n3184 & n3316 ;
  assign n3318 = ~n3021 & n3317 ;
  assign n3319 = n3318 ^ n3316 ;
  assign n3320 = n3319 ^ n3315 ;
  assign n3321 = n2993 & n3320 ;
  assign n3380 = n3261 ^ n1212 ;
  assign n3375 = n2647 ^ x98 ;
  assign n3322 = n1567 & n2638 ;
  assign n3323 = ~x122 & n3322 ;
  assign n3325 = n3323 ^ x98 ;
  assign n3376 = n3375 ^ n3325 ;
  assign n3378 = n3376 ^ n3261 ;
  assign n3381 = n3380 ^ n3376 ;
  assign n3357 = x98 & ~n3325 ;
  assign n3358 = n3381 ^ n3357 ;
  assign n3359 = n3378 ^ n3358 ;
  assign n3360 = n3359 ^ n3323 ;
  assign n3379 = n3378 ^ n3325 ;
  assign n3384 = n3381 ^ n3379 ;
  assign n3385 = n3384 ^ n3375 ;
  assign n3362 = n3385 ^ n3323 ;
  assign n3363 = ~n3360 & ~n3362 ;
  assign n3386 = n3385 ^ x98 ;
  assign n3382 = n3381 ^ n3325 ;
  assign n3346 = n3382 ^ n3376 ;
  assign n3348 = n3378 ^ n3346 ;
  assign n3366 = n3381 ^ n3348 ;
  assign n3367 = n3386 ^ n3366 ;
  assign n3368 = ~n2647 & n3367 ;
  assign n3369 = n3363 & n3368 ;
  assign n3370 = n3369 ^ n3357 ;
  assign n3371 = n3380 ^ n3370 ;
  assign n3388 = n3371 ^ n2647 ;
  assign n3389 = n3388 ^ x98 ;
  assign n3335 = n3382 ^ n3323 ;
  assign n3390 = n3389 ^ n3335 ;
  assign n3394 = x567 & n2640 ;
  assign n3395 = ~x1199 & ~n3394 ;
  assign n3396 = ~x217 & ~x588 ;
  assign n3397 = x591 & ~x1091 ;
  assign n3398 = n3396 & n3397 ;
  assign n3399 = ~n3395 & n3398 ;
  assign n3400 = ~n3019 & n3399 ;
  assign n3401 = n3308 & n3400 ;
  assign n3415 = n3394 & n3401 ;
  assign n3402 = n3237 & n3322 ;
  assign n3403 = n3402 ^ n3242 ;
  assign n3406 = n3207 & n3403 ;
  assign n3407 = n3406 ^ n3242 ;
  assign n3408 = ~n3401 & n3407 ;
  assign n3409 = ~n3236 & n3408 ;
  assign n3391 = n3390 ^ n3279 ;
  assign n3392 = n3391 ^ n3236 ;
  assign n3410 = n3409 ^ n3392 ;
  assign n3416 = n3415 ^ n3410 ;
  assign n3417 = n3390 & ~n3416 ;
  assign n3418 = n3417 ^ n3410 ;
  assign n3419 = n3418 ^ n3279 ;
  assign n3420 = n3418 ^ n3390 ;
  assign n3421 = ~n3417 & n3420 ;
  assign n3422 = ~n3419 & n3421 ;
  assign n3423 = n3422 ^ n3418 ;
  assign n3424 = n3321 & n3423 ;
  assign n3430 = ~x31 & n2985 ;
  assign n3431 = n2989 & n3430 ;
  assign n3425 = ~n3187 & n3323 ;
  assign n3426 = ~n1209 & n3425 ;
  assign n3427 = n2986 & n3426 ;
  assign n3428 = ~n2990 & ~n3313 ;
  assign n3429 = n3427 & n3428 ;
  assign n3432 = n3431 ^ n3429 ;
  assign n3433 = ~x1163 & n3432 ;
  assign n3434 = ~n3424 & ~n3433 ;
  assign n3435 = x76 & ~n1478 ;
  assign n3436 = ~n1571 & ~n3187 ;
  assign n3437 = ~x137 & ~n1551 ;
  assign n3438 = ~x50 & n3437 ;
  assign n3439 = ~n3436 & n3438 ;
  assign n3440 = n3435 & n3439 ;
  assign n3441 = x32 & ~x841 ;
  assign n3446 = ~x24 & n3441 ;
  assign n3447 = n3446 ^ x32 ;
  assign n3448 = ~n1636 & n3447 ;
  assign n3449 = ~x24 & n1259 ;
  assign n3450 = x50 & n3449 ;
  assign n3451 = ~n3448 & n3450 ;
  assign n3452 = n3451 ^ n3448 ;
  assign n3453 = ~n3440 & ~n3452 ;
  assign n3454 = n1971 & ~n3453 ;
  assign n3461 = x75 & n3246 ;
  assign n3462 = n1571 & n3461 ;
  assign n3463 = n3462 ^ n3461 ;
  assign n3464 = ~n3253 & n3463 ;
  assign n3455 = ~x252 & ~n1562 ;
  assign n3456 = n2640 ^ x129 ;
  assign n3457 = n2680 & n3456 ;
  assign n3458 = n3457 ^ x129 ;
  assign n3459 = n1210 & n3458 ;
  assign n3460 = ~n3455 & n3459 ;
  assign n3465 = n3464 ^ n3460 ;
  assign n3466 = ~x137 & ~n3252 ;
  assign n3474 = ~n1562 & n3466 ;
  assign n3475 = n3463 & n3474 ;
  assign n3476 = n3475 ^ n3463 ;
  assign n3467 = n3466 ^ x137 ;
  assign n3468 = n3467 ^ n3463 ;
  assign n3477 = n3476 ^ n3468 ;
  assign n3478 = n3465 & ~n3477 ;
  assign n3479 = n2813 & n3478 ;
  assign n3480 = ~n3454 & ~n3479 ;
  assign n3481 = x73 & n2740 ;
  assign n3482 = n1279 & n1299 ;
  assign n3483 = n3481 & n3482 ;
  assign n3486 = n1354 & n2752 ;
  assign n3484 = ~x70 & n1304 ;
  assign n3485 = n1508 & ~n3484 ;
  assign n3488 = n3486 ^ n3485 ;
  assign n3489 = ~n3483 & ~n3488 ;
  assign n3490 = ~x63 & ~x107 ;
  assign n3491 = ~x40 & n3490 ;
  assign n3501 = x954 ^ x33 ;
  assign n3492 = ~x79 & ~x118 ;
  assign n3493 = ~x33 & ~x34 ;
  assign n3494 = n3492 & n3493 ;
  assign n3495 = ~x954 & n3494 ;
  assign n3496 = ~x138 & x139 ;
  assign n3497 = n3496 ^ x138 ;
  assign n3498 = n3495 & ~n3497 ;
  assign n3499 = ~x196 & n3498 ;
  assign n3500 = ~x195 & n3499 ;
  assign n3502 = n3501 ^ n3500 ;
  assign n3503 = n3491 & n3502 ;
  assign n3504 = x186 ^ x164 ;
  assign n3505 = ~x299 & n3504 ;
  assign n3506 = n3505 ^ x164 ;
  assign n3507 = ~n1213 & n3249 ;
  assign n3508 = n3506 & n3507 ;
  assign n3509 = n3508 ^ n1213 ;
  assign n3510 = n1758 & n3509 ;
  assign n3511 = n3503 & n3510 ;
  assign n3512 = n3489 & n3511 ;
  assign n3528 = n1279 & n2742 ;
  assign n3529 = n1754 & n3528 ;
  assign n3534 = x176 ^ x154 ;
  assign n3537 = x299 & n3534 ;
  assign n3538 = n3537 ^ x176 ;
  assign n3539 = n3249 & n3538 ;
  assign n3544 = n3491 & n3539 ;
  assign n3545 = x92 & n3544 ;
  assign n3546 = n3545 ^ x92 ;
  assign n3530 = ~x39 & n3270 ;
  assign n3531 = n3503 & ~n3530 ;
  assign n3532 = n3531 ^ x92 ;
  assign n3547 = n3546 ^ n3532 ;
  assign n3548 = n3529 & n3547 ;
  assign n3549 = n3548 ^ n3531 ;
  assign n3550 = n3237 & n3270 ;
  assign n3551 = n3188 & n3550 ;
  assign n3552 = x38 & ~n3551 ;
  assign n3553 = ~x54 & ~n3552 ;
  assign n3554 = n3549 & n3553 ;
  assign n3558 = n2801 ^ n2719 ;
  assign n3559 = n2728 & n3558 ;
  assign n3560 = n3528 & n3559 ;
  assign n3561 = n3270 & n3560 ;
  assign n3564 = x39 & n3249 ;
  assign n3567 = ~n2677 & n2726 ;
  assign n3568 = ~x152 & n3567 ;
  assign n3565 = n1935 & ~n2662 ;
  assign n3566 = ~x174 & n3565 ;
  assign n3569 = n3568 ^ n3566 ;
  assign n3570 = n2801 & n3569 ;
  assign n3576 = n3570 ^ n3564 ;
  assign n3572 = x154 & n3567 ;
  assign n3571 = x176 & n3565 ;
  assign n3573 = n3572 ^ n3571 ;
  assign n3574 = n2719 & n3573 ;
  assign n3577 = n3576 ^ n3574 ;
  assign n3578 = n3564 & ~n3577 ;
  assign n3579 = n3564 ^ n3249 ;
  assign n3580 = n3579 ^ n1743 ;
  assign n3581 = n3578 & n3580 ;
  assign n3582 = n3581 ^ n3579 ;
  assign n3585 = n3561 & ~n3582 ;
  assign n3586 = n3554 & n3585 ;
  assign n3587 = n3586 ^ n3554 ;
  assign n3588 = n3587 ^ n3553 ;
  assign n3589 = n3509 & ~n3588 ;
  assign n3521 = x191 ^ x169 ;
  assign n3524 = x299 & n3521 ;
  assign n3525 = n3524 ^ x191 ;
  assign n3526 = n3249 & n3525 ;
  assign n3590 = n3589 ^ n3526 ;
  assign n3591 = ~x74 & n3590 ;
  assign n3514 = x183 ^ x178 ;
  assign n3513 = x157 ^ x149 ;
  assign n3515 = n3514 ^ n3513 ;
  assign n3518 = ~x299 & n3515 ;
  assign n3519 = n3518 ^ n3513 ;
  assign n3520 = n3249 & n3519 ;
  assign n3527 = n3526 ^ n3520 ;
  assign n3592 = n3591 ^ n3527 ;
  assign n3593 = ~n1211 & ~n3592 ;
  assign n3594 = n3593 ^ n3520 ;
  assign n3595 = n1209 & n3594 ;
  assign n3596 = ~n3512 & n3595 ;
  assign n3597 = n1216 & n3582 ;
  assign n3598 = ~x39 & n1520 ;
  assign n3599 = n1354 & n2750 ;
  assign n3635 = x193 ^ x172 ;
  assign n3638 = ~x299 & n3635 ;
  assign n3639 = n3638 ^ x172 ;
  assign n3640 = n3599 & n3639 ;
  assign n3600 = n1292 & n1300 ;
  assign n3601 = x180 ^ x158 ;
  assign n3602 = ~x299 & n3601 ;
  assign n3603 = n3602 ^ x158 ;
  assign n3604 = ~x198 & ~x299 ;
  assign n3605 = ~x841 & ~n1634 ;
  assign n3606 = n3604 & n3605 ;
  assign n3607 = n2742 & n3606 ;
  assign n3608 = ~x299 & ~n3484 ;
  assign n3609 = ~n3607 & ~n3608 ;
  assign n3610 = x183 & ~n3609 ;
  assign n3616 = ~x210 & n3441 ;
  assign n3617 = n3484 & n3616 ;
  assign n3618 = n3617 ^ n3484 ;
  assign n3623 = x149 & ~n3618 ;
  assign n3624 = x299 & n3623 ;
  assign n3625 = n3624 ^ x299 ;
  assign n3611 = x174 ^ x152 ;
  assign n3612 = ~x299 & n3611 ;
  assign n3613 = n3612 ^ x152 ;
  assign n3614 = n3613 ^ x299 ;
  assign n3626 = n3625 ^ n3614 ;
  assign n3627 = ~x73 & ~n3626 ;
  assign n3628 = n3627 ^ n3613 ;
  assign n3629 = n3610 & n3628 ;
  assign n3630 = n3629 ^ n3628 ;
  assign n3631 = n3603 & n3630 ;
  assign n3632 = n3600 & n3631 ;
  assign n3633 = n3632 ^ n3630 ;
  assign n3641 = n3640 ^ n3633 ;
  assign n3642 = n3598 & ~n3641 ;
  assign n3643 = n3642 ^ x39 ;
  assign n3644 = n3597 & n3643 ;
  assign n3645 = n3596 & ~n3644 ;
  assign n3648 = ~n1208 & n1213 ;
  assign n3653 = x164 & ~n3648 ;
  assign n3654 = n3653 ^ x169 ;
  assign n3655 = ~x74 & n3654 ;
  assign n3646 = n3513 ^ x169 ;
  assign n3656 = n3655 ^ n3646 ;
  assign n3657 = ~n1211 & n3656 ;
  assign n3658 = n3657 ^ n3513 ;
  assign n3659 = n3249 & n3658 ;
  assign n3660 = n3659 ^ n1211 ;
  assign n3661 = ~n1209 & ~n3660 ;
  assign n3662 = n1846 & ~n3648 ;
  assign n3663 = n3662 ^ n1846 ;
  assign n3664 = n3491 & n3663 ;
  assign n3667 = x149 & n3249 ;
  assign n3668 = n3667 ^ n3502 ;
  assign n3669 = n1745 & n3668 ;
  assign n3670 = n3669 ^ n3502 ;
  assign n3671 = n3664 & n3670 ;
  assign n3672 = n3661 & ~n3671 ;
  assign n3673 = ~n3645 & ~n3672 ;
  assign n3674 = ~x33 & ~x954 ;
  assign n3675 = n3674 ^ x34 ;
  assign n3676 = n3675 ^ n3500 ;
  assign n3678 = n1205 & n3530 ;
  assign n3679 = n3528 & n3678 ;
  assign n3680 = ~n1206 & ~n3679 ;
  assign n3677 = n1220 & n3489 ;
  assign n3681 = n3680 ^ n3677 ;
  assign n3682 = ~n3676 & n3681 ;
  assign n3683 = n1206 & ~n1218 ;
  assign n3684 = n2646 & n3249 ;
  assign n3686 = ~x161 & n3567 ;
  assign n3685 = ~x144 & n3565 ;
  assign n3687 = n3686 ^ n3685 ;
  assign n3688 = n3684 & n3687 ;
  assign n3689 = n3688 ^ n3249 ;
  assign n3691 = x155 & n3567 ;
  assign n3690 = x177 & n3565 ;
  assign n3692 = n3691 ^ n3690 ;
  assign n3693 = n1577 & n3692 ;
  assign n3694 = n3689 & n3693 ;
  assign n3696 = n3694 ^ n3688 ;
  assign n3697 = n3561 & ~n3696 ;
  assign n3698 = n3683 & ~n3697 ;
  assign n3699 = x39 & n3561 ;
  assign n3700 = x92 & n3529 ;
  assign n3701 = x177 ^ x155 ;
  assign n3702 = ~x299 & n3701 ;
  assign n3703 = n3702 ^ x155 ;
  assign n3708 = n3249 & n3703 ;
  assign n3709 = n3708 ^ n3676 ;
  assign n3710 = n3700 & ~n3709 ;
  assign n3711 = n3710 ^ n3676 ;
  assign n3712 = n3699 & n3711 ;
  assign n3713 = n3712 ^ n3711 ;
  assign n3714 = n3698 & ~n3713 ;
  assign n3715 = ~n3682 & ~n3714 ;
  assign n3716 = n3664 & ~n3715 ;
  assign n3729 = x162 & x299 ;
  assign n3717 = x181 ^ x159 ;
  assign n3718 = ~x299 & n3717 ;
  assign n3719 = n3718 ^ x159 ;
  assign n3720 = n2743 & n3719 ;
  assign n3721 = x73 & ~n3720 ;
  assign n3722 = x161 ^ x144 ;
  assign n3725 = ~x299 & n3722 ;
  assign n3726 = n3725 ^ x161 ;
  assign n3727 = n3721 & ~n3726 ;
  assign n3728 = n3727 ^ n3720 ;
  assign n3730 = ~n3618 & ~n3728 ;
  assign n3731 = n3729 & n3730 ;
  assign n3732 = n3731 ^ n3728 ;
  assign n3733 = ~n1554 & ~n3732 ;
  assign n3734 = n3599 & n3733 ;
  assign n3735 = n3734 ^ x140 ;
  assign n3736 = n3734 ^ n3732 ;
  assign n3737 = n1971 & ~n3736 ;
  assign n3738 = ~n3609 & n3737 ;
  assign n3739 = n3735 & n3738 ;
  assign n3740 = n3739 ^ n3737 ;
  assign n3741 = n3740 ^ n1971 ;
  assign n3770 = x145 ^ x140 ;
  assign n3768 = ~x178 & ~x183 ;
  assign n3766 = x197 ^ x162 ;
  assign n3765 = ~x149 & ~x157 ;
  assign n3767 = n3766 ^ n3765 ;
  assign n3769 = n3768 ^ n3767 ;
  assign n3771 = n3770 ^ n3769 ;
  assign n3772 = n1911 & n3771 ;
  assign n3773 = n3772 ^ n3767 ;
  assign n3748 = x148 ^ x141 ;
  assign n3749 = x299 & n3748 ;
  assign n3750 = n3749 ^ x141 ;
  assign n3742 = x188 ^ x167 ;
  assign n3745 = x299 & n3742 ;
  assign n3746 = n3745 ^ x188 ;
  assign n3747 = ~n3553 & n3746 ;
  assign n3751 = n3750 ^ n3747 ;
  assign n3752 = ~x74 & n3751 ;
  assign n3753 = n3752 ^ n3750 ;
  assign n3774 = n3773 ^ n3753 ;
  assign n3760 = x167 & ~n3648 ;
  assign n3761 = n3760 ^ x148 ;
  assign n3762 = ~x74 & n3761 ;
  assign n3754 = n3753 ^ x148 ;
  assign n3763 = n3762 ^ n3754 ;
  assign n3764 = ~n1209 & n3763 ;
  assign n3775 = n3774 ^ n3764 ;
  assign n3776 = ~n1211 & ~n3775 ;
  assign n3777 = n3776 ^ n3773 ;
  assign n3778 = n3249 & n3777 ;
  assign n3779 = ~n3741 & n3778 ;
  assign n3783 = n3779 ^ n3249 ;
  assign n3780 = n1819 & n3679 ;
  assign n3781 = x162 & n3780 ;
  assign n3782 = n3779 & n3781 ;
  assign n3784 = n3783 ^ n3782 ;
  assign n3785 = ~n3716 & ~n3784 ;
  assign n3786 = ~x55 & ~x74 ;
  assign n3787 = x24 & ~x59 ;
  assign n3788 = n3787 ^ x24 ;
  assign n3789 = n3786 & ~n3788 ;
  assign n3790 = n1763 & n3789 ;
  assign n3795 = x683 & n2644 ;
  assign n3796 = n3795 ^ x137 ;
  assign n3797 = ~n3252 & n3796 ;
  assign n3798 = n3797 ^ x137 ;
  assign n3799 = x252 & n3798 ;
  assign n3800 = n3799 ^ x252 ;
  assign n3801 = n1562 & ~n2691 ;
  assign n3802 = n1213 & ~n3801 ;
  assign n3803 = n3459 & n3802 ;
  assign n3804 = ~n3800 & n3803 ;
  assign n3829 = ~x137 & n1562 ;
  assign n3805 = x75 ^ x38 ;
  assign n3809 = n3805 ^ n3253 ;
  assign n3810 = ~n3801 & n3809 ;
  assign n3818 = x137 & n3810 ;
  assign n3819 = ~n1571 & n3818 ;
  assign n3820 = n3819 ^ n1571 ;
  assign n3811 = n3810 ^ n3801 ;
  assign n3812 = n3811 ^ n1571 ;
  assign n3821 = n3820 ^ n3812 ;
  assign n3822 = x75 & n3821 ;
  assign n3823 = n3805 & n3822 ;
  assign n3806 = n3804 ^ n3246 ;
  assign n3807 = n3806 ^ n3805 ;
  assign n3824 = n3823 ^ n3807 ;
  assign n3830 = n3829 ^ n3824 ;
  assign n3831 = n3804 & n3830 ;
  assign n3832 = n3831 ^ n3824 ;
  assign n3833 = n3832 ^ n3804 ;
  assign n3835 = n3832 ^ n3246 ;
  assign n3836 = ~n3831 & ~n3835 ;
  assign n3837 = ~n3833 & n3836 ;
  assign n3838 = n3837 ^ n3833 ;
  assign n3839 = n3838 ^ n3804 ;
  assign n3840 = n3551 & ~n3839 ;
  assign n3841 = n3840 ^ n1757 ;
  assign n3791 = n1758 & ~n3551 ;
  assign n3792 = ~n3648 & n3791 ;
  assign n3842 = n3841 ^ n3792 ;
  assign n3843 = x40 & x1082 ;
  assign n3844 = n1520 & ~n3843 ;
  assign n3846 = ~x122 & n2640 ;
  assign n3847 = ~n3436 & n3846 ;
  assign n3848 = ~n3437 & n3847 ;
  assign n3849 = x76 & n3848 ;
  assign n3850 = n3849 ^ n1608 ;
  assign n3851 = n2781 & n3850 ;
  assign n3852 = n3200 & n3851 ;
  assign n3853 = n1302 & n3852 ;
  assign n3854 = n3853 ^ n3851 ;
  assign n3855 = n3854 ^ n3850 ;
  assign n3856 = n3844 & ~n3855 ;
  assign n3857 = n3856 ^ n1520 ;
  assign n3858 = ~n3787 & ~n3857 ;
  assign n3866 = ~n2745 & n3858 ;
  assign n3867 = n1761 & n3866 ;
  assign n3868 = n3867 ^ n1761 ;
  assign n3859 = n3858 ^ n3857 ;
  assign n3860 = n3859 ^ n1761 ;
  assign n3869 = n3868 ^ n3860 ;
  assign n3870 = n3842 & n3869 ;
  assign n3871 = n3870 ^ n3840 ;
  assign n3872 = n3790 & n3871 ;
  assign n3873 = x36 & n1273 ;
  assign n3874 = ~n1478 & n3873 ;
  assign n3875 = ~n3218 & ~n3874 ;
  assign n3876 = n1277 & n2758 ;
  assign n3877 = ~n3875 & n3876 ;
  assign n3878 = ~n2640 & n3877 ;
  assign n3879 = ~x70 & ~x89 ;
  assign n3880 = x332 & n3879 ;
  assign n3881 = n3880 ^ x332 ;
  assign n3882 = n1273 & n3876 ;
  assign n3883 = ~n1478 & n3882 ;
  assign n3884 = x841 & n3883 ;
  assign n3885 = n3884 ^ n3883 ;
  assign n3894 = n3881 & n3885 ;
  assign n3886 = n1385 & n3882 ;
  assign n3887 = x64 & n3886 ;
  assign n3888 = x841 & n3887 ;
  assign n3889 = n3888 ^ n3887 ;
  assign n3890 = ~x24 & n1753 ;
  assign n3891 = n3890 ^ n1753 ;
  assign n3892 = ~n3889 & ~n3891 ;
  assign n3895 = n3894 ^ n3892 ;
  assign n3896 = ~x35 & ~x48 ;
  assign n3897 = x108 & x314 ;
  assign n3898 = x252 & ~x986 ;
  assign n3899 = n2640 & n3898 ;
  assign n3900 = n3899 ^ x252 ;
  assign n3901 = n3897 & ~n3900 ;
  assign n3906 = ~x47 & ~n3901 ;
  assign n3907 = n3906 ^ x841 ;
  assign n3908 = n3896 & n3907 ;
  assign n3909 = n3908 ^ x841 ;
  assign n3910 = n2737 & ~n3909 ;
  assign n3911 = n1635 & n1636 ;
  assign n3912 = n1220 & n3911 ;
  assign n3913 = x287 & n2942 ;
  assign n3914 = n2939 & n3913 ;
  assign n3915 = n3914 ^ n2943 ;
  assign n3916 = x835 & x984 ;
  assign n3917 = ~x979 & n3916 ;
  assign n3918 = n3917 ^ x979 ;
  assign n3919 = n2632 & ~n3918 ;
  assign n3920 = n3919 ^ n3918 ;
  assign n3921 = x835 & ~n2678 ;
  assign n3922 = ~n2667 & n3921 ;
  assign n3927 = ~x1093 & ~n2670 ;
  assign n3923 = x786 & ~x1082 ;
  assign n3924 = ~n3920 & n3923 ;
  assign n3928 = n3927 ^ n3924 ;
  assign n3929 = n3922 & ~n3928 ;
  assign n3930 = n3929 ^ n3924 ;
  assign n3931 = ~n3920 & ~n3930 ;
  assign n3932 = n3915 & n3931 ;
  assign n3933 = ~n3912 & ~n3932 ;
  assign n3934 = ~n3910 & n3933 ;
  assign n3935 = x102 ^ x40 ;
  assign n3936 = ~n3843 & n3935 ;
  assign n3937 = n1971 & n3936 ;
  assign n3962 = n1210 & ~n3272 ;
  assign n3963 = n3962 ^ n1212 ;
  assign n3964 = x228 & n3963 ;
  assign n3965 = ~n3220 & n3964 ;
  assign n3966 = ~n1296 & ~n1571 ;
  assign n3967 = ~n3210 & n3966 ;
  assign n3968 = n3967 ^ n3210 ;
  assign n3969 = n3965 & n3968 ;
  assign n3970 = x110 ^ x94 ;
  assign n3972 = ~x250 & x252 ;
  assign n3973 = x901 & ~x959 ;
  assign n3974 = n3972 & n3973 ;
  assign n3971 = ~x480 & x949 ;
  assign n3975 = n3974 ^ n3971 ;
  assign n3976 = x110 & n3975 ;
  assign n3977 = n3976 ^ n3974 ;
  assign n3978 = n3970 & n3977 ;
  assign n3979 = ~n3194 & n3978 ;
  assign n3980 = x87 & x100 ;
  assign n3981 = n3980 ^ n1792 ;
  assign n3982 = ~n1743 & n3981 ;
  assign n3983 = ~x228 & ~n3978 ;
  assign n3984 = n1215 & ~n3980 ;
  assign n3985 = n1209 & n3984 ;
  assign n3986 = ~n3983 & n3985 ;
  assign n3987 = ~n3982 & n3986 ;
  assign n3988 = ~n3257 & n3987 ;
  assign n3989 = ~n3193 & n3988 ;
  assign n3990 = ~n3979 & n3989 ;
  assign n3991 = ~n3969 & n3990 ;
  assign n3992 = ~x44 & n3991 ;
  assign n3997 = ~x101 & n3992 ;
  assign n3998 = n3997 ^ x41 ;
  assign n3999 = n2937 & ~n3998 ;
  assign n3938 = n2936 & n3249 ;
  assign n3939 = n3913 & n3938 ;
  assign n3940 = n3939 ^ n3249 ;
  assign n3941 = ~n2938 & n3940 ;
  assign n3944 = n1558 & ~n1911 ;
  assign n3945 = n3944 ^ n3940 ;
  assign n3942 = ~x166 & ~n1911 ;
  assign n3946 = n3945 ^ n3942 ;
  assign n3943 = x152 & n3942 ;
  assign n3947 = n3946 ^ n3943 ;
  assign n3948 = n3941 & n3947 ;
  assign n3951 = n1556 & n1911 ;
  assign n3949 = ~x189 & n1911 ;
  assign n3952 = n3951 ^ n3949 ;
  assign n3950 = x174 & n3949 ;
  assign n3953 = n3952 ^ n3950 ;
  assign n3954 = n3948 & ~n3953 ;
  assign n3955 = n3954 ^ n3941 ;
  assign n3956 = n3955 ^ n2938 ;
  assign n4000 = n3999 ^ n3956 ;
  assign n4001 = n2684 & n3992 ;
  assign n4002 = n2688 & n4001 ;
  assign n4003 = ~x114 & n4002 ;
  assign n4004 = n4003 ^ x42 ;
  assign n4042 = n2937 & n4004 ;
  assign n4005 = n3949 ^ n3940 ;
  assign n4006 = n3941 & ~n3942 ;
  assign n4007 = n4005 & n4006 ;
  assign n4008 = n4007 ^ n3941 ;
  assign n4009 = n4008 ^ n2938 ;
  assign n4036 = x219 ^ x199 ;
  assign n4037 = ~n1911 & n4036 ;
  assign n4038 = n4037 ^ x199 ;
  assign n4010 = ~x212 & ~x214 ;
  assign n4011 = n4010 ^ x212 ;
  assign n4012 = n4011 ^ x214 ;
  assign n4022 = x211 & ~x219 ;
  assign n4021 = x219 ^ x211 ;
  assign n4023 = n4022 ^ n4021 ;
  assign n4026 = ~n4012 & ~n4023 ;
  assign n4013 = x199 & ~x200 ;
  assign n4014 = x207 & ~x208 ;
  assign n4015 = n4014 ^ x207 ;
  assign n4016 = ~n4013 & n4015 ;
  assign n4017 = n4016 ^ x200 ;
  assign n4018 = n4017 ^ x211 ;
  assign n4027 = n4026 ^ n4018 ;
  assign n4028 = ~n1911 & n4027 ;
  assign n4029 = n4028 ^ n4017 ;
  assign n4033 = ~n1911 & ~n4022 ;
  assign n4030 = x200 ^ x199 ;
  assign n4031 = n4030 ^ n4013 ;
  assign n4032 = n1911 & ~n4031 ;
  assign n4034 = n4033 ^ n4032 ;
  assign n4035 = ~n4029 & ~n4034 ;
  assign n4039 = n4038 ^ n4035 ;
  assign n4040 = ~n4009 & n4039 ;
  assign n4043 = n4042 ^ n4040 ;
  assign n4050 = ~x42 & n4003 ;
  assign n4051 = n4050 ^ x43 ;
  assign n4052 = n2937 & n4051 ;
  assign n4044 = ~n4009 & n4029 ;
  assign n4053 = n4052 ^ n4044 ;
  assign n4054 = n3991 ^ x44 ;
  assign n4058 = n2937 & n4054 ;
  assign n4055 = n3951 ^ n3944 ;
  assign n4056 = n3941 & n4055 ;
  assign n4059 = n4058 ^ n4056 ;
  assign n4060 = x979 & n3915 ;
  assign n4062 = n1312 & n2758 ;
  assign n4063 = n1311 & n4062 ;
  assign n4064 = n1354 & n4063 ;
  assign n4065 = ~x24 & n4064 ;
  assign n4066 = n4065 ^ n4064 ;
  assign n4061 = x61 & n3885 ;
  assign n4068 = n4066 ^ n4061 ;
  assign n4079 = n2641 & n3876 ;
  assign n4069 = ~n3883 & ~n3886 ;
  assign n4070 = ~x36 & ~x88 ;
  assign n4071 = ~x104 & ~n2644 ;
  assign n4072 = n4070 & n4071 ;
  assign n4073 = n4072 ^ n2644 ;
  assign n4074 = ~n4069 & ~n4073 ;
  assign n4080 = n4079 ^ n4074 ;
  assign n4081 = ~n3875 & n4080 ;
  assign n4082 = n4081 ^ n4074 ;
  assign n4083 = x48 & n3884 ;
  assign n4140 = n3246 ^ x74 ;
  assign n4135 = n1779 ^ x49 ;
  assign n4085 = n3884 ^ x49 ;
  assign n4136 = n4135 ^ n4085 ;
  assign n4138 = n4136 ^ n3246 ;
  assign n4141 = n4140 ^ n4136 ;
  assign n4117 = ~x49 & n4085 ;
  assign n4118 = n4141 ^ n4117 ;
  assign n4119 = n4138 ^ n4118 ;
  assign n4120 = n4119 ^ n3884 ;
  assign n4139 = n4138 ^ n4085 ;
  assign n4144 = n4141 ^ n4139 ;
  assign n4145 = n4144 ^ n4135 ;
  assign n4122 = n4145 ^ n3884 ;
  assign n4123 = n4120 & ~n4122 ;
  assign n4146 = n4145 ^ x49 ;
  assign n4142 = n4141 ^ n4085 ;
  assign n4106 = n4142 ^ n4136 ;
  assign n4108 = n4138 ^ n4106 ;
  assign n4126 = n4141 ^ n4108 ;
  assign n4127 = n4146 ^ n4126 ;
  assign n4128 = n1779 & n4127 ;
  assign n4129 = n4123 & n4128 ;
  assign n4130 = n4129 ^ n4117 ;
  assign n4131 = n4140 ^ n4130 ;
  assign n4148 = n4131 ^ n1779 ;
  assign n4149 = n4148 ^ x49 ;
  assign n4095 = n4142 ^ n3884 ;
  assign n4150 = n4149 ^ n4095 ;
  assign n4151 = n1502 & n3876 ;
  assign n4152 = x24 & x50 ;
  assign n4153 = n4151 & n4152 ;
  assign n4154 = n3463 ^ n2814 ;
  assign n4155 = n3801 & n4154 ;
  assign n4156 = n2813 & n4155 ;
  assign n4157 = ~x58 & n3876 ;
  assign n4158 = ~x86 & n1262 ;
  assign n4159 = n1306 & n4158 ;
  assign n4160 = n4157 & n4159 ;
  assign n4161 = n1259 & n4160 ;
  assign n4162 = ~x94 & x110 ;
  assign n4163 = n4162 ^ n3970 ;
  assign n4164 = n4161 & n4163 ;
  assign n4165 = n3252 ^ n1571 ;
  assign n4168 = ~x252 & ~n4165 ;
  assign n4169 = n4168 ^ n1571 ;
  assign n4170 = n4164 & n4169 ;
  assign n4171 = ~n4156 & ~n4170 ;
  assign n4172 = ~n4153 & n4171 ;
  assign n4173 = n1407 & n1417 ;
  assign n4174 = n1461 & n3882 ;
  assign n4175 = n4173 & n4174 ;
  assign n4176 = n1223 & n4175 ;
  assign n4186 = n4023 ^ x211 ;
  assign n4187 = ~n4012 & ~n4186 ;
  assign n4188 = n4187 ^ n4021 ;
  assign n4189 = ~n1911 & ~n4188 ;
  assign n4183 = ~x199 & ~n4015 ;
  assign n4184 = n4183 ^ x200 ;
  assign n4185 = n4032 & n4184 ;
  assign n4190 = n4189 ^ n4185 ;
  assign n4243 = n4190 ^ n4009 ;
  assign n4238 = n4039 ^ n2937 ;
  assign n4177 = n2690 & n3991 ;
  assign n4178 = n4177 ^ x52 ;
  assign n4180 = n4178 ^ n2937 ;
  assign n4239 = n4238 ^ n4180 ;
  assign n4241 = n4239 ^ n4190 ;
  assign n4220 = ~n2937 & n4180 ;
  assign n4221 = n4239 ^ n4220 ;
  assign n4222 = n4241 ^ n4221 ;
  assign n4223 = n4222 ^ n4178 ;
  assign n4244 = n4243 ^ n4239 ;
  assign n4242 = n4241 ^ n4180 ;
  assign n4247 = n4244 ^ n4242 ;
  assign n4248 = n4247 ^ n4238 ;
  assign n4225 = n4248 ^ n4178 ;
  assign n4226 = n4223 & ~n4225 ;
  assign n4249 = n4248 ^ n2937 ;
  assign n4209 = n4244 ^ n4238 ;
  assign n4211 = n4241 ^ n4209 ;
  assign n4227 = n4244 ^ n4211 ;
  assign n4228 = n4249 ^ n4227 ;
  assign n4231 = ~n4039 & n4228 ;
  assign n4232 = n4226 & n4231 ;
  assign n4233 = n4232 ^ n4220 ;
  assign n4234 = n4243 ^ n4233 ;
  assign n4251 = n4234 ^ n4039 ;
  assign n4252 = n4251 ^ n2937 ;
  assign n4245 = n4244 ^ n4180 ;
  assign n4198 = n4245 ^ n4178 ;
  assign n4253 = n4252 ^ n4198 ;
  assign n4255 = n1266 & n4157 ;
  assign n4256 = n2607 & n4255 ;
  assign n4257 = n1316 & n4256 ;
  assign n4258 = ~x24 & n4257 ;
  assign n4259 = n4258 ^ n4257 ;
  assign n4254 = n3915 & n3917 ;
  assign n4261 = n4259 ^ n4254 ;
  assign n4265 = x106 & n3884 ;
  assign n4264 = x106 & n3883 ;
  assign n4266 = n4265 ^ n4264 ;
  assign n4262 = x24 & n1780 ;
  assign n4263 = n1758 & n4262 ;
  assign n4268 = n4266 ^ n4263 ;
  assign n4270 = x24 & n3780 ;
  assign n4269 = x45 & n3883 ;
  assign n4272 = n4270 ^ n4269 ;
  assign n4273 = x56 ^ x55 ;
  assign n4274 = ~x62 & n4273 ;
  assign n4275 = x841 ^ x24 ;
  assign n4276 = x56 & ~n4275 ;
  assign n4277 = n4276 ^ x24 ;
  assign n4278 = n4274 & ~n4277 ;
  assign n4279 = n1782 & n4278 ;
  assign n4284 = x24 & n1747 ;
  assign n4280 = ~x841 & n1785 ;
  assign n4281 = x62 & x924 ;
  assign n4282 = n4280 & n4281 ;
  assign n4283 = n4282 ^ n4280 ;
  assign n4285 = n4284 ^ n4283 ;
  assign n4286 = n1274 & n2759 ;
  assign n4287 = x841 & n4286 ;
  assign n4288 = n4287 ^ n4286 ;
  assign n4289 = ~x57 & n1206 ;
  assign n4290 = n1744 & n3788 ;
  assign n4291 = n4289 & n4290 ;
  assign n4292 = n4291 ^ n4282 ;
  assign n4293 = n3915 & n3919 ;
  assign n4294 = n1267 & n4256 ;
  assign n4295 = ~x24 & n4294 ;
  assign n4296 = n4295 ^ n4294 ;
  assign n4297 = ~n4293 & ~n4296 ;
  assign n4298 = x61 & n3884 ;
  assign n4299 = n4298 ^ n4295 ;
  assign n4300 = x62 ^ x57 ;
  assign n4305 = x62 & ~n4275 ;
  assign n4306 = n4305 ^ x24 ;
  assign n4307 = n4300 & ~n4306 ;
  assign n4308 = ~n1799 & n4307 ;
  assign n4309 = x63 & n3886 ;
  assign n4310 = ~x999 & n4309 ;
  assign n4311 = n4310 ^ n4309 ;
  assign n4312 = ~n4065 & ~n4311 ;
  assign n4313 = x107 & n3886 ;
  assign n4315 = n4313 ^ n3888 ;
  assign n4316 = ~n3922 & n3924 ;
  assign n4317 = n3915 & n4316 ;
  assign n4318 = n1355 & n3882 ;
  assign n4319 = x81 & n1250 ;
  assign n4320 = x314 & n1252 ;
  assign n4321 = n4319 & n4320 ;
  assign n4322 = n4318 & n4321 ;
  assign n4323 = x299 & n4036 ;
  assign n4324 = n4323 ^ x199 ;
  assign n4325 = n4322 & n4324 ;
  assign n4326 = ~x69 & n1455 ;
  assign n4327 = n4174 & n4326 ;
  assign n4328 = x314 & n4327 ;
  assign n4329 = x83 & ~x103 ;
  assign n4330 = n4328 & n4329 ;
  assign n4331 = n2801 & n2943 ;
  assign n4334 = n1936 & ~n2665 ;
  assign n4332 = x299 & ~n2723 ;
  assign n4333 = n1526 & n4332 ;
  assign n4335 = n4334 ^ n4333 ;
  assign n4336 = n4331 & n4335 ;
  assign n4337 = ~x71 & n3883 ;
  assign n4338 = ~x314 & n4337 ;
  assign n4339 = x69 & n4338 ;
  assign n4340 = n4339 ^ n4337 ;
  assign n4341 = n4340 ^ n3883 ;
  assign n4342 = ~x24 & x70 ;
  assign n4343 = n4342 ^ x70 ;
  assign n4344 = n2737 & n4343 ;
  assign n4345 = n2719 & n2943 ;
  assign n4346 = ~n4331 & ~n4345 ;
  assign n4349 = n1534 & ~n2665 ;
  assign n4350 = x198 & n4349 ;
  assign n4347 = n1538 & ~n2723 ;
  assign n4348 = x210 & n4347 ;
  assign n4351 = n4350 ^ n4348 ;
  assign n4352 = x589 & n4351 ;
  assign n4353 = ~n4346 & n4352 ;
  assign n4354 = x593 & n4353 ;
  assign n4355 = n4354 ^ n4353 ;
  assign n4356 = ~n3914 & ~n4355 ;
  assign n4357 = ~n4344 & n4356 ;
  assign n4363 = ~n1431 & n4174 ;
  assign n4364 = n4363 ^ n4322 ;
  assign n4358 = x85 & n1405 ;
  assign n4359 = n1444 & n4358 ;
  assign n4360 = ~n1244 & n4359 ;
  assign n4361 = ~x314 & n4360 ;
  assign n4362 = n4361 ^ n4360 ;
  assign n4365 = n4364 ^ n4362 ;
  assign n4371 = n4365 ^ n4363 ;
  assign n4366 = n4031 ^ x199 ;
  assign n4367 = n4366 ^ n4186 ;
  assign n4368 = ~x299 & n4367 ;
  assign n4369 = n4368 ^ n4186 ;
  assign n4370 = n4369 ^ n4324 ;
  assign n4372 = n4371 ^ n4370 ;
  assign n4373 = n4322 & n4372 ;
  assign n4374 = n4365 & ~n4373 ;
  assign n4375 = n4373 ^ n4371 ;
  assign n4376 = n4375 ^ n4322 ;
  assign n4377 = n4374 & n4376 ;
  assign n4378 = n4377 ^ n4375 ;
  assign n4379 = n3267 & n4331 ;
  assign n4380 = ~x38 & x88 ;
  assign n4381 = n1508 & n2645 ;
  assign n4382 = n4380 & n4381 ;
  assign n4383 = n4382 ^ x38 ;
  assign n4384 = n1220 & ~n4383 ;
  assign n4388 = x72 & n1290 ;
  assign n4393 = n4384 & n4388 ;
  assign n4394 = x24 & n4393 ;
  assign n4395 = n4394 ^ x24 ;
  assign n4385 = n4384 ^ n1220 ;
  assign n4386 = n4385 ^ x24 ;
  assign n4396 = n4395 ^ n4386 ;
  assign n4397 = ~n4379 & ~n4396 ;
  assign n4398 = x314 & x1050 ;
  assign n4399 = n4398 ^ x1050 ;
  assign n4400 = ~x39 & ~n4399 ;
  assign n4402 = n2728 & n4331 ;
  assign n4401 = x73 & n1971 ;
  assign n4404 = n4402 ^ n4401 ;
  assign n4405 = n4400 & n4404 ;
  assign n4406 = n4405 ^ n4404 ;
  assign n4407 = n1220 & ~n1571 ;
  assign n4411 = ~x479 & ~x841 ;
  assign n4408 = x479 & n1551 ;
  assign n4409 = n2640 & n4408 ;
  assign n4410 = n4409 ^ n2640 ;
  assign n4412 = n4411 ^ n4410 ;
  assign n4413 = ~x96 & n4412 ;
  assign n4414 = n4413 ^ n4411 ;
  assign n4415 = n4407 & n4414 ;
  assign n4416 = n1585 & n4415 ;
  assign n4417 = x74 & n4262 ;
  assign n4418 = ~n4416 & ~n4417 ;
  assign n4420 = x75 & n4262 ;
  assign n4419 = n1220 & n1590 ;
  assign n4422 = n4420 ^ n4419 ;
  assign n4423 = n3435 & ~n3847 ;
  assign n4430 = n3187 & n3437 ;
  assign n4424 = n4423 ^ x94 ;
  assign n4425 = n4424 ^ n3252 ;
  assign n4431 = n4430 ^ n4425 ;
  assign n4432 = n4423 & n4431 ;
  assign n4433 = n4432 ^ n4425 ;
  assign n4434 = n4433 ^ x94 ;
  assign n4435 = n4433 ^ n3252 ;
  assign n4436 = ~n4432 & ~n4435 ;
  assign n4437 = ~n4434 & n4436 ;
  assign n4438 = n4437 ^ n4433 ;
  assign n4439 = n1571 & ~n4438 ;
  assign n4440 = n3437 ^ x252 ;
  assign n4443 = x94 & n4440 ;
  assign n4444 = n4443 ^ n3437 ;
  assign n4445 = n4439 & n4444 ;
  assign n4446 = n4445 ^ n4438 ;
  assign n4447 = n1971 & ~n4446 ;
  assign n4448 = x77 & x314 ;
  assign n4449 = n4448 ^ n1263 ;
  assign n4450 = n2737 & ~n4449 ;
  assign n4451 = x232 & n2976 ;
  assign n4452 = n3270 & n3490 ;
  assign n4453 = ~x38 & n4452 ;
  assign n4454 = ~x34 & n3674 ;
  assign n4455 = n4454 ^ x79 ;
  assign n4456 = n4455 ^ n3500 ;
  assign n4457 = ~n3560 & ~n4456 ;
  assign n4458 = x39 & n3528 ;
  assign n4459 = n2801 & n3249 ;
  assign n4461 = ~x166 & n3567 ;
  assign n4460 = ~x189 & n3565 ;
  assign n4462 = n4461 ^ n4460 ;
  assign n4463 = n4459 & n4462 ;
  assign n4464 = n4463 ^ n3249 ;
  assign n4466 = x156 & n3567 ;
  assign n4465 = x179 & n3565 ;
  assign n4467 = n4466 ^ n4465 ;
  assign n4468 = n2719 & n4467 ;
  assign n4469 = n4464 & n4468 ;
  assign n4471 = n4469 ^ n4463 ;
  assign n4472 = n4458 & n4471 ;
  assign n4473 = n4472 ^ x39 ;
  assign n4474 = n4457 & n4473 ;
  assign n4475 = n4474 ^ n4473 ;
  assign n4476 = n4453 & ~n4475 ;
  assign n4477 = ~x166 & n3490 ;
  assign n4478 = n3481 & n4477 ;
  assign n4479 = ~x163 & x299 ;
  assign n4480 = ~n4478 & n4479 ;
  assign n4481 = ~n3599 & ~n4480 ;
  assign n4483 = x153 & n1330 ;
  assign n4484 = n2749 & n4483 ;
  assign n4485 = ~n1511 & n1608 ;
  assign n4486 = ~n4484 & n4485 ;
  assign n4482 = n1608 ^ x175 ;
  assign n4487 = n4486 ^ n4482 ;
  assign n4488 = x299 & n4487 ;
  assign n4489 = n4488 ^ x175 ;
  assign n4490 = ~n4481 & ~n4489 ;
  assign n4491 = x182 ^ x160 ;
  assign n4492 = ~x299 & n4491 ;
  assign n4493 = n4492 ^ x160 ;
  assign n4494 = n2744 & n3249 ;
  assign n4495 = ~n4493 & n4494 ;
  assign n4496 = n4495 ^ n3483 ;
  assign n4497 = x189 ^ x166 ;
  assign n4498 = ~x299 & n4497 ;
  assign n4499 = n4498 ^ x166 ;
  assign n4500 = n4495 ^ n3249 ;
  assign n4501 = n4499 & n4500 ;
  assign n4502 = n4496 & n4501 ;
  assign n4503 = n4502 ^ n4500 ;
  assign n4504 = ~x184 & ~n3609 ;
  assign n4505 = n4503 & n4504 ;
  assign n4506 = n4505 ^ n4503 ;
  assign n4507 = ~n4490 & n4506 ;
  assign n4508 = n4507 ^ n4456 ;
  assign n4509 = ~n3489 & ~n4508 ;
  assign n4510 = n4509 ^ n4456 ;
  assign n4511 = ~x39 & n4510 ;
  assign n4512 = n4476 & ~n4511 ;
  assign n4513 = n1848 & n3490 ;
  assign n4514 = x179 ^ x156 ;
  assign n4517 = x299 & n4514 ;
  assign n4518 = n4517 ^ x179 ;
  assign n4519 = n3249 & n4518 ;
  assign n4520 = n4519 ^ n4456 ;
  assign n4523 = n3700 & ~n4520 ;
  assign n4524 = n4523 ^ n4456 ;
  assign n4525 = n4513 & ~n4524 ;
  assign n4526 = n4525 ^ n1848 ;
  assign n4527 = ~n1750 & ~n4526 ;
  assign n4528 = ~x40 & ~n3552 ;
  assign n4529 = ~n4527 & n4528 ;
  assign n4530 = ~n4512 & n4529 ;
  assign n4543 = n3768 ^ x145 ;
  assign n4544 = n3770 & n4543 ;
  assign n4545 = n4544 ^ x140 ;
  assign n4546 = n4545 ^ x184 ;
  assign n4539 = n3765 ^ x197 ;
  assign n4540 = n3766 & n4539 ;
  assign n4541 = n4540 ^ x162 ;
  assign n4542 = n4541 ^ x163 ;
  assign n4547 = n4546 ^ n4542 ;
  assign n4548 = ~x299 & n4547 ;
  assign n4549 = n4548 ^ n4542 ;
  assign n4550 = n1211 & n3249 ;
  assign n4551 = n4549 & n4550 ;
  assign n4531 = n1847 & n3249 ;
  assign n4532 = x187 ^ x147 ;
  assign n4535 = ~x299 & n4532 ;
  assign n4536 = n4535 ^ x147 ;
  assign n4537 = n4531 & n4536 ;
  assign n4538 = n4537 ^ n1847 ;
  assign n4553 = n4551 ^ n4538 ;
  assign n4554 = ~n4530 & ~n4553 ;
  assign n4555 = n1209 & ~n4554 ;
  assign n4556 = ~x40 & ~n1206 ;
  assign n4557 = n3663 & n4556 ;
  assign n4560 = x163 & n3249 ;
  assign n4561 = n4560 ^ n4456 ;
  assign n4562 = n3679 & ~n4561 ;
  assign n4563 = n4562 ^ n4456 ;
  assign n4564 = n3490 & ~n4563 ;
  assign n4565 = n4557 & ~n4564 ;
  assign n4566 = ~n1209 & ~n3663 ;
  assign n4567 = n3249 ^ n1211 ;
  assign n4568 = n4542 ^ x74 ;
  assign n4569 = n1211 & ~n4568 ;
  assign n4570 = n4569 ^ x74 ;
  assign n4571 = n4567 & ~n4570 ;
  assign n4572 = n3249 & n4571 ;
  assign n4573 = ~x147 & n4572 ;
  assign n4574 = n4573 ^ n4571 ;
  assign n4575 = n4574 ^ n4570 ;
  assign n4576 = n4566 & ~n4575 ;
  assign n4577 = ~n4565 & ~n4576 ;
  assign n4578 = ~n4555 & n4577 ;
  assign n4579 = n2935 & n3402 ;
  assign n4580 = ~x592 & n3021 ;
  assign n4581 = n3307 & n4580 ;
  assign n4582 = n4581 ^ n3021 ;
  assign n4583 = n3323 ^ x590 ;
  assign n4584 = ~n3187 & ~n4583 ;
  assign n4585 = n4584 ^ x590 ;
  assign n4586 = x98 & ~x592 ;
  assign n4587 = x1199 & n4586 ;
  assign n4588 = n4587 ^ n3187 ;
  assign n4589 = n4588 ^ n4582 ;
  assign n4590 = ~n4585 & ~n4589 ;
  assign n4591 = n4590 ^ n3187 ;
  assign n4592 = n4582 & ~n4591 ;
  assign n4593 = ~x588 & ~x590 ;
  assign n4594 = ~n3019 & ~n4593 ;
  assign n4595 = n4592 & n4594 ;
  assign n4596 = n4595 ^ n4592 ;
  assign n4597 = n4579 & ~n4596 ;
  assign n4598 = n3240 & n4597 ;
  assign n4599 = ~x63 & n1799 ;
  assign n4600 = ~n2760 & n4599 ;
  assign n4601 = n4600 ^ n1799 ;
  assign n4602 = n4598 & ~n4601 ;
  assign n4603 = n3425 & n4582 ;
  assign n4604 = ~n4587 & n4603 ;
  assign n4605 = n4604 ^ n3425 ;
  assign n4606 = ~n4602 & ~n4605 ;
  assign n4607 = n3184 & ~n4606 ;
  assign n4608 = ~n2987 & ~n4607 ;
  assign n4609 = ~x80 & n2991 ;
  assign n4610 = ~n4608 & n4609 ;
  assign n4611 = ~x68 & ~n4069 ;
  assign n4612 = ~x314 & n4611 ;
  assign n4613 = x81 & n4612 ;
  assign n4614 = n4613 ^ n4611 ;
  assign n4615 = n4614 ^ n4069 ;
  assign n4616 = x314 ^ x66 ;
  assign n4619 = ~x69 & n4616 ;
  assign n4620 = n4619 ^ x314 ;
  assign n4621 = n3883 & n4620 ;
  assign n4625 = ~x314 & n4327 ;
  assign n4626 = n4329 & n4625 ;
  assign n4622 = ~x68 & x84 ;
  assign n4623 = n1255 & n4622 ;
  assign n4624 = n4363 & n4623 ;
  assign n4627 = n4626 ^ n4624 ;
  assign n4628 = n4322 & ~n4369 ;
  assign n4629 = ~x67 & n4363 ;
  assign n4630 = ~n4361 & n4629 ;
  assign n4631 = n4630 ^ n4363 ;
  assign n4632 = n4335 & n4345 ;
  assign n4633 = n2779 & n4328 ;
  assign n4634 = x88 & n2639 ;
  assign n4640 = n3886 & n4634 ;
  assign n4635 = x104 & n2644 ;
  assign n4636 = n3883 & n4635 ;
  assign n4637 = ~n3187 & n4636 ;
  assign n4638 = n4637 ^ n4636 ;
  assign n4641 = n4640 ^ n4638 ;
  assign n4642 = n2737 & ~n4342 ;
  assign n4643 = x89 & n4642 ;
  assign n4644 = x841 & n4643 ;
  assign n4645 = n4644 ^ n4642 ;
  assign n4646 = n4645 ^ n2737 ;
  assign n4647 = ~x1050 & n4401 ;
  assign n4648 = n4647 ^ n4287 ;
  assign n4657 = n2943 & n3268 ;
  assign n4649 = n3874 ^ x24 ;
  assign n4650 = n1577 & ~n4649 ;
  assign n4651 = n4650 ^ x24 ;
  assign n4652 = n3216 ^ n1577 ;
  assign n4653 = n4652 ^ n4157 ;
  assign n4654 = n4651 & ~n4653 ;
  assign n4655 = n4654 ^ n1577 ;
  assign n4656 = n4157 & n4655 ;
  assign n4659 = n4657 ^ n4656 ;
  assign n4662 = x92 & n4399 ;
  assign n4663 = n4662 ^ n2729 ;
  assign n4664 = ~x39 & n4663 ;
  assign n4665 = n4664 ^ n2729 ;
  assign n4666 = n1797 & n4665 ;
  assign n4668 = n1770 & n1849 ;
  assign n4669 = ~x1050 & n4668 ;
  assign n4667 = n2610 & n2737 ;
  assign n4671 = n4669 ^ n4667 ;
  assign n4689 = n3254 ^ x49 ;
  assign n4673 = n3885 ^ x49 ;
  assign n4690 = n4689 ^ n4673 ;
  assign n4701 = n4690 ^ n4164 ;
  assign n4688 = n4164 ^ n1571 ;
  assign n4691 = n4690 ^ n4688 ;
  assign n4692 = n4691 ^ n4673 ;
  assign n4704 = n4701 ^ n4692 ;
  assign n4705 = n4704 ^ n4689 ;
  assign n4706 = n4705 ^ x49 ;
  assign n4686 = ~n1571 & n4164 ;
  assign n4687 = x49 & ~n3885 ;
  assign n4693 = n4692 ^ n4687 ;
  assign n4694 = n4164 ^ n3254 ;
  assign n4695 = n4694 ^ n4687 ;
  assign n4696 = n4695 ^ n4692 ;
  assign n4697 = ~n4693 & ~n4696 ;
  assign n4698 = n4686 & n4697 ;
  assign n4699 = n4698 ^ n4695 ;
  assign n4707 = n4706 ^ n4699 ;
  assign n4708 = n4707 ^ n3254 ;
  assign n4709 = n4708 ^ x49 ;
  assign n4683 = n4692 ^ n3885 ;
  assign n4710 = n4709 ^ n4683 ;
  assign n4716 = n4349 ^ n4347 ;
  assign n4717 = ~n4346 & n4716 ;
  assign n4719 = n4717 ^ n3885 ;
  assign n4718 = n4717 ^ n4352 ;
  assign n4720 = n4719 ^ n4718 ;
  assign n4726 = n4720 ^ x89 ;
  assign n4721 = n4720 ^ x332 ;
  assign n4722 = n4721 ^ n4718 ;
  assign n4762 = n4726 ^ n4722 ;
  assign n4763 = n4762 ^ n4719 ;
  assign n4742 = ~n4717 & ~n4718 ;
  assign n4743 = n4763 ^ n4742 ;
  assign n4744 = n4743 ^ n4721 ;
  assign n4745 = n4744 ^ n4352 ;
  assign n4748 = n3885 & ~n4745 ;
  assign n4749 = n4726 ^ n4719 ;
  assign n4734 = n4719 ^ n4352 ;
  assign n4750 = n4749 ^ n4734 ;
  assign n4752 = n4762 ^ n4734 ;
  assign n4753 = ~n4750 & ~n4752 ;
  assign n4754 = n4748 & n4753 ;
  assign n4755 = n4754 ^ n4742 ;
  assign n4756 = n4755 ^ x332 ;
  assign n4735 = n4721 ^ n4719 ;
  assign n4736 = n4735 ^ n4734 ;
  assign n4757 = n4756 ^ n4736 ;
  assign n4727 = n4726 ^ n4718 ;
  assign n4728 = n4727 ^ n4722 ;
  assign n4758 = n4757 ^ n4728 ;
  assign n4771 = n4758 ^ n4734 ;
  assign n4772 = n4771 ^ n3885 ;
  assign n4773 = n4772 ^ n4352 ;
  assign n4764 = n4763 ^ n4717 ;
  assign n4774 = n4773 ^ n4764 ;
  assign n4711 = ~x32 & ~x40 ;
  assign n4712 = n1220 & n4711 ;
  assign n4713 = x95 & n4712 ;
  assign n4714 = n1300 & n4713 ;
  assign n4715 = x24 & n4714 ;
  assign n4776 = n4774 ^ n4715 ;
  assign n4777 = ~n1300 & ~n1508 ;
  assign n4778 = x96 ^ x95 ;
  assign n4781 = ~n1572 & ~n4411 ;
  assign n4782 = n4781 ^ x24 ;
  assign n4783 = x96 & ~n4782 ;
  assign n4784 = n4783 ^ x24 ;
  assign n4785 = n4778 & ~n4784 ;
  assign n4786 = n4712 & n4785 ;
  assign n4787 = ~n4777 & n4786 ;
  assign n4788 = ~n1577 & ~n4410 ;
  assign n4789 = n3876 & n4788 ;
  assign n4790 = n1580 & n4789 ;
  assign n4791 = ~n4354 & ~n4790 ;
  assign n4792 = n4668 ^ n4401 ;
  assign n4793 = n4398 & n4792 ;
  assign n4805 = n2682 & n3992 ;
  assign n4806 = n4805 ^ x99 ;
  assign n4807 = n2937 & n4806 ;
  assign n4796 = n3950 ^ n3943 ;
  assign n4795 = ~x144 & n3950 ;
  assign n4797 = n4796 ^ n4795 ;
  assign n4794 = ~x161 & n3943 ;
  assign n4798 = n4797 ^ n4794 ;
  assign n4799 = n3941 & n4798 ;
  assign n4808 = n4807 ^ n4799 ;
  assign n4809 = n2813 & ~n3253 ;
  assign n4810 = n3462 & n4809 ;
  assign n4811 = n4810 ^ n2813 ;
  assign n4812 = n3252 ^ n1562 ;
  assign n4813 = x683 & ~n3455 ;
  assign n4818 = ~n2644 & n4813 ;
  assign n4819 = n4818 ^ x252 ;
  assign n4820 = ~n4812 & ~n4819 ;
  assign n4821 = n4820 ^ n4813 ;
  assign n4822 = ~n3252 & n3458 ;
  assign n4823 = ~n4821 & n4822 ;
  assign n4824 = n4823 ^ n3458 ;
  assign n4825 = n1210 & ~n4824 ;
  assign n4826 = n4811 & n4825 ;
  assign n4828 = n4826 ^ n4810 ;
  assign n4829 = n3992 ^ x101 ;
  assign n4833 = n2937 & n4829 ;
  assign n4830 = n4795 ^ n4794 ;
  assign n4831 = n3941 & n4830 ;
  assign n4834 = n4833 ^ n4831 ;
  assign n4835 = x65 & n3886 ;
  assign n4837 = n2644 & ~n3252 ;
  assign n4838 = n4161 & n4162 ;
  assign n4839 = n4837 & n4838 ;
  assign n4840 = n4839 ^ n4838 ;
  assign n4841 = ~n4637 & ~n4840 ;
  assign n4842 = n4265 ^ n4258 ;
  assign n4844 = n3901 ^ x108 ;
  assign n4845 = ~x98 & n4151 ;
  assign n4846 = ~n4844 & n4845 ;
  assign n4847 = n4846 ^ n4151 ;
  assign n4843 = n2941 & ~n4601 ;
  assign n4849 = n4847 ^ n4843 ;
  assign n4850 = n4151 & n4448 ;
  assign n4851 = n2779 & n4175 ;
  assign n4852 = ~x314 & n4851 ;
  assign n4853 = n4852 ^ n4851 ;
  assign n4854 = ~n4839 & ~n4853 ;
  assign n4855 = ~x24 & n1220 ;
  assign n4857 = n4388 & n4855 ;
  assign n4858 = n4857 ^ n4852 ;
  assign n4859 = x124 & ~x468 ;
  assign n4864 = n2683 & n3992 ;
  assign n4865 = n4864 ^ x113 ;
  assign n4866 = n2937 & n4865 ;
  assign n4867 = n4002 ^ x114 ;
  assign n4868 = n2937 & n4867 ;
  assign n4873 = ~x116 & n4001 ;
  assign n4874 = n4873 ^ x115 ;
  assign n4875 = n2937 & n4874 ;
  assign n4876 = n4001 ^ x116 ;
  assign n4877 = n2937 & n4876 ;
  assign n4878 = x87 & n3249 ;
  assign n4879 = n4878 ^ n3249 ;
  assign n4880 = n3528 & n4879 ;
  assign n4881 = x92 ^ x39 ;
  assign n4890 = x178 ^ x157 ;
  assign n4891 = ~x299 & n4890 ;
  assign n4892 = n4891 ^ x157 ;
  assign n4887 = x157 & n2719 ;
  assign n4886 = x168 & n2801 ;
  assign n4888 = n4887 ^ n4886 ;
  assign n4889 = n3567 & n4888 ;
  assign n4893 = n4892 ^ n4889 ;
  assign n4883 = x178 & n2719 ;
  assign n4882 = x190 & n2801 ;
  assign n4884 = n4883 ^ n4882 ;
  assign n4885 = n3565 & n4884 ;
  assign n4896 = n4893 ^ n4885 ;
  assign n4897 = ~x92 & n4896 ;
  assign n4898 = n4897 ^ n4892 ;
  assign n4899 = n4881 & n4898 ;
  assign n4900 = n4880 & n4899 ;
  assign n4901 = n3491 & ~n4900 ;
  assign n4902 = n1218 & ~n3489 ;
  assign n4919 = n3249 & n3599 ;
  assign n4920 = x173 ^ x151 ;
  assign n4923 = ~x299 & n4920 ;
  assign n4924 = n4923 ^ x151 ;
  assign n4925 = n4919 & ~n4924 ;
  assign n4926 = n4925 ^ n3249 ;
  assign n4927 = ~n2744 & ~n4926 ;
  assign n4928 = ~x150 & x299 ;
  assign n4929 = ~n3618 & n4928 ;
  assign n4930 = n4929 ^ x299 ;
  assign n4932 = x73 & ~x168 ;
  assign n4933 = n4930 & n4932 ;
  assign n4934 = n4933 ^ n4929 ;
  assign n4935 = ~x185 & ~x299 ;
  assign n4936 = ~x73 & x232 ;
  assign n4937 = ~n1634 & n3618 ;
  assign n4938 = n4936 & n4937 ;
  assign n4939 = n4938 ^ n3618 ;
  assign n4940 = n4935 & ~n4939 ;
  assign n4941 = n4940 ^ x299 ;
  assign n4944 = n4940 ^ x190 ;
  assign n4945 = x73 & ~n4944 ;
  assign n4946 = ~n4941 & n4945 ;
  assign n4947 = n4946 ^ n4941 ;
  assign n4948 = n4947 ^ x299 ;
  assign n4949 = ~n4934 & ~n4948 ;
  assign n4950 = ~n4927 & n4949 ;
  assign n4903 = ~x54 & n1846 ;
  assign n4904 = ~n1755 & ~n3270 ;
  assign n4905 = n4903 & ~n4904 ;
  assign n4906 = x39 ^ x38 ;
  assign n4907 = ~x92 & n4906 ;
  assign n4908 = ~x38 & n4907 ;
  assign n4909 = ~n3559 & n4908 ;
  assign n4910 = n4909 ^ n4907 ;
  assign n4911 = n4910 ^ x92 ;
  assign n4912 = n4905 & n4911 ;
  assign n4913 = n1743 & n4912 ;
  assign n4915 = n3500 ^ x118 ;
  assign n4914 = ~x79 & n4454 ;
  assign n4916 = n4915 ^ n4914 ;
  assign n4917 = n1848 & n4916 ;
  assign n4918 = ~n4913 & ~n4917 ;
  assign n4951 = n4950 ^ n4918 ;
  assign n4952 = n4902 & n4951 ;
  assign n4953 = n4952 ^ n4918 ;
  assign n4954 = n4901 & ~n4953 ;
  assign n4955 = n1206 & ~n1911 ;
  assign n4960 = ~x163 & ~n4541 ;
  assign n4961 = n4960 ^ x150 ;
  assign n4962 = n1211 & ~n4961 ;
  assign n4963 = n4962 ^ n3662 ;
  assign n4964 = n3249 & n4963 ;
  assign n4965 = n4964 ^ n3662 ;
  assign n4966 = ~x165 & n3662 ;
  assign n4967 = ~n4965 & n4966 ;
  assign n4968 = n4967 ^ n4965 ;
  assign n4969 = n4955 & n4968 ;
  assign n4970 = n4969 ^ n3249 ;
  assign n4971 = n4969 ^ n1206 ;
  assign n4972 = n3662 & n4971 ;
  assign n4973 = ~n4970 & n4972 ;
  assign n4974 = n4973 ^ n4971 ;
  assign n4975 = ~x299 & n4550 ;
  assign n4980 = ~x184 & ~n4545 ;
  assign n4981 = n4980 ^ x185 ;
  assign n4982 = n4975 & ~n4981 ;
  assign n4983 = n4982 ^ x299 ;
  assign n4991 = ~x143 & ~n4983 ;
  assign n4992 = n1847 & n4991 ;
  assign n4993 = n4992 ^ n1847 ;
  assign n4985 = n4982 ^ n1847 ;
  assign n4994 = n4993 ^ n4985 ;
  assign n4995 = n4974 & ~n4994 ;
  assign n4996 = ~n4954 & n4995 ;
  assign n4997 = ~n1209 & ~n4968 ;
  assign n5000 = x150 & n3249 ;
  assign n5001 = n5000 ^ n4916 ;
  assign n5002 = n1745 & ~n5001 ;
  assign n5003 = n5002 ^ n4916 ;
  assign n5004 = n3664 & ~n5003 ;
  assign n5005 = n5004 ^ n3664 ;
  assign n5006 = n4997 & ~n5005 ;
  assign n5007 = ~n4996 & ~n5006 ;
  assign n5020 = n3266 & n4345 ;
  assign n5008 = n1330 & ~n1578 ;
  assign n5009 = n1328 & ~n2848 ;
  assign n5010 = n1971 & n5009 ;
  assign n5013 = n5010 ^ n1971 ;
  assign n5011 = ~x109 & n1263 ;
  assign n5012 = n5010 & n5011 ;
  assign n5014 = n5013 ^ n5012 ;
  assign n5015 = n5008 & n5014 ;
  assign n5016 = n5015 ^ n1971 ;
  assign n5017 = n1861 & n2813 ;
  assign n5018 = ~n4668 & ~n5017 ;
  assign n5019 = ~n5016 & n5018 ;
  assign n5022 = n5020 ^ n5019 ;
  assign n5023 = n5022 ^ x128 ;
  assign n5024 = ~x228 & ~n5023 ;
  assign n5025 = n5024 ^ x128 ;
  assign n5026 = ~x31 & ~x80 ;
  assign n5027 = x818 & n5026 ;
  assign n5028 = x951 & x982 ;
  assign n5029 = n2985 & n5028 ;
  assign n5030 = n2991 & n5029 ;
  assign n5031 = ~n5027 & ~n5030 ;
  assign n5032 = x1093 & ~n5031 ;
  assign n5033 = ~x120 & ~n5032 ;
  assign n5034 = n1209 & ~n3245 ;
  assign n5035 = ~n3280 & ~n3425 ;
  assign n5036 = n5034 & n5035 ;
  assign n5037 = n5036 ^ n3425 ;
  assign n5038 = ~n5033 & ~n5037 ;
  assign n5141 = ~x24 & x77 ;
  assign n5142 = n5141 ^ x77 ;
  assign n5143 = ~x86 & ~n5142 ;
  assign n5144 = ~n4448 & n5143 ;
  assign n5145 = ~x39 & ~n5144 ;
  assign n5146 = n2935 & n5145 ;
  assign n5147 = n1582 & n5146 ;
  assign n5148 = n1493 & n5147 ;
  assign n5134 = ~x24 & n4448 ;
  assign n5170 = n4519 & ~n5134 ;
  assign n5149 = x72 ^ x39 ;
  assign n5150 = n2936 & n5149 ;
  assign n5151 = x39 & ~n2802 ;
  assign n5152 = n5150 & n5151 ;
  assign n5153 = n5152 ^ n5150 ;
  assign n5156 = ~x134 & ~x135 ;
  assign n5157 = ~x136 & n5156 ;
  assign n5154 = ~x125 & ~x133 ;
  assign n5158 = ~x121 & n5154 ;
  assign n5159 = x126 & ~x132 ;
  assign n5160 = n5159 ^ x132 ;
  assign n5161 = n5158 & ~n5160 ;
  assign n5162 = ~x130 & n5161 ;
  assign n5163 = n5157 & n5162 ;
  assign n5155 = n5154 ^ x121 ;
  assign n5164 = n5163 ^ n5155 ;
  assign n5165 = ~n5153 & ~n5164 ;
  assign n5171 = n5170 ^ n5165 ;
  assign n5172 = n5148 & n5171 ;
  assign n5173 = n5172 ^ n5165 ;
  assign n5174 = n2942 & n5173 ;
  assign n5042 = ~n1911 & n3722 ;
  assign n5043 = n5042 ^ x144 ;
  assign n5463 = ~n1258 & ~n2941 ;
  assign n5044 = n5043 & n5463 ;
  assign n5045 = n5044 ^ n2942 ;
  assign n5074 = n5045 ^ n3915 ;
  assign n5065 = n5074 ^ n2799 ;
  assign n5114 = n5065 ^ n3719 ;
  assign n5051 = x184 ^ x163 ;
  assign n5052 = n1911 & n5051 ;
  assign n5053 = n5052 ^ x163 ;
  assign n5048 = n1552 & ~n1911 ;
  assign n5049 = n5048 ^ x142 ;
  assign n5050 = x51 & n5049 ;
  assign n5054 = n5053 ^ n5050 ;
  assign n5055 = ~x87 & ~n5054 ;
  assign n5056 = n5055 ^ n5053 ;
  assign n5128 = n5114 ^ n5056 ;
  assign n5100 = n2799 & n5128 ;
  assign n5076 = n3719 ^ n2799 ;
  assign n5116 = n5065 ^ n3915 ;
  assign n5057 = n5056 ^ n5045 ;
  assign n5117 = n5116 ^ n5057 ;
  assign n5087 = n5117 ^ n5045 ;
  assign n5102 = n5128 ^ n5087 ;
  assign n5105 = ~n5076 & ~n5102 ;
  assign n5106 = n5100 & n5105 ;
  assign n5107 = n5106 ^ ~n5056 ;
  assign n5115 = n5114 ^ n5057 ;
  assign n5119 = n5116 ^ n5115 ;
  assign n5066 = n5065 ^ n5057 ;
  assign n5120 = n5119 ^ n5066 ;
  assign n5075 = n5074 ^ n5057 ;
  assign n5081 = n5075 ^ n3719 ;
  assign n5082 = n5081 ^ n5057 ;
  assign n5090 = n5120 ^ n5082 ;
  assign n5108 = n5107 ^ n5090 ;
  assign n5109 = n5108 ^ n3915 ;
  assign n5077 = n5076 ^ n3915 ;
  assign n5110 = n5109 ^ n5077 ;
  assign n5111 = n5110 ^ n5087 ;
  assign n5132 = n5111 ^ n5045 ;
  assign n5133 = n5132 ^ n5128 ;
  assign n5135 = n3603 & n5134 ;
  assign n5136 = n2737 & n5135 ;
  assign n5137 = n5136 ^ n3249 ;
  assign n5138 = n3249 & n5137 ;
  assign n5139 = n5133 & n5138 ;
  assign n5140 = n5139 ^ n3249 ;
  assign n5176 = n5174 ^ n5140 ;
  assign n5177 = ~x90 & ~x111 ;
  assign n5178 = ~x72 & n5177 ;
  assign n5179 = n2777 & n5178 ;
  assign n5180 = n2737 & ~n5179 ;
  assign n5182 = ~x39 & x110 ;
  assign n5181 = x110 ^ x39 ;
  assign n5183 = n5182 ^ n5181 ;
  assign n5184 = n2954 & n5183 ;
  assign n5185 = n3249 & n4055 ;
  assign n5186 = n2644 & n5182 ;
  assign n5187 = ~n2691 & n5186 ;
  assign n5188 = ~n5185 & n5187 ;
  assign n5189 = ~n5184 & ~n5188 ;
  assign n5190 = ~n5180 & n5189 ;
  assign n5225 = ~x87 & n1209 ;
  assign n5226 = n1508 & ~n5144 ;
  assign n5227 = ~x39 & ~n4388 ;
  assign n5228 = ~n5226 & n5227 ;
  assign n5229 = n2934 & ~n5228 ;
  assign n5211 = ~x152 & ~n1258 ;
  assign n5212 = n5211 ^ x172 ;
  assign n5213 = ~x51 & n5212 ;
  assign n5214 = n5213 ^ x172 ;
  assign n5230 = x299 & n3249 ;
  assign n5231 = ~n5214 & n5230 ;
  assign n5232 = n5231 ^ n3249 ;
  assign n5235 = ~x174 & ~n1258 ;
  assign n5236 = n5235 ^ x193 ;
  assign n5237 = ~x51 & n5236 ;
  assign n5238 = n5237 ^ x193 ;
  assign n5239 = ~x299 & n5238 ;
  assign n5240 = n5239 ^ x299 ;
  assign n5241 = n5232 & n5240 ;
  assign n5203 = n5163 ^ x133 ;
  assign n5204 = n5203 ^ x125 ;
  assign n5205 = n2942 & n5204 ;
  assign n5242 = n5241 ^ n5205 ;
  assign n5243 = n5229 & ~n5242 ;
  assign n5247 = ~x287 & n3249 ;
  assign n5248 = x158 & n1523 ;
  assign n5249 = n5247 & n5248 ;
  assign n5250 = n5249 ^ n1743 ;
  assign n5251 = n1743 & n5250 ;
  assign n5252 = ~n3262 & n5251 ;
  assign n5253 = n5252 ^ n1743 ;
  assign n5254 = ~n5232 & ~n5253 ;
  assign n5255 = ~x72 & n2933 ;
  assign n5256 = ~x51 & x222 ;
  assign n5257 = ~x223 & n5256 ;
  assign n5258 = n1258 & n5257 ;
  assign n5259 = x180 & x224 ;
  assign n5260 = ~x287 & n2635 ;
  assign n5261 = n5259 & n5260 ;
  assign n5262 = n5261 ^ x224 ;
  assign n5263 = n5258 & ~n5262 ;
  assign n5264 = n5255 & n5263 ;
  assign n5265 = ~n5240 & ~n5264 ;
  assign n5266 = ~n5254 & ~n5265 ;
  assign n5271 = n5243 & ~n5266 ;
  assign n5272 = x39 & n5271 ;
  assign n5273 = n5272 ^ x39 ;
  assign n5244 = n5243 ^ n5242 ;
  assign n5245 = n5244 ^ x39 ;
  assign n5274 = n5273 ^ n5245 ;
  assign n5275 = n5225 & n5274 ;
  assign n5282 = x39 & n2934 ;
  assign n5283 = n2799 & n5282 ;
  assign n5284 = n5255 & n5283 ;
  assign n5287 = ~n5266 & n5284 ;
  assign n5288 = n5275 & n5287 ;
  assign n5289 = n5288 ^ n5275 ;
  assign n5290 = n5289 ^ n1209 ;
  assign n5293 = x162 ^ x140 ;
  assign n5294 = x299 & n5293 ;
  assign n5295 = n5294 ^ x140 ;
  assign n5296 = n4878 & n5295 ;
  assign n5297 = n5290 & n5296 ;
  assign n5206 = ~n1209 & n3249 ;
  assign n5215 = n5214 ^ x162 ;
  assign n5218 = ~x87 & n5215 ;
  assign n5219 = n5218 ^ x162 ;
  assign n5220 = n5206 & n5219 ;
  assign n5221 = n5220 ^ n1209 ;
  assign n5222 = ~n5205 & ~n5221 ;
  assign n5191 = n1218 & n5148 ;
  assign n5192 = n3249 & n5191 ;
  assign n5193 = x197 ^ x145 ;
  assign n5194 = x299 & n5193 ;
  assign n5195 = n5194 ^ x145 ;
  assign n5196 = n5195 ^ n3703 ;
  assign n5199 = n5143 & n5196 ;
  assign n5200 = n5199 ^ n3703 ;
  assign n5201 = n5192 & n5200 ;
  assign n5202 = n5201 ^ n5191 ;
  assign n5224 = n5222 ^ n5202 ;
  assign n5292 = n5290 ^ n5224 ;
  assign n5298 = n5297 ^ n5292 ;
  assign n5327 = n2942 & ~n5191 ;
  assign n5328 = n5158 ^ x126 ;
  assign n5333 = ~x130 & n5157 ;
  assign n5334 = n5333 ^ n5159 ;
  assign n5335 = ~n5160 & n5334 ;
  assign n5336 = n5328 & ~n5335 ;
  assign n5337 = n5327 & n5336 ;
  assign n5338 = n5337 ^ n5191 ;
  assign n5339 = ~n5153 & n5338 ;
  assign n5304 = x182 & n5247 ;
  assign n5305 = n5304 ^ n2799 ;
  assign n5306 = n1935 & ~n5305 ;
  assign n5307 = n5306 ^ n2799 ;
  assign n5308 = n5307 ^ x160 ;
  assign n5309 = n5308 ^ n5306 ;
  assign n5310 = n5247 ^ n2726 ;
  assign n5311 = n5306 ^ n5247 ;
  assign n5312 = ~n5310 & n5311 ;
  assign n5313 = ~n5309 & n5312 ;
  assign n5314 = n5313 ^ n5307 ;
  assign n5325 = n2943 & n5314 ;
  assign n5315 = ~n1209 & ~n2942 ;
  assign n5316 = x166 ^ x153 ;
  assign n5319 = ~x51 & ~n5316 ;
  assign n5320 = n5319 ^ x153 ;
  assign n5321 = n4879 & n5320 ;
  assign n5322 = n5315 & n5321 ;
  assign n5323 = n5322 ^ n2942 ;
  assign n5326 = n5325 ^ n5323 ;
  assign n5341 = n5339 ^ n5326 ;
  assign n5342 = n3249 & ~n5341 ;
  assign n5361 = n4892 ^ n3719 ;
  assign n5364 = ~n5143 & n5361 ;
  assign n5365 = n5364 ^ n3719 ;
  assign n5366 = n5191 & n5365 ;
  assign n5353 = x299 ^ x185 ;
  assign n5354 = n5353 ^ x150 ;
  assign n5355 = n1911 & n5354 ;
  assign n5356 = n5355 ^ x150 ;
  assign n5348 = ~n1258 & ~n4499 ;
  assign n5343 = x175 ^ x153 ;
  assign n5344 = ~x299 & n5343 ;
  assign n5345 = n5344 ^ x153 ;
  assign n5349 = n5348 ^ n5345 ;
  assign n5350 = ~x51 & n5349 ;
  assign n5351 = n5350 ^ n5345 ;
  assign n5352 = n1209 & n5351 ;
  assign n5357 = n5356 ^ n5352 ;
  assign n5358 = ~x87 & n5357 ;
  assign n5359 = n5358 ^ n5356 ;
  assign n5367 = n5366 ^ n5359 ;
  assign n5368 = n5342 & n5367 ;
  assign n5369 = n5368 ^ n5341 ;
  assign n5370 = x94 & x129 ;
  assign n5371 = n2640 ^ x127 ;
  assign n5372 = x250 & n3254 ;
  assign n5373 = n5371 & n5372 ;
  assign n5374 = n5373 ^ x127 ;
  assign n5375 = n5370 & ~n5374 ;
  assign n5376 = n5375 ^ x129 ;
  assign n5377 = ~n4601 & n5376 ;
  assign n5378 = ~x250 & n3456 ;
  assign n5386 = ~n3254 & n5378 ;
  assign n5387 = ~x100 & n5386 ;
  assign n5388 = n5387 ^ x100 ;
  assign n5379 = n5378 ^ x129 ;
  assign n5380 = n5379 ^ x100 ;
  assign n5389 = n5388 ^ n5380 ;
  assign n5390 = n1211 & ~n5389 ;
  assign n5391 = ~n1799 & ~n5390 ;
  assign n5392 = ~n1971 & ~n5391 ;
  assign n5394 = n2802 & n5247 ;
  assign n5395 = n1743 & ~n3262 ;
  assign n5396 = n5295 & n5395 ;
  assign n5397 = n5394 & n5396 ;
  assign n5398 = n5397 ^ n5395 ;
  assign n5399 = n5398 ^ n1743 ;
  assign n5400 = n5282 & ~n5399 ;
  assign n5401 = n5400 ^ n5229 ;
  assign n5403 = n5161 ^ x130 ;
  assign n5404 = n1258 & n5403 ;
  assign n5405 = n5157 & n5404 ;
  assign n5406 = n5161 & n5405 ;
  assign n5407 = n5406 ^ n5404 ;
  assign n5408 = n5407 ^ n1258 ;
  assign n5409 = ~n5284 & n5408 ;
  assign n5402 = ~n1258 & n3526 ;
  assign n5410 = n5409 ^ n5402 ;
  assign n5411 = n5225 & ~n5410 ;
  assign n5412 = ~n5401 & n5411 ;
  assign n5413 = ~n1258 & n3249 ;
  assign n5414 = x169 & n5413 ;
  assign n5415 = ~n1209 & ~n4878 ;
  assign n5416 = ~n5414 & n5415 ;
  assign n5417 = ~n5408 & n5416 ;
  assign n5418 = ~n5412 & ~n5417 ;
  assign n5419 = ~x51 & ~n5418 ;
  assign n5422 = n1911 & n3742 ;
  assign n5423 = n5422 ^ x167 ;
  assign n5424 = n4878 & n5423 ;
  assign n5425 = n5424 ^ x87 ;
  assign n5426 = ~n5419 & ~n5425 ;
  assign n5427 = n2799 & n2939 ;
  assign n5428 = n2942 & ~n5427 ;
  assign n5429 = ~n5148 & n5428 ;
  assign n5431 = x183 & n1530 ;
  assign n5430 = x149 & n2724 ;
  assign n5432 = n5431 ^ n5430 ;
  assign n5433 = n3249 & n4493 ;
  assign n5434 = n5141 & n5433 ;
  assign n5435 = n5434 ^ n5141 ;
  assign n5436 = n5432 & ~n5435 ;
  assign n5437 = n5247 & n5436 ;
  assign n5438 = n2942 & n5437 ;
  assign n5439 = ~n5429 & ~n5438 ;
  assign n5440 = x132 ^ x126 ;
  assign n5441 = n5440 ^ n5335 ;
  assign n5442 = n5441 ^ x132 ;
  assign n5445 = n5158 & ~n5442 ;
  assign n5446 = n5445 ^ x132 ;
  assign n5447 = ~n5153 & n5446 ;
  assign n5448 = ~n5439 & ~n5447 ;
  assign n5472 = n5191 & ~n5435 ;
  assign n5452 = ~n1209 & n3505 ;
  assign n5453 = n5452 ^ n3506 ;
  assign n5454 = n4878 & ~n5453 ;
  assign n5455 = n5454 ^ n3249 ;
  assign n5456 = n2940 & n5455 ;
  assign n5459 = n1911 & n4920 ;
  assign n5460 = n5459 ^ x151 ;
  assign n5461 = n5456 & ~n5460 ;
  assign n5462 = n5461 ^ n5455 ;
  assign n5464 = x190 ^ x168 ;
  assign n5467 = n1911 & n5464 ;
  assign n5468 = n5467 ^ x168 ;
  assign n5469 = n5463 & n5468 ;
  assign n5470 = n5469 ^ n2941 ;
  assign n5471 = n5462 & n5470 ;
  assign n5474 = n5472 ^ n5471 ;
  assign n5475 = ~n5448 & ~n5474 ;
  assign n5482 = x183 ^ x149 ;
  assign n5485 = ~n1911 & n5482 ;
  assign n5486 = n5485 ^ x183 ;
  assign n5487 = n4878 & n5486 ;
  assign n5477 = ~x86 & n3449 ;
  assign n5478 = ~n3539 & n5477 ;
  assign n5479 = n5478 ^ n3539 ;
  assign n5476 = n5203 & n5428 ;
  assign n5480 = n5479 ^ n5476 ;
  assign n5489 = n5487 ^ n5480 ;
  assign n5490 = ~n5191 & n5489 ;
  assign n5491 = n5490 ^ n5479 ;
  assign n5492 = ~n4601 & ~n5491 ;
  assign n5493 = ~x72 & ~n3262 ;
  assign n5494 = n5149 & n5493 ;
  assign n5495 = n5394 & n5494 ;
  assign n5496 = n5195 & n5495 ;
  assign n5497 = n5496 ^ n5494 ;
  assign n5498 = n5497 ^ n5149 ;
  assign n5499 = n5492 & n5498 ;
  assign n5500 = n5499 ^ n5491 ;
  assign n5501 = ~n2941 & ~n5148 ;
  assign n5514 = x192 ^ x171 ;
  assign n5517 = ~n1911 & n5514 ;
  assign n5518 = n5517 ^ x192 ;
  assign n5519 = n3249 & n5518 ;
  assign n5509 = n5163 ^ x134 ;
  assign n5507 = ~x136 & n5162 ;
  assign n5508 = ~x135 & n5507 ;
  assign n5510 = n5509 ^ n5508 ;
  assign n5511 = ~n5153 & ~n5510 ;
  assign n5527 = n5247 & n5427 ;
  assign n5504 = n3506 & n5527 ;
  assign n5502 = n5150 & n5493 ;
  assign n5505 = n5504 ^ n5502 ;
  assign n5506 = n5505 ^ n5150 ;
  assign n5513 = n5511 ^ n5506 ;
  assign n5520 = n5519 ^ n5513 ;
  assign n5521 = ~n1258 & n5520 ;
  assign n5522 = n5521 ^ n5513 ;
  assign n5523 = n5501 & ~n5522 ;
  assign n5525 = x185 & n1530 ;
  assign n5524 = x150 & n2724 ;
  assign n5526 = n5525 ^ n5524 ;
  assign n5528 = n5526 & n5527 ;
  assign n5529 = n5528 ^ n5427 ;
  assign n5530 = n1258 & ~n5529 ;
  assign n5531 = n5163 ^ x135 ;
  assign n5532 = n5531 ^ n5507 ;
  assign n5533 = ~n5153 & n5532 ;
  assign n5534 = n5530 & ~n5533 ;
  assign n5535 = x194 ^ x170 ;
  assign n5540 = n1911 & n5535 ;
  assign n5541 = n5540 ^ x170 ;
  assign n5542 = n5413 & n5541 ;
  assign n5543 = ~n5534 & ~n5542 ;
  assign n5544 = n5501 & n5543 ;
  assign n5546 = x184 & n1530 ;
  assign n5545 = x163 & n2724 ;
  assign n5547 = n5546 ^ n5545 ;
  assign n5548 = ~n3262 & n5247 ;
  assign n5549 = n5547 & n5548 ;
  assign n5550 = n5549 ^ n3262 ;
  assign n5551 = n5255 & n5550 ;
  assign n5552 = x39 & n1258 ;
  assign n5553 = ~n5551 & n5552 ;
  assign n5554 = n3249 & n3750 ;
  assign n5555 = ~n1258 & n2935 ;
  assign n5556 = ~n5554 & n5555 ;
  assign n5557 = n5556 ^ n2935 ;
  assign n5558 = ~n5553 & n5557 ;
  assign n5559 = ~n5228 & n5558 ;
  assign n5566 = n5162 ^ x136 ;
  assign n5567 = n1258 & ~n5157 ;
  assign n5568 = n5566 & n5567 ;
  assign n5562 = n1911 & n3748 ;
  assign n5563 = n5562 ^ x148 ;
  assign n5564 = n5413 & n5563 ;
  assign n5565 = n5564 ^ n1258 ;
  assign n5569 = n5568 ^ n5565 ;
  assign n5570 = ~n2941 & ~n5427 ;
  assign n5571 = n5569 & n5570 ;
  assign n5572 = n5571 ^ n2941 ;
  assign n5573 = ~n5559 & ~n5572 ;
  assign n5575 = ~x210 & n3944 ;
  assign n5574 = ~x198 & n3951 ;
  assign n5576 = n5575 ^ n5574 ;
  assign n5577 = n3249 & n4009 ;
  assign n5578 = n5576 & n5577 ;
  assign n5579 = n5578 ^ x137 ;
  assign n5580 = x39 & n5579 ;
  assign n5581 = n5580 ^ x137 ;
  assign n5582 = n1206 & n3270 ;
  assign n5587 = n2729 & n3528 ;
  assign n5588 = n5587 ^ n3488 ;
  assign n5589 = x39 & n5588 ;
  assign n5590 = n5589 ^ n3488 ;
  assign n5591 = n5582 & n5590 ;
  assign n5592 = n1781 & n3664 ;
  assign n5593 = ~n5591 & n5592 ;
  assign n5599 = ~x195 & ~x196 ;
  assign n5600 = n5599 ^ n3496 ;
  assign n5601 = ~n3497 & n5600 ;
  assign n5594 = x139 ^ x138 ;
  assign n5602 = n5601 ^ n5594 ;
  assign n5603 = n5602 ^ x138 ;
  assign n5606 = n3495 & ~n5603 ;
  assign n5607 = n5606 ^ x138 ;
  assign n5608 = n5593 & n5607 ;
  assign n5609 = n5608 ^ n5554 ;
  assign n5610 = ~n4404 & ~n5609 ;
  assign n5611 = n5610 ^ n5554 ;
  assign n5612 = n3500 ^ n3495 ;
  assign n5613 = n5612 ^ x139 ;
  assign n5614 = n5593 & n5613 ;
  assign n5615 = n5614 ^ n3526 ;
  assign n5616 = n4404 & ~n5615 ;
  assign n5617 = n5616 ^ n5614 ;
  assign n5618 = ~n2647 & n3911 ;
  assign n5619 = ~x841 & n1275 ;
  assign n5620 = n1301 & n5619 ;
  assign n5621 = ~x45 & ~x47 ;
  assign n5622 = ~x102 & n5621 ;
  assign n5623 = ~n3897 & n5622 ;
  assign n5624 = ~n5620 & n5623 ;
  assign n5625 = ~x47 & ~x252 ;
  assign n5626 = ~n1255 & n5625 ;
  assign n5627 = n5626 ^ x252 ;
  assign n5628 = ~n5624 & n5627 ;
  assign n5629 = ~x40 & ~n5628 ;
  assign n5630 = ~n5618 & n5629 ;
  assign n5631 = ~n4383 & n5630 ;
  assign n5632 = ~n4601 & ~n5631 ;
  assign n5638 = ~x120 & ~x287 ;
  assign n5639 = n3920 & n5638 ;
  assign n5640 = n5639 ^ x120 ;
  assign n5653 = n2943 & n5640 ;
  assign n5656 = n5640 ^ n2679 ;
  assign n5654 = ~n3266 & ~n4346 ;
  assign n5655 = n5654 ^ n2943 ;
  assign n5657 = n5656 ^ n5655 ;
  assign n5658 = n5657 ^ n4346 ;
  assign n5660 = n5656 & n5658 ;
  assign n5661 = n5653 & n5660 ;
  assign n5662 = n5661 ^ n5657 ;
  assign n5634 = n3266 ^ n2943 ;
  assign n5652 = n5634 ^ n4346 ;
  assign n5663 = n5662 ^ n5652 ;
  assign n5671 = n5663 ^ n2943 ;
  assign n5672 = n5671 ^ n4346 ;
  assign n5633 = n4346 ^ n3266 ;
  assign n5635 = n5634 ^ n5633 ;
  assign n5644 = n5640 ^ n5635 ;
  assign n5636 = n5635 ^ n2679 ;
  assign n5637 = n5636 ^ n5633 ;
  assign n5666 = n5644 ^ n5637 ;
  assign n5667 = n5666 ^ n5634 ;
  assign n5668 = n5667 ^ n3266 ;
  assign n5673 = n5672 ^ n5668 ;
  assign n5674 = ~n5632 & n5673 ;
  assign n5675 = n2985 & ~n5674 ;
  assign n5676 = x832 & n2985 ;
  assign n5677 = ~n5675 & ~n5676 ;
  assign n5781 = x761 ^ x140 ;
  assign n5678 = x621 & x1091 ;
  assign n5679 = x1157 ^ x630 ;
  assign n5680 = x1158 ^ x626 ;
  assign n5708 = x1154 ^ x618 ;
  assign n5681 = x1155 ^ x609 ;
  assign n5682 = x1156 ^ x629 ;
  assign n5684 = x789 ^ x778 ;
  assign n5683 = x1153 ^ x608 ;
  assign n5685 = n5684 ^ n5683 ;
  assign n5687 = x1159 ^ x619 ;
  assign n5688 = n5687 ^ n5684 ;
  assign n5689 = n5688 ^ n5685 ;
  assign n5690 = x789 & ~n5689 ;
  assign n5691 = n5685 & ~n5690 ;
  assign n5692 = n5685 ^ x778 ;
  assign n5693 = n5692 ^ n5690 ;
  assign n5694 = n5693 ^ x789 ;
  assign n5695 = n5691 & n5694 ;
  assign n5696 = n5695 ^ n5693 ;
  assign n5697 = x792 & ~n5696 ;
  assign n5698 = n5682 & n5697 ;
  assign n5699 = n5698 ^ n5696 ;
  assign n5700 = x1160 ^ x644 ;
  assign n5701 = x603 & x790 ;
  assign n5702 = n5700 & n5701 ;
  assign n5703 = n5702 ^ x603 ;
  assign n5704 = ~n5699 & n5703 ;
  assign n5705 = x785 & n5704 ;
  assign n5706 = n5681 & n5705 ;
  assign n5707 = n5706 ^ n5704 ;
  assign n5709 = x781 & n5707 ;
  assign n5710 = n5708 & n5709 ;
  assign n5711 = n5710 ^ n5707 ;
  assign n5712 = x788 & n5711 ;
  assign n5713 = n5680 & n5712 ;
  assign n5714 = n5713 ^ n5711 ;
  assign n5715 = x787 & n5714 ;
  assign n5716 = n5679 & n5715 ;
  assign n5717 = n5716 ^ n5714 ;
  assign n5718 = n5678 & n5717 ;
  assign n5719 = n5718 ^ n5717 ;
  assign n5722 = x665 & x1091 ;
  assign n5770 = x1154 ^ x627 ;
  assign n5723 = x1157 ^ x647 ;
  assign n5743 = x1155 ^ x660 ;
  assign n5724 = x1153 ^ x625 ;
  assign n5726 = x790 ^ x788 ;
  assign n5725 = x1158 ^ x641 ;
  assign n5727 = n5726 ^ n5725 ;
  assign n5729 = x1160 ^ x715 ;
  assign n5730 = n5729 ^ n5726 ;
  assign n5731 = n5730 ^ n5727 ;
  assign n5732 = x790 & ~n5731 ;
  assign n5733 = n5727 & ~n5732 ;
  assign n5734 = n5727 ^ x788 ;
  assign n5735 = n5734 ^ n5732 ;
  assign n5736 = n5735 ^ x790 ;
  assign n5737 = n5733 & n5736 ;
  assign n5738 = n5737 ^ n5735 ;
  assign n5739 = x680 & ~n5738 ;
  assign n5740 = x778 & n5739 ;
  assign n5741 = n5724 & n5740 ;
  assign n5742 = n5741 ^ n5739 ;
  assign n5744 = x785 & n5742 ;
  assign n5745 = n5743 & n5744 ;
  assign n5746 = n5745 ^ n5742 ;
  assign n5747 = x787 & n5746 ;
  assign n5748 = n5723 & n5747 ;
  assign n5749 = n5748 ^ n5746 ;
  assign n5755 = x1156 ^ x628 ;
  assign n5751 = x792 ^ x789 ;
  assign n5756 = n5755 ^ n5751 ;
  assign n5750 = x1159 ^ x648 ;
  assign n5752 = n5751 ^ n5750 ;
  assign n5757 = n5756 ^ n5752 ;
  assign n5758 = x792 & ~n5757 ;
  assign n5753 = n5752 ^ x789 ;
  assign n5759 = n5758 ^ n5753 ;
  assign n5760 = n5759 ^ x792 ;
  assign n5765 = n5752 & ~n5758 ;
  assign n5766 = n5760 & n5765 ;
  assign n5767 = n5766 ^ n5760 ;
  assign n5768 = n5767 ^ x792 ;
  assign n5769 = n5749 & ~n5768 ;
  assign n5771 = x781 & n5769 ;
  assign n5772 = n5770 & n5771 ;
  assign n5773 = n5772 ^ n5769 ;
  assign n5774 = n5722 & n5773 ;
  assign n5775 = n5774 ^ n5773 ;
  assign n5778 = ~x738 & n5775 ;
  assign n5779 = n5778 ^ x761 ;
  assign n5780 = ~n5719 & ~n5779 ;
  assign n5782 = n5781 ^ n5780 ;
  assign n5783 = ~n5677 & n5782 ;
  assign n5784 = n5783 ^ x140 ;
  assign n5792 = x749 ^ x141 ;
  assign n5789 = x706 & n5775 ;
  assign n5790 = n5789 ^ x749 ;
  assign n5791 = ~n5719 & n5790 ;
  assign n5793 = n5792 ^ n5791 ;
  assign n5794 = ~n5677 & ~n5793 ;
  assign n5795 = n5794 ^ x141 ;
  assign n5803 = x743 ^ x142 ;
  assign n5800 = x735 & n5775 ;
  assign n5801 = n5800 ^ x743 ;
  assign n5802 = ~n5719 & n5801 ;
  assign n5804 = n5803 ^ n5802 ;
  assign n5805 = ~n5677 & n5804 ;
  assign n5806 = n5805 ^ x142 ;
  assign n5814 = x774 ^ x143 ;
  assign n5811 = x687 & n5775 ;
  assign n5812 = n5811 ^ x774 ;
  assign n5813 = ~n5719 & ~n5812 ;
  assign n5815 = n5814 ^ n5813 ;
  assign n5816 = ~n5677 & n5815 ;
  assign n5817 = n5816 ^ x143 ;
  assign n5825 = x758 ^ x144 ;
  assign n5822 = x736 & n5775 ;
  assign n5823 = n5822 ^ x758 ;
  assign n5824 = ~n5719 & n5823 ;
  assign n5826 = n5825 ^ n5824 ;
  assign n5827 = ~n5677 & n5826 ;
  assign n5828 = n5827 ^ x144 ;
  assign n5836 = x767 ^ x145 ;
  assign n5833 = ~x698 & n5775 ;
  assign n5834 = n5833 ^ x767 ;
  assign n5835 = ~n5719 & ~n5834 ;
  assign n5837 = n5836 ^ n5835 ;
  assign n5838 = ~n5677 & n5837 ;
  assign n5839 = n5838 ^ x145 ;
  assign n5845 = x743 ^ x146 ;
  assign n5842 = x735 & x907 ;
  assign n5843 = n5842 ^ x743 ;
  assign n5844 = ~x947 & n5843 ;
  assign n5846 = n5845 ^ n5844 ;
  assign n5847 = ~n5677 & n5846 ;
  assign n5848 = n5847 ^ x146 ;
  assign n5856 = x770 ^ x147 ;
  assign n5853 = x726 & x907 ;
  assign n5854 = n5853 ^ x770 ;
  assign n5855 = ~x947 & ~n5854 ;
  assign n5857 = n5856 ^ n5855 ;
  assign n5858 = ~n5677 & n5857 ;
  assign n5859 = n5858 ^ x147 ;
  assign n5865 = x749 ^ x148 ;
  assign n5862 = x706 & x907 ;
  assign n5863 = n5862 ^ x749 ;
  assign n5864 = ~x947 & n5863 ;
  assign n5866 = n5865 ^ n5864 ;
  assign n5867 = ~n5677 & ~n5866 ;
  assign n5868 = n5867 ^ x148 ;
  assign n5892 = ~x149 & n5677 ;
  assign n5869 = n2985 & ~n5632 ;
  assign n5870 = n3263 & n3558 ;
  assign n5871 = n2943 & ~n5870 ;
  assign n5872 = n1537 & n2668 ;
  assign n5873 = n5871 & n5872 ;
  assign n5874 = n5873 ^ n5871 ;
  assign n5878 = n5874 ^ n2943 ;
  assign n5875 = n5640 & n5874 ;
  assign n5876 = n5870 ^ n2670 ;
  assign n5877 = n5875 & ~n5876 ;
  assign n5879 = n5878 ^ n5877 ;
  assign n5880 = n5869 & ~n5879 ;
  assign n5881 = n5880 ^ n2985 ;
  assign n5882 = ~n5676 & ~n5881 ;
  assign n5887 = ~x725 & x907 ;
  assign n5888 = n5887 ^ x755 ;
  assign n5889 = ~x947 & ~n5888 ;
  assign n5890 = n5889 ^ x755 ;
  assign n5891 = ~n5882 & ~n5890 ;
  assign n5894 = n5892 ^ n5891 ;
  assign n5904 = ~x150 & n5677 ;
  assign n5899 = ~x701 & x907 ;
  assign n5900 = n5899 ^ x751 ;
  assign n5901 = ~x947 & ~n5900 ;
  assign n5902 = n5901 ^ x751 ;
  assign n5903 = ~n5882 & ~n5902 ;
  assign n5906 = n5904 ^ n5903 ;
  assign n5914 = x745 ^ x151 ;
  assign n5911 = ~x723 & x907 ;
  assign n5912 = n5911 ^ x745 ;
  assign n5913 = ~x947 & ~n5912 ;
  assign n5915 = n5914 ^ n5913 ;
  assign n5916 = ~n5677 & n5915 ;
  assign n5917 = n5916 ^ x151 ;
  assign n5925 = x759 ^ x152 ;
  assign n5922 = x696 & x907 ;
  assign n5923 = n5922 ^ x759 ;
  assign n5924 = ~x947 & n5923 ;
  assign n5926 = n5925 ^ n5924 ;
  assign n5927 = ~n5677 & n5926 ;
  assign n5928 = n5927 ^ x152 ;
  assign n5936 = x766 ^ x153 ;
  assign n5933 = x700 & x907 ;
  assign n5934 = n5933 ^ x766 ;
  assign n5935 = ~x947 & n5934 ;
  assign n5937 = n5936 ^ n5935 ;
  assign n5938 = ~n5677 & ~n5937 ;
  assign n5939 = n5938 ^ x153 ;
  assign n5949 = ~x154 & n5677 ;
  assign n5944 = ~x704 & x907 ;
  assign n5945 = n5944 ^ x742 ;
  assign n5946 = ~x947 & ~n5945 ;
  assign n5947 = n5946 ^ x742 ;
  assign n5948 = ~n5882 & ~n5947 ;
  assign n5951 = n5949 ^ n5948 ;
  assign n5961 = ~x155 & n5677 ;
  assign n5956 = ~x686 & x907 ;
  assign n5957 = n5956 ^ x757 ;
  assign n5958 = ~x947 & ~n5957 ;
  assign n5959 = n5958 ^ x757 ;
  assign n5960 = ~n5882 & ~n5959 ;
  assign n5963 = n5961 ^ n5960 ;
  assign n5973 = ~x156 & n5677 ;
  assign n5968 = ~x724 & x907 ;
  assign n5969 = n5968 ^ x741 ;
  assign n5970 = ~x947 & ~n5969 ;
  assign n5971 = n5970 ^ x741 ;
  assign n5972 = ~n5882 & ~n5971 ;
  assign n5975 = n5973 ^ n5972 ;
  assign n5983 = x760 ^ x157 ;
  assign n5980 = ~x688 & x907 ;
  assign n5981 = n5980 ^ x760 ;
  assign n5982 = ~x947 & ~n5981 ;
  assign n5984 = n5983 ^ n5982 ;
  assign n5985 = ~n5677 & n5984 ;
  assign n5986 = n5985 ^ x157 ;
  assign n5996 = ~x158 & n5677 ;
  assign n5991 = ~x702 & x907 ;
  assign n5992 = n5991 ^ x753 ;
  assign n5993 = ~x947 & ~n5992 ;
  assign n5994 = n5993 ^ x753 ;
  assign n5995 = ~n5882 & ~n5994 ;
  assign n5998 = n5996 ^ n5995 ;
  assign n6006 = x754 ^ x159 ;
  assign n6003 = ~x709 & x907 ;
  assign n6004 = n6003 ^ x754 ;
  assign n6005 = ~x947 & ~n6004 ;
  assign n6007 = n6006 ^ n6005 ;
  assign n6008 = ~n5677 & n6007 ;
  assign n6009 = n6008 ^ x159 ;
  assign n6017 = x756 ^ x160 ;
  assign n6014 = ~x734 & x907 ;
  assign n6015 = n6014 ^ x756 ;
  assign n6016 = ~x947 & ~n6015 ;
  assign n6018 = n6017 ^ n6016 ;
  assign n6019 = ~n5677 & n6018 ;
  assign n6020 = n6019 ^ x160 ;
  assign n6026 = x758 ^ x161 ;
  assign n6023 = x736 & x907 ;
  assign n6024 = n6023 ^ x758 ;
  assign n6025 = ~x947 & n6024 ;
  assign n6027 = n6026 ^ n6025 ;
  assign n6028 = ~n5677 & n6027 ;
  assign n6029 = n6028 ^ x161 ;
  assign n6035 = x761 ^ x162 ;
  assign n6032 = ~x738 & x907 ;
  assign n6033 = n6032 ^ x761 ;
  assign n6034 = ~x947 & ~n6033 ;
  assign n6036 = n6035 ^ n6034 ;
  assign n6037 = ~n5677 & n6036 ;
  assign n6038 = n6037 ^ x162 ;
  assign n6046 = x777 ^ x163 ;
  assign n6043 = ~x737 & x907 ;
  assign n6044 = n6043 ^ x777 ;
  assign n6045 = ~x947 & ~n6044 ;
  assign n6047 = n6046 ^ n6045 ;
  assign n6048 = ~n5677 & n6047 ;
  assign n6049 = n6048 ^ x163 ;
  assign n6057 = x752 ^ x164 ;
  assign n6054 = x703 & x907 ;
  assign n6055 = n6054 ^ x752 ;
  assign n6056 = ~x947 & ~n6055 ;
  assign n6058 = n6057 ^ n6056 ;
  assign n6059 = ~n5677 & n6058 ;
  assign n6060 = n6059 ^ x164 ;
  assign n6068 = ~x165 & n5677 ;
  assign n6063 = x687 & x907 ;
  assign n6064 = n6063 ^ x774 ;
  assign n6065 = ~x947 & ~n6064 ;
  assign n6066 = n6065 ^ x774 ;
  assign n6067 = ~n5882 & ~n6066 ;
  assign n6070 = n6068 ^ n6067 ;
  assign n6078 = x772 ^ x166 ;
  assign n6075 = x727 & x907 ;
  assign n6076 = n6075 ^ x772 ;
  assign n6077 = ~x947 & n6076 ;
  assign n6079 = n6078 ^ n6077 ;
  assign n6080 = ~n5677 & n6079 ;
  assign n6081 = n6080 ^ x166 ;
  assign n6089 = x768 ^ x167 ;
  assign n6086 = x705 & x907 ;
  assign n6087 = n6086 ^ x768 ;
  assign n6088 = ~x947 & ~n6087 ;
  assign n6090 = n6089 ^ n6088 ;
  assign n6091 = ~n5677 & n6090 ;
  assign n6092 = n6091 ^ x167 ;
  assign n6100 = x763 ^ x168 ;
  assign n6097 = x699 & x907 ;
  assign n6098 = n6097 ^ x763 ;
  assign n6099 = ~x947 & n6098 ;
  assign n6101 = n6100 ^ n6099 ;
  assign n6102 = ~n5677 & ~n6101 ;
  assign n6103 = n6102 ^ x168 ;
  assign n6111 = x746 ^ x169 ;
  assign n6108 = x729 & x907 ;
  assign n6109 = n6108 ^ x746 ;
  assign n6110 = ~x947 & n6109 ;
  assign n6112 = n6111 ^ n6110 ;
  assign n6113 = ~n5677 & ~n6112 ;
  assign n6114 = n6113 ^ x169 ;
  assign n6122 = x748 ^ x170 ;
  assign n6119 = x730 & x907 ;
  assign n6120 = n6119 ^ x748 ;
  assign n6121 = ~x947 & n6120 ;
  assign n6123 = n6122 ^ n6121 ;
  assign n6124 = ~n5677 & ~n6123 ;
  assign n6125 = n6124 ^ x170 ;
  assign n6133 = x764 ^ x171 ;
  assign n6130 = x691 & x907 ;
  assign n6131 = n6130 ^ x764 ;
  assign n6132 = ~x947 & n6131 ;
  assign n6134 = n6133 ^ n6132 ;
  assign n6135 = ~n5677 & ~n6134 ;
  assign n6136 = n6135 ^ x171 ;
  assign n6144 = x739 ^ x172 ;
  assign n6141 = x690 & x907 ;
  assign n6142 = n6141 ^ x739 ;
  assign n6143 = ~x947 & n6142 ;
  assign n6145 = n6144 ^ n6143 ;
  assign n6146 = ~n5677 & ~n6145 ;
  assign n6147 = n6146 ^ x172 ;
  assign n6153 = x745 ^ x173 ;
  assign n6150 = ~x723 & n5775 ;
  assign n6151 = n6150 ^ x745 ;
  assign n6152 = ~n5719 & ~n6151 ;
  assign n6154 = n6153 ^ n6152 ;
  assign n6155 = ~n5677 & n6154 ;
  assign n6156 = n6155 ^ x173 ;
  assign n6162 = x759 ^ x174 ;
  assign n6159 = x696 & n5775 ;
  assign n6160 = n6159 ^ x759 ;
  assign n6161 = ~n5719 & n6160 ;
  assign n6163 = n6162 ^ n6161 ;
  assign n6164 = ~n5677 & n6163 ;
  assign n6165 = n6164 ^ x174 ;
  assign n6171 = x766 ^ x175 ;
  assign n6168 = x700 & n5775 ;
  assign n6169 = n6168 ^ x766 ;
  assign n6170 = ~n5719 & n6169 ;
  assign n6172 = n6171 ^ n6170 ;
  assign n6173 = ~n5677 & ~n6172 ;
  assign n6174 = n6173 ^ x175 ;
  assign n6180 = x742 ^ x176 ;
  assign n6177 = ~x704 & n5775 ;
  assign n6178 = n6177 ^ x742 ;
  assign n6179 = ~n5719 & ~n6178 ;
  assign n6181 = n6180 ^ n6179 ;
  assign n6182 = ~n5677 & n6181 ;
  assign n6183 = n6182 ^ x176 ;
  assign n6189 = x757 ^ x177 ;
  assign n6186 = ~x686 & n5775 ;
  assign n6187 = n6186 ^ x757 ;
  assign n6188 = ~n5719 & ~n6187 ;
  assign n6190 = n6189 ^ n6188 ;
  assign n6191 = ~n5677 & n6190 ;
  assign n6192 = n6191 ^ x177 ;
  assign n6198 = x760 ^ x178 ;
  assign n6195 = ~x688 & n5775 ;
  assign n6196 = n6195 ^ x760 ;
  assign n6197 = ~n5719 & ~n6196 ;
  assign n6199 = n6198 ^ n6197 ;
  assign n6200 = ~n5677 & n6199 ;
  assign n6201 = n6200 ^ x178 ;
  assign n6207 = x741 ^ x179 ;
  assign n6204 = ~x724 & n5775 ;
  assign n6205 = n6204 ^ x741 ;
  assign n6206 = ~n5719 & ~n6205 ;
  assign n6208 = n6207 ^ n6206 ;
  assign n6209 = ~n5677 & n6208 ;
  assign n6210 = n6209 ^ x179 ;
  assign n6216 = x753 ^ x180 ;
  assign n6213 = ~x702 & n5775 ;
  assign n6214 = n6213 ^ x753 ;
  assign n6215 = ~n5719 & ~n6214 ;
  assign n6217 = n6216 ^ n6215 ;
  assign n6218 = ~n5677 & n6217 ;
  assign n6219 = n6218 ^ x180 ;
  assign n6225 = x754 ^ x181 ;
  assign n6222 = ~x709 & n5775 ;
  assign n6223 = n6222 ^ x754 ;
  assign n6224 = ~n5719 & ~n6223 ;
  assign n6226 = n6225 ^ n6224 ;
  assign n6227 = ~n5677 & n6226 ;
  assign n6228 = n6227 ^ x181 ;
  assign n6234 = x756 ^ x182 ;
  assign n6231 = ~x734 & n5775 ;
  assign n6232 = n6231 ^ x756 ;
  assign n6233 = ~n5719 & ~n6232 ;
  assign n6235 = n6234 ^ n6233 ;
  assign n6236 = ~n5677 & n6235 ;
  assign n6237 = n6236 ^ x182 ;
  assign n6243 = x755 ^ x183 ;
  assign n6240 = ~x725 & n5775 ;
  assign n6241 = n6240 ^ x755 ;
  assign n6242 = ~n5719 & ~n6241 ;
  assign n6244 = n6243 ^ n6242 ;
  assign n6245 = ~n5677 & n6244 ;
  assign n6246 = n6245 ^ x183 ;
  assign n6252 = x777 ^ x184 ;
  assign n6249 = ~x737 & n5775 ;
  assign n6250 = n6249 ^ x777 ;
  assign n6251 = ~n5719 & ~n6250 ;
  assign n6253 = n6252 ^ n6251 ;
  assign n6254 = ~n5677 & n6253 ;
  assign n6255 = n6254 ^ x184 ;
  assign n6261 = x751 ^ x185 ;
  assign n6258 = ~x701 & n5775 ;
  assign n6259 = n6258 ^ x751 ;
  assign n6260 = ~n5719 & ~n6259 ;
  assign n6262 = n6261 ^ n6260 ;
  assign n6263 = ~n5677 & n6262 ;
  assign n6264 = n6263 ^ x185 ;
  assign n6270 = x752 ^ x186 ;
  assign n6267 = x703 & n5775 ;
  assign n6268 = n6267 ^ x752 ;
  assign n6269 = ~n5719 & ~n6268 ;
  assign n6271 = n6270 ^ n6269 ;
  assign n6272 = ~n5677 & n6271 ;
  assign n6273 = n6272 ^ x186 ;
  assign n6279 = x770 ^ x187 ;
  assign n6276 = x726 & n5775 ;
  assign n6277 = n6276 ^ x770 ;
  assign n6278 = ~n5719 & ~n6277 ;
  assign n6280 = n6279 ^ n6278 ;
  assign n6281 = ~n5677 & n6280 ;
  assign n6282 = n6281 ^ x187 ;
  assign n6288 = x768 ^ x188 ;
  assign n6285 = x705 & n5775 ;
  assign n6286 = n6285 ^ x768 ;
  assign n6287 = ~n5719 & ~n6286 ;
  assign n6289 = n6288 ^ n6287 ;
  assign n6290 = ~n5677 & n6289 ;
  assign n6291 = n6290 ^ x188 ;
  assign n6297 = x772 ^ x189 ;
  assign n6294 = x727 & n5775 ;
  assign n6295 = n6294 ^ x772 ;
  assign n6296 = ~n5719 & n6295 ;
  assign n6298 = n6297 ^ n6296 ;
  assign n6299 = ~n5677 & n6298 ;
  assign n6300 = n6299 ^ x189 ;
  assign n6306 = x763 ^ x190 ;
  assign n6303 = x699 & n5775 ;
  assign n6304 = n6303 ^ x763 ;
  assign n6305 = ~n5719 & n6304 ;
  assign n6307 = n6306 ^ n6305 ;
  assign n6308 = ~n5677 & ~n6307 ;
  assign n6309 = n6308 ^ x190 ;
  assign n6315 = x746 ^ x191 ;
  assign n6312 = x729 & n5775 ;
  assign n6313 = n6312 ^ x746 ;
  assign n6314 = ~n5719 & n6313 ;
  assign n6316 = n6315 ^ n6314 ;
  assign n6317 = ~n5677 & ~n6316 ;
  assign n6318 = n6317 ^ x191 ;
  assign n6324 = x764 ^ x192 ;
  assign n6321 = x691 & n5775 ;
  assign n6322 = n6321 ^ x764 ;
  assign n6323 = ~n5719 & n6322 ;
  assign n6325 = n6324 ^ n6323 ;
  assign n6326 = ~n5677 & ~n6325 ;
  assign n6327 = n6326 ^ x192 ;
  assign n6333 = x739 ^ x193 ;
  assign n6330 = x690 & n5775 ;
  assign n6331 = n6330 ^ x739 ;
  assign n6332 = ~n5719 & n6331 ;
  assign n6334 = n6333 ^ n6332 ;
  assign n6335 = ~n5677 & ~n6334 ;
  assign n6336 = n6335 ^ x193 ;
  assign n6342 = x748 ^ x194 ;
  assign n6339 = x730 & n5775 ;
  assign n6340 = n6339 ^ x748 ;
  assign n6341 = ~n5719 & n6340 ;
  assign n6343 = n6342 ^ n6341 ;
  assign n6344 = ~n5677 & ~n6343 ;
  assign n6345 = n6344 ^ x194 ;
  assign n6353 = n3499 ^ x195 ;
  assign n6354 = n6353 ^ n3500 ;
  assign n6359 = ~n5593 & n6354 ;
  assign n6350 = ~x299 & n5514 ;
  assign n6351 = n6350 ^ x171 ;
  assign n6352 = n3249 & n6351 ;
  assign n6355 = n6354 ^ n6352 ;
  assign n6360 = n6359 ^ n6355 ;
  assign n6361 = ~n4404 & ~n6360 ;
  assign n6362 = n6361 ^ n6352 ;
  assign n6368 = n3500 ^ n3498 ;
  assign n6369 = n6368 ^ x196 ;
  assign n6370 = n5593 & n6369 ;
  assign n6365 = x299 & n5535 ;
  assign n6366 = n6365 ^ x194 ;
  assign n6367 = n3249 & n6366 ;
  assign n6371 = n6370 ^ n6367 ;
  assign n6372 = n4404 & ~n6371 ;
  assign n6373 = n6372 ^ n6370 ;
  assign n6379 = x767 ^ x197 ;
  assign n6376 = ~x698 & x907 ;
  assign n6377 = n6376 ^ x767 ;
  assign n6378 = ~x947 & ~n6377 ;
  assign n6380 = n6379 ^ n6378 ;
  assign n6381 = ~n5677 & n6380 ;
  assign n6382 = n6381 ^ x197 ;
  assign n6390 = x633 ^ x198 ;
  assign n6387 = x634 & n5775 ;
  assign n6388 = n6387 ^ x633 ;
  assign n6389 = ~n5719 & n6388 ;
  assign n6391 = n6390 ^ n6389 ;
  assign n6392 = n5675 & n6391 ;
  assign n6393 = n6392 ^ x198 ;
  assign n6401 = x617 ^ x199 ;
  assign n6398 = x637 & n5775 ;
  assign n6399 = n6398 ^ x617 ;
  assign n6400 = ~n5719 & n6399 ;
  assign n6402 = n6401 ^ n6400 ;
  assign n6403 = n5675 & n6402 ;
  assign n6404 = n6403 ^ x199 ;
  assign n6412 = x606 ^ x200 ;
  assign n6409 = x643 & n5775 ;
  assign n6410 = n6409 ^ x606 ;
  assign n6411 = ~n5719 & n6410 ;
  assign n6413 = n6412 ^ n6411 ;
  assign n6414 = n5675 & n6413 ;
  assign n6415 = n6414 ^ x200 ;
  assign n6416 = n1268 & n4151 ;
  assign n6417 = ~x332 & ~n1767 ;
  assign n6418 = ~n6416 & n6417 ;
  assign n6419 = x70 ^ x32 ;
  assign n6420 = x841 ^ x96 ;
  assign n6421 = x70 & ~n6420 ;
  assign n6422 = n6421 ^ x841 ;
  assign n6423 = n1549 & ~n1911 ;
  assign n6424 = n6423 ^ x198 ;
  assign n6425 = n6424 ^ x70 ;
  assign n6426 = n6425 ^ n6419 ;
  assign n6427 = ~n6422 & n6426 ;
  assign n6428 = n6427 ^ x70 ;
  assign n6429 = n6419 & n6428 ;
  assign n6430 = ~x233 & n6429 ;
  assign n6431 = n6430 ^ n6429 ;
  assign n6432 = ~x237 & n6431 ;
  assign n6433 = n6432 ^ n6431 ;
  assign n6434 = n6418 & ~n6433 ;
  assign n6435 = x947 ^ x587 ;
  assign n6436 = n1911 & n2635 ;
  assign n6437 = n6435 & n6436 ;
  assign n6438 = n6437 ^ n2860 ;
  assign n6439 = ~x332 & ~n6438 ;
  assign n6440 = x96 & n6424 ;
  assign n6441 = ~x237 & n6440 ;
  assign n6442 = n6441 ^ n6440 ;
  assign n6443 = ~x233 & n6438 ;
  assign n6444 = n6443 ^ n6438 ;
  assign n6445 = n6442 & n6444 ;
  assign n6446 = ~x201 & ~n6445 ;
  assign n6447 = ~n6439 & n6446 ;
  assign n6448 = ~n6434 & n6447 ;
  assign n6449 = n6448 ^ n6446 ;
  assign n6450 = n6449 ^ n6445 ;
  assign n6451 = ~x237 & n6430 ;
  assign n6452 = n6451 ^ n6430 ;
  assign n6453 = n6418 & ~n6452 ;
  assign n6454 = n6442 & n6443 ;
  assign n6455 = ~x202 & ~n6454 ;
  assign n6456 = ~n6453 & n6455 ;
  assign n6457 = ~n6439 & n6456 ;
  assign n6458 = n6457 ^ n6455 ;
  assign n6459 = n6458 ^ n6454 ;
  assign n6460 = n6418 & ~n6451 ;
  assign n6461 = n6441 & n6443 ;
  assign n6462 = ~x203 & ~n6461 ;
  assign n6463 = ~n6460 & n6462 ;
  assign n6464 = ~n6439 & n6463 ;
  assign n6465 = n6464 ^ n6462 ;
  assign n6466 = n6465 ^ n6461 ;
  assign n6468 = n2654 ^ x602 ;
  assign n6467 = n2654 ^ x907 ;
  assign n6469 = n6468 ^ n6467 ;
  assign n6472 = n1911 & n6469 ;
  assign n6473 = n6472 ^ n6467 ;
  assign n6474 = n2635 & n6473 ;
  assign n6475 = n6474 ^ n2654 ;
  assign n6476 = ~x332 & ~n6475 ;
  assign n6477 = n6442 & n6475 ;
  assign n6478 = ~x233 & n6477 ;
  assign n6479 = n6478 ^ n6477 ;
  assign n6480 = ~x204 & ~n6479 ;
  assign n6481 = ~n6476 & n6480 ;
  assign n6482 = ~n6434 & n6481 ;
  assign n6483 = n6482 ^ n6480 ;
  assign n6484 = n6483 ^ n6479 ;
  assign n6485 = ~x205 & ~n6478 ;
  assign n6486 = ~n6476 & n6485 ;
  assign n6487 = ~n6453 & n6486 ;
  assign n6488 = n6487 ^ n6485 ;
  assign n6489 = n6488 ^ n6478 ;
  assign n6490 = n6418 & ~n6432 ;
  assign n6491 = n6441 & n6475 ;
  assign n6492 = ~x233 & n6491 ;
  assign n6493 = n6492 ^ n6491 ;
  assign n6494 = ~x206 & ~n6493 ;
  assign n6495 = ~n6490 & n6494 ;
  assign n6496 = ~n6476 & n6495 ;
  assign n6497 = n6496 ^ n6494 ;
  assign n6498 = n6497 ^ n6493 ;
  assign n6506 = x623 ^ x207 ;
  assign n6503 = x710 & n5775 ;
  assign n6504 = n6503 ^ x623 ;
  assign n6505 = ~n5719 & n6504 ;
  assign n6507 = n6506 ^ n6505 ;
  assign n6508 = n5675 & ~n6507 ;
  assign n6509 = n6508 ^ x207 ;
  assign n6517 = x607 ^ x208 ;
  assign n6514 = x638 & n5775 ;
  assign n6515 = n6514 ^ x607 ;
  assign n6516 = ~n5719 & n6515 ;
  assign n6518 = n6517 ^ n6516 ;
  assign n6519 = n5675 & ~n6518 ;
  assign n6520 = n6519 ^ x208 ;
  assign n6528 = x622 ^ x209 ;
  assign n6525 = x639 & n5775 ;
  assign n6526 = n6525 ^ x622 ;
  assign n6527 = ~n5719 & n6526 ;
  assign n6529 = n6528 ^ n6527 ;
  assign n6530 = n5675 & ~n6529 ;
  assign n6531 = n6530 ^ x209 ;
  assign n6537 = x633 ^ x210 ;
  assign n6534 = x634 & x907 ;
  assign n6535 = n6534 ^ x633 ;
  assign n6536 = ~x947 & n6535 ;
  assign n6538 = n6537 ^ n6536 ;
  assign n6539 = n5675 & n6538 ;
  assign n6540 = n6539 ^ x210 ;
  assign n6546 = x606 ^ x211 ;
  assign n6543 = x643 & x907 ;
  assign n6544 = n6543 ^ x606 ;
  assign n6545 = ~x947 & n6544 ;
  assign n6547 = n6546 ^ n6545 ;
  assign n6548 = n5675 & n6547 ;
  assign n6549 = n6548 ^ x211 ;
  assign n6557 = ~x212 & ~n5675 ;
  assign n6552 = x638 & x907 ;
  assign n6553 = n6552 ^ x607 ;
  assign n6554 = ~x947 & n6553 ;
  assign n6555 = n6554 ^ x607 ;
  assign n6556 = n5881 & n6555 ;
  assign n6559 = n6557 ^ n6556 ;
  assign n6567 = ~x213 & ~n5675 ;
  assign n6562 = x639 & x907 ;
  assign n6563 = n6562 ^ x622 ;
  assign n6564 = ~x947 & n6563 ;
  assign n6565 = n6564 ^ x622 ;
  assign n6566 = n5881 & n6565 ;
  assign n6569 = n6567 ^ n6566 ;
  assign n6575 = x623 ^ x214 ;
  assign n6572 = x710 & x907 ;
  assign n6573 = n6572 ^ x623 ;
  assign n6574 = ~x947 & n6573 ;
  assign n6576 = n6575 ^ n6574 ;
  assign n6577 = n5675 & ~n6576 ;
  assign n6578 = n6577 ^ x214 ;
  assign n6586 = x642 ^ x215 ;
  assign n6583 = x681 & x907 ;
  assign n6584 = n6583 ^ x642 ;
  assign n6585 = ~x947 & n6584 ;
  assign n6587 = n6586 ^ n6585 ;
  assign n6588 = n5675 & n6587 ;
  assign n6589 = n6588 ^ x215 ;
  assign n6597 = x614 ^ x216 ;
  assign n6594 = x662 & x907 ;
  assign n6595 = n6594 ^ x614 ;
  assign n6596 = ~x947 & n6595 ;
  assign n6598 = n6597 ^ n6596 ;
  assign n6599 = n5675 & n6598 ;
  assign n6600 = n6599 ^ x216 ;
  assign n6608 = x612 ^ x217 ;
  assign n6605 = ~x695 & n5775 ;
  assign n6606 = n6605 ^ x612 ;
  assign n6607 = ~n5719 & n6606 ;
  assign n6609 = n6608 ^ n6607 ;
  assign n6610 = n5675 & ~n6609 ;
  assign n6611 = n6610 ^ x217 ;
  assign n6612 = ~x218 & ~n6492 ;
  assign n6613 = ~n6476 & n6612 ;
  assign n6614 = ~n6460 & n6613 ;
  assign n6615 = n6614 ^ n6612 ;
  assign n6616 = n6615 ^ n6492 ;
  assign n6624 = x219 & ~n5675 ;
  assign n6619 = x637 & x907 ;
  assign n6620 = n6619 ^ x617 ;
  assign n6621 = ~x947 & n6620 ;
  assign n6622 = n6621 ^ x617 ;
  assign n6623 = n5881 & n6622 ;
  assign n6626 = n6624 ^ n6623 ;
  assign n6627 = n6441 & n6444 ;
  assign n6628 = ~x220 & ~n6627 ;
  assign n6629 = ~n6490 & n6628 ;
  assign n6630 = ~n6439 & n6629 ;
  assign n6631 = n6630 ^ n6628 ;
  assign n6632 = n6631 ^ n6627 ;
  assign n6640 = x616 ^ x221 ;
  assign n6637 = x661 & x907 ;
  assign n6638 = n6637 ^ x616 ;
  assign n6639 = ~x947 & n6638 ;
  assign n6641 = n6640 ^ n6639 ;
  assign n6642 = n5675 & n6641 ;
  assign n6643 = n6642 ^ x221 ;
  assign n6649 = x616 ^ x222 ;
  assign n6646 = x661 & n5775 ;
  assign n6647 = n6646 ^ x616 ;
  assign n6648 = ~n5719 & n6647 ;
  assign n6650 = n6649 ^ n6648 ;
  assign n6651 = n5675 & n6650 ;
  assign n6652 = n6651 ^ x222 ;
  assign n6658 = x642 ^ x223 ;
  assign n6655 = x681 & n5775 ;
  assign n6656 = n6655 ^ x642 ;
  assign n6657 = ~n5719 & n6656 ;
  assign n6659 = n6658 ^ n6657 ;
  assign n6660 = n5675 & n6659 ;
  assign n6661 = n6660 ^ x223 ;
  assign n6667 = x614 ^ x224 ;
  assign n6664 = x662 & n5775 ;
  assign n6665 = n6664 ^ x614 ;
  assign n6666 = ~n5719 & n6665 ;
  assign n6668 = n6667 ^ n6666 ;
  assign n6669 = n5675 & n6668 ;
  assign n6670 = n6669 ^ x224 ;
  assign n6671 = n1220 & n1627 ;
  assign n6672 = ~n1639 & n1971 ;
  assign n6673 = x70 & n6672 ;
  assign n6674 = x332 & n6673 ;
  assign n6675 = n6674 ^ n6672 ;
  assign n6676 = n6675 ^ n1971 ;
  assign n6677 = ~x55 & ~x137 ;
  assign n6678 = ~n1799 & n6677 ;
  assign n6686 = n1563 & n6678 ;
  assign n6687 = n5017 & n6686 ;
  assign n6688 = n6687 ^ n5017 ;
  assign n6679 = n6678 ^ n1799 ;
  assign n6680 = n6679 ^ n5017 ;
  assign n6689 = n6688 ^ n6680 ;
  assign n6690 = ~n6676 & n6689 ;
  assign n6691 = ~n6671 & n6690 ;
  assign n6697 = n1971 & n2623 ;
  assign n6694 = n1780 & ~n1786 ;
  assign n6692 = x479 & n4714 ;
  assign n6693 = n6692 ^ n1798 ;
  assign n6696 = n6694 ^ n6693 ;
  assign n6699 = n6697 ^ n6696 ;
  assign n6700 = n6699 ^ x231 ;
  assign n6701 = ~x228 & n6700 ;
  assign n6702 = n6701 ^ x231 ;
  assign n6703 = x1093 & n3874 ;
  assign n6704 = n1337 & n1614 ;
  assign n6705 = ~x58 & n6704 ;
  assign n6706 = n6705 ^ x72 ;
  assign n6707 = ~x72 & ~n6706 ;
  assign n6708 = n4073 & n6707 ;
  assign n6709 = ~n6703 & n6708 ;
  assign n6710 = n1971 & ~n6709 ;
  assign n6711 = ~n4379 & ~n6710 ;
  assign n6712 = x36 & n1571 ;
  assign n6713 = ~n6711 & ~n6712 ;
  assign n6714 = n1209 & n1216 ;
  assign n6715 = n1576 ^ n1566 ;
  assign n6716 = n6714 & n6715 ;
  assign n6717 = n1585 & n6716 ;
  assign n6718 = ~x228 & ~n6717 ;
  assign n6719 = ~x39 & ~n6718 ;
  assign n6720 = x1091 & n4717 ;
  assign n6721 = ~n6719 & ~n6720 ;
  assign n6722 = ~x47 & ~n2640 ;
  assign n6723 = n1259 & n6722 ;
  assign n6724 = ~n3528 & n6723 ;
  assign n6725 = ~n5674 & ~n6724 ;
  assign n6726 = ~x64 & n3490 ;
  assign n6727 = x102 ^ x65 ;
  assign n6728 = n6726 & n6727 ;
  assign n6729 = n1372 & n6728 ;
  assign n6730 = ~n3843 & ~n6729 ;
  assign n6731 = ~n2760 & n6730 ;
  assign n6732 = ~n1799 & ~n4317 ;
  assign n6733 = ~n6731 & ~n6732 ;
  assign n6734 = x209 & n1911 ;
  assign n6735 = n6734 ^ n1911 ;
  assign n6759 = x1155 & ~n4366 ;
  assign n6758 = x1153 & n4013 ;
  assign n6760 = n6759 ^ n6758 ;
  assign n6757 = x1154 & n4031 ;
  assign n6761 = n6760 ^ n6757 ;
  assign n6762 = x208 & n6761 ;
  assign n6736 = x1156 ^ x1155 ;
  assign n6737 = x200 & n6736 ;
  assign n6738 = n6737 ^ x1155 ;
  assign n6748 = n6738 ^ n6736 ;
  assign n6749 = ~x199 & n6748 ;
  assign n6747 = x1154 & n4013 ;
  assign n6750 = n6749 ^ n6747 ;
  assign n6743 = ~x200 & x1157 ;
  assign n6744 = n6743 ^ n6738 ;
  assign n6745 = ~n4030 & n6744 ;
  assign n6746 = n6745 ^ n6738 ;
  assign n6751 = n6750 ^ n6746 ;
  assign n6752 = x207 & n6751 ;
  assign n6753 = n6752 ^ n6750 ;
  assign n6763 = n6762 ^ n6753 ;
  assign n6830 = n4014 ^ x208 ;
  assign n7061 = n6830 ^ n4015 ;
  assign n6764 = n6763 & ~n7061 ;
  assign n6765 = n6764 ^ n6753 ;
  assign n6766 = n6735 & n6765 ;
  assign n6767 = n6766 ^ n6735 ;
  assign n6820 = x1142 & ~n4183 ;
  assign n6821 = n7061 ^ x200 ;
  assign n6822 = x1144 ^ x1143 ;
  assign n6823 = n6821 & n6822 ;
  assign n6824 = n6823 ^ x1143 ;
  assign n6825 = n6824 & ~n7061 ;
  assign n6826 = x208 & n6825 ;
  assign n6827 = ~x200 & n6826 ;
  assign n6828 = n6827 ^ n6825 ;
  assign n6829 = n6828 ^ n6824 ;
  assign n6840 = n4366 & ~n6829 ;
  assign n6841 = n6820 & n6840 ;
  assign n6831 = ~x200 & n6830 ;
  assign n6832 = n6831 ^ n6829 ;
  assign n6835 = ~x1142 & ~n6832 ;
  assign n6836 = n6835 ^ n6831 ;
  assign n6837 = x199 & ~n6836 ;
  assign n6838 = n6837 ^ n6829 ;
  assign n6842 = n6841 ^ n6838 ;
  assign n6843 = n6734 & ~n6842 ;
  assign n6768 = x213 & ~n1911 ;
  assign n6769 = n6768 ^ n1911 ;
  assign n6777 = ~x219 & x1156 ;
  assign n6770 = x1157 ^ x1155 ;
  assign n6771 = ~x219 & n6770 ;
  assign n6772 = n6771 ^ x1155 ;
  assign n6778 = n6777 ^ n6772 ;
  assign n6779 = x211 & n6778 ;
  assign n6780 = n6779 ^ n6772 ;
  assign n6781 = ~n4011 & n6780 ;
  assign n6782 = ~n6769 & n6781 ;
  assign n6783 = n6782 ^ n6769 ;
  assign n6793 = x1155 ^ x1154 ;
  assign n6796 = ~x214 & n6793 ;
  assign n6797 = n6796 ^ x1154 ;
  assign n6798 = ~x219 & n6797 ;
  assign n6787 = x1156 ^ x1154 ;
  assign n6788 = ~x219 & n6787 ;
  assign n6789 = n6788 ^ x1154 ;
  assign n6784 = x1155 ^ x1153 ;
  assign n6785 = ~x219 & n6784 ;
  assign n6786 = n6785 ^ x1153 ;
  assign n6790 = n6789 ^ n6786 ;
  assign n6791 = x214 & n6790 ;
  assign n6792 = n6791 ^ n6789 ;
  assign n6799 = n6798 ^ n6792 ;
  assign n6800 = x211 & n6799 ;
  assign n6801 = n6800 ^ n6792 ;
  assign n6802 = x212 & n6801 ;
  assign n6803 = ~n6783 & n6802 ;
  assign n6804 = n6803 ^ n6783 ;
  assign n6805 = x214 ^ x212 ;
  assign n6806 = ~x219 & n6805 ;
  assign n6807 = x211 & n6806 ;
  assign n6814 = n6807 ^ n6806 ;
  assign n6815 = x1144 & n6814 ;
  assign n6811 = ~n4010 & n4023 ;
  assign n6810 = ~n4012 & n4022 ;
  assign n6812 = n6811 ^ n6810 ;
  assign n6813 = x1142 & n6812 ;
  assign n6816 = n6815 ^ n6813 ;
  assign n6808 = n6807 ^ n4187 ;
  assign n6809 = x1143 & n6808 ;
  assign n6817 = n6816 ^ n6809 ;
  assign n6818 = n6804 & ~n6817 ;
  assign n6819 = n6768 & n6818 ;
  assign n6844 = n6843 ^ n6819 ;
  assign n6845 = n6844 ^ n6804 ;
  assign n6846 = ~n6767 & n6845 ;
  assign n6847 = n6846 ^ x233 ;
  assign n6848 = x230 & ~n6847 ;
  assign n6849 = n6848 ^ x233 ;
  assign n6869 = x1156 & n6768 ;
  assign n6870 = n6814 & n6869 ;
  assign n6871 = n6870 ^ x1155 ;
  assign n6872 = n6870 ^ n6768 ;
  assign n6882 = n6808 & n6872 ;
  assign n6883 = n6871 & n6882 ;
  assign n6884 = n6883 ^ n6872 ;
  assign n6875 = x208 & n6759 ;
  assign n6876 = n6875 ^ n6749 ;
  assign n6877 = n6876 & ~n7061 ;
  assign n6878 = n6877 ^ n6749 ;
  assign n6879 = n6734 & n6878 ;
  assign n6880 = n6879 ^ n6734 ;
  assign n6885 = n6884 ^ n6880 ;
  assign n6896 = n6885 ^ x234 ;
  assign n6867 = n6768 ^ n6734 ;
  assign n6897 = n6896 ^ n6867 ;
  assign n6850 = n6830 ^ n4010 ;
  assign n6851 = n1911 & ~n6850 ;
  assign n6852 = n6851 ^ n4010 ;
  assign n6862 = ~n4190 & ~n6852 ;
  assign n6863 = n4039 & n6862 ;
  assign n6864 = x1152 & n6863 ;
  assign n6853 = ~n4039 & ~n6852 ;
  assign n6854 = x1154 ^ x1153 ;
  assign n6859 = n4190 & n6854 ;
  assign n6860 = n6859 ^ x1153 ;
  assign n6861 = n6853 & n6860 ;
  assign n6866 = n6864 ^ n6861 ;
  assign n6898 = n6897 ^ n6866 ;
  assign n6891 = x1154 & n6863 ;
  assign n6868 = n6867 ^ n6866 ;
  assign n6892 = n6891 ^ n6868 ;
  assign n6893 = n6885 & ~n6892 ;
  assign n6899 = n6898 ^ n6893 ;
  assign n6886 = n6885 ^ n6867 ;
  assign n6895 = ~n6868 & n6886 ;
  assign n6900 = n6899 ^ n6895 ;
  assign n6901 = x230 & n6900 ;
  assign n6902 = n6901 ^ x234 ;
  assign n6910 = ~x211 & n6805 ;
  assign n6903 = ~n1911 & n6810 ;
  assign n6906 = ~x213 & n6784 ;
  assign n6907 = n6906 ^ x1155 ;
  assign n6908 = n6903 & n6907 ;
  assign n6909 = n6908 ^ n1911 ;
  assign n6911 = n6786 ^ n6772 ;
  assign n6914 = ~x213 & n6911 ;
  assign n6915 = n6914 ^ n6772 ;
  assign n6916 = ~n6909 & n6915 ;
  assign n6917 = n6910 & n6916 ;
  assign n6918 = n6917 ^ n6909 ;
  assign n6919 = n6808 & ~n6918 ;
  assign n6922 = ~x213 & n6787 ;
  assign n6923 = n6922 ^ x1156 ;
  assign n6924 = n6919 & n6923 ;
  assign n6925 = n6924 ^ n6918 ;
  assign n6926 = n1911 & n4015 ;
  assign n6929 = ~x200 & n6854 ;
  assign n6930 = n6929 ^ x1153 ;
  assign n6931 = ~x199 & n6930 ;
  assign n6932 = n6931 ^ n6749 ;
  assign n6935 = ~x209 & n6932 ;
  assign n6936 = n6935 ^ n6749 ;
  assign n6937 = n6926 & n6936 ;
  assign n6938 = n6937 ^ n1911 ;
  assign n6939 = n6938 & n7061 ;
  assign n6940 = n6761 ^ n6746 ;
  assign n6943 = x209 & n6940 ;
  assign n6944 = n6943 ^ n6761 ;
  assign n6945 = n6939 & n6944 ;
  assign n6946 = n6945 ^ n6938 ;
  assign n6947 = n6925 & ~n6946 ;
  assign n6948 = n6947 ^ x235 ;
  assign n6949 = x230 & n6948 ;
  assign n6950 = n6949 ^ x235 ;
  assign n6969 = x208 & n6750 ;
  assign n6958 = ~x200 & x1158 ;
  assign n6951 = x1157 ^ x1156 ;
  assign n6952 = x200 & n6951 ;
  assign n6953 = n6952 ^ x1156 ;
  assign n6959 = n6958 ^ n6953 ;
  assign n6960 = ~n4030 & n6959 ;
  assign n6961 = n6960 ^ n6953 ;
  assign n6962 = n6961 ^ n6746 ;
  assign n6963 = ~x208 & n6962 ;
  assign n6964 = n6963 ^ n6746 ;
  assign n6970 = n6969 ^ n6964 ;
  assign n6971 = n6970 & ~n7061 ;
  assign n6972 = n6971 ^ n6964 ;
  assign n6973 = x230 & n6735 ;
  assign n6974 = n6972 & n6973 ;
  assign n6975 = n6974 ^ n6768 ;
  assign n6979 = x1143 & n6812 ;
  assign n6977 = x1145 & n6814 ;
  assign n6976 = x1144 & n6808 ;
  assign n6978 = n6977 ^ n6976 ;
  assign n6980 = n6979 ^ n6978 ;
  assign n6981 = n6974 ^ x230 ;
  assign n6982 = n6980 & n6981 ;
  assign n6983 = n6975 & n6982 ;
  assign n6984 = n6983 ^ n6981 ;
  assign n7007 = ~x219 & n6951 ;
  assign n6998 = x1158 ^ x1156 ;
  assign n6999 = n6998 ^ n6951 ;
  assign n7000 = n6999 ^ x1156 ;
  assign n7003 = ~x219 & n7000 ;
  assign n7004 = n7003 ^ x1156 ;
  assign n7005 = ~n4021 & n7004 ;
  assign n6990 = n6789 ^ n6772 ;
  assign n6991 = x214 & n6990 ;
  assign n6992 = n6991 ^ n6772 ;
  assign n6987 = ~x214 & n6736 ;
  assign n6988 = n6987 ^ x1155 ;
  assign n6989 = ~x219 & n6988 ;
  assign n6993 = n6992 ^ n6989 ;
  assign n6994 = x211 & n6993 ;
  assign n6995 = n6994 ^ n6992 ;
  assign n6996 = n6995 ^ x1156 ;
  assign n7006 = n7005 ^ n6996 ;
  assign n7008 = n7007 ^ n7006 ;
  assign n7009 = n7008 ^ n6995 ;
  assign n7012 = x214 & n7009 ;
  assign n7013 = n7012 ^ n6995 ;
  assign n7014 = ~x212 & n7013 ;
  assign n7015 = n7014 ^ n6995 ;
  assign n7016 = ~n6769 & n7015 ;
  assign n7017 = n6984 & n7016 ;
  assign n7018 = n7017 ^ n6984 ;
  assign n7019 = n7018 ^ x230 ;
  assign n7039 = n7061 ^ n6831 ;
  assign n7040 = ~x199 & x1144 ;
  assign n7041 = n7039 & n7040 ;
  assign n7029 = ~x199 & n4015 ;
  assign n7030 = n7029 ^ n6831 ;
  assign n7031 = x1145 ^ x1143 ;
  assign n7033 = n4183 & n7031 ;
  assign n7034 = n7033 ^ x1145 ;
  assign n7035 = n7034 ^ n7031 ;
  assign n7036 = ~n7030 & n7035 ;
  assign n7037 = n7036 ^ n7033 ;
  assign n7038 = n7037 ^ x1143 ;
  assign n7042 = n7041 ^ n7038 ;
  assign n7045 = n6734 & n7042 ;
  assign n7020 = n7019 ^ x237 ;
  assign n7046 = n7045 ^ n7020 ;
  assign n7047 = n7018 & ~n7046 ;
  assign n7048 = n7047 ^ n7020 ;
  assign n7049 = n7048 ^ x230 ;
  assign n7051 = n7019 & ~n7049 ;
  assign n7052 = n7051 ^ n7048 ;
  assign n7078 = x1151 & n6863 ;
  assign n7074 = x1153 ^ x1152 ;
  assign n7075 = ~n4190 & n7074 ;
  assign n7076 = n7075 ^ x1153 ;
  assign n7077 = n6853 & n7076 ;
  assign n7080 = n7078 ^ n7077 ;
  assign n7081 = ~n6867 & ~n7080 ;
  assign n7058 = n6734 & n6761 ;
  assign n7063 = n4015 & ~n6758 ;
  assign n7064 = n7063 ^ n6830 ;
  assign n7065 = n7058 & n7064 ;
  assign n7066 = n7065 ^ n6734 ;
  assign n7067 = n4015 & n6931 ;
  assign n7068 = n7066 & n7067 ;
  assign n7069 = n7068 ^ n7066 ;
  assign n7072 = n7069 ^ x238 ;
  assign n7055 = x1154 & n6808 ;
  assign n7054 = x1155 & n6814 ;
  assign n7056 = n7055 ^ n7054 ;
  assign n7053 = x1153 & n6812 ;
  assign n7057 = n7056 ^ n7053 ;
  assign n7071 = n6768 & ~n7057 ;
  assign n7073 = n7072 ^ n7071 ;
  assign n7082 = n7081 ^ n7073 ;
  assign n7083 = x230 & ~n7082 ;
  assign n7084 = n7083 ^ x238 ;
  assign n7085 = n1911 & n4014 ;
  assign n7086 = n6961 ^ n6750 ;
  assign n7087 = x209 & n7086 ;
  assign n7088 = n7087 ^ n6750 ;
  assign n7089 = n7085 & n7088 ;
  assign n7090 = ~n1911 & ~n4011 ;
  assign n7091 = x213 & n7008 ;
  assign n7092 = n7091 ^ n6995 ;
  assign n7093 = n7090 & n7092 ;
  assign n7094 = ~n7089 & ~n7093 ;
  assign n7095 = n7094 ^ x239 ;
  assign n7096 = x230 & ~n7095 ;
  assign n7097 = n7096 ^ x239 ;
  assign n7116 = x1147 & n6863 ;
  assign n7110 = x1149 ^ x1148 ;
  assign n7113 = ~n4190 & n7110 ;
  assign n7114 = n7113 ^ x1149 ;
  assign n7115 = n6853 & n7114 ;
  assign n7118 = n7116 ^ n7115 ;
  assign n7119 = n7118 ^ x240 ;
  assign n7104 = x1145 & n6863 ;
  assign n7098 = x1147 ^ x1146 ;
  assign n7101 = ~n4190 & n7098 ;
  assign n7102 = n7101 ^ x1147 ;
  assign n7103 = n6853 & n7102 ;
  assign n7106 = n7104 ^ n7103 ;
  assign n7107 = n7106 ^ x240 ;
  assign n7120 = n7119 ^ n7107 ;
  assign n7121 = n6867 & n7120 ;
  assign n7122 = n7121 ^ n7107 ;
  assign n7123 = x230 & n7122 ;
  assign n7124 = n7123 ^ x240 ;
  assign n7134 = x1149 & n6863 ;
  assign n7128 = x1151 ^ x1150 ;
  assign n7131 = ~n4190 & n7128 ;
  assign n7132 = n7131 ^ x1151 ;
  assign n7133 = n6853 & n7132 ;
  assign n7136 = n7134 ^ n7133 ;
  assign n7137 = n7136 ^ x241 ;
  assign n7125 = n7080 ^ x241 ;
  assign n7138 = n7137 ^ n7125 ;
  assign n7139 = ~n6867 & n7138 ;
  assign n7140 = n7139 ^ n7125 ;
  assign n7141 = x230 & n7140 ;
  assign n7142 = n7141 ^ x241 ;
  assign n7154 = n6735 & ~n6842 ;
  assign n7150 = x1144 & n6863 ;
  assign n7144 = x1146 ^ x1145 ;
  assign n7147 = ~n4190 & n7144 ;
  assign n7148 = n7147 ^ x1146 ;
  assign n7149 = n6853 & n7148 ;
  assign n7152 = n7150 ^ n7149 ;
  assign n7153 = n6867 & ~n7152 ;
  assign n7155 = n7154 ^ n7153 ;
  assign n7156 = n7155 ^ x242 ;
  assign n7143 = ~n6769 & ~n6817 ;
  assign n7157 = n7156 ^ n7143 ;
  assign n7158 = x230 & ~n7157 ;
  assign n7159 = n7158 ^ x242 ;
  assign n7160 = ~x230 & ~x1091 ;
  assign n7185 = n4038 ^ n4034 ;
  assign n7186 = x1155 & n7185 ;
  assign n7181 = n4023 ^ n4013 ;
  assign n7182 = n1911 & n7181 ;
  assign n7183 = n7182 ^ n4023 ;
  assign n7184 = x1157 & n7183 ;
  assign n7187 = n7186 ^ n7184 ;
  assign n7162 = ~x83 & ~x85 ;
  assign n7163 = x314 & n7162 ;
  assign n7165 = x81 & ~n4038 ;
  assign n7166 = n7163 & n7165 ;
  assign n7164 = n7163 ^ x314 ;
  assign n7167 = n7166 ^ n7164 ;
  assign n7168 = x802 & n7167 ;
  assign n7169 = x276 & n7168 ;
  assign n7170 = x271 & n7169 ;
  assign n7171 = x273 & n7170 ;
  assign n7172 = x283 & n7171 ;
  assign n7173 = x272 & n7172 ;
  assign n7174 = x275 & n7173 ;
  assign n7175 = x268 & n7174 ;
  assign n7176 = x253 & n7175 ;
  assign n7177 = x254 & n7176 ;
  assign n7178 = x267 & n7177 ;
  assign n7179 = ~x263 & n7178 ;
  assign n7180 = n7179 ^ x243 ;
  assign n7188 = n7187 ^ n7180 ;
  assign n7161 = x1156 & ~n4034 ;
  assign n7189 = n7188 ^ n7161 ;
  assign n7190 = ~n7160 & ~n7189 ;
  assign n7191 = n7190 ^ n7180 ;
  assign n7194 = ~n6769 & ~n6980 ;
  assign n7193 = n6867 & ~n7106 ;
  assign n7195 = n7194 ^ n7193 ;
  assign n7196 = n7195 ^ x244 ;
  assign n7192 = n6735 & ~n7042 ;
  assign n7197 = n7196 ^ n7192 ;
  assign n7198 = x230 & ~n7197 ;
  assign n7199 = n7198 ^ x244 ;
  assign n7209 = x1146 & n6863 ;
  assign n7203 = x1148 ^ x1147 ;
  assign n7206 = ~n4190 & n7203 ;
  assign n7207 = n7206 ^ x1148 ;
  assign n7208 = n6853 & n7207 ;
  assign n7211 = n7209 ^ n7208 ;
  assign n7212 = n7211 ^ x245 ;
  assign n7200 = n7152 ^ x245 ;
  assign n7213 = n7212 ^ n7200 ;
  assign n7214 = n6867 & n7213 ;
  assign n7215 = n7214 ^ n7200 ;
  assign n7216 = x230 & n7215 ;
  assign n7217 = n7216 ^ x245 ;
  assign n7227 = x1148 & n6863 ;
  assign n7221 = x1150 ^ x1149 ;
  assign n7224 = ~n4190 & n7221 ;
  assign n7225 = n7224 ^ x1150 ;
  assign n7226 = n6853 & n7225 ;
  assign n7229 = n7227 ^ n7226 ;
  assign n7230 = n7229 ^ x246 ;
  assign n7218 = n7211 ^ x246 ;
  assign n7231 = n7230 ^ n7218 ;
  assign n7232 = n6867 & n7231 ;
  assign n7233 = n7232 ^ n7218 ;
  assign n7234 = x230 & n7233 ;
  assign n7235 = n7234 ^ x246 ;
  assign n7239 = n7136 ^ x247 ;
  assign n7236 = n7118 ^ x247 ;
  assign n7240 = n7239 ^ n7236 ;
  assign n7241 = n6867 & n7240 ;
  assign n7242 = n7241 ^ n7236 ;
  assign n7243 = x230 & n7242 ;
  assign n7244 = n7243 ^ x247 ;
  assign n7254 = x1150 & n6863 ;
  assign n7248 = x1152 ^ x1151 ;
  assign n7251 = ~n4190 & n7248 ;
  assign n7252 = n7251 ^ x1152 ;
  assign n7253 = n6853 & n7252 ;
  assign n7256 = n7254 ^ n7253 ;
  assign n7257 = n7256 ^ x248 ;
  assign n7245 = n7229 ^ x248 ;
  assign n7258 = n7257 ^ n7245 ;
  assign n7259 = n6867 & n7258 ;
  assign n7260 = n7259 ^ n7245 ;
  assign n7261 = x230 & n7260 ;
  assign n7262 = n7261 ^ x248 ;
  assign n7266 = n7256 ^ x249 ;
  assign n7263 = n6866 ^ x249 ;
  assign n7267 = n7266 ^ n7263 ;
  assign n7268 = ~n6867 & n7267 ;
  assign n7269 = n7268 ^ n7263 ;
  assign n7270 = x230 & n7269 ;
  assign n7271 = n7270 ^ x249 ;
  assign n7272 = ~x250 & ~n4164 ;
  assign n7273 = ~n5017 & n7272 ;
  assign n7274 = n7273 ^ x250 ;
  assign n7275 = x1053 ^ x1039 ;
  assign n7276 = ~x200 & n7275 ;
  assign n7277 = n7276 ^ x1039 ;
  assign n7278 = n7277 ^ x251 ;
  assign n7279 = x897 ^ x476 ;
  assign n7280 = ~x200 & ~n7279 ;
  assign n7281 = n7280 ^ x476 ;
  assign n7282 = ~x199 & ~n7281 ;
  assign n7283 = n7278 & n7282 ;
  assign n7284 = n7283 ^ x251 ;
  assign n7285 = n2668 & ~n2678 ;
  assign n7286 = n2943 & n7285 ;
  assign n7287 = x1093 & ~n2991 ;
  assign n7288 = x252 & x1092 ;
  assign n7289 = ~n7287 & n7288 ;
  assign n7290 = ~n7286 & ~n7289 ;
  assign n7294 = x1151 & n7185 ;
  assign n7293 = x1153 & n7183 ;
  assign n7295 = n7294 ^ n7293 ;
  assign n7292 = n7175 ^ x253 ;
  assign n7296 = n7295 ^ n7292 ;
  assign n7291 = x1152 & ~n4034 ;
  assign n7297 = n7296 ^ n7291 ;
  assign n7298 = ~n7160 & n7297 ;
  assign n7299 = n7298 ^ n7292 ;
  assign n7303 = x1154 & n7183 ;
  assign n7302 = x1152 & n7185 ;
  assign n7304 = n7303 ^ n7302 ;
  assign n7301 = n7176 ^ x254 ;
  assign n7305 = n7304 ^ n7301 ;
  assign n7300 = x1153 & ~n4034 ;
  assign n7306 = n7305 ^ n7300 ;
  assign n7307 = ~n7160 & n7306 ;
  assign n7308 = n7307 ^ n7301 ;
  assign n7309 = x1049 ^ x1036 ;
  assign n7310 = ~x200 & n7309 ;
  assign n7311 = n7310 ^ x1036 ;
  assign n7312 = n7311 ^ x255 ;
  assign n7313 = n7282 & n7312 ;
  assign n7314 = n7313 ^ x255 ;
  assign n7315 = x1070 ^ x1048 ;
  assign n7316 = x200 & n7315 ;
  assign n7317 = n7316 ^ x1048 ;
  assign n7318 = n7317 ^ x256 ;
  assign n7319 = n7282 & n7318 ;
  assign n7320 = n7319 ^ x256 ;
  assign n7321 = x1084 ^ x1065 ;
  assign n7322 = ~x200 & n7321 ;
  assign n7323 = n7322 ^ x1065 ;
  assign n7324 = n7323 ^ x257 ;
  assign n7325 = n7282 & n7324 ;
  assign n7326 = n7325 ^ x257 ;
  assign n7327 = x1072 ^ x1062 ;
  assign n7328 = ~x200 & n7327 ;
  assign n7329 = n7328 ^ x1062 ;
  assign n7330 = n7329 ^ x258 ;
  assign n7331 = n7282 & n7330 ;
  assign n7332 = n7331 ^ x258 ;
  assign n7333 = x1069 ^ x1059 ;
  assign n7334 = x200 & n7333 ;
  assign n7335 = n7334 ^ x1059 ;
  assign n7336 = n7335 ^ x259 ;
  assign n7337 = n7282 & n7336 ;
  assign n7338 = n7337 ^ x259 ;
  assign n7339 = x1067 ^ x1044 ;
  assign n7340 = x200 & n7339 ;
  assign n7341 = n7340 ^ x1044 ;
  assign n7342 = n7341 ^ x260 ;
  assign n7343 = n7282 & n7342 ;
  assign n7344 = n7343 ^ x260 ;
  assign n7345 = x1040 ^ x1037 ;
  assign n7346 = x200 & n7345 ;
  assign n7347 = n7346 ^ x1037 ;
  assign n7348 = n7347 ^ x261 ;
  assign n7349 = n7282 & n7348 ;
  assign n7350 = n7349 ^ x261 ;
  assign n7351 = x1093 ^ x123 ;
  assign n7352 = ~x228 & ~n7351 ;
  assign n7353 = n7352 ^ x123 ;
  assign n7358 = x1142 & n6853 ;
  assign n7359 = n7358 ^ x262 ;
  assign n7360 = ~n7353 & ~n7359 ;
  assign n7361 = n7360 ^ x262 ;
  assign n7365 = x1154 & n7185 ;
  assign n7364 = x1156 & n7183 ;
  assign n7366 = n7365 ^ n7364 ;
  assign n7363 = n7178 ^ x263 ;
  assign n7367 = n7366 ^ n7363 ;
  assign n7362 = x1155 & ~n4034 ;
  assign n7368 = n7367 ^ n7362 ;
  assign n7369 = ~n7160 & ~n7368 ;
  assign n7370 = n7369 ^ n7363 ;
  assign n7376 = x1143 & n7183 ;
  assign n7375 = x1141 & n7185 ;
  assign n7377 = n7376 ^ n7375 ;
  assign n7372 = x796 ^ x264 ;
  assign n7373 = n7167 & ~n7372 ;
  assign n7374 = n7373 ^ x264 ;
  assign n7378 = n7377 ^ n7374 ;
  assign n7371 = x1142 & ~n4034 ;
  assign n7379 = n7378 ^ n7371 ;
  assign n7380 = ~n7160 & ~n7379 ;
  assign n7381 = n7380 ^ n7374 ;
  assign n7387 = x1144 & n7183 ;
  assign n7386 = x1142 & n7185 ;
  assign n7388 = n7387 ^ n7386 ;
  assign n7383 = x819 ^ x265 ;
  assign n7384 = n7167 & ~n7383 ;
  assign n7385 = n7384 ^ x265 ;
  assign n7389 = n7388 ^ n7385 ;
  assign n7382 = x1143 & ~n4034 ;
  assign n7390 = n7389 ^ n7382 ;
  assign n7391 = ~n7160 & ~n7390 ;
  assign n7392 = n7391 ^ n7385 ;
  assign n7398 = x1136 & n7183 ;
  assign n7397 = x1134 & n7185 ;
  assign n7399 = n7398 ^ n7397 ;
  assign n7394 = x948 ^ x266 ;
  assign n7395 = n7167 & n7394 ;
  assign n7396 = n7395 ^ x266 ;
  assign n7400 = n7399 ^ n7396 ;
  assign n7393 = x1135 & ~n4034 ;
  assign n7401 = n7400 ^ n7393 ;
  assign n7402 = ~n7160 & n7401 ;
  assign n7403 = n7402 ^ n7396 ;
  assign n7407 = x1155 & n7183 ;
  assign n7406 = x1153 & n7185 ;
  assign n7408 = n7407 ^ n7406 ;
  assign n7405 = n7177 ^ x267 ;
  assign n7409 = n7408 ^ n7405 ;
  assign n7404 = x1154 & ~n4034 ;
  assign n7410 = n7409 ^ n7404 ;
  assign n7411 = ~n7160 & n7410 ;
  assign n7412 = n7411 ^ n7405 ;
  assign n7416 = x1150 & n7185 ;
  assign n7415 = x1152 & n7183 ;
  assign n7417 = n7416 ^ n7415 ;
  assign n7414 = n7174 ^ x268 ;
  assign n7418 = n7417 ^ n7414 ;
  assign n7413 = x1151 & ~n4034 ;
  assign n7419 = n7418 ^ n7413 ;
  assign n7420 = ~n7160 & n7419 ;
  assign n7421 = n7420 ^ n7414 ;
  assign n7427 = x1138 & n7183 ;
  assign n7426 = x1136 & n7185 ;
  assign n7428 = n7427 ^ n7426 ;
  assign n7423 = x817 ^ x269 ;
  assign n7424 = n7167 & ~n7423 ;
  assign n7425 = n7424 ^ x269 ;
  assign n7429 = n7428 ^ n7425 ;
  assign n7422 = x1137 & ~n4034 ;
  assign n7430 = n7429 ^ n7422 ;
  assign n7431 = ~n7160 & ~n7430 ;
  assign n7432 = n7431 ^ n7425 ;
  assign n7438 = x1141 & n7183 ;
  assign n7437 = x1139 & n7185 ;
  assign n7439 = n7438 ^ n7437 ;
  assign n7434 = x805 ^ x270 ;
  assign n7435 = n7167 & ~n7434 ;
  assign n7436 = n7435 ^ x270 ;
  assign n7440 = n7439 ^ n7436 ;
  assign n7433 = x1140 & ~n4034 ;
  assign n7441 = n7440 ^ n7433 ;
  assign n7442 = ~n7160 & ~n7441 ;
  assign n7443 = n7442 ^ n7436 ;
  assign n7447 = x1147 & n7183 ;
  assign n7446 = x1145 & n7185 ;
  assign n7448 = n7447 ^ n7446 ;
  assign n7445 = n7169 ^ x271 ;
  assign n7449 = n7448 ^ n7445 ;
  assign n7444 = x1146 & ~n4034 ;
  assign n7450 = n7449 ^ n7444 ;
  assign n7451 = ~n7160 & n7450 ;
  assign n7452 = n7451 ^ n7445 ;
  assign n7456 = x1148 & n7185 ;
  assign n7455 = x1150 & n7183 ;
  assign n7457 = n7456 ^ n7455 ;
  assign n7454 = n7172 ^ x272 ;
  assign n7458 = n7457 ^ n7454 ;
  assign n7453 = x1149 & ~n4034 ;
  assign n7459 = n7458 ^ n7453 ;
  assign n7460 = ~n7160 & n7459 ;
  assign n7461 = n7460 ^ n7454 ;
  assign n7465 = x1148 & n7183 ;
  assign n7464 = x1146 & n7185 ;
  assign n7466 = n7465 ^ n7464 ;
  assign n7463 = n7170 ^ x273 ;
  assign n7467 = n7466 ^ n7463 ;
  assign n7462 = x1147 & ~n4034 ;
  assign n7468 = n7467 ^ n7462 ;
  assign n7469 = ~n7160 & n7468 ;
  assign n7470 = n7469 ^ n7463 ;
  assign n7476 = x1143 & n7185 ;
  assign n7475 = x1145 & n7183 ;
  assign n7477 = n7476 ^ n7475 ;
  assign n7472 = x659 ^ x274 ;
  assign n7473 = n7167 & ~n7472 ;
  assign n7474 = n7473 ^ x274 ;
  assign n7478 = n7477 ^ n7474 ;
  assign n7471 = x1144 & ~n4034 ;
  assign n7479 = n7478 ^ n7471 ;
  assign n7480 = ~n7160 & ~n7479 ;
  assign n7481 = n7480 ^ n7474 ;
  assign n7485 = x1149 & n7185 ;
  assign n7484 = x1151 & n7183 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7483 = n7173 ^ x275 ;
  assign n7487 = n7486 ^ n7483 ;
  assign n7482 = x1150 & ~n4034 ;
  assign n7488 = n7487 ^ n7482 ;
  assign n7489 = ~n7160 & n7488 ;
  assign n7490 = n7489 ^ n7483 ;
  assign n7494 = x1144 & n7185 ;
  assign n7493 = x1146 & n7183 ;
  assign n7495 = n7494 ^ n7493 ;
  assign n7492 = n7168 ^ x276 ;
  assign n7496 = n7495 ^ n7492 ;
  assign n7491 = x1145 & ~n4034 ;
  assign n7497 = n7496 ^ n7491 ;
  assign n7498 = ~n7160 & n7497 ;
  assign n7499 = n7498 ^ n7492 ;
  assign n7505 = x1142 & n7183 ;
  assign n7504 = x1140 & n7185 ;
  assign n7506 = n7505 ^ n7504 ;
  assign n7501 = x820 ^ x277 ;
  assign n7502 = n7167 & ~n7501 ;
  assign n7503 = n7502 ^ x277 ;
  assign n7507 = n7506 ^ n7503 ;
  assign n7500 = x1141 & ~n4034 ;
  assign n7508 = n7507 ^ n7500 ;
  assign n7509 = ~n7160 & ~n7508 ;
  assign n7510 = n7509 ^ n7503 ;
  assign n7518 = x1133 & ~n4034 ;
  assign n7516 = x1134 & n7183 ;
  assign n7514 = x1132 & n7185 ;
  assign n7511 = x976 ^ x278 ;
  assign n7512 = n7167 & n7511 ;
  assign n7513 = n7512 ^ x278 ;
  assign n7515 = n7514 ^ n7513 ;
  assign n7517 = n7516 ^ n7515 ;
  assign n7519 = n7518 ^ n7517 ;
  assign n7520 = ~n7160 & n7519 ;
  assign n7521 = n7520 ^ n7513 ;
  assign n7527 = x1135 & n7183 ;
  assign n7526 = x1133 & n7185 ;
  assign n7528 = n7527 ^ n7526 ;
  assign n7523 = x958 ^ x279 ;
  assign n7524 = n7167 & n7523 ;
  assign n7525 = n7524 ^ x279 ;
  assign n7529 = n7528 ^ n7525 ;
  assign n7522 = x1134 & ~n4034 ;
  assign n7530 = n7529 ^ n7522 ;
  assign n7531 = ~n7160 & n7530 ;
  assign n7532 = n7531 ^ n7525 ;
  assign n7538 = x1137 & n7183 ;
  assign n7537 = x1135 & n7185 ;
  assign n7539 = n7538 ^ n7537 ;
  assign n7534 = x914 ^ x280 ;
  assign n7535 = n7167 & ~n7534 ;
  assign n7536 = n7535 ^ x280 ;
  assign n7540 = n7539 ^ n7536 ;
  assign n7533 = x1136 & ~n4034 ;
  assign n7541 = n7540 ^ n7533 ;
  assign n7542 = ~n7160 & ~n7541 ;
  assign n7543 = n7542 ^ n7536 ;
  assign n7549 = x1139 & n7183 ;
  assign n7548 = x1137 & n7185 ;
  assign n7550 = n7549 ^ n7548 ;
  assign n7545 = x830 ^ x281 ;
  assign n7546 = n7167 & ~n7545 ;
  assign n7547 = n7546 ^ x281 ;
  assign n7551 = n7550 ^ n7547 ;
  assign n7544 = x1138 & ~n4034 ;
  assign n7552 = n7551 ^ n7544 ;
  assign n7553 = ~n7160 & ~n7552 ;
  assign n7554 = n7553 ^ n7547 ;
  assign n7560 = x1140 & n7183 ;
  assign n7559 = x1138 & n7185 ;
  assign n7561 = n7560 ^ n7559 ;
  assign n7556 = x836 ^ x282 ;
  assign n7557 = n7167 & ~n7556 ;
  assign n7558 = n7557 ^ x282 ;
  assign n7562 = n7561 ^ n7558 ;
  assign n7555 = x1139 & ~n4034 ;
  assign n7563 = n7562 ^ n7555 ;
  assign n7564 = ~n7160 & ~n7563 ;
  assign n7565 = n7564 ^ n7558 ;
  assign n7569 = x1147 & n7185 ;
  assign n7568 = x1149 & n7183 ;
  assign n7570 = n7569 ^ n7568 ;
  assign n7567 = n7171 ^ x283 ;
  assign n7571 = n7570 ^ n7567 ;
  assign n7566 = x1148 & ~n4034 ;
  assign n7572 = n7571 ^ n7566 ;
  assign n7573 = ~n7160 & n7572 ;
  assign n7574 = n7573 ^ n7567 ;
  assign n7581 = x1143 & n6853 ;
  assign n7582 = n4190 & n7581 ;
  assign n7583 = n7582 ^ n4190 ;
  assign n7575 = n4190 ^ x284 ;
  assign n7584 = n7583 ^ n7575 ;
  assign n7585 = ~n7353 & ~n7584 ;
  assign n7586 = n7585 ^ x284 ;
  assign n7587 = n3978 & n4161 ;
  assign n7588 = ~n3323 & n7587 ;
  assign n7589 = x289 & n7588 ;
  assign n7590 = x286 & x288 ;
  assign n7591 = n7589 & n7590 ;
  assign n7592 = n7591 ^ x285 ;
  assign n7593 = ~x288 & n3323 ;
  assign n7594 = ~n7587 & n7593 ;
  assign n7595 = x285 & n3186 ;
  assign n7596 = n7594 & n7595 ;
  assign n7597 = ~x793 & ~n7596 ;
  assign n7598 = n7592 & n7597 ;
  assign n7599 = x288 & n7588 ;
  assign n7600 = n7599 ^ x286 ;
  assign n7601 = n7600 ^ n7594 ;
  assign n7602 = ~x793 & n7601 ;
  assign n7604 = n3187 & n7602 ;
  assign n7605 = n7604 ^ n7602 ;
  assign n7606 = ~x287 & ~x332 ;
  assign n7607 = x457 & n7606 ;
  assign n7608 = n7607 ^ x332 ;
  assign n7609 = n3425 ^ x288 ;
  assign n7610 = n7609 ^ n7587 ;
  assign n7611 = ~x793 & n7610 ;
  assign n7615 = ~x286 & n7594 ;
  assign n7616 = x289 & n7615 ;
  assign n7613 = n7596 ^ x289 ;
  assign n7617 = n7616 ^ n7613 ;
  assign n7612 = n7590 & n7599 ;
  assign n7618 = n7617 ^ n7612 ;
  assign n7619 = ~x793 & n7618 ;
  assign n7620 = x1048 ^ x290 ;
  assign n7621 = ~x476 & n7620 ;
  assign n7622 = n7621 ^ x290 ;
  assign n7623 = x1049 ^ x291 ;
  assign n7624 = ~x476 & n7623 ;
  assign n7625 = n7624 ^ x291 ;
  assign n7626 = x1084 ^ x292 ;
  assign n7627 = ~x476 & n7626 ;
  assign n7628 = n7627 ^ x292 ;
  assign n7629 = x1059 ^ x293 ;
  assign n7630 = ~x476 & n7629 ;
  assign n7631 = n7630 ^ x293 ;
  assign n7632 = x1072 ^ x294 ;
  assign n7633 = ~x476 & n7632 ;
  assign n7634 = n7633 ^ x294 ;
  assign n7635 = x1053 ^ x295 ;
  assign n7636 = ~x476 & n7635 ;
  assign n7637 = n7636 ^ x295 ;
  assign n7638 = x1037 ^ x296 ;
  assign n7639 = ~x476 & n7638 ;
  assign n7640 = n7639 ^ x296 ;
  assign n7641 = x1044 ^ x297 ;
  assign n7642 = ~x476 & n7641 ;
  assign n7643 = n7642 ^ x297 ;
  assign n7644 = x1044 ^ x298 ;
  assign n7645 = ~x478 & n7644 ;
  assign n7646 = n7645 ^ x298 ;
  assign n7647 = n1209 & n1767 ;
  assign n7648 = x39 & n3917 ;
  assign n7649 = ~x287 & n7648 ;
  assign n7650 = n7649 ^ n4257 ;
  assign n7652 = ~n4264 & ~n7650 ;
  assign n7653 = ~n7647 & n7652 ;
  assign n7654 = ~x24 & n1746 ;
  assign n7659 = ~x312 & n7654 ;
  assign n7660 = n7659 ^ x300 ;
  assign n7661 = ~x55 & ~n7660 ;
  assign n7662 = ~x300 & ~x312 ;
  assign n7667 = n7654 & n7662 ;
  assign n7668 = n7667 ^ x301 ;
  assign n7669 = ~x55 & ~n7668 ;
  assign n7675 = n7674 ^ n1968 ;
  assign n7676 = ~x237 & n7675 ;
  assign n7670 = n1931 ^ n1663 ;
  assign n7671 = n1911 & n7670 ;
  assign n7672 = n7671 ^ n1663 ;
  assign n7673 = x937 & n7672 ;
  assign n7677 = n7676 ^ n7673 ;
  assign n7682 = x1148 & n2591 ;
  assign n7678 = n1936 ^ n1526 ;
  assign n7679 = n1911 & n7678 ;
  assign n7680 = n7679 ^ n1526 ;
  assign n7681 = x273 & n7680 ;
  assign n7683 = n7682 ^ n7681 ;
  assign n7684 = ~n7677 & ~n7683 ;
  assign n7685 = x1049 ^ x303 ;
  assign n7686 = ~x478 & n7685 ;
  assign n7687 = n7686 ^ x303 ;
  assign n7688 = x1048 ^ x304 ;
  assign n7689 = ~x478 & n7688 ;
  assign n7690 = n7689 ^ x304 ;
  assign n7691 = x1084 ^ x305 ;
  assign n7692 = ~x478 & n7691 ;
  assign n7693 = n7692 ^ x305 ;
  assign n7694 = x1059 ^ x306 ;
  assign n7695 = ~x478 & n7694 ;
  assign n7696 = n7695 ^ x306 ;
  assign n7697 = x1053 ^ x307 ;
  assign n7698 = ~x478 & n7697 ;
  assign n7699 = n7698 ^ x307 ;
  assign n7700 = x1037 ^ x308 ;
  assign n7701 = ~x478 & n7700 ;
  assign n7702 = n7701 ^ x308 ;
  assign n7703 = x1072 ^ x309 ;
  assign n7704 = ~x478 & n7703 ;
  assign n7705 = n7704 ^ x309 ;
  assign n7707 = ~x233 & n7675 ;
  assign n7706 = x271 & n7680 ;
  assign n7708 = n7707 ^ n7706 ;
  assign n7710 = x934 & n7672 ;
  assign n7709 = x1147 & n2591 ;
  assign n7711 = n7710 ^ n7709 ;
  assign n7712 = ~n7708 & ~n7711 ;
  assign n7713 = x301 & n7662 ;
  assign n7718 = n7654 & n7713 ;
  assign n7719 = n7718 ^ x311 ;
  assign n7720 = ~x55 & ~n7719 ;
  assign n7721 = n7654 ^ x312 ;
  assign n7722 = ~x55 & n7721 ;
  assign n7723 = n4851 ^ n2640 ;
  assign n7724 = n4838 ^ x314 ;
  assign n7727 = ~n4851 & n7724 ;
  assign n7728 = n7727 ^ x314 ;
  assign n7729 = n7723 & ~n7728 ;
  assign n7730 = n7729 ^ n2640 ;
  assign n7731 = n7730 ^ x313 ;
  assign n7732 = ~x954 & ~n7731 ;
  assign n7733 = n7732 ^ x313 ;
  assign n7734 = n5163 & n5429 ;
  assign n7735 = ~x340 & n7587 ;
  assign n7736 = x1080 ^ x315 ;
  assign n7737 = n7735 & n7736 ;
  assign n7738 = n7737 ^ x315 ;
  assign n7739 = x1047 ^ x316 ;
  assign n7740 = n7735 & n7739 ;
  assign n7741 = n7740 ^ x316 ;
  assign n7742 = ~x330 & n7587 ;
  assign n7743 = x1078 ^ x317 ;
  assign n7744 = n7742 & n7743 ;
  assign n7745 = n7744 ^ x317 ;
  assign n7746 = ~x341 & n7587 ;
  assign n7747 = x1074 ^ x318 ;
  assign n7748 = n7746 & n7747 ;
  assign n7749 = n7748 ^ x318 ;
  assign n7750 = x1072 ^ x319 ;
  assign n7751 = n7746 & n7750 ;
  assign n7752 = n7751 ^ x319 ;
  assign n7753 = x1048 ^ x320 ;
  assign n7754 = n7735 & n7753 ;
  assign n7755 = n7754 ^ x320 ;
  assign n7756 = x1058 ^ x321 ;
  assign n7757 = n7735 & n7756 ;
  assign n7758 = n7757 ^ x321 ;
  assign n7759 = x1051 ^ x322 ;
  assign n7760 = n7735 & n7759 ;
  assign n7761 = n7760 ^ x322 ;
  assign n7762 = x1065 ^ x323 ;
  assign n7763 = n7735 & n7762 ;
  assign n7764 = n7763 ^ x323 ;
  assign n7765 = x1086 ^ x324 ;
  assign n7766 = n7746 & n7765 ;
  assign n7767 = n7766 ^ x324 ;
  assign n7768 = x1063 ^ x325 ;
  assign n7769 = n7746 & n7768 ;
  assign n7770 = n7769 ^ x325 ;
  assign n7771 = x1057 ^ x326 ;
  assign n7772 = n7746 & n7771 ;
  assign n7773 = n7772 ^ x326 ;
  assign n7774 = x1040 ^ x327 ;
  assign n7775 = n7735 & n7774 ;
  assign n7776 = n7775 ^ x327 ;
  assign n7777 = x1058 ^ x328 ;
  assign n7778 = n7746 & n7777 ;
  assign n7779 = n7778 ^ x328 ;
  assign n7780 = x1043 ^ x329 ;
  assign n7781 = n7746 & n7780 ;
  assign n7782 = n7781 ^ x329 ;
  assign n7783 = x1091 & n2985 ;
  assign n7784 = n7783 ^ x1092 ;
  assign n7785 = n7742 ^ n7735 ;
  assign n7786 = n7785 ^ x330 ;
  assign n7787 = n7784 & ~n7786 ;
  assign n7789 = ~x331 & n7587 ;
  assign n7788 = n7746 ^ x331 ;
  assign n7790 = n7789 ^ n7788 ;
  assign n7791 = n7784 & ~n7790 ;
  assign n7792 = n1971 & n3881 ;
  assign n7793 = ~n3914 & ~n4064 ;
  assign n7794 = ~n1753 & n7793 ;
  assign n7795 = ~n7792 & n7794 ;
  assign n7796 = x1040 ^ x333 ;
  assign n7797 = n7746 & n7796 ;
  assign n7798 = n7797 ^ x333 ;
  assign n7799 = x1065 ^ x334 ;
  assign n7800 = n7746 & n7799 ;
  assign n7801 = n7800 ^ x334 ;
  assign n7802 = x1069 ^ x335 ;
  assign n7803 = n7746 & n7802 ;
  assign n7804 = n7803 ^ x335 ;
  assign n7805 = x1070 ^ x336 ;
  assign n7806 = n7742 & n7805 ;
  assign n7807 = n7806 ^ x336 ;
  assign n7808 = x1044 ^ x337 ;
  assign n7809 = n7742 & n7808 ;
  assign n7810 = n7809 ^ x337 ;
  assign n7811 = x1072 ^ x338 ;
  assign n7812 = n7742 & n7811 ;
  assign n7813 = n7812 ^ x338 ;
  assign n7814 = x1086 ^ x339 ;
  assign n7815 = n7742 & n7814 ;
  assign n7816 = n7815 ^ x339 ;
  assign n7817 = n7735 ^ x340 ;
  assign n7818 = n7817 ^ n7789 ;
  assign n7819 = n7784 & n7818 ;
  assign n7820 = n7746 ^ n7742 ;
  assign n7821 = n7820 ^ x341 ;
  assign n7822 = n7784 & ~n7821 ;
  assign n7823 = x1049 ^ x342 ;
  assign n7824 = n7735 & n7823 ;
  assign n7825 = n7824 ^ x342 ;
  assign n7826 = x1062 ^ x343 ;
  assign n7827 = n7735 & n7826 ;
  assign n7828 = n7827 ^ x343 ;
  assign n7829 = x1069 ^ x344 ;
  assign n7830 = n7735 & n7829 ;
  assign n7831 = n7830 ^ x344 ;
  assign n7832 = x1039 ^ x345 ;
  assign n7833 = n7735 & n7832 ;
  assign n7834 = n7833 ^ x345 ;
  assign n7835 = x1067 ^ x346 ;
  assign n7836 = n7735 & n7835 ;
  assign n7837 = n7836 ^ x346 ;
  assign n7838 = x1055 ^ x347 ;
  assign n7839 = n7735 & n7838 ;
  assign n7840 = n7839 ^ x347 ;
  assign n7841 = x1087 ^ x348 ;
  assign n7842 = n7735 & n7841 ;
  assign n7843 = n7842 ^ x348 ;
  assign n7844 = x1043 ^ x349 ;
  assign n7845 = n7735 & n7844 ;
  assign n7846 = n7845 ^ x349 ;
  assign n7847 = x1035 ^ x350 ;
  assign n7848 = n7735 & n7847 ;
  assign n7849 = n7848 ^ x350 ;
  assign n7850 = x1079 ^ x351 ;
  assign n7851 = n7735 & n7850 ;
  assign n7852 = n7851 ^ x351 ;
  assign n7853 = x1078 ^ x352 ;
  assign n7854 = n7735 & n7853 ;
  assign n7855 = n7854 ^ x352 ;
  assign n7856 = x1063 ^ x353 ;
  assign n7857 = n7735 & n7856 ;
  assign n7858 = n7857 ^ x353 ;
  assign n7859 = x1045 ^ x354 ;
  assign n7860 = n7735 & n7859 ;
  assign n7861 = n7860 ^ x354 ;
  assign n7862 = x1084 ^ x355 ;
  assign n7863 = n7735 & n7862 ;
  assign n7864 = n7863 ^ x355 ;
  assign n7865 = x1081 ^ x356 ;
  assign n7866 = n7735 & n7865 ;
  assign n7867 = n7866 ^ x356 ;
  assign n7868 = x1076 ^ x357 ;
  assign n7869 = n7735 & n7868 ;
  assign n7870 = n7869 ^ x357 ;
  assign n7871 = x1071 ^ x358 ;
  assign n7872 = n7735 & n7871 ;
  assign n7873 = n7872 ^ x358 ;
  assign n7874 = x1068 ^ x359 ;
  assign n7875 = n7735 & n7874 ;
  assign n7876 = n7875 ^ x359 ;
  assign n7877 = x1042 ^ x360 ;
  assign n7878 = n7735 & n7877 ;
  assign n7879 = n7878 ^ x360 ;
  assign n7880 = x1059 ^ x361 ;
  assign n7881 = n7735 & n7880 ;
  assign n7882 = n7881 ^ x361 ;
  assign n7883 = x1070 ^ x362 ;
  assign n7884 = n7735 & n7883 ;
  assign n7885 = n7884 ^ x362 ;
  assign n7886 = x1049 ^ x363 ;
  assign n7887 = n7742 & n7886 ;
  assign n7888 = n7887 ^ x363 ;
  assign n7889 = x1062 ^ x364 ;
  assign n7890 = n7742 & n7889 ;
  assign n7891 = n7890 ^ x364 ;
  assign n7892 = x1065 ^ x365 ;
  assign n7893 = n7742 & n7892 ;
  assign n7894 = n7893 ^ x365 ;
  assign n7895 = x1069 ^ x366 ;
  assign n7896 = n7742 & n7895 ;
  assign n7897 = n7896 ^ x366 ;
  assign n7898 = x1039 ^ x367 ;
  assign n7899 = n7742 & n7898 ;
  assign n7900 = n7899 ^ x367 ;
  assign n7901 = x1067 ^ x368 ;
  assign n7902 = n7742 & n7901 ;
  assign n7903 = n7902 ^ x368 ;
  assign n7904 = x1080 ^ x369 ;
  assign n7905 = n7742 & n7904 ;
  assign n7906 = n7905 ^ x369 ;
  assign n7907 = x1055 ^ x370 ;
  assign n7908 = n7742 & n7907 ;
  assign n7909 = n7908 ^ x370 ;
  assign n7910 = x1051 ^ x371 ;
  assign n7911 = n7742 & n7910 ;
  assign n7912 = n7911 ^ x371 ;
  assign n7913 = x1048 ^ x372 ;
  assign n7914 = n7742 & n7913 ;
  assign n7915 = n7914 ^ x372 ;
  assign n7916 = x1087 ^ x373 ;
  assign n7917 = n7742 & n7916 ;
  assign n7918 = n7917 ^ x373 ;
  assign n7919 = x1035 ^ x374 ;
  assign n7920 = n7742 & n7919 ;
  assign n7921 = n7920 ^ x374 ;
  assign n7922 = x1047 ^ x375 ;
  assign n7923 = n7742 & n7922 ;
  assign n7924 = n7923 ^ x375 ;
  assign n7925 = x1079 ^ x376 ;
  assign n7926 = n7742 & n7925 ;
  assign n7927 = n7926 ^ x376 ;
  assign n7928 = x1074 ^ x377 ;
  assign n7929 = n7742 & n7928 ;
  assign n7930 = n7929 ^ x377 ;
  assign n7931 = x1063 ^ x378 ;
  assign n7932 = n7742 & n7931 ;
  assign n7933 = n7932 ^ x378 ;
  assign n7934 = x1045 ^ x379 ;
  assign n7935 = n7742 & n7934 ;
  assign n7936 = n7935 ^ x379 ;
  assign n7937 = x1084 ^ x380 ;
  assign n7938 = n7742 & n7937 ;
  assign n7939 = n7938 ^ x380 ;
  assign n7940 = x1081 ^ x381 ;
  assign n7941 = n7742 & n7940 ;
  assign n7942 = n7941 ^ x381 ;
  assign n7943 = x1076 ^ x382 ;
  assign n7944 = n7742 & n7943 ;
  assign n7945 = n7944 ^ x382 ;
  assign n7946 = x1071 ^ x383 ;
  assign n7947 = n7742 & n7946 ;
  assign n7948 = n7947 ^ x383 ;
  assign n7949 = x1068 ^ x384 ;
  assign n7950 = n7742 & n7949 ;
  assign n7951 = n7950 ^ x384 ;
  assign n7952 = x1042 ^ x385 ;
  assign n7953 = n7742 & n7952 ;
  assign n7954 = n7953 ^ x385 ;
  assign n7955 = x1059 ^ x386 ;
  assign n7956 = n7742 & n7955 ;
  assign n7957 = n7956 ^ x386 ;
  assign n7958 = x1053 ^ x387 ;
  assign n7959 = n7742 & n7958 ;
  assign n7960 = n7959 ^ x387 ;
  assign n7961 = x1037 ^ x388 ;
  assign n7962 = n7742 & n7961 ;
  assign n7963 = n7962 ^ x388 ;
  assign n7964 = x1036 ^ x389 ;
  assign n7965 = n7742 & n7964 ;
  assign n7966 = n7965 ^ x389 ;
  assign n7967 = x1049 ^ x390 ;
  assign n7968 = n7746 & n7967 ;
  assign n7969 = n7968 ^ x390 ;
  assign n7970 = x1062 ^ x391 ;
  assign n7971 = n7746 & n7970 ;
  assign n7972 = n7971 ^ x391 ;
  assign n7973 = x1039 ^ x392 ;
  assign n7974 = n7746 & n7973 ;
  assign n7975 = n7974 ^ x392 ;
  assign n7976 = x1067 ^ x393 ;
  assign n7977 = n7746 & n7976 ;
  assign n7978 = n7977 ^ x393 ;
  assign n7979 = x1080 ^ x394 ;
  assign n7980 = n7746 & n7979 ;
  assign n7981 = n7980 ^ x394 ;
  assign n7982 = x1055 ^ x395 ;
  assign n7983 = n7746 & n7982 ;
  assign n7984 = n7983 ^ x395 ;
  assign n7985 = x1051 ^ x396 ;
  assign n7986 = n7746 & n7985 ;
  assign n7987 = n7986 ^ x396 ;
  assign n7988 = x1048 ^ x397 ;
  assign n7989 = n7746 & n7988 ;
  assign n7990 = n7989 ^ x397 ;
  assign n7991 = x1087 ^ x398 ;
  assign n7992 = n7746 & n7991 ;
  assign n7993 = n7992 ^ x398 ;
  assign n7994 = x1047 ^ x399 ;
  assign n7995 = n7746 & n7994 ;
  assign n7996 = n7995 ^ x399 ;
  assign n7997 = x1035 ^ x400 ;
  assign n7998 = n7746 & n7997 ;
  assign n7999 = n7998 ^ x400 ;
  assign n8000 = x1079 ^ x401 ;
  assign n8001 = n7746 & n8000 ;
  assign n8002 = n8001 ^ x401 ;
  assign n8003 = x1078 ^ x402 ;
  assign n8004 = n7746 & n8003 ;
  assign n8005 = n8004 ^ x402 ;
  assign n8006 = x1045 ^ x403 ;
  assign n8007 = n7746 & n8006 ;
  assign n8008 = n8007 ^ x403 ;
  assign n8009 = x1084 ^ x404 ;
  assign n8010 = n7746 & n8009 ;
  assign n8011 = n8010 ^ x404 ;
  assign n8012 = x1081 ^ x405 ;
  assign n8013 = n7746 & n8012 ;
  assign n8014 = n8013 ^ x405 ;
  assign n8015 = x1076 ^ x406 ;
  assign n8016 = n7746 & n8015 ;
  assign n8017 = n8016 ^ x406 ;
  assign n8018 = x1071 ^ x407 ;
  assign n8019 = n7746 & n8018 ;
  assign n8020 = n8019 ^ x407 ;
  assign n8021 = x1068 ^ x408 ;
  assign n8022 = n7746 & n8021 ;
  assign n8023 = n8022 ^ x408 ;
  assign n8024 = x1042 ^ x409 ;
  assign n8025 = n7746 & n8024 ;
  assign n8026 = n8025 ^ x409 ;
  assign n8027 = x1059 ^ x410 ;
  assign n8028 = n7746 & n8027 ;
  assign n8029 = n8028 ^ x410 ;
  assign n8030 = x1053 ^ x411 ;
  assign n8031 = n7746 & n8030 ;
  assign n8032 = n8031 ^ x411 ;
  assign n8033 = x1037 ^ x412 ;
  assign n8034 = n7746 & n8033 ;
  assign n8035 = n8034 ^ x412 ;
  assign n8036 = x1036 ^ x413 ;
  assign n8037 = n7746 & n8036 ;
  assign n8038 = n8037 ^ x413 ;
  assign n8039 = x1049 ^ x414 ;
  assign n8040 = n7789 & n8039 ;
  assign n8041 = n8040 ^ x414 ;
  assign n8042 = x1062 ^ x415 ;
  assign n8043 = n7789 & n8042 ;
  assign n8044 = n8043 ^ x415 ;
  assign n8045 = x1069 ^ x416 ;
  assign n8046 = n7789 & n8045 ;
  assign n8047 = n8046 ^ x416 ;
  assign n8048 = x1039 ^ x417 ;
  assign n8049 = n7789 & n8048 ;
  assign n8050 = n8049 ^ x417 ;
  assign n8051 = x1067 ^ x418 ;
  assign n8052 = n7789 & n8051 ;
  assign n8053 = n8052 ^ x418 ;
  assign n8054 = x1080 ^ x419 ;
  assign n8055 = n7789 & n8054 ;
  assign n8056 = n8055 ^ x419 ;
  assign n8057 = x1055 ^ x420 ;
  assign n8058 = n7789 & n8057 ;
  assign n8059 = n8058 ^ x420 ;
  assign n8060 = x1051 ^ x421 ;
  assign n8061 = n7789 & n8060 ;
  assign n8062 = n8061 ^ x421 ;
  assign n8063 = x1048 ^ x422 ;
  assign n8064 = n7789 & n8063 ;
  assign n8065 = n8064 ^ x422 ;
  assign n8066 = x1087 ^ x423 ;
  assign n8067 = n7789 & n8066 ;
  assign n8068 = n8067 ^ x423 ;
  assign n8069 = x1047 ^ x424 ;
  assign n8070 = n7789 & n8069 ;
  assign n8071 = n8070 ^ x424 ;
  assign n8072 = x1035 ^ x425 ;
  assign n8073 = n7789 & n8072 ;
  assign n8074 = n8073 ^ x425 ;
  assign n8075 = x1079 ^ x426 ;
  assign n8076 = n7789 & n8075 ;
  assign n8077 = n8076 ^ x426 ;
  assign n8078 = x1078 ^ x427 ;
  assign n8079 = n7789 & n8078 ;
  assign n8080 = n8079 ^ x427 ;
  assign n8081 = x1045 ^ x428 ;
  assign n8082 = n7789 & n8081 ;
  assign n8083 = n8082 ^ x428 ;
  assign n8084 = x1084 ^ x429 ;
  assign n8085 = n7789 & n8084 ;
  assign n8086 = n8085 ^ x429 ;
  assign n8087 = x1076 ^ x430 ;
  assign n8088 = n7789 & n8087 ;
  assign n8089 = n8088 ^ x430 ;
  assign n8090 = x1071 ^ x431 ;
  assign n8091 = n7789 & n8090 ;
  assign n8092 = n8091 ^ x431 ;
  assign n8093 = x1068 ^ x432 ;
  assign n8094 = n7789 & n8093 ;
  assign n8095 = n8094 ^ x432 ;
  assign n8096 = x1042 ^ x433 ;
  assign n8097 = n7789 & n8096 ;
  assign n8098 = n8097 ^ x433 ;
  assign n8099 = x1059 ^ x434 ;
  assign n8100 = n7789 & n8099 ;
  assign n8101 = n8100 ^ x434 ;
  assign n8102 = x1053 ^ x435 ;
  assign n8103 = n7789 & n8102 ;
  assign n8104 = n8103 ^ x435 ;
  assign n8105 = x1037 ^ x436 ;
  assign n8106 = n7789 & n8105 ;
  assign n8107 = n8106 ^ x436 ;
  assign n8108 = x1070 ^ x437 ;
  assign n8109 = n7789 & n8108 ;
  assign n8110 = n8109 ^ x437 ;
  assign n8111 = x1036 ^ x438 ;
  assign n8112 = n7789 & n8111 ;
  assign n8113 = n8112 ^ x438 ;
  assign n8114 = x1057 ^ x439 ;
  assign n8115 = n7742 & n8114 ;
  assign n8116 = n8115 ^ x439 ;
  assign n8117 = x1043 ^ x440 ;
  assign n8118 = n7742 & n8117 ;
  assign n8119 = n8118 ^ x440 ;
  assign n8120 = x1044 ^ x441 ;
  assign n8121 = n7735 & n8120 ;
  assign n8122 = n8121 ^ x441 ;
  assign n8123 = x1058 ^ x442 ;
  assign n8124 = n7742 & n8123 ;
  assign n8125 = n8124 ^ x442 ;
  assign n8126 = x1044 ^ x443 ;
  assign n8127 = n7789 & n8126 ;
  assign n8128 = n8127 ^ x443 ;
  assign n8129 = x1072 ^ x444 ;
  assign n8130 = n7789 & n8129 ;
  assign n8131 = n8130 ^ x444 ;
  assign n8132 = x1081 ^ x445 ;
  assign n8133 = n7789 & n8132 ;
  assign n8134 = n8133 ^ x445 ;
  assign n8135 = x1086 ^ x446 ;
  assign n8136 = n7789 & n8135 ;
  assign n8137 = n8136 ^ x446 ;
  assign n8138 = x1040 ^ x447 ;
  assign n8139 = n7742 & n8138 ;
  assign n8140 = n8139 ^ x447 ;
  assign n8141 = x1074 ^ x448 ;
  assign n8142 = n7789 & n8141 ;
  assign n8143 = n8142 ^ x448 ;
  assign n8144 = x1057 ^ x449 ;
  assign n8145 = n7789 & n8144 ;
  assign n8146 = n8145 ^ x449 ;
  assign n8147 = x1036 ^ x450 ;
  assign n8148 = n7735 & n8147 ;
  assign n8149 = n8148 ^ x450 ;
  assign n8150 = x1063 ^ x451 ;
  assign n8151 = n7789 & n8150 ;
  assign n8152 = n8151 ^ x451 ;
  assign n8153 = x1053 ^ x452 ;
  assign n8154 = n7735 & n8153 ;
  assign n8155 = n8154 ^ x452 ;
  assign n8156 = x1040 ^ x453 ;
  assign n8157 = n7789 & n8156 ;
  assign n8158 = n8157 ^ x453 ;
  assign n8159 = x1043 ^ x454 ;
  assign n8160 = n7789 & n8159 ;
  assign n8161 = n8160 ^ x454 ;
  assign n8162 = x1037 ^ x455 ;
  assign n8163 = n7735 & n8162 ;
  assign n8164 = n8163 ^ x455 ;
  assign n8165 = x1044 ^ x456 ;
  assign n8166 = n7746 & n8165 ;
  assign n8167 = n8166 ^ x456 ;
  assign n8168 = x594 & x600 ;
  assign n8169 = x597 & x601 ;
  assign n8170 = n8168 & n8169 ;
  assign n8171 = n8170 ^ x804 ;
  assign n8172 = n8171 ^ x595 ;
  assign n8175 = x804 ^ x596 ;
  assign n8176 = n8175 ^ x810 ;
  assign n8177 = x815 ^ x804 ;
  assign n8178 = n8177 ^ n8176 ;
  assign n8179 = x815 ^ x810 ;
  assign n8180 = n8179 ^ n8176 ;
  assign n8181 = x810 ^ x599 ;
  assign n8182 = n8181 ^ x804 ;
  assign n8183 = n8180 & n8182 ;
  assign n8184 = n8178 & n8183 ;
  assign n8185 = n8184 ^ x810 ;
  assign n8186 = n8185 ^ x804 ;
  assign n8187 = n8176 & n8186 ;
  assign n8188 = x804 & n8187 ;
  assign n8173 = x810 ^ x804 ;
  assign n8189 = n8188 ^ n8173 ;
  assign n8190 = n8172 & n8189 ;
  assign n8191 = n8190 ^ x804 ;
  assign n8192 = n8170 & ~n8191 ;
  assign n8193 = x600 & x804 ;
  assign n8194 = ~x810 & n8193 ;
  assign n8195 = n8194 ^ x804 ;
  assign n8196 = ~x601 & ~x815 ;
  assign n8204 = ~x804 & n8196 ;
  assign n8205 = ~x810 & n8204 ;
  assign n8206 = n8205 ^ x810 ;
  assign n8197 = n8196 ^ x815 ;
  assign n8198 = n8197 ^ x810 ;
  assign n8207 = n8206 ^ n8198 ;
  assign n8208 = ~n8195 & ~n8207 ;
  assign n8209 = ~n8192 & ~n8208 ;
  assign n8210 = x605 & ~n8209 ;
  assign n8211 = ~x815 & x990 ;
  assign n8212 = n8168 & n8211 ;
  assign n8213 = n8195 & n8212 ;
  assign n8214 = ~n8210 & ~n8213 ;
  assign n8215 = x821 & ~n8214 ;
  assign n8216 = x1072 ^ x458 ;
  assign n8217 = n7735 & n8216 ;
  assign n8218 = n8217 ^ x458 ;
  assign n8219 = x1058 ^ x459 ;
  assign n8220 = n7789 & n8219 ;
  assign n8221 = n8220 ^ x459 ;
  assign n8222 = x1086 ^ x460 ;
  assign n8223 = n7735 & n8222 ;
  assign n8224 = n8223 ^ x460 ;
  assign n8225 = x1057 ^ x461 ;
  assign n8226 = n7735 & n8225 ;
  assign n8227 = n8226 ^ x461 ;
  assign n8228 = x1074 ^ x462 ;
  assign n8229 = n7735 & n8228 ;
  assign n8230 = n8229 ^ x462 ;
  assign n8231 = x1070 ^ x463 ;
  assign n8232 = n7746 & n8231 ;
  assign n8233 = n8232 ^ x463 ;
  assign n8234 = x1065 ^ x464 ;
  assign n8235 = n7789 & n8234 ;
  assign n8236 = n8235 ^ x464 ;
  assign n8239 = x1157 & n2591 ;
  assign n8238 = ~x243 & n7680 ;
  assign n8240 = n8239 ^ n8238 ;
  assign n8237 = x926 & n7672 ;
  assign n8241 = n8240 ^ n8237 ;
  assign n8244 = x1151 & n2591 ;
  assign n8243 = x275 & n7680 ;
  assign n8245 = n8244 ^ n8243 ;
  assign n8242 = x943 & n7672 ;
  assign n8246 = n8245 ^ n8242 ;
  assign n8247 = n4318 & n6729 ;
  assign n8248 = x40 & x1001 ;
  assign n8249 = n2631 & n8248 ;
  assign n8250 = n2647 & n8249 ;
  assign n8251 = ~n8247 & ~n8250 ;
  assign n8252 = x468 & ~n3890 ;
  assign n8253 = ~n4293 & n8252 ;
  assign n8254 = n8253 ^ n4293 ;
  assign n8257 = x1156 & n2591 ;
  assign n8256 = ~x263 & n7680 ;
  assign n8258 = n8257 ^ n8256 ;
  assign n8255 = x942 & n7672 ;
  assign n8259 = n8258 ^ n8255 ;
  assign n8262 = x1155 & n2591 ;
  assign n8261 = x267 & n7680 ;
  assign n8263 = n8262 ^ n8261 ;
  assign n8260 = x925 & n7672 ;
  assign n8264 = n8263 ^ n8260 ;
  assign n8267 = x1153 & n2591 ;
  assign n8266 = x253 & n7680 ;
  assign n8268 = n8267 ^ n8266 ;
  assign n8265 = x941 & n7672 ;
  assign n8269 = n8268 ^ n8265 ;
  assign n8272 = x1154 & n2591 ;
  assign n8271 = x254 & n7680 ;
  assign n8273 = n8272 ^ n8271 ;
  assign n8270 = x923 & n7672 ;
  assign n8274 = n8273 ^ n8270 ;
  assign n8277 = x1152 & n2591 ;
  assign n8276 = x268 & n7680 ;
  assign n8278 = n8277 ^ n8276 ;
  assign n8275 = x922 & n7672 ;
  assign n8279 = n8278 ^ n8275 ;
  assign n8282 = x1150 & n2591 ;
  assign n8281 = x272 & n7680 ;
  assign n8283 = n8282 ^ n8281 ;
  assign n8280 = x931 & n7672 ;
  assign n8284 = n8283 ^ n8280 ;
  assign n8287 = x1149 & n2591 ;
  assign n8286 = x283 & n7680 ;
  assign n8288 = n8287 ^ n8286 ;
  assign n8285 = x936 & n7672 ;
  assign n8289 = n8288 ^ n8285 ;
  assign n8290 = x71 & ~n4034 ;
  assign n8292 = n8290 ^ n4624 ;
  assign n8293 = x71 & n7185 ;
  assign n8294 = x481 ^ x248 ;
  assign n8295 = ~n6445 & n8294 ;
  assign n8296 = n8295 ^ x248 ;
  assign n8297 = x482 ^ x249 ;
  assign n8298 = ~n6461 & n8297 ;
  assign n8299 = n8298 ^ x249 ;
  assign n8300 = x483 ^ x242 ;
  assign n8301 = ~n6493 & n8300 ;
  assign n8302 = n8301 ^ x242 ;
  assign n8303 = x484 ^ x249 ;
  assign n8304 = ~n6493 & n8303 ;
  assign n8305 = n8304 ^ x249 ;
  assign n8306 = x485 ^ x234 ;
  assign n8307 = ~n6492 & n8306 ;
  assign n8308 = n8307 ^ x234 ;
  assign n8309 = x486 ^ x244 ;
  assign n8310 = ~n6492 & n8309 ;
  assign n8311 = n8310 ^ x244 ;
  assign n8312 = x487 ^ x246 ;
  assign n8313 = ~n6445 & n8312 ;
  assign n8314 = n8313 ^ x246 ;
  assign n8315 = x488 ^ x239 ;
  assign n8316 = ~n6445 & ~n8315 ;
  assign n8317 = n8316 ^ x239 ;
  assign n8318 = x489 ^ x242 ;
  assign n8319 = ~n6492 & n8318 ;
  assign n8320 = n8319 ^ x242 ;
  assign n8321 = x490 ^ x241 ;
  assign n8322 = ~n6493 & n8321 ;
  assign n8323 = n8322 ^ x241 ;
  assign n8324 = x491 ^ x238 ;
  assign n8325 = ~n6493 & n8324 ;
  assign n8326 = n8325 ^ x238 ;
  assign n8327 = x492 ^ x240 ;
  assign n8328 = ~n6493 & n8327 ;
  assign n8329 = n8328 ^ x240 ;
  assign n8330 = x493 ^ x244 ;
  assign n8331 = ~n6493 & n8330 ;
  assign n8332 = n8331 ^ x244 ;
  assign n8333 = x494 ^ x239 ;
  assign n8334 = ~n6493 & ~n8333 ;
  assign n8335 = n8334 ^ x239 ;
  assign n8336 = x495 ^ x235 ;
  assign n8337 = ~n6493 & n8336 ;
  assign n8338 = n8337 ^ x235 ;
  assign n8339 = x496 ^ x249 ;
  assign n8340 = ~n6478 & n8339 ;
  assign n8341 = n8340 ^ x249 ;
  assign n8342 = x497 ^ x239 ;
  assign n8343 = ~n6478 & ~n8342 ;
  assign n8344 = n8343 ^ x239 ;
  assign n8345 = x498 ^ x238 ;
  assign n8346 = ~n6461 & n8345 ;
  assign n8347 = n8346 ^ x238 ;
  assign n8348 = x499 ^ x246 ;
  assign n8349 = ~n6478 & n8348 ;
  assign n8350 = n8349 ^ x246 ;
  assign n8351 = x500 ^ x241 ;
  assign n8352 = ~n6478 & n8351 ;
  assign n8353 = n8352 ^ x241 ;
  assign n8354 = x501 ^ x248 ;
  assign n8355 = ~n6478 & n8354 ;
  assign n8356 = n8355 ^ x248 ;
  assign n8357 = x502 ^ x247 ;
  assign n8358 = ~n6478 & n8357 ;
  assign n8359 = n8358 ^ x247 ;
  assign n8360 = x503 ^ x245 ;
  assign n8361 = ~n6478 & n8360 ;
  assign n8362 = n8361 ^ x245 ;
  assign n8363 = x504 ^ x242 ;
  assign n8364 = ~n6479 & n8363 ;
  assign n8365 = n8364 ^ x242 ;
  assign n8366 = x505 ^ x234 ;
  assign n8367 = ~n6478 & n8366 ;
  assign n8368 = n8367 ^ x234 ;
  assign n8369 = x506 ^ x241 ;
  assign n8370 = ~n6479 & n8369 ;
  assign n8371 = n8370 ^ x241 ;
  assign n8372 = x507 ^ x238 ;
  assign n8373 = ~n6479 & n8372 ;
  assign n8374 = n8373 ^ x238 ;
  assign n8375 = x508 ^ x247 ;
  assign n8376 = ~n6479 & n8375 ;
  assign n8377 = n8376 ^ x247 ;
  assign n8378 = x509 ^ x245 ;
  assign n8379 = ~n6479 & n8378 ;
  assign n8380 = n8379 ^ x245 ;
  assign n8381 = x510 ^ x242 ;
  assign n8382 = ~n6445 & n8381 ;
  assign n8383 = n8382 ^ x242 ;
  assign n8384 = x511 ^ x234 ;
  assign n8385 = ~n6445 & n8384 ;
  assign n8386 = n8385 ^ x234 ;
  assign n8387 = x512 ^ x235 ;
  assign n8388 = ~n6445 & n8387 ;
  assign n8389 = n8388 ^ x235 ;
  assign n8390 = x513 ^ x244 ;
  assign n8391 = ~n6445 & n8390 ;
  assign n8392 = n8391 ^ x244 ;
  assign n8393 = x514 ^ x245 ;
  assign n8394 = ~n6445 & n8393 ;
  assign n8395 = n8394 ^ x245 ;
  assign n8396 = x515 ^ x240 ;
  assign n8397 = ~n6445 & n8396 ;
  assign n8398 = n8397 ^ x240 ;
  assign n8399 = x516 ^ x247 ;
  assign n8400 = ~n6445 & n8399 ;
  assign n8401 = n8400 ^ x247 ;
  assign n8402 = x517 ^ x238 ;
  assign n8403 = ~n6445 & n8402 ;
  assign n8404 = n8403 ^ x238 ;
  assign n8405 = x518 ^ x234 ;
  assign n8406 = ~n6454 & n8405 ;
  assign n8407 = n8406 ^ x234 ;
  assign n8408 = x519 ^ x239 ;
  assign n8409 = ~n6454 & ~n8408 ;
  assign n8410 = n8409 ^ x239 ;
  assign n8411 = x520 ^ x246 ;
  assign n8412 = ~n6454 & n8411 ;
  assign n8413 = n8412 ^ x246 ;
  assign n8414 = x521 ^ x248 ;
  assign n8415 = ~n6454 & n8414 ;
  assign n8416 = n8415 ^ x248 ;
  assign n8417 = x522 ^ x238 ;
  assign n8418 = ~n6454 & n8417 ;
  assign n8419 = n8418 ^ x238 ;
  assign n8420 = x523 ^ x234 ;
  assign n8421 = ~n6627 & n8420 ;
  assign n8422 = n8421 ^ x234 ;
  assign n8423 = x524 ^ x239 ;
  assign n8424 = ~n6627 & ~n8423 ;
  assign n8425 = n8424 ^ x239 ;
  assign n8426 = x525 ^ x245 ;
  assign n8427 = ~n6627 & n8426 ;
  assign n8428 = n8427 ^ x245 ;
  assign n8429 = x526 ^ x246 ;
  assign n8430 = ~n6627 & n8429 ;
  assign n8431 = n8430 ^ x246 ;
  assign n8432 = x527 ^ x247 ;
  assign n8433 = ~n6627 & n8432 ;
  assign n8434 = n8433 ^ x247 ;
  assign n8435 = x528 ^ x249 ;
  assign n8436 = ~n6627 & n8435 ;
  assign n8437 = n8436 ^ x249 ;
  assign n8438 = x529 ^ x238 ;
  assign n8439 = ~n6627 & n8438 ;
  assign n8440 = n8439 ^ x238 ;
  assign n8441 = x530 ^ x240 ;
  assign n8442 = ~n6627 & n8441 ;
  assign n8443 = n8442 ^ x240 ;
  assign n8444 = x531 ^ x235 ;
  assign n8445 = ~n6461 & n8444 ;
  assign n8446 = n8445 ^ x235 ;
  assign n8447 = x532 ^ x247 ;
  assign n8448 = ~n6461 & n8447 ;
  assign n8449 = n8448 ^ x247 ;
  assign n8450 = x533 ^ x235 ;
  assign n8451 = ~n6479 & n8450 ;
  assign n8452 = n8451 ^ x235 ;
  assign n8453 = x534 ^ x239 ;
  assign n8454 = ~n6479 & ~n8453 ;
  assign n8455 = n8454 ^ x239 ;
  assign n8456 = x535 ^ x240 ;
  assign n8457 = ~n6479 & n8456 ;
  assign n8458 = n8457 ^ x240 ;
  assign n8459 = x536 ^ x246 ;
  assign n8460 = ~n6479 & n8459 ;
  assign n8461 = n8460 ^ x246 ;
  assign n8462 = x537 ^ x248 ;
  assign n8463 = ~n6479 & n8462 ;
  assign n8464 = n8463 ^ x248 ;
  assign n8465 = x538 ^ x249 ;
  assign n8466 = ~n6479 & n8465 ;
  assign n8467 = n8466 ^ x249 ;
  assign n8468 = x539 ^ x242 ;
  assign n8469 = ~n6478 & n8468 ;
  assign n8470 = n8469 ^ x242 ;
  assign n8471 = x540 ^ x235 ;
  assign n8472 = ~n6478 & n8471 ;
  assign n8473 = n8472 ^ x235 ;
  assign n8474 = x541 ^ x244 ;
  assign n8475 = ~n6478 & n8474 ;
  assign n8476 = n8475 ^ x244 ;
  assign n8477 = x542 ^ x240 ;
  assign n8478 = ~n6478 & n8477 ;
  assign n8479 = n8478 ^ x240 ;
  assign n8480 = x543 ^ x238 ;
  assign n8481 = ~n6478 & n8480 ;
  assign n8482 = n8481 ^ x238 ;
  assign n8483 = x544 ^ x234 ;
  assign n8484 = ~n6493 & n8483 ;
  assign n8485 = n8484 ^ x234 ;
  assign n8486 = x545 ^ x245 ;
  assign n8487 = ~n6493 & n8486 ;
  assign n8488 = n8487 ^ x245 ;
  assign n8489 = x546 ^ x246 ;
  assign n8490 = ~n6493 & n8489 ;
  assign n8491 = n8490 ^ x246 ;
  assign n8492 = x547 ^ x247 ;
  assign n8493 = ~n6493 & n8492 ;
  assign n8494 = n8493 ^ x247 ;
  assign n8495 = x548 ^ x248 ;
  assign n8496 = ~n6493 & n8495 ;
  assign n8497 = n8496 ^ x248 ;
  assign n8498 = x549 ^ x235 ;
  assign n8499 = ~n6492 & n8498 ;
  assign n8500 = n8499 ^ x235 ;
  assign n8501 = x550 ^ x239 ;
  assign n8502 = ~n6492 & ~n8501 ;
  assign n8503 = n8502 ^ x239 ;
  assign n8504 = x551 ^ x240 ;
  assign n8505 = ~n6492 & n8504 ;
  assign n8506 = n8505 ^ x240 ;
  assign n8507 = x552 ^ x247 ;
  assign n8508 = ~n6492 & n8507 ;
  assign n8509 = n8508 ^ x247 ;
  assign n8510 = x553 ^ x241 ;
  assign n8511 = ~n6492 & n8510 ;
  assign n8512 = n8511 ^ x241 ;
  assign n8513 = x554 ^ x248 ;
  assign n8514 = ~n6492 & n8513 ;
  assign n8515 = n8514 ^ x248 ;
  assign n8516 = x555 ^ x249 ;
  assign n8517 = ~n6492 & n8516 ;
  assign n8518 = n8517 ^ x249 ;
  assign n8519 = x556 ^ x242 ;
  assign n8520 = ~n6461 & n8519 ;
  assign n8521 = n8520 ^ x242 ;
  assign n8522 = x557 ^ x234 ;
  assign n8523 = ~n6479 & n8522 ;
  assign n8524 = n8523 ^ x234 ;
  assign n8525 = x558 ^ x244 ;
  assign n8526 = ~n6479 & n8525 ;
  assign n8527 = n8526 ^ x244 ;
  assign n8528 = x559 ^ x241 ;
  assign n8529 = ~n6445 & n8528 ;
  assign n8530 = n8529 ^ x241 ;
  assign n8531 = x560 ^ x240 ;
  assign n8532 = ~n6461 & n8531 ;
  assign n8533 = n8532 ^ x240 ;
  assign n8534 = x561 ^ x247 ;
  assign n8535 = ~n6454 & n8534 ;
  assign n8536 = n8535 ^ x247 ;
  assign n8537 = x562 ^ x241 ;
  assign n8538 = ~n6461 & n8537 ;
  assign n8539 = n8538 ^ x241 ;
  assign n8540 = x563 ^ x246 ;
  assign n8541 = ~n6492 & n8540 ;
  assign n8542 = n8541 ^ x246 ;
  assign n8543 = x564 ^ x246 ;
  assign n8544 = ~n6461 & n8543 ;
  assign n8545 = n8544 ^ x246 ;
  assign n8546 = x565 ^ x248 ;
  assign n8547 = ~n6461 & n8546 ;
  assign n8548 = n8547 ^ x248 ;
  assign n8549 = x566 ^ x244 ;
  assign n8550 = ~n6461 & n8549 ;
  assign n8551 = n8550 ^ x244 ;
  assign n8552 = x230 & x1093 ;
  assign n8556 = n5774 ^ x567 ;
  assign n8553 = n5774 ^ x1091 ;
  assign n8554 = x621 & n5717 ;
  assign n8555 = n8553 & n8554 ;
  assign n8557 = n8556 ^ n8555 ;
  assign n8558 = n8552 & ~n8557 ;
  assign n8559 = n8558 ^ x567 ;
  assign n8560 = x1092 & ~n8559 ;
  assign n8561 = x568 ^ x245 ;
  assign n8562 = ~n6461 & n8561 ;
  assign n8563 = n8562 ^ x245 ;
  assign n8564 = x569 ^ x239 ;
  assign n8565 = ~n6461 & ~n8564 ;
  assign n8566 = n8565 ^ x239 ;
  assign n8567 = x570 ^ x234 ;
  assign n8568 = ~n6461 & n8567 ;
  assign n8569 = n8568 ^ x234 ;
  assign n8570 = x571 ^ x241 ;
  assign n8571 = ~n6627 & n8570 ;
  assign n8572 = n8571 ^ x241 ;
  assign n8573 = x572 ^ x244 ;
  assign n8574 = ~n6627 & n8573 ;
  assign n8575 = n8574 ^ x244 ;
  assign n8576 = x573 ^ x242 ;
  assign n8577 = ~n6627 & n8576 ;
  assign n8578 = n8577 ^ x242 ;
  assign n8579 = x574 ^ x241 ;
  assign n8580 = ~n6454 & n8579 ;
  assign n8581 = n8580 ^ x241 ;
  assign n8582 = x575 ^ x235 ;
  assign n8583 = ~n6627 & n8582 ;
  assign n8584 = n8583 ^ x235 ;
  assign n8585 = x576 ^ x248 ;
  assign n8586 = ~n6627 & n8585 ;
  assign n8587 = n8586 ^ x248 ;
  assign n8588 = x577 ^ x238 ;
  assign n8589 = ~n6492 & n8588 ;
  assign n8590 = n8589 ^ x238 ;
  assign n8591 = x578 ^ x249 ;
  assign n8592 = ~n6454 & n8591 ;
  assign n8593 = n8592 ^ x249 ;
  assign n8594 = x579 ^ x249 ;
  assign n8595 = ~n6445 & n8594 ;
  assign n8596 = n8595 ^ x249 ;
  assign n8597 = x580 ^ x245 ;
  assign n8598 = ~n6492 & n8597 ;
  assign n8599 = n8598 ^ x245 ;
  assign n8600 = x581 ^ x235 ;
  assign n8601 = ~n6454 & n8600 ;
  assign n8602 = n8601 ^ x235 ;
  assign n8603 = x582 ^ x240 ;
  assign n8604 = ~n6454 & n8603 ;
  assign n8605 = n8604 ^ x240 ;
  assign n8606 = x584 ^ x245 ;
  assign n8607 = ~n6454 & n8606 ;
  assign n8608 = n8607 ^ x245 ;
  assign n8609 = x585 ^ x244 ;
  assign n8610 = ~n6454 & n8609 ;
  assign n8611 = n8610 ^ x244 ;
  assign n8612 = x586 ^ x242 ;
  assign n8613 = ~n6454 & n8612 ;
  assign n8614 = n8613 ^ x242 ;
  assign n8615 = n5719 ^ x587 ;
  assign n8616 = x230 & n8615 ;
  assign n8617 = n8616 ^ x587 ;
  assign n8618 = x591 ^ x588 ;
  assign n8619 = ~x123 & x824 ;
  assign n8620 = x950 & n8619 ;
  assign n8623 = n8618 & ~n8620 ;
  assign n8624 = n8623 ^ x591 ;
  assign n8625 = n7784 & n8624 ;
  assign n8626 = x218 ^ x205 ;
  assign n8627 = ~x237 & n8626 ;
  assign n8628 = n8627 ^ x205 ;
  assign n8630 = n8628 ^ x204 ;
  assign n8629 = n8628 ^ x206 ;
  assign n8631 = n8630 ^ n8629 ;
  assign n8634 = x237 & n8631 ;
  assign n8635 = n8634 ^ n8629 ;
  assign n8636 = x233 & n8635 ;
  assign n8637 = n8636 ^ n8628 ;
  assign n8638 = n6475 & ~n8637 ;
  assign n8639 = x203 ^ x202 ;
  assign n8640 = ~x237 & n8639 ;
  assign n8641 = n8640 ^ x202 ;
  assign n8643 = n8641 ^ x201 ;
  assign n8642 = n8641 ^ x220 ;
  assign n8644 = n8643 ^ n8642 ;
  assign n8647 = x237 & n8644 ;
  assign n8648 = n8647 ^ n8642 ;
  assign n8649 = x233 & n8648 ;
  assign n8650 = n8649 ^ n8641 ;
  assign n8651 = n6438 & ~n8650 ;
  assign n8652 = ~n8638 & n8651 ;
  assign n8653 = n8652 ^ n8638 ;
  assign n8654 = x590 ^ x588 ;
  assign n8657 = n8620 & n8654 ;
  assign n8658 = n8657 ^ x590 ;
  assign n8659 = n7784 & ~n8658 ;
  assign n8660 = x592 ^ x591 ;
  assign n8663 = n8620 & n8660 ;
  assign n8664 = n8663 ^ x591 ;
  assign n8665 = n7784 & n8664 ;
  assign n8666 = x592 ^ x590 ;
  assign n8669 = n8620 & n8666 ;
  assign n8670 = n8669 ^ x592 ;
  assign n8671 = n7784 & n8670 ;
  assign n8699 = ~n8540 & ~n8588 ;
  assign n8700 = ~n8306 & ~n8597 ;
  assign n8701 = n8699 & n8700 ;
  assign n8702 = ~n8498 & ~n8516 ;
  assign n8703 = n8501 & ~n8510 ;
  assign n8704 = n8702 & n8703 ;
  assign n8705 = n8701 & n8704 ;
  assign n8706 = ~x233 & ~n8507 ;
  assign n8707 = ~n8318 & n8706 ;
  assign n8708 = ~n8309 & ~n8513 ;
  assign n8709 = ~n8504 & n8708 ;
  assign n8710 = n8707 & n8709 ;
  assign n8711 = n8705 & n8710 ;
  assign n8712 = ~n8303 & ~n8489 ;
  assign n8713 = ~n8330 & ~n8495 ;
  assign n8714 = n8712 & n8713 ;
  assign n8715 = ~n8327 & ~n8483 ;
  assign n8716 = n8333 & ~n8336 ;
  assign n8717 = n8715 & n8716 ;
  assign n8718 = n8714 & n8717 ;
  assign n8719 = x233 & ~n8486 ;
  assign n8720 = ~n8321 & n8719 ;
  assign n8721 = ~n8300 & ~n8492 ;
  assign n8722 = ~n8324 & n8721 ;
  assign n8723 = n8720 & n8722 ;
  assign n8724 = n8718 & n8723 ;
  assign n8725 = ~n8711 & ~n8724 ;
  assign n8672 = ~n8456 & ~n8522 ;
  assign n8673 = ~n8369 & ~n8525 ;
  assign n8674 = n8672 & n8673 ;
  assign n8675 = ~n8378 & ~n8462 ;
  assign n8676 = n8453 & ~n8459 ;
  assign n8677 = n8675 & n8676 ;
  assign n8678 = n8674 & n8677 ;
  assign n8679 = x233 & ~n8450 ;
  assign n8680 = ~n8372 & n8679 ;
  assign n8681 = ~n8363 & ~n8465 ;
  assign n8682 = ~n8375 & n8681 ;
  assign n8683 = n8680 & n8682 ;
  assign n8684 = n8678 & n8683 ;
  assign n8685 = ~n8354 & ~n8480 ;
  assign n8686 = ~n8357 & ~n8471 ;
  assign n8687 = n8685 & n8686 ;
  assign n8688 = ~n8366 & ~n8474 ;
  assign n8689 = n8342 & ~n8477 ;
  assign n8690 = n8688 & n8689 ;
  assign n8691 = n8687 & n8690 ;
  assign n8692 = ~x233 & ~n8351 ;
  assign n8693 = ~n8339 & n8692 ;
  assign n8694 = ~n8360 & ~n8468 ;
  assign n8695 = n8693 & n8694 ;
  assign n8696 = ~n8348 & n8695 ;
  assign n8697 = n8691 & n8696 ;
  assign n8698 = ~n8684 & ~n8697 ;
  assign n8726 = n8725 ^ n8698 ;
  assign n8727 = x237 & n8726 ;
  assign n8728 = n8727 ^ n8725 ;
  assign n8729 = n6475 & ~n8728 ;
  assign n8730 = ~n8384 & ~n8390 ;
  assign n8731 = ~n8381 & ~n8396 ;
  assign n8732 = n8730 & n8731 ;
  assign n8733 = n8315 & ~n8387 ;
  assign n8734 = ~n8312 & ~n8402 ;
  assign n8735 = n8733 & n8734 ;
  assign n8736 = n8732 & n8735 ;
  assign n8737 = x233 & ~n8528 ;
  assign n8738 = ~n8393 & n8737 ;
  assign n8739 = ~n8294 & ~n8594 ;
  assign n8740 = ~n8399 & n8739 ;
  assign n8741 = n8738 & n8740 ;
  assign n8742 = n8736 & n8741 ;
  assign n8743 = x237 & ~n8742 ;
  assign n8744 = n8408 & ~n8606 ;
  assign n8745 = ~n8405 & ~n8411 ;
  assign n8746 = n8744 & n8745 ;
  assign n8747 = ~n8534 & ~n8612 ;
  assign n8748 = ~n8600 & ~n8603 ;
  assign n8749 = n8747 & n8748 ;
  assign n8750 = n8746 & n8749 ;
  assign n8751 = ~x233 & ~n8591 ;
  assign n8752 = ~n8417 & n8751 ;
  assign n8753 = ~n8414 & ~n8609 ;
  assign n8754 = ~n8579 & n8753 ;
  assign n8755 = n8752 & n8754 ;
  assign n8756 = n8750 & n8755 ;
  assign n8757 = n8743 & ~n8756 ;
  assign n8758 = n6438 & ~n8757 ;
  assign n8759 = n8423 & ~n8426 ;
  assign n8760 = ~n8435 & ~n8438 ;
  assign n8761 = n8759 & n8760 ;
  assign n8762 = ~n8429 & ~n8582 ;
  assign n8763 = ~n8420 & ~n8576 ;
  assign n8764 = n8762 & n8763 ;
  assign n8765 = n8761 & n8764 ;
  assign n8766 = x244 & ~x572 ;
  assign n8767 = n8766 ^ n8573 ;
  assign n8768 = x247 & ~x527 ;
  assign n8769 = n8768 ^ n8432 ;
  assign n8770 = ~n8767 & ~n8769 ;
  assign n8771 = ~n8585 & n8770 ;
  assign n8772 = x233 & ~n8768 ;
  assign n8773 = ~n8570 & n8772 ;
  assign n8774 = n8771 & n8773 ;
  assign n8775 = n8765 & n8774 ;
  assign n8776 = ~n8441 & ~n8766 ;
  assign n8777 = n8775 & n8776 ;
  assign n8778 = ~n8546 & ~n8567 ;
  assign n8779 = ~n8531 & ~n8543 ;
  assign n8780 = n8778 & n8779 ;
  assign n8781 = ~n8447 & ~n8561 ;
  assign n8782 = ~n8345 & n8564 ;
  assign n8783 = n8781 & n8782 ;
  assign n8784 = n8780 & n8783 ;
  assign n8785 = x249 & ~x482 ;
  assign n8786 = n8785 ^ n8297 ;
  assign n8787 = ~x233 & ~n8786 ;
  assign n8788 = ~n8537 & n8787 ;
  assign n8789 = ~n8444 & ~n8549 ;
  assign n8790 = n8788 & n8789 ;
  assign n8791 = n8784 & n8790 ;
  assign n8792 = ~n8519 & ~n8785 ;
  assign n8793 = n8791 & n8792 ;
  assign n8794 = ~n8777 & ~n8793 ;
  assign n8795 = ~x237 & n8794 ;
  assign n8796 = n8758 & ~n8795 ;
  assign n8797 = ~n8729 & ~n8796 ;
  assign n8798 = ~x806 & x990 ;
  assign n8803 = x600 & n8798 ;
  assign n8804 = n8803 ^ x594 ;
  assign n8805 = ~x332 & n8804 ;
  assign n8812 = ~x806 & n8170 ;
  assign n8813 = x605 & n8812 ;
  assign n8814 = n8813 ^ x605 ;
  assign n8806 = x605 ^ x595 ;
  assign n8815 = n8814 ^ n8806 ;
  assign n8816 = ~x332 & n8815 ;
  assign n8817 = n8168 & n8798 ;
  assign n8818 = x595 & x597 ;
  assign n8819 = n8817 & n8818 ;
  assign n8820 = n8819 ^ x596 ;
  assign n8821 = ~x332 & n8820 ;
  assign n8822 = n8817 ^ x597 ;
  assign n8823 = ~x332 & n8822 ;
  assign n8824 = x780 ^ x598 ;
  assign n8889 = n8824 ^ n2651 ;
  assign n8825 = ~x882 & n1209 ;
  assign n8826 = x947 & n8825 ;
  assign n8827 = n8826 ^ x598 ;
  assign n8890 = n8889 ^ n8827 ;
  assign n8830 = n8824 ^ x740 ;
  assign n8892 = n8890 ^ n8830 ;
  assign n8888 = n8827 ^ n8824 ;
  assign n8893 = n8892 ^ n8888 ;
  assign n8894 = n8893 ^ n8826 ;
  assign n8852 = ~x598 & ~n8827 ;
  assign n8831 = n8830 ^ n8827 ;
  assign n8853 = n8852 ^ n8831 ;
  assign n8832 = n8831 ^ n8824 ;
  assign n8838 = n8832 ^ n8826 ;
  assign n8842 = n8838 ^ n8827 ;
  assign n8854 = n8853 ^ n8842 ;
  assign n8855 = n8854 ^ n8826 ;
  assign n8883 = n8893 ^ n8827 ;
  assign n8857 = n8883 ^ n8826 ;
  assign n8858 = ~n8855 & n8857 ;
  assign n8880 = n8893 ^ x780 ;
  assign n8881 = n8880 ^ n8827 ;
  assign n8859 = n8893 ^ n8881 ;
  assign n8860 = n8894 ^ n8859 ;
  assign n8861 = n8893 ^ n8831 ;
  assign n8862 = n8894 ^ n8861 ;
  assign n8863 = ~n8860 & ~n8862 ;
  assign n8864 = n8858 & n8863 ;
  assign n8865 = n8864 ^ n8852 ;
  assign n8848 = n8881 ^ n8831 ;
  assign n8866 = n8865 ^ n8848 ;
  assign n8867 = n8866 ^ x740 ;
  assign n8887 = n8867 ^ x598 ;
  assign n8895 = n8894 ^ n8887 ;
  assign n8900 = x596 & n8819 ;
  assign n8901 = n8900 ^ x599 ;
  assign n8902 = ~x332 & n8901 ;
  assign n8903 = n8798 ^ x600 ;
  assign n8904 = ~x332 & n8903 ;
  assign n8905 = x989 ^ x601 ;
  assign n8906 = ~x806 & n8905 ;
  assign n8907 = n8906 ^ x601 ;
  assign n8908 = ~x332 & n8907 ;
  assign n8909 = n5775 ^ x602 ;
  assign n8910 = x230 & n8909 ;
  assign n8911 = n8910 ^ x602 ;
  assign n8925 = ~x871 & ~x872 ;
  assign n8912 = x1100 ^ x603 ;
  assign n8913 = x832 & ~x980 ;
  assign n8914 = x1060 & n8913 ;
  assign n8915 = x1038 & ~x1061 ;
  assign n8916 = n8914 & n8915 ;
  assign n8917 = ~x952 & n8916 ;
  assign n8918 = n8917 ^ n8916 ;
  assign n8919 = n8912 & n8918 ;
  assign n8920 = n8919 ^ x603 ;
  assign n8926 = n8925 ^ n8920 ;
  assign n8927 = x966 & ~n8926 ;
  assign n8928 = n8927 ^ n8920 ;
  assign n8931 = ~x299 & x983 ;
  assign n8932 = x907 & n8931 ;
  assign n8933 = x604 & n8932 ;
  assign n8929 = x779 ^ x604 ;
  assign n8934 = n8933 ^ n8929 ;
  assign n8937 = n8934 ^ x779 ;
  assign n8935 = x823 & n2653 ;
  assign n8936 = ~n8934 & n8935 ;
  assign n8938 = n8937 ^ n8936 ;
  assign n8939 = x806 ^ x605 ;
  assign n8940 = ~x332 & ~n8939 ;
  assign n8944 = x1104 ^ x837 ;
  assign n8941 = x837 ^ x606 ;
  assign n8945 = n8944 ^ n8941 ;
  assign n8946 = n8918 & n8945 ;
  assign n8947 = n8946 ^ n8941 ;
  assign n8948 = ~x966 & n8947 ;
  assign n8949 = n8948 ^ x837 ;
  assign n8950 = x1107 ^ x607 ;
  assign n8953 = n8918 & n8950 ;
  assign n8954 = n8953 ^ x607 ;
  assign n8955 = ~x966 & n8954 ;
  assign n8956 = x1116 ^ x608 ;
  assign n8959 = n8918 & n8956 ;
  assign n8960 = n8959 ^ x608 ;
  assign n8961 = ~x966 & n8960 ;
  assign n8962 = x1118 ^ x609 ;
  assign n8965 = n8918 & n8962 ;
  assign n8966 = n8965 ^ x609 ;
  assign n8967 = ~x966 & n8966 ;
  assign n8968 = x1113 ^ x610 ;
  assign n8971 = n8918 & n8968 ;
  assign n8972 = n8971 ^ x610 ;
  assign n8973 = ~x966 & n8972 ;
  assign n8974 = x1114 ^ x611 ;
  assign n8977 = n8918 & n8974 ;
  assign n8978 = n8977 ^ x611 ;
  assign n8979 = ~x966 & n8978 ;
  assign n8980 = x1111 ^ x612 ;
  assign n8983 = n8918 & n8980 ;
  assign n8984 = n8983 ^ x612 ;
  assign n8985 = ~x966 & n8984 ;
  assign n8986 = x1115 ^ x613 ;
  assign n8989 = n8918 & n8986 ;
  assign n8990 = n8989 ^ x613 ;
  assign n8991 = ~x966 & n8990 ;
  assign n8995 = x1102 ^ x871 ;
  assign n8992 = x871 ^ x614 ;
  assign n8996 = n8995 ^ n8992 ;
  assign n8997 = n8918 & n8996 ;
  assign n8998 = n8997 ^ n8992 ;
  assign n8999 = ~x966 & n8998 ;
  assign n9000 = n8999 ^ x871 ;
  assign n9001 = x907 & n8825 ;
  assign n9003 = n9001 ^ x797 ;
  assign n9002 = n9001 ^ x615 ;
  assign n9004 = n9003 ^ n9002 ;
  assign n9011 = n9004 ^ x779 ;
  assign n9043 = n9011 ^ n9002 ;
  assign n9008 = n9004 ^ n2654 ;
  assign n9042 = n9008 ^ n9002 ;
  assign n9044 = n9043 ^ n9042 ;
  assign n9024 = x615 & n9002 ;
  assign n9025 = n9042 ^ n9024 ;
  assign n9026 = n9025 ^ n9003 ;
  assign n9027 = n9026 ^ n9001 ;
  assign n9046 = n9042 ^ x779 ;
  assign n9029 = n9046 ^ n9001 ;
  assign n9030 = ~n9027 & n9029 ;
  assign n9058 = n9042 ^ n9011 ;
  assign n9059 = n9058 ^ n9003 ;
  assign n9060 = n9059 ^ n9001 ;
  assign n9051 = n9046 ^ n9011 ;
  assign n9032 = n9060 ^ n9051 ;
  assign n9033 = n9059 ^ n9042 ;
  assign n9034 = n9060 ^ n9033 ;
  assign n9035 = ~n9032 & ~n9034 ;
  assign n9036 = n9030 & n9035 ;
  assign n9037 = n9036 ^ n9024 ;
  assign n9038 = n9044 ^ n9037 ;
  assign n9063 = n9038 ^ x797 ;
  assign n9064 = n9063 ^ x615 ;
  assign n9065 = n9064 ^ n9060 ;
  assign n9069 = x1101 ^ x872 ;
  assign n9066 = x872 ^ x616 ;
  assign n9070 = n9069 ^ n9066 ;
  assign n9071 = n8918 & n9070 ;
  assign n9072 = n9071 ^ n9066 ;
  assign n9073 = ~x966 & n9072 ;
  assign n9074 = n9073 ^ x872 ;
  assign n9078 = x1105 ^ x850 ;
  assign n9075 = x850 ^ x617 ;
  assign n9079 = n9078 ^ n9075 ;
  assign n9080 = n8918 & n9079 ;
  assign n9081 = n9080 ^ n9075 ;
  assign n9082 = ~x966 & n9081 ;
  assign n9083 = n9082 ^ x850 ;
  assign n9084 = x1117 ^ x618 ;
  assign n9087 = n8918 & n9084 ;
  assign n9088 = n9087 ^ x618 ;
  assign n9089 = ~x966 & n9088 ;
  assign n9090 = x1122 ^ x619 ;
  assign n9093 = n8918 & n9090 ;
  assign n9094 = n9093 ^ x619 ;
  assign n9095 = ~x966 & n9094 ;
  assign n9096 = x1112 ^ x620 ;
  assign n9099 = n8918 & n9096 ;
  assign n9100 = n9099 ^ x620 ;
  assign n9101 = ~x966 & n9100 ;
  assign n9102 = x1108 ^ x621 ;
  assign n9105 = n8918 & n9102 ;
  assign n9106 = n9105 ^ x621 ;
  assign n9107 = ~x966 & n9106 ;
  assign n9108 = x1109 ^ x622 ;
  assign n9111 = n8918 & n9108 ;
  assign n9112 = n9111 ^ x622 ;
  assign n9113 = ~x966 & n9112 ;
  assign n9114 = x1106 ^ x623 ;
  assign n9117 = n8918 & n9114 ;
  assign n9118 = n9117 ^ x623 ;
  assign n9119 = ~x966 & n9118 ;
  assign n9122 = x947 & n8931 ;
  assign n9123 = x624 & n9122 ;
  assign n9120 = x780 ^ x624 ;
  assign n9124 = n9123 ^ n9120 ;
  assign n9127 = n9124 ^ x780 ;
  assign n9125 = x831 & n2650 ;
  assign n9126 = ~n9124 & n9125 ;
  assign n9128 = n9127 ^ n9126 ;
  assign n9129 = x1116 ^ x625 ;
  assign n9130 = x1066 & x1088 ;
  assign n9131 = ~x973 & ~x1054 ;
  assign n9132 = n9130 & n9131 ;
  assign n9133 = x832 & n9132 ;
  assign n9134 = x953 & n9133 ;
  assign n9135 = n9134 ^ n9133 ;
  assign n9138 = n9129 & n9135 ;
  assign n9139 = n9138 ^ x625 ;
  assign n9140 = ~x962 & n9139 ;
  assign n9141 = x1121 ^ x626 ;
  assign n9144 = n8918 & n9141 ;
  assign n9145 = n9144 ^ x626 ;
  assign n9146 = ~x966 & n9145 ;
  assign n9147 = x1117 ^ x627 ;
  assign n9150 = n9135 & n9147 ;
  assign n9151 = n9150 ^ x627 ;
  assign n9152 = ~x962 & n9151 ;
  assign n9153 = x1119 ^ x628 ;
  assign n9156 = n9135 & n9153 ;
  assign n9157 = n9156 ^ x628 ;
  assign n9158 = ~x962 & n9157 ;
  assign n9159 = x1119 ^ x629 ;
  assign n9162 = n8918 & n9159 ;
  assign n9163 = n9162 ^ x629 ;
  assign n9164 = ~x966 & n9163 ;
  assign n9165 = x1120 ^ x630 ;
  assign n9168 = n8918 & n9165 ;
  assign n9169 = n9168 ^ x630 ;
  assign n9170 = ~x966 & n9169 ;
  assign n9171 = x1113 ^ x631 ;
  assign n9174 = n9135 & ~n9171 ;
  assign n9175 = n9174 ^ x631 ;
  assign n9176 = ~x962 & ~n9175 ;
  assign n9177 = x1115 ^ x632 ;
  assign n9180 = n9135 & ~n9177 ;
  assign n9181 = n9180 ^ x632 ;
  assign n9182 = ~x962 & ~n9181 ;
  assign n9183 = x1110 ^ x633 ;
  assign n9186 = n8918 & n9183 ;
  assign n9187 = n9186 ^ x633 ;
  assign n9188 = ~x966 & n9187 ;
  assign n9189 = x1110 ^ x634 ;
  assign n9192 = n9135 & n9189 ;
  assign n9193 = n9192 ^ x634 ;
  assign n9194 = ~x962 & n9193 ;
  assign n9195 = x1112 ^ x635 ;
  assign n9198 = n9135 & ~n9195 ;
  assign n9199 = n9198 ^ x635 ;
  assign n9200 = ~x962 & ~n9199 ;
  assign n9201 = x1127 ^ x636 ;
  assign n9204 = n8918 & n9201 ;
  assign n9205 = n9204 ^ x636 ;
  assign n9206 = ~x966 & n9205 ;
  assign n9207 = x1105 ^ x637 ;
  assign n9210 = n9135 & n9207 ;
  assign n9211 = n9210 ^ x637 ;
  assign n9212 = ~x962 & n9211 ;
  assign n9213 = x1107 ^ x638 ;
  assign n9216 = n9135 & n9213 ;
  assign n9217 = n9216 ^ x638 ;
  assign n9218 = ~x962 & n9217 ;
  assign n9219 = x1109 ^ x639 ;
  assign n9222 = n9135 & n9219 ;
  assign n9223 = n9222 ^ x639 ;
  assign n9224 = ~x962 & n9223 ;
  assign n9225 = x1128 ^ x640 ;
  assign n9228 = n8918 & n9225 ;
  assign n9229 = n9228 ^ x640 ;
  assign n9230 = ~x966 & n9229 ;
  assign n9231 = x1121 ^ x641 ;
  assign n9234 = n9135 & n9231 ;
  assign n9235 = n9234 ^ x641 ;
  assign n9236 = ~x962 & n9235 ;
  assign n9237 = x1103 ^ x642 ;
  assign n9240 = n8918 & n9237 ;
  assign n9241 = n9240 ^ x642 ;
  assign n9242 = ~x966 & n9241 ;
  assign n9243 = x1104 ^ x643 ;
  assign n9246 = n9135 & n9243 ;
  assign n9247 = n9246 ^ x643 ;
  assign n9248 = ~x962 & n9247 ;
  assign n9249 = x1123 ^ x644 ;
  assign n9252 = n8918 & n9249 ;
  assign n9253 = n9252 ^ x644 ;
  assign n9254 = ~x966 & n9253 ;
  assign n9255 = x1125 ^ x645 ;
  assign n9258 = n8918 & n9255 ;
  assign n9259 = n9258 ^ x645 ;
  assign n9260 = ~x966 & n9259 ;
  assign n9261 = x1114 ^ x646 ;
  assign n9264 = n9135 & ~n9261 ;
  assign n9265 = n9264 ^ x646 ;
  assign n9266 = ~x962 & ~n9265 ;
  assign n9267 = x1120 ^ x647 ;
  assign n9270 = n9135 & n9267 ;
  assign n9271 = n9270 ^ x647 ;
  assign n9272 = ~x962 & n9271 ;
  assign n9273 = x1122 ^ x648 ;
  assign n9276 = n9135 & n9273 ;
  assign n9277 = n9276 ^ x648 ;
  assign n9278 = ~x962 & n9277 ;
  assign n9279 = x1126 ^ x649 ;
  assign n9282 = n9135 & ~n9279 ;
  assign n9283 = n9282 ^ x649 ;
  assign n9284 = ~x962 & ~n9283 ;
  assign n9285 = x1127 ^ x650 ;
  assign n9288 = n9135 & ~n9285 ;
  assign n9289 = n9288 ^ x650 ;
  assign n9290 = ~x962 & ~n9289 ;
  assign n9291 = x1130 ^ x651 ;
  assign n9294 = n8918 & n9291 ;
  assign n9295 = n9294 ^ x651 ;
  assign n9296 = ~x966 & n9295 ;
  assign n9297 = x1131 ^ x652 ;
  assign n9300 = n8918 & n9297 ;
  assign n9301 = n9300 ^ x652 ;
  assign n9302 = ~x966 & n9301 ;
  assign n9303 = x1129 ^ x653 ;
  assign n9306 = n8918 & n9303 ;
  assign n9307 = n9306 ^ x653 ;
  assign n9308 = ~x966 & n9307 ;
  assign n9309 = x1130 ^ x654 ;
  assign n9312 = n9135 & ~n9309 ;
  assign n9313 = n9312 ^ x654 ;
  assign n9314 = ~x962 & ~n9313 ;
  assign n9315 = x1124 ^ x655 ;
  assign n9318 = n9135 & ~n9315 ;
  assign n9319 = n9318 ^ x655 ;
  assign n9320 = ~x962 & ~n9319 ;
  assign n9321 = x1126 ^ x656 ;
  assign n9324 = n8918 & n9321 ;
  assign n9325 = n9324 ^ x656 ;
  assign n9326 = ~x966 & n9325 ;
  assign n9327 = x1131 ^ x657 ;
  assign n9330 = n9135 & ~n9327 ;
  assign n9331 = n9330 ^ x657 ;
  assign n9332 = ~x962 & ~n9331 ;
  assign n9333 = x1124 ^ x658 ;
  assign n9336 = n8918 & n9333 ;
  assign n9337 = n9336 ^ x658 ;
  assign n9338 = ~x966 & n9337 ;
  assign n9339 = x266 & x992 ;
  assign n9340 = ~x280 & n9339 ;
  assign n9341 = ~x269 & n9340 ;
  assign n9342 = ~x281 & ~x282 ;
  assign n9343 = n9341 & n9342 ;
  assign n9344 = ~x270 & ~x277 ;
  assign n9345 = ~x264 & n9344 ;
  assign n9346 = n9343 & n9345 ;
  assign n9347 = ~x265 & n9346 ;
  assign n9348 = n9347 ^ x274 ;
  assign n9349 = x1118 ^ x660 ;
  assign n9352 = n9135 & n9349 ;
  assign n9353 = n9352 ^ x660 ;
  assign n9354 = ~x962 & n9353 ;
  assign n9355 = x1101 ^ x661 ;
  assign n9358 = n9135 & n9355 ;
  assign n9359 = n9358 ^ x661 ;
  assign n9360 = ~x962 & n9359 ;
  assign n9361 = x1102 ^ x662 ;
  assign n9364 = n9135 & n9361 ;
  assign n9365 = n9364 ^ x662 ;
  assign n9366 = ~x962 & n9365 ;
  assign n9471 = ~x1137 & ~x1138 ;
  assign n9472 = ~n2991 & n9471 ;
  assign n9482 = x815 ^ x633 ;
  assign n9483 = ~x1136 & n9482 ;
  assign n9484 = n9483 ^ x633 ;
  assign n9486 = n9484 ^ x766 ;
  assign n9485 = n9484 ^ x855 ;
  assign n9487 = n9486 ^ n9485 ;
  assign n9490 = x1136 & n9487 ;
  assign n9491 = n9490 ^ n9485 ;
  assign n9492 = x1134 & n9491 ;
  assign n9493 = n9492 ^ n9484 ;
  assign n9474 = x1135 ^ x1134 ;
  assign n9475 = x700 ^ x634 ;
  assign n9476 = n9475 ^ x784 ;
  assign n9479 = x1136 & n9476 ;
  assign n9480 = n9479 ^ x784 ;
  assign n9481 = n9474 & n9480 ;
  assign n9494 = n9493 ^ n9481 ;
  assign n9473 = x700 & x1136 ;
  assign n9495 = n9494 ^ n9473 ;
  assign n9496 = x1135 & n9495 ;
  assign n9497 = n9496 ^ n9493 ;
  assign n9498 = n9472 & n9497 ;
  assign n9367 = ~x223 & ~x224 ;
  assign n9369 = ~x588 & ~n3076 ;
  assign n9368 = n3076 ^ x588 ;
  assign n9370 = n9369 ^ n9368 ;
  assign n9371 = n9370 ^ n8660 ;
  assign n9372 = n9371 ^ x334 ;
  assign n9373 = n9372 ^ x365 ;
  assign n9374 = n9373 ^ n9371 ;
  assign n9375 = x592 & n9374 ;
  assign n9376 = n9375 ^ n9372 ;
  assign n9400 = n9376 ^ x464 ;
  assign n9401 = n9400 ^ n9370 ;
  assign n9378 = n9370 ^ x464 ;
  assign n9381 = n9378 ^ n9371 ;
  assign n9382 = n9381 ^ n4593 ;
  assign n9383 = n9382 ^ n9378 ;
  assign n9448 = n9401 ^ n9383 ;
  assign n9449 = n9448 ^ n9371 ;
  assign n9437 = n9449 ^ n9383 ;
  assign n9438 = n9437 ^ x464 ;
  assign n9416 = ~x464 & ~n9378 ;
  assign n9417 = n9438 ^ n9416 ;
  assign n9396 = n9448 ^ n9370 ;
  assign n9406 = n9396 ^ n9378 ;
  assign n9418 = n9417 ^ n9406 ;
  assign n9419 = n9418 ^ n9370 ;
  assign n9393 = n9376 ^ n4593 ;
  assign n9421 = n9393 ^ n9370 ;
  assign n9422 = ~n9419 & n9421 ;
  assign n9450 = n9449 ^ n9370 ;
  assign n9423 = n9449 ^ n9376 ;
  assign n9424 = n9450 ^ n9423 ;
  assign n9425 = n9449 ^ n9438 ;
  assign n9426 = n9450 ^ n9425 ;
  assign n9427 = ~n9424 & n9426 ;
  assign n9428 = n9422 & n9427 ;
  assign n9429 = n9428 ^ n9416 ;
  assign n9430 = n9429 ^ n8660 ;
  assign n9408 = n9449 ^ n9406 ;
  assign n9410 = n9450 ^ n9408 ;
  assign n9431 = n9430 ^ n9410 ;
  assign n9454 = n9431 ^ x464 ;
  assign n9455 = n9454 ^ n9450 ;
  assign n9456 = n9367 & n9455 ;
  assign n9457 = n2991 & ~n9367 ;
  assign n9458 = x1065 ^ x257 ;
  assign n9461 = x199 & n9458 ;
  assign n9462 = n9461 ^ x257 ;
  assign n9463 = n9457 & ~n9462 ;
  assign n9464 = n9463 ^ n2991 ;
  assign n9465 = n9456 & n9464 ;
  assign n9469 = n9465 ^ n9464 ;
  assign n9466 = n3109 & n9369 ;
  assign n9467 = x323 & n9466 ;
  assign n9468 = n9465 & n9467 ;
  assign n9470 = n9469 ^ n9468 ;
  assign n9500 = n9498 ^ n9470 ;
  assign n9606 = x811 ^ x614 ;
  assign n9607 = ~x1136 & n9606 ;
  assign n9608 = n9607 ^ x614 ;
  assign n9610 = n9608 ^ x772 ;
  assign n9609 = n9608 ^ x872 ;
  assign n9611 = n9610 ^ n9609 ;
  assign n9614 = x1136 & n9611 ;
  assign n9615 = n9614 ^ n9609 ;
  assign n9616 = x1134 & n9615 ;
  assign n9617 = n9616 ^ n9608 ;
  assign n9599 = x727 ^ x662 ;
  assign n9600 = n9599 ^ x785 ;
  assign n9603 = x1136 & n9600 ;
  assign n9604 = n9603 ^ x785 ;
  assign n9605 = n9474 & n9604 ;
  assign n9618 = n9617 ^ n9605 ;
  assign n9598 = x727 & x1136 ;
  assign n9619 = n9618 ^ n9598 ;
  assign n9620 = x1135 & n9619 ;
  assign n9621 = n9620 ^ n9617 ;
  assign n9622 = n9472 & n9621 ;
  assign n9501 = x355 & n9466 ;
  assign n9504 = x199 & n7626 ;
  assign n9505 = n9504 ^ x292 ;
  assign n9506 = n9457 & ~n9505 ;
  assign n9507 = n9506 ^ n2991 ;
  assign n9508 = n9371 ^ x380 ;
  assign n9509 = n9508 ^ x404 ;
  assign n9510 = n9509 ^ n9371 ;
  assign n9511 = ~x592 & n9510 ;
  assign n9512 = n9511 ^ n9508 ;
  assign n9536 = n9512 ^ x429 ;
  assign n9537 = n9536 ^ n9370 ;
  assign n9514 = n9370 ^ x429 ;
  assign n9517 = n9514 ^ n9371 ;
  assign n9518 = n9517 ^ n4593 ;
  assign n9519 = n9518 ^ n9514 ;
  assign n9584 = n9537 ^ n9519 ;
  assign n9585 = n9584 ^ n9371 ;
  assign n9573 = n9585 ^ n9519 ;
  assign n9574 = n9573 ^ x429 ;
  assign n9552 = ~x429 & ~n9514 ;
  assign n9553 = n9574 ^ n9552 ;
  assign n9532 = n9584 ^ n9370 ;
  assign n9542 = n9532 ^ n9514 ;
  assign n9554 = n9553 ^ n9542 ;
  assign n9555 = n9554 ^ n9370 ;
  assign n9529 = n9512 ^ n4593 ;
  assign n9557 = n9529 ^ n9370 ;
  assign n9558 = ~n9555 & n9557 ;
  assign n9586 = n9585 ^ n9370 ;
  assign n9559 = n9585 ^ n9512 ;
  assign n9560 = n9586 ^ n9559 ;
  assign n9561 = n9585 ^ n9574 ;
  assign n9562 = n9586 ^ n9561 ;
  assign n9563 = ~n9560 & n9562 ;
  assign n9564 = n9558 & n9563 ;
  assign n9565 = n9564 ^ n9552 ;
  assign n9566 = n9565 ^ n8660 ;
  assign n9544 = n9585 ^ n9542 ;
  assign n9546 = n9586 ^ n9544 ;
  assign n9567 = n9566 ^ n9546 ;
  assign n9590 = n9567 ^ x429 ;
  assign n9591 = n9590 ^ n9586 ;
  assign n9592 = n9367 & n9591 ;
  assign n9593 = n9507 & n9592 ;
  assign n9596 = n9501 & n9593 ;
  assign n9594 = n9593 ^ n9507 ;
  assign n9597 = n9596 ^ n9594 ;
  assign n9624 = n9622 ^ n9597 ;
  assign n9625 = x1108 ^ x665 ;
  assign n9628 = n9135 & n9625 ;
  assign n9629 = n9628 ^ x665 ;
  assign n9630 = ~x962 & n9629 ;
  assign n9736 = x799 ^ x607 ;
  assign n9737 = ~x1136 & ~n9736 ;
  assign n9738 = n9737 ^ x607 ;
  assign n9740 = n9738 ^ x764 ;
  assign n9739 = n9738 ^ x873 ;
  assign n9741 = n9740 ^ n9739 ;
  assign n9744 = x1136 & n9741 ;
  assign n9745 = n9744 ^ n9739 ;
  assign n9746 = x1134 & n9745 ;
  assign n9747 = n9746 ^ n9738 ;
  assign n9729 = x691 ^ x638 ;
  assign n9730 = n9729 ^ x790 ;
  assign n9733 = x1136 & n9730 ;
  assign n9734 = n9733 ^ x790 ;
  assign n9735 = n9474 & n9734 ;
  assign n9748 = n9747 ^ n9735 ;
  assign n9728 = x691 & x1136 ;
  assign n9749 = n9748 ^ n9728 ;
  assign n9750 = x1135 & n9749 ;
  assign n9751 = n9750 ^ n9747 ;
  assign n9752 = n9472 & n9751 ;
  assign n9631 = x441 & n9466 ;
  assign n9634 = x199 & n7641 ;
  assign n9635 = n9634 ^ x297 ;
  assign n9636 = n9457 & ~n9635 ;
  assign n9637 = n9636 ^ n2991 ;
  assign n9638 = n9371 ^ x337 ;
  assign n9639 = n9638 ^ x456 ;
  assign n9640 = n9639 ^ n9371 ;
  assign n9641 = ~x592 & n9640 ;
  assign n9642 = n9641 ^ n9638 ;
  assign n9666 = n9642 ^ x443 ;
  assign n9667 = n9666 ^ n9370 ;
  assign n9644 = n9370 ^ x443 ;
  assign n9647 = n9644 ^ n9371 ;
  assign n9648 = n9647 ^ n4593 ;
  assign n9649 = n9648 ^ n9644 ;
  assign n9714 = n9667 ^ n9649 ;
  assign n9715 = n9714 ^ n9371 ;
  assign n9703 = n9715 ^ n9649 ;
  assign n9704 = n9703 ^ x443 ;
  assign n9682 = ~x443 & ~n9644 ;
  assign n9683 = n9704 ^ n9682 ;
  assign n9662 = n9714 ^ n9370 ;
  assign n9672 = n9662 ^ n9644 ;
  assign n9684 = n9683 ^ n9672 ;
  assign n9685 = n9684 ^ n9370 ;
  assign n9659 = n9642 ^ n4593 ;
  assign n9687 = n9659 ^ n9370 ;
  assign n9688 = ~n9685 & n9687 ;
  assign n9716 = n9715 ^ n9370 ;
  assign n9689 = n9715 ^ n9642 ;
  assign n9690 = n9716 ^ n9689 ;
  assign n9691 = n9715 ^ n9704 ;
  assign n9692 = n9716 ^ n9691 ;
  assign n9693 = ~n9690 & n9692 ;
  assign n9694 = n9688 & n9693 ;
  assign n9695 = n9694 ^ n9682 ;
  assign n9696 = n9695 ^ n8660 ;
  assign n9674 = n9715 ^ n9672 ;
  assign n9676 = n9716 ^ n9674 ;
  assign n9697 = n9696 ^ n9676 ;
  assign n9720 = n9697 ^ x443 ;
  assign n9721 = n9720 ^ n9716 ;
  assign n9722 = n9367 & n9721 ;
  assign n9723 = n9637 & n9722 ;
  assign n9726 = n9631 & n9723 ;
  assign n9724 = n9723 ^ n9637 ;
  assign n9727 = n9726 ^ n9724 ;
  assign n9754 = n9752 ^ n9727 ;
  assign n9858 = x809 ^ x642 ;
  assign n9859 = ~x1136 & ~n9858 ;
  assign n9860 = n9859 ^ x642 ;
  assign n9862 = n9860 ^ x763 ;
  assign n9861 = n9860 ^ x871 ;
  assign n9863 = n9862 ^ n9861 ;
  assign n9866 = x1136 & n9863 ;
  assign n9867 = n9866 ^ n9861 ;
  assign n9868 = x1134 & n9867 ;
  assign n9869 = n9868 ^ n9860 ;
  assign n9851 = x699 ^ x681 ;
  assign n9852 = n9851 ^ x792 ;
  assign n9855 = x1136 & n9852 ;
  assign n9856 = n9855 ^ x792 ;
  assign n9857 = n9474 & n9856 ;
  assign n9870 = n9869 ^ n9857 ;
  assign n9850 = x699 & x1136 ;
  assign n9871 = n9870 ^ n9850 ;
  assign n9872 = x1135 & n9871 ;
  assign n9873 = n9872 ^ n9869 ;
  assign n9874 = n9471 & n9873 ;
  assign n9756 = n9371 ^ x319 ;
  assign n9757 = n9756 ^ x338 ;
  assign n9758 = n9757 ^ n9371 ;
  assign n9759 = x592 & n9758 ;
  assign n9760 = n9759 ^ n9756 ;
  assign n9784 = n9760 ^ x444 ;
  assign n9785 = n9784 ^ n9370 ;
  assign n9762 = n9370 ^ x444 ;
  assign n9765 = n9762 ^ n9371 ;
  assign n9766 = n9765 ^ n4593 ;
  assign n9767 = n9766 ^ n9762 ;
  assign n9832 = n9785 ^ n9767 ;
  assign n9833 = n9832 ^ n9371 ;
  assign n9821 = n9833 ^ n9767 ;
  assign n9822 = n9821 ^ x444 ;
  assign n9800 = ~x444 & ~n9762 ;
  assign n9801 = n9822 ^ n9800 ;
  assign n9780 = n9832 ^ n9370 ;
  assign n9790 = n9780 ^ n9762 ;
  assign n9802 = n9801 ^ n9790 ;
  assign n9803 = n9802 ^ n9370 ;
  assign n9777 = n9760 ^ n4593 ;
  assign n9805 = n9777 ^ n9370 ;
  assign n9806 = ~n9803 & n9805 ;
  assign n9834 = n9833 ^ n9370 ;
  assign n9807 = n9833 ^ n9760 ;
  assign n9808 = n9834 ^ n9807 ;
  assign n9809 = n9833 ^ n9822 ;
  assign n9810 = n9834 ^ n9809 ;
  assign n9811 = ~n9808 & n9810 ;
  assign n9812 = n9806 & n9811 ;
  assign n9813 = n9812 ^ n9800 ;
  assign n9814 = n9813 ^ n8660 ;
  assign n9792 = n9833 ^ n9790 ;
  assign n9794 = n9834 ^ n9792 ;
  assign n9815 = n9814 ^ n9794 ;
  assign n9838 = n9815 ^ x444 ;
  assign n9839 = n9838 ^ n9834 ;
  assign n9755 = x458 & n9466 ;
  assign n9841 = n9839 ^ n9755 ;
  assign n9875 = n9874 ^ n9841 ;
  assign n9847 = x199 & n7632 ;
  assign n9843 = n9841 ^ x294 ;
  assign n9848 = n9847 ^ n9843 ;
  assign n9849 = ~n9367 & ~n9848 ;
  assign n9876 = n9875 ^ n9849 ;
  assign n9877 = n2991 & ~n9876 ;
  assign n9878 = n9877 ^ n9874 ;
  assign n9982 = x981 ^ x603 ;
  assign n9983 = ~x1136 & n9982 ;
  assign n9984 = n9983 ^ x603 ;
  assign n9986 = n9984 ^ x759 ;
  assign n9985 = n9984 ^ x837 ;
  assign n9987 = n9986 ^ n9985 ;
  assign n9990 = x1136 & n9987 ;
  assign n9991 = n9990 ^ n9985 ;
  assign n9992 = x1134 & n9991 ;
  assign n9993 = n9992 ^ n9984 ;
  assign n9975 = x696 ^ x680 ;
  assign n9976 = n9975 ^ x778 ;
  assign n9979 = x1136 & n9976 ;
  assign n9980 = n9979 ^ x778 ;
  assign n9981 = n9474 & n9980 ;
  assign n9994 = n9993 ^ n9981 ;
  assign n9974 = x696 & x1136 ;
  assign n9995 = n9994 ^ n9974 ;
  assign n9996 = x1135 & n9995 ;
  assign n9997 = n9996 ^ n9993 ;
  assign n9998 = n9471 & n9997 ;
  assign n9880 = n9371 ^ x363 ;
  assign n9881 = n9880 ^ x390 ;
  assign n9882 = n9881 ^ n9371 ;
  assign n9883 = ~x592 & n9882 ;
  assign n9884 = n9883 ^ n9880 ;
  assign n9908 = n9884 ^ x414 ;
  assign n9909 = n9908 ^ n9370 ;
  assign n9886 = n9370 ^ x414 ;
  assign n9889 = n9886 ^ n9371 ;
  assign n9890 = n9889 ^ n4593 ;
  assign n9891 = n9890 ^ n9886 ;
  assign n9956 = n9909 ^ n9891 ;
  assign n9957 = n9956 ^ n9371 ;
  assign n9945 = n9957 ^ n9891 ;
  assign n9946 = n9945 ^ x414 ;
  assign n9924 = ~x414 & ~n9886 ;
  assign n9925 = n9946 ^ n9924 ;
  assign n9904 = n9956 ^ n9370 ;
  assign n9914 = n9904 ^ n9886 ;
  assign n9926 = n9925 ^ n9914 ;
  assign n9927 = n9926 ^ n9370 ;
  assign n9901 = n9884 ^ n4593 ;
  assign n9929 = n9901 ^ n9370 ;
  assign n9930 = ~n9927 & n9929 ;
  assign n9958 = n9957 ^ n9370 ;
  assign n9931 = n9957 ^ n9884 ;
  assign n9932 = n9958 ^ n9931 ;
  assign n9933 = n9957 ^ n9946 ;
  assign n9934 = n9958 ^ n9933 ;
  assign n9935 = ~n9932 & n9934 ;
  assign n9936 = n9930 & n9935 ;
  assign n9937 = n9936 ^ n9924 ;
  assign n9938 = n9937 ^ n8660 ;
  assign n9916 = n9957 ^ n9914 ;
  assign n9918 = n9958 ^ n9916 ;
  assign n9939 = n9938 ^ n9918 ;
  assign n9962 = n9939 ^ x414 ;
  assign n9963 = n9962 ^ n9958 ;
  assign n9879 = x342 & n9466 ;
  assign n9965 = n9963 ^ n9879 ;
  assign n9999 = n9998 ^ n9965 ;
  assign n9971 = x199 & n7623 ;
  assign n9967 = n9965 ^ x291 ;
  assign n9972 = n9971 ^ n9967 ;
  assign n9973 = ~n9367 & ~n9972 ;
  assign n10000 = n9999 ^ n9973 ;
  assign n10001 = n2991 & ~n10000 ;
  assign n10002 = n10001 ^ n9998 ;
  assign n10003 = x1125 ^ x669 ;
  assign n10006 = n9135 & ~n10003 ;
  assign n10007 = n10006 ^ x669 ;
  assign n10008 = ~x962 & ~n10007 ;
  assign n5907 = x745 ^ x723 ;
  assign n10009 = ~x1135 & n5907 ;
  assign n10010 = n10009 ^ x723 ;
  assign n10012 = n10010 ^ x612 ;
  assign n10011 = n10010 ^ x695 ;
  assign n10013 = n10012 ^ n10011 ;
  assign n10016 = ~x1135 & ~n10013 ;
  assign n10017 = n10016 ^ n10011 ;
  assign n10018 = ~x1134 & n10017 ;
  assign n10019 = n10018 ^ n10010 ;
  assign n10020 = x1136 & n9472 ;
  assign n10021 = ~n10019 & n10020 ;
  assign n10022 = n10021 ^ n9472 ;
  assign n10023 = ~x1135 & ~x1136 ;
  assign n10024 = x1134 & n10023 ;
  assign n10025 = x852 & n10024 ;
  assign n10026 = n10022 & n10025 ;
  assign n10028 = n10026 ^ n10021 ;
  assign n10029 = x1062 ^ x258 ;
  assign n10032 = x199 & n10029 ;
  assign n10033 = n10032 ^ x258 ;
  assign n10034 = n9457 & ~n10033 ;
  assign n10035 = n10034 ^ n2991 ;
  assign n10036 = x391 & ~x590 ;
  assign n10037 = ~x592 & n10036 ;
  assign n10038 = n10037 ^ x364 ;
  assign n10041 = n10037 ^ x590 ;
  assign n10042 = ~x591 & ~n10041 ;
  assign n10043 = n10038 & n10042 ;
  assign n10044 = n10043 ^ n10038 ;
  assign n10045 = n10044 ^ x364 ;
  assign n10046 = n9369 & ~n10045 ;
  assign n10054 = x343 & n10046 ;
  assign n10055 = n3109 & n10054 ;
  assign n10056 = n10055 ^ n3109 ;
  assign n10047 = n10046 ^ n9369 ;
  assign n10048 = n10047 ^ n3109 ;
  assign n10057 = n10056 ^ n10048 ;
  assign n10058 = n9367 & ~n10057 ;
  assign n10059 = n10035 & n10058 ;
  assign n10067 = x415 & n10059 ;
  assign n10068 = ~n9370 & n10067 ;
  assign n10069 = n10068 ^ n9370 ;
  assign n10060 = n10059 ^ n10035 ;
  assign n10061 = n10060 ^ n9370 ;
  assign n10070 = n10069 ^ n10061 ;
  assign n10071 = ~n10028 & ~n10070 ;
  assign n10072 = n9371 ^ x333 ;
  assign n10073 = n10072 ^ x447 ;
  assign n10074 = n10073 ^ n9371 ;
  assign n10075 = x592 & n10074 ;
  assign n10076 = n10075 ^ n10072 ;
  assign n10100 = n10076 ^ x453 ;
  assign n10101 = n10100 ^ n9370 ;
  assign n10078 = n9370 ^ x453 ;
  assign n10081 = n10078 ^ n9371 ;
  assign n10082 = n10081 ^ n4593 ;
  assign n10083 = n10082 ^ n10078 ;
  assign n10148 = n10101 ^ n10083 ;
  assign n10149 = n10148 ^ n9371 ;
  assign n10137 = n10149 ^ n10083 ;
  assign n10138 = n10137 ^ x453 ;
  assign n10116 = ~x453 & ~n10078 ;
  assign n10117 = n10138 ^ n10116 ;
  assign n10096 = n10148 ^ n9370 ;
  assign n10106 = n10096 ^ n10078 ;
  assign n10118 = n10117 ^ n10106 ;
  assign n10119 = n10118 ^ n9370 ;
  assign n10093 = n10076 ^ n4593 ;
  assign n10121 = n10093 ^ n9370 ;
  assign n10122 = ~n10119 & n10121 ;
  assign n10150 = n10149 ^ n9370 ;
  assign n10123 = n10149 ^ n10076 ;
  assign n10124 = n10150 ^ n10123 ;
  assign n10125 = n10149 ^ n10138 ;
  assign n10126 = n10150 ^ n10125 ;
  assign n10127 = ~n10124 & n10126 ;
  assign n10128 = n10122 & n10127 ;
  assign n10129 = n10128 ^ n10116 ;
  assign n10130 = n10129 ^ n8660 ;
  assign n10108 = n10149 ^ n10106 ;
  assign n10110 = n10150 ^ n10108 ;
  assign n10131 = n10130 ^ n10110 ;
  assign n10154 = n10131 ^ x453 ;
  assign n10155 = n10154 ^ n10150 ;
  assign n10156 = n9367 & n10155 ;
  assign n10157 = x327 & n9466 ;
  assign n10158 = n10156 & ~n10157 ;
  assign n10159 = x1040 ^ x261 ;
  assign n10162 = x199 & n10159 ;
  assign n10163 = n10162 ^ x261 ;
  assign n10164 = n9457 & ~n10163 ;
  assign n10165 = n10164 ^ n2991 ;
  assign n10166 = ~n10158 & n10165 ;
  assign n5966 = x741 ^ x724 ;
  assign n10167 = ~x1135 & n5966 ;
  assign n10168 = n10167 ^ x724 ;
  assign n10170 = n10168 ^ x611 ;
  assign n10169 = n10168 ^ x646 ;
  assign n10171 = n10170 ^ n10169 ;
  assign n10174 = ~x1135 & ~n10171 ;
  assign n10175 = n10174 ^ n10169 ;
  assign n10176 = ~x1134 & n10175 ;
  assign n10177 = n10176 ^ n10168 ;
  assign n10178 = n10020 & ~n10177 ;
  assign n10179 = n10178 ^ n9472 ;
  assign n10181 = x865 & n10024 ;
  assign n10182 = n10179 & n10181 ;
  assign n10183 = n10182 ^ n10178 ;
  assign n10184 = ~n10166 & ~n10183 ;
  assign n10288 = x808 ^ x616 ;
  assign n10289 = ~x1136 & n10288 ;
  assign n10290 = n10289 ^ x616 ;
  assign n10292 = n10290 ^ x758 ;
  assign n10291 = n10290 ^ x850 ;
  assign n10293 = n10292 ^ n10291 ;
  assign n10296 = x1136 & n10293 ;
  assign n10297 = n10296 ^ n10291 ;
  assign n10298 = x1134 & n10297 ;
  assign n10299 = n10298 ^ n10290 ;
  assign n10281 = x736 ^ x661 ;
  assign n10282 = n10281 ^ x781 ;
  assign n10285 = x1136 & n10282 ;
  assign n10286 = n10285 ^ x781 ;
  assign n10287 = n9474 & n10286 ;
  assign n10300 = n10299 ^ n10287 ;
  assign n10280 = x736 & x1136 ;
  assign n10301 = n10300 ^ n10280 ;
  assign n10302 = x1135 & n10301 ;
  assign n10303 = n10302 ^ n10299 ;
  assign n10304 = n9471 & n10303 ;
  assign n10186 = n9371 ^ x372 ;
  assign n10187 = n10186 ^ x397 ;
  assign n10188 = n10187 ^ n9371 ;
  assign n10189 = ~x592 & n10188 ;
  assign n10190 = n10189 ^ n10186 ;
  assign n10214 = n10190 ^ x422 ;
  assign n10215 = n10214 ^ n9370 ;
  assign n10192 = n9370 ^ x422 ;
  assign n10195 = n10192 ^ n9371 ;
  assign n10196 = n10195 ^ n4593 ;
  assign n10197 = n10196 ^ n10192 ;
  assign n10262 = n10215 ^ n10197 ;
  assign n10263 = n10262 ^ n9371 ;
  assign n10251 = n10263 ^ n10197 ;
  assign n10252 = n10251 ^ x422 ;
  assign n10230 = ~x422 & ~n10192 ;
  assign n10231 = n10252 ^ n10230 ;
  assign n10210 = n10262 ^ n9370 ;
  assign n10220 = n10210 ^ n10192 ;
  assign n10232 = n10231 ^ n10220 ;
  assign n10233 = n10232 ^ n9370 ;
  assign n10207 = n10190 ^ n4593 ;
  assign n10235 = n10207 ^ n9370 ;
  assign n10236 = ~n10233 & n10235 ;
  assign n10264 = n10263 ^ n9370 ;
  assign n10237 = n10263 ^ n10190 ;
  assign n10238 = n10264 ^ n10237 ;
  assign n10239 = n10263 ^ n10252 ;
  assign n10240 = n10264 ^ n10239 ;
  assign n10241 = ~n10238 & n10240 ;
  assign n10242 = n10236 & n10241 ;
  assign n10243 = n10242 ^ n10230 ;
  assign n10244 = n10243 ^ n8660 ;
  assign n10222 = n10263 ^ n10220 ;
  assign n10224 = n10264 ^ n10222 ;
  assign n10245 = n10244 ^ n10224 ;
  assign n10268 = n10245 ^ x422 ;
  assign n10269 = n10268 ^ n10264 ;
  assign n10185 = x320 & n9466 ;
  assign n10271 = n10269 ^ n10185 ;
  assign n10305 = n10304 ^ n10271 ;
  assign n10277 = x199 & n7620 ;
  assign n10273 = n10271 ^ x290 ;
  assign n10278 = n10277 ^ n10273 ;
  assign n10279 = ~n9367 & ~n10278 ;
  assign n10306 = n10305 ^ n10279 ;
  assign n10307 = n2991 & ~n10306 ;
  assign n10308 = n10307 ^ n10304 ;
  assign n10414 = x866 ^ x749 ;
  assign n10415 = ~x1136 & n10414 ;
  assign n10416 = n10415 ^ x749 ;
  assign n10418 = n10416 ^ x617 ;
  assign n10417 = n10416 ^ x814 ;
  assign n10419 = n10418 ^ n10417 ;
  assign n10422 = x1136 & ~n10419 ;
  assign n10423 = n10422 ^ n10417 ;
  assign n10424 = ~x1134 & ~n10423 ;
  assign n10425 = n10424 ^ n10416 ;
  assign n10407 = x706 ^ x637 ;
  assign n10408 = n10407 ^ x788 ;
  assign n10411 = x1136 & n10408 ;
  assign n10412 = n10411 ^ x788 ;
  assign n10413 = n9474 & n10412 ;
  assign n10426 = n10425 ^ n10413 ;
  assign n10406 = x706 & x1136 ;
  assign n10427 = n10426 ^ n10406 ;
  assign n10428 = x1135 & n10427 ;
  assign n10429 = n10428 ^ n10425 ;
  assign n10430 = n9472 & n10429 ;
  assign n10309 = x452 & n9466 ;
  assign n10312 = x199 & n7635 ;
  assign n10313 = n10312 ^ x295 ;
  assign n10314 = n9457 & ~n10313 ;
  assign n10315 = n10314 ^ n2991 ;
  assign n10316 = n9371 ^ x387 ;
  assign n10317 = n10316 ^ x411 ;
  assign n10318 = n10317 ^ n9371 ;
  assign n10319 = ~x592 & n10318 ;
  assign n10320 = n10319 ^ n10316 ;
  assign n10344 = n10320 ^ x435 ;
  assign n10345 = n10344 ^ n9370 ;
  assign n10322 = n9370 ^ x435 ;
  assign n10325 = n10322 ^ n9371 ;
  assign n10326 = n10325 ^ n4593 ;
  assign n10327 = n10326 ^ n10322 ;
  assign n10392 = n10345 ^ n10327 ;
  assign n10393 = n10392 ^ n9371 ;
  assign n10381 = n10393 ^ n10327 ;
  assign n10382 = n10381 ^ x435 ;
  assign n10360 = ~x435 & ~n10322 ;
  assign n10361 = n10382 ^ n10360 ;
  assign n10340 = n10392 ^ n9370 ;
  assign n10350 = n10340 ^ n10322 ;
  assign n10362 = n10361 ^ n10350 ;
  assign n10363 = n10362 ^ n9370 ;
  assign n10337 = n10320 ^ n4593 ;
  assign n10365 = n10337 ^ n9370 ;
  assign n10366 = ~n10363 & n10365 ;
  assign n10394 = n10393 ^ n9370 ;
  assign n10367 = n10393 ^ n10320 ;
  assign n10368 = n10394 ^ n10367 ;
  assign n10369 = n10393 ^ n10382 ;
  assign n10370 = n10394 ^ n10369 ;
  assign n10371 = ~n10368 & n10370 ;
  assign n10372 = n10366 & n10371 ;
  assign n10373 = n10372 ^ n10360 ;
  assign n10374 = n10373 ^ n8660 ;
  assign n10352 = n10393 ^ n10350 ;
  assign n10354 = n10394 ^ n10352 ;
  assign n10375 = n10374 ^ n10354 ;
  assign n10398 = n10375 ^ x435 ;
  assign n10399 = n10398 ^ n10394 ;
  assign n10400 = n9367 & n10399 ;
  assign n10401 = n10315 & n10400 ;
  assign n10404 = n10309 & n10401 ;
  assign n10402 = n10401 ^ n10315 ;
  assign n10405 = n10404 ^ n10402 ;
  assign n10432 = n10430 ^ n10405 ;
  assign n10536 = x804 ^ x622 ;
  assign n10537 = ~x1136 & n10536 ;
  assign n10538 = n10537 ^ x622 ;
  assign n10540 = n10538 ^ x743 ;
  assign n10539 = n10538 ^ x859 ;
  assign n10541 = n10540 ^ n10539 ;
  assign n10544 = x1136 & n10541 ;
  assign n10545 = n10544 ^ n10539 ;
  assign n10546 = x1134 & n10545 ;
  assign n10547 = n10546 ^ n10538 ;
  assign n10529 = x735 ^ x639 ;
  assign n10530 = n10529 ^ x783 ;
  assign n10533 = x1136 & n10530 ;
  assign n10534 = n10533 ^ x783 ;
  assign n10535 = n9474 & n10534 ;
  assign n10548 = n10547 ^ n10535 ;
  assign n10528 = x735 & x1136 ;
  assign n10549 = n10548 ^ n10528 ;
  assign n10550 = x1135 & n10549 ;
  assign n10551 = n10550 ^ n10547 ;
  assign n10552 = n9471 & n10551 ;
  assign n10434 = n9371 ^ x336 ;
  assign n10435 = n10434 ^ x463 ;
  assign n10436 = n10435 ^ n9371 ;
  assign n10437 = ~x592 & n10436 ;
  assign n10438 = n10437 ^ n10434 ;
  assign n10462 = n10438 ^ x437 ;
  assign n10463 = n10462 ^ n9370 ;
  assign n10440 = n9370 ^ x437 ;
  assign n10443 = n10440 ^ n9371 ;
  assign n10444 = n10443 ^ n4593 ;
  assign n10445 = n10444 ^ n10440 ;
  assign n10510 = n10463 ^ n10445 ;
  assign n10511 = n10510 ^ n9371 ;
  assign n10499 = n10511 ^ n10445 ;
  assign n10500 = n10499 ^ x437 ;
  assign n10478 = ~x437 & ~n10440 ;
  assign n10479 = n10500 ^ n10478 ;
  assign n10458 = n10510 ^ n9370 ;
  assign n10468 = n10458 ^ n10440 ;
  assign n10480 = n10479 ^ n10468 ;
  assign n10481 = n10480 ^ n9370 ;
  assign n10455 = n10438 ^ n4593 ;
  assign n10483 = n10455 ^ n9370 ;
  assign n10484 = ~n10481 & n10483 ;
  assign n10512 = n10511 ^ n9370 ;
  assign n10485 = n10511 ^ n10438 ;
  assign n10486 = n10512 ^ n10485 ;
  assign n10487 = n10511 ^ n10500 ;
  assign n10488 = n10512 ^ n10487 ;
  assign n10489 = ~n10486 & n10488 ;
  assign n10490 = n10484 & n10489 ;
  assign n10491 = n10490 ^ n10478 ;
  assign n10492 = n10491 ^ n8660 ;
  assign n10470 = n10511 ^ n10468 ;
  assign n10472 = n10512 ^ n10470 ;
  assign n10493 = n10492 ^ n10472 ;
  assign n10516 = n10493 ^ x437 ;
  assign n10517 = n10516 ^ n10512 ;
  assign n10433 = x362 & n9466 ;
  assign n10519 = n10517 ^ n10433 ;
  assign n10553 = n10552 ^ n10519 ;
  assign n10521 = n10519 ^ x256 ;
  assign n10520 = n10519 ^ x1070 ;
  assign n10522 = n10521 ^ n10520 ;
  assign n10525 = x199 & n10522 ;
  assign n10526 = n10525 ^ n10521 ;
  assign n10527 = ~n9367 & ~n10526 ;
  assign n10554 = n10553 ^ n10527 ;
  assign n10555 = n2991 & ~n10554 ;
  assign n10556 = n10555 ^ n10552 ;
  assign n10662 = x803 ^ x623 ;
  assign n10663 = ~x1136 & ~n10662 ;
  assign n10664 = n10663 ^ x623 ;
  assign n10666 = n10664 ^ x748 ;
  assign n10665 = n10664 ^ x876 ;
  assign n10667 = n10666 ^ n10665 ;
  assign n10670 = x1136 & n10667 ;
  assign n10671 = n10670 ^ n10665 ;
  assign n10672 = x1134 & n10671 ;
  assign n10673 = n10672 ^ n10664 ;
  assign n10655 = x730 ^ x710 ;
  assign n10656 = n10655 ^ x789 ;
  assign n10659 = x1136 & n10656 ;
  assign n10660 = n10659 ^ x789 ;
  assign n10661 = n9474 & n10660 ;
  assign n10674 = n10673 ^ n10661 ;
  assign n10654 = x730 & x1136 ;
  assign n10675 = n10674 ^ n10654 ;
  assign n10676 = x1135 & n10675 ;
  assign n10677 = n10676 ^ n10673 ;
  assign n10678 = n9472 & n10677 ;
  assign n10557 = x455 & n9466 ;
  assign n10560 = x199 & n7638 ;
  assign n10561 = n10560 ^ x296 ;
  assign n10562 = n9457 & ~n10561 ;
  assign n10563 = n10562 ^ n2991 ;
  assign n10564 = n9371 ^ x388 ;
  assign n10565 = n10564 ^ x412 ;
  assign n10566 = n10565 ^ n9371 ;
  assign n10567 = ~x592 & n10566 ;
  assign n10568 = n10567 ^ n10564 ;
  assign n10592 = n10568 ^ x436 ;
  assign n10593 = n10592 ^ n9370 ;
  assign n10570 = n9370 ^ x436 ;
  assign n10573 = n10570 ^ n9371 ;
  assign n10574 = n10573 ^ n4593 ;
  assign n10575 = n10574 ^ n10570 ;
  assign n10640 = n10593 ^ n10575 ;
  assign n10641 = n10640 ^ n9371 ;
  assign n10629 = n10641 ^ n10575 ;
  assign n10630 = n10629 ^ x436 ;
  assign n10608 = ~x436 & ~n10570 ;
  assign n10609 = n10630 ^ n10608 ;
  assign n10588 = n10640 ^ n9370 ;
  assign n10598 = n10588 ^ n10570 ;
  assign n10610 = n10609 ^ n10598 ;
  assign n10611 = n10610 ^ n9370 ;
  assign n10585 = n10568 ^ n4593 ;
  assign n10613 = n10585 ^ n9370 ;
  assign n10614 = ~n10611 & n10613 ;
  assign n10642 = n10641 ^ n9370 ;
  assign n10615 = n10641 ^ n10568 ;
  assign n10616 = n10642 ^ n10615 ;
  assign n10617 = n10641 ^ n10630 ;
  assign n10618 = n10642 ^ n10617 ;
  assign n10619 = ~n10616 & n10618 ;
  assign n10620 = n10614 & n10619 ;
  assign n10621 = n10620 ^ n10608 ;
  assign n10622 = n10621 ^ n8660 ;
  assign n10600 = n10641 ^ n10598 ;
  assign n10602 = n10642 ^ n10600 ;
  assign n10623 = n10622 ^ n10602 ;
  assign n10646 = n10623 ^ x436 ;
  assign n10647 = n10646 ^ n10642 ;
  assign n10648 = n9367 & n10647 ;
  assign n10649 = n10563 & n10648 ;
  assign n10652 = n10557 & n10649 ;
  assign n10650 = n10649 ^ n10563 ;
  assign n10653 = n10652 ^ n10650 ;
  assign n10680 = n10678 ^ n10653 ;
  assign n10784 = x881 ^ x746 ;
  assign n10785 = ~x1136 & n10784 ;
  assign n10786 = n10785 ^ x746 ;
  assign n10788 = n10786 ^ x606 ;
  assign n10787 = n10786 ^ x812 ;
  assign n10789 = n10788 ^ n10787 ;
  assign n10792 = x1136 & ~n10789 ;
  assign n10793 = n10792 ^ n10787 ;
  assign n10794 = ~x1134 & ~n10793 ;
  assign n10795 = n10794 ^ n10786 ;
  assign n10777 = x729 ^ x643 ;
  assign n10778 = n10777 ^ x787 ;
  assign n10781 = x1136 & n10778 ;
  assign n10782 = n10781 ^ x787 ;
  assign n10783 = n9474 & n10782 ;
  assign n10796 = n10795 ^ n10783 ;
  assign n10776 = x729 & x1136 ;
  assign n10797 = n10796 ^ n10776 ;
  assign n10798 = x1135 & n10797 ;
  assign n10799 = n10798 ^ n10795 ;
  assign n10800 = n9471 & n10799 ;
  assign n10682 = n9371 ^ x386 ;
  assign n10683 = n10682 ^ x410 ;
  assign n10684 = n10683 ^ n9371 ;
  assign n10685 = ~x592 & n10684 ;
  assign n10686 = n10685 ^ n10682 ;
  assign n10710 = n10686 ^ x434 ;
  assign n10711 = n10710 ^ n9370 ;
  assign n10688 = n9370 ^ x434 ;
  assign n10691 = n10688 ^ n9371 ;
  assign n10692 = n10691 ^ n4593 ;
  assign n10693 = n10692 ^ n10688 ;
  assign n10758 = n10711 ^ n10693 ;
  assign n10759 = n10758 ^ n9371 ;
  assign n10747 = n10759 ^ n10693 ;
  assign n10748 = n10747 ^ x434 ;
  assign n10726 = ~x434 & ~n10688 ;
  assign n10727 = n10748 ^ n10726 ;
  assign n10706 = n10758 ^ n9370 ;
  assign n10716 = n10706 ^ n10688 ;
  assign n10728 = n10727 ^ n10716 ;
  assign n10729 = n10728 ^ n9370 ;
  assign n10703 = n10686 ^ n4593 ;
  assign n10731 = n10703 ^ n9370 ;
  assign n10732 = ~n10729 & n10731 ;
  assign n10760 = n10759 ^ n9370 ;
  assign n10733 = n10759 ^ n10686 ;
  assign n10734 = n10760 ^ n10733 ;
  assign n10735 = n10759 ^ n10748 ;
  assign n10736 = n10760 ^ n10735 ;
  assign n10737 = ~n10734 & n10736 ;
  assign n10738 = n10732 & n10737 ;
  assign n10739 = n10738 ^ n10726 ;
  assign n10740 = n10739 ^ n8660 ;
  assign n10718 = n10759 ^ n10716 ;
  assign n10720 = n10760 ^ n10718 ;
  assign n10741 = n10740 ^ n10720 ;
  assign n10764 = n10741 ^ x434 ;
  assign n10765 = n10764 ^ n10760 ;
  assign n10681 = x361 & n9466 ;
  assign n10767 = n10765 ^ n10681 ;
  assign n10801 = n10800 ^ n10767 ;
  assign n10773 = x199 & n7629 ;
  assign n10769 = n10767 ^ x293 ;
  assign n10774 = n10773 ^ n10769 ;
  assign n10775 = ~n9367 & ~n10774 ;
  assign n10802 = n10801 ^ n10775 ;
  assign n10803 = n2991 & ~n10802 ;
  assign n10804 = n10803 ^ n10800 ;
  assign n10822 = n9371 ^ x335 ;
  assign n10823 = n10822 ^ x366 ;
  assign n10824 = n10823 ^ n9371 ;
  assign n10825 = x592 & n10824 ;
  assign n10826 = n10825 ^ n10822 ;
  assign n10850 = n10826 ^ x416 ;
  assign n10851 = n10850 ^ n9370 ;
  assign n10828 = n9370 ^ x416 ;
  assign n10831 = n10828 ^ n9371 ;
  assign n10832 = n10831 ^ n4593 ;
  assign n10833 = n10832 ^ n10828 ;
  assign n10898 = n10851 ^ n10833 ;
  assign n10899 = n10898 ^ n9371 ;
  assign n10887 = n10899 ^ n10833 ;
  assign n10888 = n10887 ^ x416 ;
  assign n10866 = ~x416 & ~n10828 ;
  assign n10867 = n10888 ^ n10866 ;
  assign n10846 = n10898 ^ n9370 ;
  assign n10856 = n10846 ^ n10828 ;
  assign n10868 = n10867 ^ n10856 ;
  assign n10869 = n10868 ^ n9370 ;
  assign n10843 = n10826 ^ n4593 ;
  assign n10871 = n10843 ^ n9370 ;
  assign n10872 = ~n10869 & n10871 ;
  assign n10900 = n10899 ^ n9370 ;
  assign n10873 = n10899 ^ n10826 ;
  assign n10874 = n10900 ^ n10873 ;
  assign n10875 = n10899 ^ n10888 ;
  assign n10876 = n10900 ^ n10875 ;
  assign n10877 = ~n10874 & n10876 ;
  assign n10878 = n10872 & n10877 ;
  assign n10879 = n10878 ^ n10866 ;
  assign n10880 = n10879 ^ n8660 ;
  assign n10858 = n10899 ^ n10856 ;
  assign n10860 = n10900 ^ n10858 ;
  assign n10881 = n10880 ^ n10860 ;
  assign n10904 = n10881 ^ x416 ;
  assign n10905 = n10904 ^ n10900 ;
  assign n10821 = x344 & n9466 ;
  assign n10907 = n10905 ^ n10821 ;
  assign n10909 = n10907 ^ x259 ;
  assign n10908 = n10907 ^ x1069 ;
  assign n10910 = n10909 ^ n10908 ;
  assign n10913 = x199 & n10910 ;
  assign n10914 = n10913 ^ n10909 ;
  assign n10915 = ~n9367 & ~n10914 ;
  assign n10916 = n10915 ^ n10907 ;
  assign n5942 = x742 ^ x704 ;
  assign n10805 = ~x1135 & n5942 ;
  assign n10806 = n10805 ^ x704 ;
  assign n10808 = n10806 ^ x620 ;
  assign n10807 = n10806 ^ x635 ;
  assign n10809 = n10808 ^ n10807 ;
  assign n10812 = ~x1135 & ~n10809 ;
  assign n10813 = n10812 ^ n10807 ;
  assign n10814 = ~x1134 & n10813 ;
  assign n10815 = n10814 ^ n10806 ;
  assign n10816 = x1136 & n9471 ;
  assign n10817 = ~n10815 & n10816 ;
  assign n10918 = n10916 ^ n10817 ;
  assign n10818 = n10817 ^ n9471 ;
  assign n10819 = x870 & n10024 ;
  assign n10820 = n10818 & n10819 ;
  assign n10919 = n10918 ^ n10820 ;
  assign n10920 = ~n2991 & ~n10919 ;
  assign n10921 = n10920 ^ n10916 ;
  assign n5976 = x760 ^ x688 ;
  assign n10922 = ~x1135 & n5976 ;
  assign n10923 = n10922 ^ x688 ;
  assign n10925 = n10923 ^ x613 ;
  assign n10924 = n10923 ^ x632 ;
  assign n10926 = n10925 ^ n10924 ;
  assign n10929 = ~x1135 & ~n10926 ;
  assign n10930 = n10929 ^ n10924 ;
  assign n10931 = ~x1134 & n10930 ;
  assign n10932 = n10931 ^ n10923 ;
  assign n10933 = n10020 & ~n10932 ;
  assign n10934 = n10933 ^ n9472 ;
  assign n10936 = x856 & n10024 ;
  assign n10937 = n10934 & n10936 ;
  assign n10938 = n10937 ^ n10933 ;
  assign n10939 = x1067 ^ x260 ;
  assign n10942 = x199 & n10939 ;
  assign n10943 = n10942 ^ x260 ;
  assign n10944 = n9457 & ~n10943 ;
  assign n10945 = n10944 ^ n2991 ;
  assign n10946 = x393 & n3022 ;
  assign n10947 = x368 & ~x590 ;
  assign n10948 = ~x591 & n9369 ;
  assign n10949 = n10947 & n10948 ;
  assign n10950 = n10949 ^ n9369 ;
  assign n10951 = n10946 & n10950 ;
  assign n10952 = n10951 ^ n10950 ;
  assign n10960 = x346 & n10952 ;
  assign n10961 = n3109 & n10960 ;
  assign n10962 = n10961 ^ n3109 ;
  assign n10953 = n10952 ^ n9369 ;
  assign n10954 = n10953 ^ n3109 ;
  assign n10963 = n10962 ^ n10954 ;
  assign n10964 = n9367 & ~n10963 ;
  assign n10965 = n10945 & n10964 ;
  assign n10973 = ~n9370 & n10965 ;
  assign n10974 = x418 & n10973 ;
  assign n10975 = n10974 ^ x418 ;
  assign n10966 = n10965 ^ n10945 ;
  assign n10967 = n10966 ^ x418 ;
  assign n10976 = n10975 ^ n10967 ;
  assign n10977 = ~n10938 & ~n10976 ;
  assign n10978 = n9371 ^ x389 ;
  assign n10979 = n10978 ^ x413 ;
  assign n10980 = n10979 ^ n9371 ;
  assign n10981 = ~x592 & n10980 ;
  assign n10982 = n10981 ^ n10978 ;
  assign n11006 = n10982 ^ x438 ;
  assign n11007 = n11006 ^ n9370 ;
  assign n10984 = n9370 ^ x438 ;
  assign n10987 = n10984 ^ n9371 ;
  assign n10988 = n10987 ^ n4593 ;
  assign n10989 = n10988 ^ n10984 ;
  assign n11054 = n11007 ^ n10989 ;
  assign n11055 = n11054 ^ n9371 ;
  assign n11043 = n11055 ^ n10989 ;
  assign n11044 = n11043 ^ x438 ;
  assign n11022 = ~x438 & ~n10984 ;
  assign n11023 = n11044 ^ n11022 ;
  assign n11002 = n11054 ^ n9370 ;
  assign n11012 = n11002 ^ n10984 ;
  assign n11024 = n11023 ^ n11012 ;
  assign n11025 = n11024 ^ n9370 ;
  assign n10999 = n10982 ^ n4593 ;
  assign n11027 = n10999 ^ n9370 ;
  assign n11028 = ~n11025 & n11027 ;
  assign n11056 = n11055 ^ n9370 ;
  assign n11029 = n11055 ^ n10982 ;
  assign n11030 = n11056 ^ n11029 ;
  assign n11031 = n11055 ^ n11044 ;
  assign n11032 = n11056 ^ n11031 ;
  assign n11033 = ~n11030 & n11032 ;
  assign n11034 = n11028 & n11033 ;
  assign n11035 = n11034 ^ n11022 ;
  assign n11036 = n11035 ^ n8660 ;
  assign n11014 = n11055 ^ n11012 ;
  assign n11016 = n11056 ^ n11014 ;
  assign n11037 = n11036 ^ n11016 ;
  assign n11060 = n11037 ^ x438 ;
  assign n11061 = n11060 ^ n11056 ;
  assign n11062 = n9367 & n11061 ;
  assign n11063 = x450 & n9466 ;
  assign n11064 = n11062 & ~n11063 ;
  assign n11065 = x1036 ^ x255 ;
  assign n11068 = x199 & n11065 ;
  assign n11069 = n11068 ^ x255 ;
  assign n11070 = n9457 & ~n11069 ;
  assign n11071 = n11070 ^ n2991 ;
  assign n11072 = ~n11064 & n11071 ;
  assign n11081 = x810 ^ x621 ;
  assign n11082 = ~x1136 & n11081 ;
  assign n11083 = n11082 ^ x621 ;
  assign n11085 = n11083 ^ x739 ;
  assign n11084 = n11083 ^ x874 ;
  assign n11086 = n11085 ^ n11084 ;
  assign n11089 = x1136 & n11086 ;
  assign n11090 = n11089 ^ n11084 ;
  assign n11091 = x1134 & n11090 ;
  assign n11092 = n11091 ^ n11083 ;
  assign n11074 = x690 ^ x665 ;
  assign n11075 = n11074 ^ x791 ;
  assign n11078 = x1136 & n11075 ;
  assign n11079 = n11078 ^ x791 ;
  assign n11080 = n9474 & n11079 ;
  assign n11093 = n11092 ^ n11080 ;
  assign n11073 = x690 & x1136 ;
  assign n11094 = n11093 ^ n11073 ;
  assign n11095 = x1135 & n11094 ;
  assign n11096 = n11095 ^ n11092 ;
  assign n11097 = n9472 & n11096 ;
  assign n11098 = ~n11072 & ~n11097 ;
  assign n11099 = x1100 ^ x680 ;
  assign n11102 = n9135 & n11099 ;
  assign n11103 = n11102 ^ x680 ;
  assign n11104 = ~x962 & n11103 ;
  assign n11105 = x1103 ^ x681 ;
  assign n11108 = n9135 & n11105 ;
  assign n11109 = n11108 ^ x681 ;
  assign n11110 = ~x962 & n11109 ;
  assign n11111 = n9371 ^ x367 ;
  assign n11112 = n11111 ^ x392 ;
  assign n11113 = n11112 ^ n9371 ;
  assign n11114 = ~x592 & n11113 ;
  assign n11115 = n11114 ^ n11111 ;
  assign n11139 = n11115 ^ x417 ;
  assign n11140 = n11139 ^ n9370 ;
  assign n11117 = n9370 ^ x417 ;
  assign n11120 = n11117 ^ n9371 ;
  assign n11121 = n11120 ^ n4593 ;
  assign n11122 = n11121 ^ n11117 ;
  assign n11187 = n11140 ^ n11122 ;
  assign n11188 = n11187 ^ n9371 ;
  assign n11176 = n11188 ^ n11122 ;
  assign n11177 = n11176 ^ x417 ;
  assign n11155 = ~x417 & ~n11117 ;
  assign n11156 = n11177 ^ n11155 ;
  assign n11135 = n11187 ^ n9370 ;
  assign n11145 = n11135 ^ n11117 ;
  assign n11157 = n11156 ^ n11145 ;
  assign n11158 = n11157 ^ n9370 ;
  assign n11132 = n11115 ^ n4593 ;
  assign n11160 = n11132 ^ n9370 ;
  assign n11161 = ~n11158 & n11160 ;
  assign n11189 = n11188 ^ n9370 ;
  assign n11162 = n11188 ^ n11115 ;
  assign n11163 = n11189 ^ n11162 ;
  assign n11164 = n11188 ^ n11177 ;
  assign n11165 = n11189 ^ n11164 ;
  assign n11166 = ~n11163 & n11165 ;
  assign n11167 = n11161 & n11166 ;
  assign n11168 = n11167 ^ n11155 ;
  assign n11169 = n11168 ^ n8660 ;
  assign n11147 = n11188 ^ n11145 ;
  assign n11149 = n11189 ^ n11147 ;
  assign n11170 = n11169 ^ n11149 ;
  assign n11193 = n11170 ^ x417 ;
  assign n11194 = n11193 ^ n11189 ;
  assign n11195 = n9367 & n11194 ;
  assign n11196 = x345 & n9466 ;
  assign n11197 = n11195 & ~n11196 ;
  assign n11198 = x1039 ^ x251 ;
  assign n11201 = x199 & n11198 ;
  assign n11202 = n11201 ^ x251 ;
  assign n11203 = n9457 & ~n11202 ;
  assign n11204 = n11203 ^ n2991 ;
  assign n11205 = ~n11197 & n11204 ;
  assign n5954 = x757 ^ x686 ;
  assign n11206 = ~x1135 & n5954 ;
  assign n11207 = n11206 ^ x686 ;
  assign n11209 = n11207 ^ x610 ;
  assign n11208 = n11207 ^ x631 ;
  assign n11210 = n11209 ^ n11208 ;
  assign n11213 = ~x1135 & ~n11210 ;
  assign n11214 = n11213 ^ n11208 ;
  assign n11215 = ~x1134 & n11214 ;
  assign n11216 = n11215 ^ n11207 ;
  assign n11217 = n10020 & ~n11216 ;
  assign n11218 = n11217 ^ n9472 ;
  assign n11220 = x848 & n10024 ;
  assign n11221 = n11218 & n11220 ;
  assign n11222 = n11221 ^ n11217 ;
  assign n11223 = ~n11205 & ~n11222 ;
  assign n11224 = x1130 ^ x684 ;
  assign n11227 = n9134 & ~n11224 ;
  assign n11228 = n11227 ^ x684 ;
  assign n11229 = ~x962 & ~n11228 ;
  assign n11230 = n9371 ^ x382 ;
  assign n11231 = n11230 ^ x406 ;
  assign n11232 = n11231 ^ n9371 ;
  assign n11233 = ~x592 & n11232 ;
  assign n11234 = n11233 ^ n11230 ;
  assign n11258 = n11234 ^ x430 ;
  assign n11259 = n11258 ^ n9370 ;
  assign n11236 = n9370 ^ x430 ;
  assign n11239 = n11236 ^ n9371 ;
  assign n11240 = n11239 ^ n4593 ;
  assign n11241 = n11240 ^ n11236 ;
  assign n11306 = n11259 ^ n11241 ;
  assign n11307 = n11306 ^ n9371 ;
  assign n11295 = n11307 ^ n11241 ;
  assign n11296 = n11295 ^ x430 ;
  assign n11274 = ~x430 & ~n11236 ;
  assign n11275 = n11296 ^ n11274 ;
  assign n11254 = n11306 ^ n9370 ;
  assign n11264 = n11254 ^ n11236 ;
  assign n11276 = n11275 ^ n11264 ;
  assign n11277 = n11276 ^ n9370 ;
  assign n11251 = n11234 ^ n4593 ;
  assign n11279 = n11251 ^ n9370 ;
  assign n11280 = ~n11277 & n11279 ;
  assign n11308 = n11307 ^ n9370 ;
  assign n11281 = n11307 ^ n11234 ;
  assign n11282 = n11308 ^ n11281 ;
  assign n11283 = n11307 ^ n11296 ;
  assign n11284 = n11308 ^ n11283 ;
  assign n11285 = ~n11282 & n11284 ;
  assign n11286 = n11280 & n11285 ;
  assign n11287 = n11286 ^ n11274 ;
  assign n11288 = n11287 ^ n8660 ;
  assign n11266 = n11307 ^ n11264 ;
  assign n11268 = n11308 ^ n11266 ;
  assign n11289 = n11288 ^ n11268 ;
  assign n11312 = n11289 ^ x430 ;
  assign n11313 = n11312 ^ n11308 ;
  assign n11314 = n9367 & n11313 ;
  assign n11315 = x357 & n9466 ;
  assign n11316 = n11314 & ~n11315 ;
  assign n11317 = n7341 ^ x1076 ;
  assign n11320 = ~x199 & n11317 ;
  assign n11321 = n11320 ^ x1076 ;
  assign n11322 = n9457 & ~n11321 ;
  assign n11323 = n11322 ^ n2991 ;
  assign n11324 = ~n11316 & n11323 ;
  assign n11331 = x744 ^ x728 ;
  assign n11332 = ~x1135 & n11331 ;
  assign n11333 = n11332 ^ x728 ;
  assign n11335 = n11333 ^ x652 ;
  assign n11334 = n11333 ^ x657 ;
  assign n11336 = n11335 ^ n11334 ;
  assign n11339 = ~x1135 & ~n11336 ;
  assign n11340 = n11339 ^ n11334 ;
  assign n11341 = ~x1134 & n11340 ;
  assign n11342 = n11341 ^ n11333 ;
  assign n11325 = x860 ^ x813 ;
  assign n11328 = ~x1134 & n11325 ;
  assign n11329 = n11328 ^ x860 ;
  assign n11330 = ~x1135 & n11329 ;
  assign n11343 = n11342 ^ n11330 ;
  assign n11344 = ~x1136 & ~n11343 ;
  assign n11345 = n11344 ^ n11342 ;
  assign n11346 = n9472 & ~n11345 ;
  assign n11347 = ~n11324 & ~n11346 ;
  assign n11348 = x1113 ^ x686 ;
  assign n11351 = n9134 & ~n11348 ;
  assign n11352 = n11351 ^ x686 ;
  assign n11353 = ~x962 & ~n11352 ;
  assign n11354 = x1127 ^ x687 ;
  assign n11357 = n9134 & n11354 ;
  assign n11358 = n11357 ^ x687 ;
  assign n11359 = ~x962 & n11358 ;
  assign n11360 = x1115 ^ x688 ;
  assign n11363 = n9134 & ~n11360 ;
  assign n11364 = n11363 ^ x688 ;
  assign n11365 = ~x962 & ~n11364 ;
  assign n6050 = x752 ^ x703 ;
  assign n11467 = ~x1135 & ~n6050 ;
  assign n11468 = n11467 ^ x703 ;
  assign n11470 = n11468 ^ x655 ;
  assign n11469 = n11468 ^ x658 ;
  assign n11471 = n11470 ^ n11469 ;
  assign n11474 = x1135 & ~n11471 ;
  assign n11475 = n11474 ^ n11469 ;
  assign n11476 = ~x1134 & n11475 ;
  assign n11477 = n11476 ^ n11468 ;
  assign n11461 = x843 ^ x798 ;
  assign n11464 = ~x1134 & n11461 ;
  assign n11465 = n11464 ^ x843 ;
  assign n11466 = ~x1135 & n11465 ;
  assign n11478 = n11477 ^ n11466 ;
  assign n11479 = ~x1136 & n11478 ;
  assign n11480 = n11479 ^ n11477 ;
  assign n11481 = n9471 & n11480 ;
  assign n11367 = n9371 ^ x376 ;
  assign n11368 = n11367 ^ x401 ;
  assign n11369 = n11368 ^ n9371 ;
  assign n11370 = ~x592 & n11369 ;
  assign n11371 = n11370 ^ n11367 ;
  assign n11395 = n11371 ^ x426 ;
  assign n11396 = n11395 ^ n9370 ;
  assign n11373 = n9370 ^ x426 ;
  assign n11376 = n11373 ^ n9371 ;
  assign n11377 = n11376 ^ n4593 ;
  assign n11378 = n11377 ^ n11373 ;
  assign n11443 = n11396 ^ n11378 ;
  assign n11444 = n11443 ^ n9371 ;
  assign n11432 = n11444 ^ n11378 ;
  assign n11433 = n11432 ^ x426 ;
  assign n11411 = ~x426 & ~n11373 ;
  assign n11412 = n11433 ^ n11411 ;
  assign n11391 = n11443 ^ n9370 ;
  assign n11401 = n11391 ^ n11373 ;
  assign n11413 = n11412 ^ n11401 ;
  assign n11414 = n11413 ^ n9370 ;
  assign n11388 = n11371 ^ n4593 ;
  assign n11416 = n11388 ^ n9370 ;
  assign n11417 = ~n11414 & n11416 ;
  assign n11445 = n11444 ^ n9370 ;
  assign n11418 = n11444 ^ n11371 ;
  assign n11419 = n11445 ^ n11418 ;
  assign n11420 = n11444 ^ n11433 ;
  assign n11421 = n11445 ^ n11420 ;
  assign n11422 = ~n11419 & n11421 ;
  assign n11423 = n11417 & n11422 ;
  assign n11424 = n11423 ^ n11411 ;
  assign n11425 = n11424 ^ n8660 ;
  assign n11403 = n11444 ^ n11401 ;
  assign n11405 = n11445 ^ n11403 ;
  assign n11426 = n11425 ^ n11405 ;
  assign n11449 = n11426 ^ x426 ;
  assign n11450 = n11449 ^ n11445 ;
  assign n11366 = x351 & n9466 ;
  assign n11452 = n11450 ^ n11366 ;
  assign n11482 = n11481 ^ n11452 ;
  assign n11454 = n11452 ^ x1079 ;
  assign n11453 = n11452 ^ n7311 ;
  assign n11455 = n11454 ^ n11453 ;
  assign n11458 = ~x199 & n11455 ;
  assign n11459 = n11458 ^ n11454 ;
  assign n11460 = ~n9367 & ~n11459 ;
  assign n11483 = n11482 ^ n11460 ;
  assign n11484 = n2991 & ~n11483 ;
  assign n11485 = n11484 ^ n11481 ;
  assign n11486 = x1108 ^ x690 ;
  assign n11489 = n9134 & n11486 ;
  assign n11490 = n11489 ^ x690 ;
  assign n11491 = ~x962 & n11490 ;
  assign n11492 = x1107 ^ x691 ;
  assign n11495 = n9134 & n11492 ;
  assign n11496 = n11495 ^ x691 ;
  assign n11497 = ~x962 & n11496 ;
  assign n11498 = n9371 ^ x317 ;
  assign n11499 = n11498 ^ x402 ;
  assign n11500 = n11499 ^ n9371 ;
  assign n11501 = ~x592 & n11500 ;
  assign n11502 = n11501 ^ n11498 ;
  assign n11526 = n11502 ^ x427 ;
  assign n11527 = n11526 ^ n9370 ;
  assign n11504 = n9370 ^ x427 ;
  assign n11507 = n11504 ^ n9371 ;
  assign n11508 = n11507 ^ n4593 ;
  assign n11509 = n11508 ^ n11504 ;
  assign n11574 = n11527 ^ n11509 ;
  assign n11575 = n11574 ^ n9371 ;
  assign n11563 = n11575 ^ n11509 ;
  assign n11564 = n11563 ^ x427 ;
  assign n11542 = ~x427 & ~n11504 ;
  assign n11543 = n11564 ^ n11542 ;
  assign n11522 = n11574 ^ n9370 ;
  assign n11532 = n11522 ^ n11504 ;
  assign n11544 = n11543 ^ n11532 ;
  assign n11545 = n11544 ^ n9370 ;
  assign n11519 = n11502 ^ n4593 ;
  assign n11547 = n11519 ^ n9370 ;
  assign n11548 = ~n11545 & n11547 ;
  assign n11576 = n11575 ^ n9370 ;
  assign n11549 = n11575 ^ n11502 ;
  assign n11550 = n11576 ^ n11549 ;
  assign n11551 = n11575 ^ n11564 ;
  assign n11552 = n11576 ^ n11551 ;
  assign n11553 = ~n11550 & n11552 ;
  assign n11554 = n11548 & n11553 ;
  assign n11555 = n11554 ^ n11542 ;
  assign n11556 = n11555 ^ n8660 ;
  assign n11534 = n11575 ^ n11532 ;
  assign n11536 = n11576 ^ n11534 ;
  assign n11557 = n11556 ^ n11536 ;
  assign n11580 = n11557 ^ x427 ;
  assign n11581 = n11580 ^ n11576 ;
  assign n11582 = n9367 & n11581 ;
  assign n11583 = x352 & n9466 ;
  assign n11584 = n11582 & ~n11583 ;
  assign n11585 = n7323 ^ x1078 ;
  assign n11588 = ~x199 & n11585 ;
  assign n11589 = n11588 ^ x1078 ;
  assign n11590 = n9457 & ~n11589 ;
  assign n11591 = n11590 ^ n2991 ;
  assign n11592 = ~n11584 & n11591 ;
  assign n5849 = x770 ^ x726 ;
  assign n11599 = ~x1135 & ~n5849 ;
  assign n11600 = n11599 ^ x726 ;
  assign n11602 = n11600 ^ x649 ;
  assign n11601 = n11600 ^ x656 ;
  assign n11603 = n11602 ^ n11601 ;
  assign n11606 = x1135 & ~n11603 ;
  assign n11607 = n11606 ^ n11601 ;
  assign n11608 = ~x1134 & n11607 ;
  assign n11609 = n11608 ^ n11600 ;
  assign n11593 = x844 ^ x801 ;
  assign n11596 = ~x1134 & n11593 ;
  assign n11597 = n11596 ^ x844 ;
  assign n11598 = ~x1135 & n11597 ;
  assign n11610 = n11609 ^ n11598 ;
  assign n11611 = ~x1136 & n11610 ;
  assign n11612 = n11611 ^ n11609 ;
  assign n11613 = n9472 & n11612 ;
  assign n11614 = ~n11592 & ~n11613 ;
  assign n11615 = x1129 ^ x693 ;
  assign n11618 = n9135 & ~n11615 ;
  assign n11619 = n11618 ^ x693 ;
  assign n11620 = ~x962 & ~n11619 ;
  assign n11621 = x1128 ^ x694 ;
  assign n11624 = n9134 & ~n11621 ;
  assign n11625 = n11624 ^ x694 ;
  assign n11626 = ~x962 & ~n11625 ;
  assign n11627 = x1111 ^ x695 ;
  assign n11630 = n9135 & ~n11627 ;
  assign n11631 = n11630 ^ x695 ;
  assign n11632 = ~x962 & ~n11631 ;
  assign n11633 = x1100 ^ x696 ;
  assign n11636 = n9134 & n11633 ;
  assign n11637 = n11636 ^ x696 ;
  assign n11638 = ~x962 & n11637 ;
  assign n11639 = x1129 ^ x697 ;
  assign n11642 = n9134 & ~n11639 ;
  assign n11643 = n11642 ^ x697 ;
  assign n11644 = ~x962 & ~n11643 ;
  assign n11645 = x1116 ^ x698 ;
  assign n11648 = n9134 & ~n11645 ;
  assign n11649 = n11648 ^ x698 ;
  assign n11650 = ~x962 & ~n11649 ;
  assign n11651 = x1103 ^ x699 ;
  assign n11654 = n9134 & n11651 ;
  assign n11655 = n11654 ^ x699 ;
  assign n11656 = ~x962 & n11655 ;
  assign n11657 = x1110 ^ x700 ;
  assign n11660 = n9134 & n11657 ;
  assign n11661 = n11660 ^ x700 ;
  assign n11662 = ~x962 & n11661 ;
  assign n11663 = x1123 ^ x701 ;
  assign n11666 = n9134 & ~n11663 ;
  assign n11667 = n11666 ^ x701 ;
  assign n11668 = ~x962 & ~n11667 ;
  assign n11669 = x1117 ^ x702 ;
  assign n11672 = n9134 & ~n11669 ;
  assign n11673 = n11672 ^ x702 ;
  assign n11674 = ~x962 & ~n11673 ;
  assign n11675 = x1124 ^ x703 ;
  assign n11678 = n9134 & n11675 ;
  assign n11679 = n11678 ^ x703 ;
  assign n11680 = ~x962 & n11679 ;
  assign n11681 = x1112 ^ x704 ;
  assign n11684 = n9134 & ~n11681 ;
  assign n11685 = n11684 ^ x704 ;
  assign n11686 = ~x962 & ~n11685 ;
  assign n11687 = x1125 ^ x705 ;
  assign n11690 = n9134 & n11687 ;
  assign n11691 = n11690 ^ x705 ;
  assign n11692 = ~x962 & n11691 ;
  assign n11693 = x1105 ^ x706 ;
  assign n11696 = n9134 & n11693 ;
  assign n11697 = n11696 ^ x706 ;
  assign n11698 = ~x962 & n11697 ;
  assign n11699 = n9371 ^ x370 ;
  assign n11700 = n11699 ^ x395 ;
  assign n11701 = n11700 ^ n9371 ;
  assign n11702 = ~x592 & n11701 ;
  assign n11703 = n11702 ^ n11699 ;
  assign n11727 = n11703 ^ x420 ;
  assign n11728 = n11727 ^ n9370 ;
  assign n11705 = n9370 ^ x420 ;
  assign n11708 = n11705 ^ n9371 ;
  assign n11709 = n11708 ^ n4593 ;
  assign n11710 = n11709 ^ n11705 ;
  assign n11775 = n11728 ^ n11710 ;
  assign n11776 = n11775 ^ n9371 ;
  assign n11764 = n11776 ^ n11710 ;
  assign n11765 = n11764 ^ x420 ;
  assign n11743 = ~x420 & ~n11705 ;
  assign n11744 = n11765 ^ n11743 ;
  assign n11723 = n11775 ^ n9370 ;
  assign n11733 = n11723 ^ n11705 ;
  assign n11745 = n11744 ^ n11733 ;
  assign n11746 = n11745 ^ n9370 ;
  assign n11720 = n11703 ^ n4593 ;
  assign n11748 = n11720 ^ n9370 ;
  assign n11749 = ~n11746 & n11748 ;
  assign n11777 = n11776 ^ n9370 ;
  assign n11750 = n11776 ^ n11703 ;
  assign n11751 = n11777 ^ n11750 ;
  assign n11752 = n11776 ^ n11765 ;
  assign n11753 = n11777 ^ n11752 ;
  assign n11754 = ~n11751 & n11753 ;
  assign n11755 = n11749 & n11754 ;
  assign n11756 = n11755 ^ n11743 ;
  assign n11757 = n11756 ^ n8660 ;
  assign n11735 = n11776 ^ n11733 ;
  assign n11737 = n11777 ^ n11735 ;
  assign n11758 = n11757 ^ n11737 ;
  assign n11781 = n11758 ^ x420 ;
  assign n11782 = n11781 ^ n11777 ;
  assign n11783 = n9367 & n11782 ;
  assign n11784 = x347 & n9466 ;
  assign n11785 = n11783 & ~n11784 ;
  assign n11791 = x200 & n7688 ;
  assign n11787 = x1055 ^ x304 ;
  assign n11792 = n11791 ^ n11787 ;
  assign n11793 = ~x199 & n11792 ;
  assign n11794 = n11793 ^ x1055 ;
  assign n11795 = n9457 & ~n11794 ;
  assign n11796 = n11795 ^ n2991 ;
  assign n11797 = ~n11785 & n11796 ;
  assign n5989 = x753 ^ x702 ;
  assign n11798 = ~x1135 & n5989 ;
  assign n11799 = n11798 ^ x702 ;
  assign n11801 = n11799 ^ x618 ;
  assign n11800 = n11799 ^ x627 ;
  assign n11802 = n11801 ^ n11800 ;
  assign n11805 = ~x1135 & n11802 ;
  assign n11806 = n11805 ^ n11800 ;
  assign n11807 = ~x1134 & ~n11806 ;
  assign n11808 = n11807 ^ n11799 ;
  assign n11809 = n10020 & ~n11808 ;
  assign n11810 = n11809 ^ n9472 ;
  assign n11812 = x847 & n10024 ;
  assign n11813 = n11810 & n11812 ;
  assign n11814 = n11813 ^ n11809 ;
  assign n11815 = ~n11797 & ~n11814 ;
  assign n11840 = n9371 ^ x328 ;
  assign n11841 = n11840 ^ x442 ;
  assign n11842 = n11841 ^ n9371 ;
  assign n11843 = x592 & n11842 ;
  assign n11844 = n11843 ^ n11840 ;
  assign n11868 = n11844 ^ x459 ;
  assign n11869 = n11868 ^ n9370 ;
  assign n11846 = n9370 ^ x459 ;
  assign n11849 = n11846 ^ n9371 ;
  assign n11850 = n11849 ^ n4593 ;
  assign n11851 = n11850 ^ n11846 ;
  assign n11916 = n11869 ^ n11851 ;
  assign n11917 = n11916 ^ n9371 ;
  assign n11905 = n11917 ^ n11851 ;
  assign n11906 = n11905 ^ x459 ;
  assign n11884 = ~x459 & ~n11846 ;
  assign n11885 = n11906 ^ n11884 ;
  assign n11864 = n11916 ^ n9370 ;
  assign n11874 = n11864 ^ n11846 ;
  assign n11886 = n11885 ^ n11874 ;
  assign n11887 = n11886 ^ n9370 ;
  assign n11861 = n11844 ^ n4593 ;
  assign n11889 = n11861 ^ n9370 ;
  assign n11890 = ~n11887 & n11889 ;
  assign n11918 = n11917 ^ n9370 ;
  assign n11891 = n11917 ^ n11844 ;
  assign n11892 = n11918 ^ n11891 ;
  assign n11893 = n11917 ^ n11906 ;
  assign n11894 = n11918 ^ n11893 ;
  assign n11895 = ~n11892 & n11894 ;
  assign n11896 = n11890 & n11895 ;
  assign n11897 = n11896 ^ n11884 ;
  assign n11898 = n11897 ^ n8660 ;
  assign n11876 = n11917 ^ n11874 ;
  assign n11878 = n11918 ^ n11876 ;
  assign n11899 = n11898 ^ n11878 ;
  assign n11922 = n11899 ^ x459 ;
  assign n11923 = n11922 ^ n11918 ;
  assign n11839 = x321 & n9466 ;
  assign n11925 = n11923 ^ n11839 ;
  assign n11926 = n11925 ^ x1058 ;
  assign n11836 = x200 & n7691 ;
  assign n11832 = x1058 ^ x305 ;
  assign n11837 = n11836 ^ n11832 ;
  assign n11838 = ~x199 & n11837 ;
  assign n11927 = n11926 ^ n11838 ;
  assign n11928 = ~n9367 & ~n11927 ;
  assign n11929 = n11928 ^ n11925 ;
  assign n5999 = x754 ^ x709 ;
  assign n11816 = ~x1135 & n5999 ;
  assign n11817 = n11816 ^ x709 ;
  assign n11819 = n11817 ^ x609 ;
  assign n11818 = n11817 ^ x660 ;
  assign n11820 = n11819 ^ n11818 ;
  assign n11823 = ~x1135 & n11820 ;
  assign n11824 = n11823 ^ n11818 ;
  assign n11825 = ~x1134 & ~n11824 ;
  assign n11826 = n11825 ^ n11817 ;
  assign n11827 = n10816 & ~n11826 ;
  assign n11931 = n11929 ^ n11827 ;
  assign n11828 = n11827 ^ n9471 ;
  assign n11829 = x857 & n10024 ;
  assign n11830 = n11828 & n11829 ;
  assign n11932 = n11931 ^ n11830 ;
  assign n11933 = ~n2991 & ~n11932 ;
  assign n11934 = n11933 ^ n11929 ;
  assign n11935 = x1118 ^ x709 ;
  assign n11938 = n9134 & ~n11935 ;
  assign n11939 = n11938 ^ x709 ;
  assign n11940 = ~x962 & ~n11939 ;
  assign n11941 = x1106 ^ x710 ;
  assign n11944 = n9135 & n11941 ;
  assign n11945 = n11944 ^ x710 ;
  assign n11946 = ~x962 & n11945 ;
  assign n11947 = n9371 ^ x373 ;
  assign n11948 = n11947 ^ x398 ;
  assign n11949 = n11948 ^ n9371 ;
  assign n11950 = ~x592 & n11949 ;
  assign n11951 = n11950 ^ n11947 ;
  assign n11975 = n11951 ^ x423 ;
  assign n11976 = n11975 ^ n9370 ;
  assign n11953 = n9370 ^ x423 ;
  assign n11956 = n11953 ^ n9371 ;
  assign n11957 = n11956 ^ n4593 ;
  assign n11958 = n11957 ^ n11953 ;
  assign n12023 = n11976 ^ n11958 ;
  assign n12024 = n12023 ^ n9371 ;
  assign n12012 = n12024 ^ n11958 ;
  assign n12013 = n12012 ^ x423 ;
  assign n11991 = ~x423 & ~n11953 ;
  assign n11992 = n12013 ^ n11991 ;
  assign n11971 = n12023 ^ n9370 ;
  assign n11981 = n11971 ^ n11953 ;
  assign n11993 = n11992 ^ n11981 ;
  assign n11994 = n11993 ^ n9370 ;
  assign n11968 = n11951 ^ n4593 ;
  assign n11996 = n11968 ^ n9370 ;
  assign n11997 = ~n11994 & n11996 ;
  assign n12025 = n12024 ^ n9370 ;
  assign n11998 = n12024 ^ n11951 ;
  assign n11999 = n12025 ^ n11998 ;
  assign n12000 = n12024 ^ n12013 ;
  assign n12001 = n12025 ^ n12000 ;
  assign n12002 = ~n11999 & n12001 ;
  assign n12003 = n11997 & n12002 ;
  assign n12004 = n12003 ^ n11991 ;
  assign n12005 = n12004 ^ n8660 ;
  assign n11983 = n12024 ^ n11981 ;
  assign n11985 = n12025 ^ n11983 ;
  assign n12006 = n12005 ^ n11985 ;
  assign n12029 = n12006 ^ x423 ;
  assign n12030 = n12029 ^ n12025 ;
  assign n12031 = n9367 & n12030 ;
  assign n12032 = x348 & n9466 ;
  assign n12033 = n12031 & ~n12032 ;
  assign n12039 = x200 & n7694 ;
  assign n12035 = x1087 ^ x306 ;
  assign n12040 = n12039 ^ n12035 ;
  assign n12041 = ~x199 & n12040 ;
  assign n12042 = n12041 ^ x1087 ;
  assign n12043 = n9457 & ~n12042 ;
  assign n12044 = n12043 ^ n2991 ;
  assign n12045 = ~n12033 & n12044 ;
  assign n5885 = x755 ^ x725 ;
  assign n12046 = ~x1135 & n5885 ;
  assign n12047 = n12046 ^ x725 ;
  assign n12049 = n12047 ^ x630 ;
  assign n12048 = n12047 ^ x647 ;
  assign n12050 = n12049 ^ n12048 ;
  assign n12053 = ~x1135 & n12050 ;
  assign n12054 = n12053 ^ n12048 ;
  assign n12055 = ~x1134 & ~n12054 ;
  assign n12056 = n12055 ^ n12047 ;
  assign n12057 = n10020 & ~n12056 ;
  assign n12058 = n12057 ^ n9472 ;
  assign n12060 = x858 & n10024 ;
  assign n12061 = n12058 & n12060 ;
  assign n12062 = n12061 ^ n12057 ;
  assign n12063 = ~n12045 & ~n12062 ;
  assign n12064 = n9371 ^ x374 ;
  assign n12065 = n12064 ^ x400 ;
  assign n12066 = n12065 ^ n9371 ;
  assign n12067 = ~x592 & n12066 ;
  assign n12068 = n12067 ^ n12064 ;
  assign n12092 = n12068 ^ x425 ;
  assign n12093 = n12092 ^ n9370 ;
  assign n12070 = n9370 ^ x425 ;
  assign n12073 = n12070 ^ n9371 ;
  assign n12074 = n12073 ^ n4593 ;
  assign n12075 = n12074 ^ n12070 ;
  assign n12140 = n12093 ^ n12075 ;
  assign n12141 = n12140 ^ n9371 ;
  assign n12129 = n12141 ^ n12075 ;
  assign n12130 = n12129 ^ x425 ;
  assign n12108 = ~x425 & ~n12070 ;
  assign n12109 = n12130 ^ n12108 ;
  assign n12088 = n12140 ^ n9370 ;
  assign n12098 = n12088 ^ n12070 ;
  assign n12110 = n12109 ^ n12098 ;
  assign n12111 = n12110 ^ n9370 ;
  assign n12085 = n12068 ^ n4593 ;
  assign n12113 = n12085 ^ n9370 ;
  assign n12114 = ~n12111 & n12113 ;
  assign n12142 = n12141 ^ n9370 ;
  assign n12115 = n12141 ^ n12068 ;
  assign n12116 = n12142 ^ n12115 ;
  assign n12117 = n12141 ^ n12130 ;
  assign n12118 = n12142 ^ n12117 ;
  assign n12119 = ~n12116 & n12118 ;
  assign n12120 = n12114 & n12119 ;
  assign n12121 = n12120 ^ n12108 ;
  assign n12122 = n12121 ^ n8660 ;
  assign n12100 = n12141 ^ n12098 ;
  assign n12102 = n12142 ^ n12100 ;
  assign n12123 = n12122 ^ n12102 ;
  assign n12146 = n12123 ^ x425 ;
  assign n12147 = n12146 ^ n12142 ;
  assign n12148 = n9367 & n12147 ;
  assign n12149 = x350 & n9466 ;
  assign n12150 = n12148 & ~n12149 ;
  assign n12156 = x200 & n7644 ;
  assign n12152 = x1035 ^ x298 ;
  assign n12157 = n12156 ^ n12152 ;
  assign n12158 = ~x199 & n12157 ;
  assign n12159 = n12158 ^ x1035 ;
  assign n12160 = n9457 & ~n12159 ;
  assign n12161 = n12160 ^ n2991 ;
  assign n12162 = ~n12150 & n12161 ;
  assign n5897 = x751 ^ x701 ;
  assign n12163 = ~x1135 & n5897 ;
  assign n12164 = n12163 ^ x701 ;
  assign n12166 = n12164 ^ x644 ;
  assign n12165 = n12164 ^ x715 ;
  assign n12167 = n12166 ^ n12165 ;
  assign n12170 = ~x1135 & n12167 ;
  assign n12171 = n12170 ^ n12165 ;
  assign n12172 = ~x1134 & ~n12171 ;
  assign n12173 = n12172 ^ n12164 ;
  assign n12174 = n10020 & ~n12173 ;
  assign n12175 = n12174 ^ n9472 ;
  assign n12177 = x842 & n10024 ;
  assign n12178 = n12175 & n12177 ;
  assign n12179 = n12178 ^ n12174 ;
  assign n12180 = ~n12162 & ~n12179 ;
  assign n12181 = n9371 ^ x371 ;
  assign n12182 = n12181 ^ x396 ;
  assign n12183 = n12182 ^ n9371 ;
  assign n12184 = ~x592 & n12183 ;
  assign n12185 = n12184 ^ n12181 ;
  assign n12209 = n12185 ^ x421 ;
  assign n12210 = n12209 ^ n9370 ;
  assign n12187 = n9370 ^ x421 ;
  assign n12190 = n12187 ^ n9371 ;
  assign n12191 = n12190 ^ n4593 ;
  assign n12192 = n12191 ^ n12187 ;
  assign n12257 = n12210 ^ n12192 ;
  assign n12258 = n12257 ^ n9371 ;
  assign n12246 = n12258 ^ n12192 ;
  assign n12247 = n12246 ^ x421 ;
  assign n12225 = ~x421 & ~n12187 ;
  assign n12226 = n12247 ^ n12225 ;
  assign n12205 = n12257 ^ n9370 ;
  assign n12215 = n12205 ^ n12187 ;
  assign n12227 = n12226 ^ n12215 ;
  assign n12228 = n12227 ^ n9370 ;
  assign n12202 = n12185 ^ n4593 ;
  assign n12230 = n12202 ^ n9370 ;
  assign n12231 = ~n12228 & n12230 ;
  assign n12259 = n12258 ^ n9370 ;
  assign n12232 = n12258 ^ n12185 ;
  assign n12233 = n12259 ^ n12232 ;
  assign n12234 = n12258 ^ n12247 ;
  assign n12235 = n12259 ^ n12234 ;
  assign n12236 = ~n12233 & n12235 ;
  assign n12237 = n12231 & n12236 ;
  assign n12238 = n12237 ^ n12225 ;
  assign n12239 = n12238 ^ n8660 ;
  assign n12217 = n12258 ^ n12215 ;
  assign n12219 = n12259 ^ n12217 ;
  assign n12240 = n12239 ^ n12219 ;
  assign n12263 = n12240 ^ x421 ;
  assign n12264 = n12263 ^ n12259 ;
  assign n12265 = n9367 & n12264 ;
  assign n12266 = x322 & n9466 ;
  assign n12267 = n12265 & ~n12266 ;
  assign n12273 = x200 & n7703 ;
  assign n12269 = x1051 ^ x309 ;
  assign n12274 = n12273 ^ n12269 ;
  assign n12275 = ~x199 & n12274 ;
  assign n12276 = n12275 ^ x1051 ;
  assign n12277 = n9457 & ~n12276 ;
  assign n12278 = n12277 ^ n2991 ;
  assign n12279 = ~n12267 & n12278 ;
  assign n6010 = x756 ^ x734 ;
  assign n12280 = ~x1135 & n6010 ;
  assign n12281 = n12280 ^ x734 ;
  assign n12283 = n12281 ^ x628 ;
  assign n12282 = n12281 ^ x629 ;
  assign n12284 = n12283 ^ n12282 ;
  assign n12287 = x1135 & n12284 ;
  assign n12288 = n12287 ^ n12282 ;
  assign n12289 = ~x1134 & ~n12288 ;
  assign n12290 = n12289 ^ n12281 ;
  assign n12291 = n10020 & ~n12290 ;
  assign n12292 = n12291 ^ n9472 ;
  assign n12294 = x854 & n10024 ;
  assign n12295 = n12292 & n12294 ;
  assign n12296 = n12295 ^ n12291 ;
  assign n12297 = ~n12279 & ~n12296 ;
  assign n12399 = x762 ^ x697 ;
  assign n12400 = ~x1135 & n12399 ;
  assign n12401 = n12400 ^ x697 ;
  assign n12403 = n12401 ^ x653 ;
  assign n12402 = n12401 ^ x693 ;
  assign n12404 = n12403 ^ n12402 ;
  assign n12407 = ~x1135 & ~n12404 ;
  assign n12408 = n12407 ^ n12402 ;
  assign n12409 = ~x1134 & n12408 ;
  assign n12410 = n12409 ^ n12401 ;
  assign n12393 = x867 ^ x816 ;
  assign n12396 = ~x1134 & n12393 ;
  assign n12397 = n12396 ^ x867 ;
  assign n12398 = ~x1135 & n12397 ;
  assign n12411 = n12410 ^ n12398 ;
  assign n12412 = ~x1136 & ~n12411 ;
  assign n12413 = n12412 ^ n12410 ;
  assign n12414 = n9471 & ~n12413 ;
  assign n12299 = n9371 ^ x326 ;
  assign n12300 = n12299 ^ x439 ;
  assign n12301 = n12300 ^ n9371 ;
  assign n12302 = x592 & n12301 ;
  assign n12303 = n12302 ^ n12299 ;
  assign n12327 = n12303 ^ x449 ;
  assign n12328 = n12327 ^ n9370 ;
  assign n12305 = n9370 ^ x449 ;
  assign n12308 = n12305 ^ n9371 ;
  assign n12309 = n12308 ^ n4593 ;
  assign n12310 = n12309 ^ n12305 ;
  assign n12375 = n12328 ^ n12310 ;
  assign n12376 = n12375 ^ n9371 ;
  assign n12364 = n12376 ^ n12310 ;
  assign n12365 = n12364 ^ x449 ;
  assign n12343 = ~x449 & ~n12305 ;
  assign n12344 = n12365 ^ n12343 ;
  assign n12323 = n12375 ^ n9370 ;
  assign n12333 = n12323 ^ n12305 ;
  assign n12345 = n12344 ^ n12333 ;
  assign n12346 = n12345 ^ n9370 ;
  assign n12320 = n12303 ^ n4593 ;
  assign n12348 = n12320 ^ n9370 ;
  assign n12349 = ~n12346 & n12348 ;
  assign n12377 = n12376 ^ n9370 ;
  assign n12350 = n12376 ^ n12303 ;
  assign n12351 = n12377 ^ n12350 ;
  assign n12352 = n12376 ^ n12365 ;
  assign n12353 = n12377 ^ n12352 ;
  assign n12354 = ~n12351 & n12353 ;
  assign n12355 = n12349 & n12354 ;
  assign n12356 = n12355 ^ n12343 ;
  assign n12357 = n12356 ^ n8660 ;
  assign n12335 = n12376 ^ n12333 ;
  assign n12337 = n12377 ^ n12335 ;
  assign n12358 = n12357 ^ n12337 ;
  assign n12381 = n12358 ^ x449 ;
  assign n12382 = n12381 ^ n12377 ;
  assign n12298 = x461 & n9466 ;
  assign n12384 = n12382 ^ n12298 ;
  assign n12415 = n12414 ^ n12384 ;
  assign n12386 = n12384 ^ x1057 ;
  assign n12385 = n12384 ^ n7277 ;
  assign n12387 = n12386 ^ n12385 ;
  assign n12390 = ~x199 & n12387 ;
  assign n12391 = n12390 ^ n12386 ;
  assign n12392 = ~n9367 & ~n12391 ;
  assign n12416 = n12415 ^ n12392 ;
  assign n12417 = n2991 & ~n12416 ;
  assign n12418 = n12417 ^ n12414 ;
  assign n12419 = x1123 ^ x715 ;
  assign n12422 = n9135 & n12419 ;
  assign n12423 = n12422 ^ x715 ;
  assign n12424 = ~x962 & n12423 ;
  assign n12430 = x200 & n7697 ;
  assign n12426 = x1043 ^ x307 ;
  assign n12431 = n12430 ^ n12426 ;
  assign n12432 = ~x199 & n12431 ;
  assign n12433 = n12432 ^ x1043 ;
  assign n12434 = n9457 & ~n12433 ;
  assign n12435 = n12434 ^ n2991 ;
  assign n12437 = x591 ^ x329 ;
  assign n12438 = n12437 ^ n9466 ;
  assign n12436 = x591 ^ x440 ;
  assign n12439 = n12438 ^ n12436 ;
  assign n12440 = n12439 ^ n9466 ;
  assign n12441 = x592 & ~n12440 ;
  assign n12442 = n12441 ^ n12438 ;
  assign n12445 = x349 & n9466 ;
  assign n12443 = n8660 ^ n4593 ;
  assign n12444 = n12443 ^ n12442 ;
  assign n12446 = n12445 ^ n12444 ;
  assign n12454 = ~n12442 & ~n12446 ;
  assign n12455 = n8660 & n12454 ;
  assign n12456 = n12455 ^ n8660 ;
  assign n12448 = n12445 ^ n8660 ;
  assign n12457 = n12456 ^ n12448 ;
  assign n12458 = n9367 & ~n12457 ;
  assign n12459 = n12435 & n12458 ;
  assign n12461 = x454 & ~n9370 ;
  assign n12462 = n12459 & n12461 ;
  assign n12460 = n12459 ^ n12435 ;
  assign n12463 = n12462 ^ n12460 ;
  assign n5720 = x761 ^ x738 ;
  assign n12464 = ~x1135 & n5720 ;
  assign n12465 = n12464 ^ x738 ;
  assign n12467 = n12465 ^ x626 ;
  assign n12466 = n12465 ^ x641 ;
  assign n12468 = n12467 ^ n12466 ;
  assign n12471 = ~x1135 & n12468 ;
  assign n12472 = n12471 ^ n12466 ;
  assign n12473 = ~x1134 & ~n12472 ;
  assign n12474 = n12473 ^ n12465 ;
  assign n12475 = n10020 & ~n12474 ;
  assign n12476 = n12475 ^ n9472 ;
  assign n12484 = x845 & n12476 ;
  assign n12485 = n10024 & n12484 ;
  assign n12486 = n12485 ^ n10024 ;
  assign n12478 = n12475 ^ n10024 ;
  assign n12487 = n12486 ^ n12478 ;
  assign n12488 = ~n12463 & ~n12487 ;
  assign n6082 = x768 ^ x705 ;
  assign n12590 = ~x1135 & ~n6082 ;
  assign n12591 = n12590 ^ x705 ;
  assign n12593 = n12591 ^ x645 ;
  assign n12592 = n12591 ^ x669 ;
  assign n12594 = n12593 ^ n12592 ;
  assign n12597 = ~x1135 & ~n12594 ;
  assign n12598 = n12597 ^ n12592 ;
  assign n12599 = ~x1134 & ~n12598 ;
  assign n12600 = n12599 ^ n12591 ;
  assign n12584 = x839 ^ x800 ;
  assign n12587 = ~x1134 & n12584 ;
  assign n12588 = n12587 ^ x839 ;
  assign n12589 = ~x1135 & n12588 ;
  assign n12601 = n12600 ^ n12589 ;
  assign n12602 = ~x1136 & n12601 ;
  assign n12603 = n12602 ^ n12600 ;
  assign n12604 = n9471 & n12603 ;
  assign n12490 = n9371 ^ x318 ;
  assign n12491 = n12490 ^ x377 ;
  assign n12492 = n12491 ^ n9371 ;
  assign n12493 = x592 & n12492 ;
  assign n12494 = n12493 ^ n12490 ;
  assign n12518 = n12494 ^ x448 ;
  assign n12519 = n12518 ^ n9370 ;
  assign n12496 = n9370 ^ x448 ;
  assign n12499 = n12496 ^ n9371 ;
  assign n12500 = n12499 ^ n4593 ;
  assign n12501 = n12500 ^ n12496 ;
  assign n12566 = n12519 ^ n12501 ;
  assign n12567 = n12566 ^ n9371 ;
  assign n12555 = n12567 ^ n12501 ;
  assign n12556 = n12555 ^ x448 ;
  assign n12534 = ~x448 & ~n12496 ;
  assign n12535 = n12556 ^ n12534 ;
  assign n12514 = n12566 ^ n9370 ;
  assign n12524 = n12514 ^ n12496 ;
  assign n12536 = n12535 ^ n12524 ;
  assign n12537 = n12536 ^ n9370 ;
  assign n12511 = n12494 ^ n4593 ;
  assign n12539 = n12511 ^ n9370 ;
  assign n12540 = ~n12537 & n12539 ;
  assign n12568 = n12567 ^ n9370 ;
  assign n12541 = n12567 ^ n12494 ;
  assign n12542 = n12568 ^ n12541 ;
  assign n12543 = n12567 ^ n12556 ;
  assign n12544 = n12568 ^ n12543 ;
  assign n12545 = ~n12542 & n12544 ;
  assign n12546 = n12540 & n12545 ;
  assign n12547 = n12546 ^ n12534 ;
  assign n12548 = n12547 ^ n8660 ;
  assign n12526 = n12567 ^ n12524 ;
  assign n12528 = n12568 ^ n12526 ;
  assign n12549 = n12548 ^ n12528 ;
  assign n12572 = n12549 ^ x448 ;
  assign n12573 = n12572 ^ n12568 ;
  assign n12489 = x462 & n9466 ;
  assign n12575 = n12573 ^ n12489 ;
  assign n12605 = n12604 ^ n12575 ;
  assign n12577 = n12575 ^ x1074 ;
  assign n12576 = n12575 ^ n7317 ;
  assign n12578 = n12577 ^ n12576 ;
  assign n12581 = ~x199 & n12578 ;
  assign n12582 = n12581 ^ n12577 ;
  assign n12583 = ~n9367 & ~n12582 ;
  assign n12606 = n12605 ^ n12583 ;
  assign n12607 = n2991 & ~n12606 ;
  assign n12608 = n12607 ^ n12604 ;
  assign n12610 = x419 & ~n9370 ;
  assign n12609 = x315 & n9466 ;
  assign n12611 = n12610 ^ n12609 ;
  assign n12612 = n4593 & n8660 ;
  assign n12613 = x394 ^ x369 ;
  assign n12616 = x592 & n12613 ;
  assign n12617 = n12616 ^ x394 ;
  assign n12618 = n9367 & n12617 ;
  assign n12619 = n12612 & n12618 ;
  assign n12620 = n12619 ^ n9367 ;
  assign n12621 = ~n12611 & n12620 ;
  assign n12627 = x200 & n7685 ;
  assign n12623 = x1080 ^ x303 ;
  assign n12628 = n12627 ^ n12623 ;
  assign n12629 = ~x199 & n12628 ;
  assign n12630 = n12629 ^ x1080 ;
  assign n12631 = n9457 & ~n12630 ;
  assign n12632 = n12631 ^ n2991 ;
  assign n12633 = n12621 & n12632 ;
  assign n12634 = n12633 ^ n12632 ;
  assign n5829 = x767 ^ x698 ;
  assign n12635 = ~x1135 & n5829 ;
  assign n12636 = n12635 ^ x698 ;
  assign n12638 = n12636 ^ x608 ;
  assign n12637 = n12636 ^ x625 ;
  assign n12639 = n12638 ^ n12637 ;
  assign n12642 = ~x1135 & n12639 ;
  assign n12643 = n12642 ^ n12637 ;
  assign n12644 = ~x1134 & ~n12643 ;
  assign n12645 = n12644 ^ n12636 ;
  assign n12646 = n10020 & ~n12645 ;
  assign n12647 = n12646 ^ n9472 ;
  assign n12655 = x853 & n12647 ;
  assign n12656 = n10024 & n12655 ;
  assign n12657 = n12656 ^ n10024 ;
  assign n12649 = n12646 ^ n10024 ;
  assign n12658 = n12657 ^ n12649 ;
  assign n12659 = ~n12634 & ~n12658 ;
  assign n5807 = x774 ^ x687 ;
  assign n12761 = ~x1135 & ~n5807 ;
  assign n12762 = n12761 ^ x687 ;
  assign n12764 = n12762 ^ x636 ;
  assign n12763 = n12762 ^ x650 ;
  assign n12765 = n12764 ^ n12763 ;
  assign n12768 = ~x1135 & ~n12765 ;
  assign n12769 = n12768 ^ n12763 ;
  assign n12770 = ~x1134 & ~n12769 ;
  assign n12771 = n12770 ^ n12762 ;
  assign n12755 = x868 ^ x807 ;
  assign n12758 = ~x1134 & n12755 ;
  assign n12759 = n12758 ^ x868 ;
  assign n12760 = ~x1135 & n12759 ;
  assign n12772 = n12771 ^ n12760 ;
  assign n12773 = ~x1136 & n12772 ;
  assign n12774 = n12773 ^ n12771 ;
  assign n12775 = n9471 & n12774 ;
  assign n12661 = n9371 ^ x325 ;
  assign n12662 = n12661 ^ x378 ;
  assign n12663 = n12662 ^ n9371 ;
  assign n12664 = x592 & n12663 ;
  assign n12665 = n12664 ^ n12661 ;
  assign n12689 = n12665 ^ x451 ;
  assign n12690 = n12689 ^ n9370 ;
  assign n12667 = n9370 ^ x451 ;
  assign n12670 = n12667 ^ n9371 ;
  assign n12671 = n12670 ^ n4593 ;
  assign n12672 = n12671 ^ n12667 ;
  assign n12737 = n12690 ^ n12672 ;
  assign n12738 = n12737 ^ n9371 ;
  assign n12726 = n12738 ^ n12672 ;
  assign n12727 = n12726 ^ x451 ;
  assign n12705 = ~x451 & ~n12667 ;
  assign n12706 = n12727 ^ n12705 ;
  assign n12685 = n12737 ^ n9370 ;
  assign n12695 = n12685 ^ n12667 ;
  assign n12707 = n12706 ^ n12695 ;
  assign n12708 = n12707 ^ n9370 ;
  assign n12682 = n12665 ^ n4593 ;
  assign n12710 = n12682 ^ n9370 ;
  assign n12711 = ~n12708 & n12710 ;
  assign n12739 = n12738 ^ n9370 ;
  assign n12712 = n12738 ^ n12665 ;
  assign n12713 = n12739 ^ n12712 ;
  assign n12714 = n12738 ^ n12727 ;
  assign n12715 = n12739 ^ n12714 ;
  assign n12716 = ~n12713 & n12715 ;
  assign n12717 = n12711 & n12716 ;
  assign n12718 = n12717 ^ n12705 ;
  assign n12719 = n12718 ^ n8660 ;
  assign n12697 = n12738 ^ n12695 ;
  assign n12699 = n12739 ^ n12697 ;
  assign n12720 = n12719 ^ n12699 ;
  assign n12743 = n12720 ^ x451 ;
  assign n12744 = n12743 ^ n12739 ;
  assign n12660 = x353 & n9466 ;
  assign n12746 = n12744 ^ n12660 ;
  assign n12776 = n12775 ^ n12746 ;
  assign n12748 = n12746 ^ x1063 ;
  assign n12747 = n12746 ^ n7329 ;
  assign n12749 = n12748 ^ n12747 ;
  assign n12752 = ~x199 & n12749 ;
  assign n12753 = n12752 ^ n12748 ;
  assign n12754 = ~n9367 & ~n12753 ;
  assign n12777 = n12776 ^ n12754 ;
  assign n12778 = n2991 & ~n12777 ;
  assign n12779 = n12778 ^ n12775 ;
  assign n12881 = x750 ^ x684 ;
  assign n12882 = ~x1135 & n12881 ;
  assign n12883 = n12882 ^ x684 ;
  assign n12885 = n12883 ^ x651 ;
  assign n12884 = n12883 ^ x654 ;
  assign n12886 = n12885 ^ n12884 ;
  assign n12889 = ~x1135 & ~n12886 ;
  assign n12890 = n12889 ^ n12884 ;
  assign n12891 = ~x1134 & n12890 ;
  assign n12892 = n12891 ^ n12883 ;
  assign n12875 = x880 ^ x794 ;
  assign n12878 = ~x1134 & n12875 ;
  assign n12879 = n12878 ^ x880 ;
  assign n12880 = ~x1135 & n12879 ;
  assign n12893 = n12892 ^ n12880 ;
  assign n12894 = ~x1136 & ~n12893 ;
  assign n12895 = n12894 ^ n12892 ;
  assign n12896 = n9471 & ~n12895 ;
  assign n12781 = n9371 ^ x381 ;
  assign n12782 = n12781 ^ x405 ;
  assign n12783 = n12782 ^ n9371 ;
  assign n12784 = ~x592 & n12783 ;
  assign n12785 = n12784 ^ n12781 ;
  assign n12809 = n12785 ^ x445 ;
  assign n12810 = n12809 ^ n9370 ;
  assign n12787 = n9370 ^ x445 ;
  assign n12790 = n12787 ^ n9371 ;
  assign n12791 = n12790 ^ n4593 ;
  assign n12792 = n12791 ^ n12787 ;
  assign n12857 = n12810 ^ n12792 ;
  assign n12858 = n12857 ^ n9371 ;
  assign n12846 = n12858 ^ n12792 ;
  assign n12847 = n12846 ^ x445 ;
  assign n12825 = ~x445 & ~n12787 ;
  assign n12826 = n12847 ^ n12825 ;
  assign n12805 = n12857 ^ n9370 ;
  assign n12815 = n12805 ^ n12787 ;
  assign n12827 = n12826 ^ n12815 ;
  assign n12828 = n12827 ^ n9370 ;
  assign n12802 = n12785 ^ n4593 ;
  assign n12830 = n12802 ^ n9370 ;
  assign n12831 = ~n12828 & n12830 ;
  assign n12859 = n12858 ^ n9370 ;
  assign n12832 = n12858 ^ n12785 ;
  assign n12833 = n12859 ^ n12832 ;
  assign n12834 = n12858 ^ n12847 ;
  assign n12835 = n12859 ^ n12834 ;
  assign n12836 = ~n12833 & n12835 ;
  assign n12837 = n12831 & n12836 ;
  assign n12838 = n12837 ^ n12825 ;
  assign n12839 = n12838 ^ n8660 ;
  assign n12817 = n12858 ^ n12815 ;
  assign n12819 = n12859 ^ n12817 ;
  assign n12840 = n12839 ^ n12819 ;
  assign n12863 = n12840 ^ x445 ;
  assign n12864 = n12863 ^ n12859 ;
  assign n12780 = x356 & n9466 ;
  assign n12866 = n12864 ^ n12780 ;
  assign n12897 = n12896 ^ n12866 ;
  assign n12868 = n12866 ^ x1081 ;
  assign n12867 = n12866 ^ n7347 ;
  assign n12869 = n12868 ^ n12867 ;
  assign n12872 = ~x199 & n12869 ;
  assign n12873 = n12872 ^ n12868 ;
  assign n12874 = ~n9367 & ~n12873 ;
  assign n12898 = n12897 ^ n12874 ;
  assign n12899 = n2991 & ~n12898 ;
  assign n12900 = n12899 ^ n12896 ;
  assign n12901 = x798 ^ x765 ;
  assign n12902 = x800 ^ x771 ;
  assign n12903 = ~n12901 & ~n12902 ;
  assign n12904 = x807 ^ x747 ;
  assign n12905 = x816 ^ x775 ;
  assign n12906 = ~n12904 & ~n12905 ;
  assign n12907 = n12903 & n12906 ;
  assign n12908 = x794 ^ x769 ;
  assign n12909 = x801 ^ x773 ;
  assign n12910 = ~n12908 & ~n12909 ;
  assign n12911 = x813 ^ x721 ;
  assign n12912 = x795 ^ x731 ;
  assign n12913 = ~n12911 & ~n12912 ;
  assign n12914 = n12910 & n12913 ;
  assign n12915 = n12907 & n12914 ;
  assign n12916 = x747 & x773 ;
  assign n12917 = x731 & ~x945 ;
  assign n12918 = n12916 & n12917 ;
  assign n12919 = x775 & x988 ;
  assign n12920 = n12918 & n12919 ;
  assign n12925 = x769 & n12920 ;
  assign n12926 = n12925 ^ x721 ;
  assign n12927 = ~n12915 & n12926 ;
  assign n12928 = n9371 ^ x379 ;
  assign n12929 = n12928 ^ x403 ;
  assign n12930 = n12929 ^ n9371 ;
  assign n12931 = ~x592 & n12930 ;
  assign n12932 = n12931 ^ n12928 ;
  assign n12956 = n12932 ^ x428 ;
  assign n12957 = n12956 ^ n9370 ;
  assign n12934 = n9370 ^ x428 ;
  assign n12937 = n12934 ^ n9371 ;
  assign n12938 = n12937 ^ n4593 ;
  assign n12939 = n12938 ^ n12934 ;
  assign n13004 = n12957 ^ n12939 ;
  assign n13005 = n13004 ^ n9371 ;
  assign n12993 = n13005 ^ n12939 ;
  assign n12994 = n12993 ^ x428 ;
  assign n12972 = ~x428 & ~n12934 ;
  assign n12973 = n12994 ^ n12972 ;
  assign n12952 = n13004 ^ n9370 ;
  assign n12962 = n12952 ^ n12934 ;
  assign n12974 = n12973 ^ n12962 ;
  assign n12975 = n12974 ^ n9370 ;
  assign n12949 = n12932 ^ n4593 ;
  assign n12977 = n12949 ^ n9370 ;
  assign n12978 = ~n12975 & n12977 ;
  assign n13006 = n13005 ^ n9370 ;
  assign n12979 = n13005 ^ n12932 ;
  assign n12980 = n13006 ^ n12979 ;
  assign n12981 = n13005 ^ n12994 ;
  assign n12982 = n13006 ^ n12981 ;
  assign n12983 = ~n12980 & n12982 ;
  assign n12984 = n12978 & n12983 ;
  assign n12985 = n12984 ^ n12972 ;
  assign n12986 = n12985 ^ n8660 ;
  assign n12964 = n13005 ^ n12962 ;
  assign n12966 = n13006 ^ n12964 ;
  assign n12987 = n12986 ^ n12966 ;
  assign n13010 = n12987 ^ x428 ;
  assign n13011 = n13010 ^ n13006 ;
  assign n13012 = n9367 & n13011 ;
  assign n13013 = x354 & n9466 ;
  assign n13014 = n13012 & ~n13013 ;
  assign n13015 = n7335 ^ x1045 ;
  assign n13018 = ~x199 & n13015 ;
  assign n13019 = n13018 ^ x1045 ;
  assign n13020 = n9457 & ~n13019 ;
  assign n13021 = n13020 ^ n2991 ;
  assign n13022 = ~n13014 & n13021 ;
  assign n13029 = x776 ^ x694 ;
  assign n13030 = ~x1135 & n13029 ;
  assign n13031 = n13030 ^ x694 ;
  assign n13033 = n13031 ^ x640 ;
  assign n13032 = n13031 ^ x732 ;
  assign n13034 = n13033 ^ n13032 ;
  assign n13037 = ~x1135 & ~n13034 ;
  assign n13038 = n13037 ^ n13032 ;
  assign n13039 = ~x1134 & n13038 ;
  assign n13040 = n13039 ^ n13031 ;
  assign n13023 = x851 ^ x795 ;
  assign n13026 = ~x1134 & n13023 ;
  assign n13027 = n13026 ^ x851 ;
  assign n13028 = ~x1135 & n13027 ;
  assign n13041 = n13040 ^ n13028 ;
  assign n13042 = ~x1136 & ~n13041 ;
  assign n13043 = n13042 ^ n13040 ;
  assign n13044 = n9472 & ~n13043 ;
  assign n13045 = ~n13022 & ~n13044 ;
  assign n13046 = x1111 ^ x723 ;
  assign n13049 = n9134 & ~n13046 ;
  assign n13050 = n13049 ^ x723 ;
  assign n13051 = ~x962 & ~n13050 ;
  assign n13052 = x1114 ^ x724 ;
  assign n13055 = n9134 & ~n13052 ;
  assign n13056 = n13055 ^ x724 ;
  assign n13057 = ~x962 & ~n13056 ;
  assign n13058 = x1120 ^ x725 ;
  assign n13061 = n9134 & ~n13058 ;
  assign n13062 = n13061 ^ x725 ;
  assign n13063 = ~x962 & ~n13062 ;
  assign n13064 = x1126 ^ x726 ;
  assign n13067 = n9134 & n13064 ;
  assign n13068 = n13067 ^ x726 ;
  assign n13069 = ~x962 & n13068 ;
  assign n13070 = x1102 ^ x727 ;
  assign n13073 = n9134 & n13070 ;
  assign n13074 = n13073 ^ x727 ;
  assign n13075 = ~x962 & n13074 ;
  assign n13076 = x1131 ^ x728 ;
  assign n13079 = n9134 & ~n13076 ;
  assign n13080 = n13079 ^ x728 ;
  assign n13081 = ~x962 & ~n13080 ;
  assign n13082 = x1104 ^ x729 ;
  assign n13085 = n9134 & n13082 ;
  assign n13086 = n13085 ^ x729 ;
  assign n13087 = ~x962 & n13086 ;
  assign n13088 = x1106 ^ x730 ;
  assign n13091 = n9134 & n13088 ;
  assign n13092 = n13091 ^ x730 ;
  assign n13093 = ~x962 & n13092 ;
  assign n13094 = ~x945 & x988 ;
  assign n13099 = n12916 & n13094 ;
  assign n13100 = n13099 ^ x731 ;
  assign n13101 = ~n12915 & n13100 ;
  assign n13102 = x1128 ^ x732 ;
  assign n13105 = n9135 & ~n13102 ;
  assign n13106 = n13105 ^ x732 ;
  assign n13107 = ~x962 & ~n13106 ;
  assign n13132 = n9371 ^ x375 ;
  assign n13133 = n13132 ^ x399 ;
  assign n13134 = n13133 ^ n9371 ;
  assign n13135 = ~x592 & n13134 ;
  assign n13136 = n13135 ^ n13132 ;
  assign n13160 = n13136 ^ x424 ;
  assign n13161 = n13160 ^ n9370 ;
  assign n13138 = n9370 ^ x424 ;
  assign n13141 = n13138 ^ n9371 ;
  assign n13142 = n13141 ^ n4593 ;
  assign n13143 = n13142 ^ n13138 ;
  assign n13208 = n13161 ^ n13143 ;
  assign n13209 = n13208 ^ n9371 ;
  assign n13197 = n13209 ^ n13143 ;
  assign n13198 = n13197 ^ x424 ;
  assign n13176 = ~x424 & ~n13138 ;
  assign n13177 = n13198 ^ n13176 ;
  assign n13156 = n13208 ^ n9370 ;
  assign n13166 = n13156 ^ n13138 ;
  assign n13178 = n13177 ^ n13166 ;
  assign n13179 = n13178 ^ n9370 ;
  assign n13153 = n13136 ^ n4593 ;
  assign n13181 = n13153 ^ n9370 ;
  assign n13182 = ~n13179 & n13181 ;
  assign n13210 = n13209 ^ n9370 ;
  assign n13183 = n13209 ^ n13136 ;
  assign n13184 = n13210 ^ n13183 ;
  assign n13185 = n13209 ^ n13198 ;
  assign n13186 = n13210 ^ n13185 ;
  assign n13187 = ~n13184 & n13186 ;
  assign n13188 = n13182 & n13187 ;
  assign n13189 = n13188 ^ n13176 ;
  assign n13190 = n13189 ^ n8660 ;
  assign n13168 = n13209 ^ n13166 ;
  assign n13170 = n13210 ^ n13168 ;
  assign n13191 = n13190 ^ n13170 ;
  assign n13214 = n13191 ^ x424 ;
  assign n13215 = n13214 ^ n13210 ;
  assign n13131 = x316 & n9466 ;
  assign n13217 = n13215 ^ n13131 ;
  assign n13218 = n13217 ^ x1047 ;
  assign n13128 = x200 & n7700 ;
  assign n13124 = x1047 ^ x308 ;
  assign n13129 = n13128 ^ n13124 ;
  assign n13130 = ~x199 & n13129 ;
  assign n13219 = n13218 ^ n13130 ;
  assign n13220 = ~n9367 & ~n13219 ;
  assign n13221 = n13220 ^ n13217 ;
  assign n6039 = x777 ^ x737 ;
  assign n13108 = ~x1135 & n6039 ;
  assign n13109 = n13108 ^ x737 ;
  assign n13111 = n13109 ^ x619 ;
  assign n13110 = n13109 ^ x648 ;
  assign n13112 = n13111 ^ n13110 ;
  assign n13115 = ~x1135 & n13112 ;
  assign n13116 = n13115 ^ n13110 ;
  assign n13117 = ~x1134 & ~n13116 ;
  assign n13118 = n13117 ^ n13109 ;
  assign n13119 = n10816 & ~n13118 ;
  assign n13223 = n13221 ^ n13119 ;
  assign n13120 = n13119 ^ n9471 ;
  assign n13121 = x838 & n10024 ;
  assign n13122 = n13120 & n13121 ;
  assign n13224 = n13223 ^ n13122 ;
  assign n13225 = ~n2991 & ~n13224 ;
  assign n13226 = n13225 ^ n13221 ;
  assign n13227 = x1119 ^ x734 ;
  assign n13230 = n9134 & ~n13227 ;
  assign n13231 = n13230 ^ x734 ;
  assign n13232 = ~x962 & ~n13231 ;
  assign n13233 = x1109 ^ x735 ;
  assign n13236 = n9134 & n13233 ;
  assign n13237 = n13236 ^ x735 ;
  assign n13238 = ~x962 & n13237 ;
  assign n13239 = x1101 ^ x736 ;
  assign n13242 = n9134 & n13239 ;
  assign n13243 = n13242 ^ x736 ;
  assign n13244 = ~x962 & n13243 ;
  assign n13245 = x1122 ^ x737 ;
  assign n13248 = n9134 & ~n13245 ;
  assign n13249 = n13248 ^ x737 ;
  assign n13250 = ~x962 & ~n13249 ;
  assign n13251 = x1121 ^ x738 ;
  assign n13254 = n9134 & ~n13251 ;
  assign n13255 = n13254 ^ x738 ;
  assign n13256 = ~x962 & ~n13255 ;
  assign n13257 = x1108 ^ x739 ;
  assign n13260 = n8917 & n13257 ;
  assign n13261 = n13260 ^ x739 ;
  assign n13262 = ~x966 & ~n13261 ;
  assign n13263 = x1114 ^ x741 ;
  assign n13266 = n8917 & ~n13263 ;
  assign n13267 = n13266 ^ x741 ;
  assign n13268 = ~x966 & n13267 ;
  assign n13269 = x1112 ^ x742 ;
  assign n13272 = n8917 & ~n13269 ;
  assign n13273 = n13272 ^ x742 ;
  assign n13274 = ~x966 & n13273 ;
  assign n13275 = x1109 ^ x743 ;
  assign n13278 = n8917 & n13275 ;
  assign n13279 = n13278 ^ x743 ;
  assign n13280 = ~x966 & ~n13279 ;
  assign n13281 = x1131 ^ x744 ;
  assign n13284 = n8917 & ~n13281 ;
  assign n13285 = n13284 ^ x744 ;
  assign n13286 = ~x966 & n13285 ;
  assign n13287 = x1111 ^ x745 ;
  assign n13290 = n8917 & ~n13287 ;
  assign n13291 = n13290 ^ x745 ;
  assign n13292 = ~x966 & n13291 ;
  assign n13293 = x1104 ^ x746 ;
  assign n13296 = n8917 & n13293 ;
  assign n13297 = n13296 ^ x746 ;
  assign n13298 = ~x966 & ~n13297 ;
  assign n13303 = x773 & n13094 ;
  assign n13304 = n13303 ^ x747 ;
  assign n13305 = ~n12915 & n13304 ;
  assign n13306 = x1106 ^ x748 ;
  assign n13309 = n8917 & n13306 ;
  assign n13310 = n13309 ^ x748 ;
  assign n13311 = ~x966 & ~n13310 ;
  assign n13312 = x1105 ^ x749 ;
  assign n13315 = n8917 & n13312 ;
  assign n13316 = n13315 ^ x749 ;
  assign n13317 = ~x966 & ~n13316 ;
  assign n13318 = x1130 ^ x750 ;
  assign n13321 = n8917 & ~n13318 ;
  assign n13322 = n13321 ^ x750 ;
  assign n13323 = ~x966 & n13322 ;
  assign n13324 = x1123 ^ x751 ;
  assign n13327 = n8917 & ~n13324 ;
  assign n13328 = n13327 ^ x751 ;
  assign n13329 = ~x966 & n13328 ;
  assign n13330 = x1124 ^ x752 ;
  assign n13333 = n8917 & ~n13330 ;
  assign n13334 = n13333 ^ x752 ;
  assign n13335 = ~x966 & n13334 ;
  assign n13336 = x1117 ^ x753 ;
  assign n13339 = n8917 & ~n13336 ;
  assign n13340 = n13339 ^ x753 ;
  assign n13341 = ~x966 & n13340 ;
  assign n13342 = x1118 ^ x754 ;
  assign n13345 = n8917 & ~n13342 ;
  assign n13346 = n13345 ^ x754 ;
  assign n13347 = ~x966 & n13346 ;
  assign n13348 = x1120 ^ x755 ;
  assign n13351 = n8917 & ~n13348 ;
  assign n13352 = n13351 ^ x755 ;
  assign n13353 = ~x966 & n13352 ;
  assign n13354 = x1119 ^ x756 ;
  assign n13357 = n8917 & ~n13354 ;
  assign n13358 = n13357 ^ x756 ;
  assign n13359 = ~x966 & n13358 ;
  assign n13360 = x1113 ^ x757 ;
  assign n13363 = n8917 & ~n13360 ;
  assign n13364 = n13363 ^ x757 ;
  assign n13365 = ~x966 & n13364 ;
  assign n13366 = x1101 ^ x758 ;
  assign n13369 = n8917 & n13366 ;
  assign n13370 = n13369 ^ x758 ;
  assign n13371 = ~x966 & ~n13370 ;
  assign n13372 = x1100 ^ x759 ;
  assign n13375 = n8917 & n13372 ;
  assign n13376 = n13375 ^ x759 ;
  assign n13377 = ~x966 & ~n13376 ;
  assign n13378 = x1115 ^ x760 ;
  assign n13381 = n8917 & ~n13378 ;
  assign n13382 = n13381 ^ x760 ;
  assign n13383 = ~x966 & n13382 ;
  assign n13384 = x1121 ^ x761 ;
  assign n13387 = n8917 & ~n13384 ;
  assign n13388 = n13387 ^ x761 ;
  assign n13389 = ~x966 & n13388 ;
  assign n13390 = x1129 ^ x762 ;
  assign n13393 = n8917 & ~n13390 ;
  assign n13394 = n13393 ^ x762 ;
  assign n13395 = ~x966 & n13394 ;
  assign n13396 = x1103 ^ x763 ;
  assign n13399 = n8917 & n13396 ;
  assign n13400 = n13399 ^ x763 ;
  assign n13401 = ~x966 & ~n13400 ;
  assign n13402 = x1107 ^ x764 ;
  assign n13405 = n8917 & n13402 ;
  assign n13406 = n13405 ^ x764 ;
  assign n13407 = ~x966 & ~n13406 ;
  assign n13408 = ~x773 & ~x794 ;
  assign n13409 = ~x795 & ~x816 ;
  assign n13410 = n13408 & n13409 ;
  assign n13411 = ~x721 & ~x747 ;
  assign n13413 = x765 & x771 ;
  assign n13412 = x771 ^ x765 ;
  assign n13414 = n13413 ^ n13412 ;
  assign n13415 = n13411 & ~n13414 ;
  assign n13416 = n13410 & n13415 ;
  assign n13417 = n12915 & ~n13416 ;
  assign n13418 = x945 ^ x765 ;
  assign n13419 = ~n13417 & ~n13418 ;
  assign n13420 = x1110 ^ x766 ;
  assign n13423 = n8917 & n13420 ;
  assign n13424 = n13423 ^ x766 ;
  assign n13425 = ~x966 & ~n13424 ;
  assign n13426 = x1116 ^ x767 ;
  assign n13429 = n8917 & ~n13426 ;
  assign n13430 = n13429 ^ x767 ;
  assign n13431 = ~x966 & n13430 ;
  assign n13432 = x1125 ^ x768 ;
  assign n13435 = n8917 & ~n13432 ;
  assign n13436 = n13435 ^ x768 ;
  assign n13437 = ~x966 & n13436 ;
  assign n13438 = n12920 ^ x769 ;
  assign n13439 = ~n12915 & n13438 ;
  assign n13440 = x1126 ^ x770 ;
  assign n13443 = n8917 & ~n13440 ;
  assign n13444 = n13443 ^ x770 ;
  assign n13445 = ~x966 & n13444 ;
  assign n13446 = x987 ^ x771 ;
  assign n13447 = ~x945 & n13446 ;
  assign n13448 = n13447 ^ x771 ;
  assign n13449 = ~n13417 & n13448 ;
  assign n13450 = x1102 ^ x772 ;
  assign n13453 = n8917 & n13450 ;
  assign n13454 = n13453 ^ x772 ;
  assign n13455 = ~x966 & ~n13454 ;
  assign n13456 = n13094 ^ x773 ;
  assign n13457 = ~n13417 & n13456 ;
  assign n13458 = x1127 ^ x774 ;
  assign n13461 = n8917 & ~n13458 ;
  assign n13462 = n13461 ^ x774 ;
  assign n13463 = ~x966 & n13462 ;
  assign n13468 = n12918 & n13413 ;
  assign n13469 = n13468 ^ x775 ;
  assign n13470 = ~n12915 & n13469 ;
  assign n13471 = x1128 ^ x776 ;
  assign n13474 = n8917 & ~n13471 ;
  assign n13475 = n13474 ^ x776 ;
  assign n13476 = ~x966 & n13475 ;
  assign n13477 = x1122 ^ x777 ;
  assign n13480 = n8917 & ~n13477 ;
  assign n13481 = n13480 ^ x777 ;
  assign n13482 = ~x966 & n13481 ;
  assign n13483 = x1100 ^ x778 ;
  assign n13484 = x832 & x956 ;
  assign n13485 = ~x1083 & x1085 ;
  assign n13486 = n13484 & n13485 ;
  assign n13487 = ~x1046 & n13486 ;
  assign n13488 = x968 & n13487 ;
  assign n13489 = n13488 ^ n13487 ;
  assign n13490 = n13483 & n13489 ;
  assign n13491 = n13490 ^ x778 ;
  assign n13492 = x779 & ~n9001 ;
  assign n13493 = x780 & ~n8826 ;
  assign n13494 = x1101 ^ x781 ;
  assign n13495 = n13489 & n13494 ;
  assign n13496 = n13495 ^ x781 ;
  assign n13497 = ~n2630 & ~n8931 ;
  assign n13498 = ~n8825 & n13497 ;
  assign n13499 = x1109 ^ x783 ;
  assign n13500 = n13489 & n13499 ;
  assign n13501 = n13500 ^ x783 ;
  assign n13502 = x1110 ^ x784 ;
  assign n13503 = n13489 & n13502 ;
  assign n13504 = n13503 ^ x784 ;
  assign n13505 = x1102 ^ x785 ;
  assign n13506 = n13489 & n13505 ;
  assign n13507 = n13506 ^ x785 ;
  assign n13508 = x786 ^ x24 ;
  assign n13509 = x954 & n13508 ;
  assign n13510 = n13509 ^ x24 ;
  assign n13511 = x1104 ^ x787 ;
  assign n13512 = n13489 & n13511 ;
  assign n13513 = n13512 ^ x787 ;
  assign n13514 = x1105 ^ x788 ;
  assign n13515 = n13489 & n13514 ;
  assign n13516 = n13515 ^ x788 ;
  assign n13517 = x1106 ^ x789 ;
  assign n13518 = n13489 & n13517 ;
  assign n13519 = n13518 ^ x789 ;
  assign n13520 = x1107 ^ x790 ;
  assign n13521 = n13489 & n13520 ;
  assign n13522 = n13521 ^ x790 ;
  assign n13523 = x1108 ^ x791 ;
  assign n13524 = n13489 & n13523 ;
  assign n13525 = n13524 ^ x791 ;
  assign n13526 = x1103 ^ x792 ;
  assign n13527 = n13489 & n13526 ;
  assign n13528 = n13527 ^ x792 ;
  assign n13529 = x1130 ^ x794 ;
  assign n13530 = n13488 & n13529 ;
  assign n13531 = n13530 ^ x794 ;
  assign n13532 = x1128 ^ x795 ;
  assign n13533 = n13488 & n13532 ;
  assign n13534 = n13533 ^ x795 ;
  assign n13535 = x266 & ~x269 ;
  assign n13536 = x279 & n13535 ;
  assign n13537 = x278 & ~x280 ;
  assign n13538 = n13536 & n13537 ;
  assign n13539 = n9342 & n9344 ;
  assign n13540 = n13538 & n13539 ;
  assign n13541 = n13540 ^ x264 ;
  assign n13542 = x1124 ^ x798 ;
  assign n13543 = n13488 & n13542 ;
  assign n13544 = n13543 ^ x798 ;
  assign n13545 = x1107 ^ x799 ;
  assign n13546 = n13488 & ~n13545 ;
  assign n13547 = n13546 ^ x799 ;
  assign n13548 = x1125 ^ x800 ;
  assign n13549 = n13488 & n13548 ;
  assign n13550 = n13549 ^ x800 ;
  assign n13551 = x1126 ^ x801 ;
  assign n13552 = n13488 & n13551 ;
  assign n13553 = n13552 ^ x801 ;
  assign n13554 = ~x274 & n9347 ;
  assign n13555 = x1106 ^ x803 ;
  assign n13556 = n13488 & ~n13555 ;
  assign n13557 = n13556 ^ x803 ;
  assign n13558 = x1109 ^ x804 ;
  assign n13559 = n13488 & n13558 ;
  assign n13560 = n13559 ^ x804 ;
  assign n13561 = n9343 ^ x270 ;
  assign n13562 = x1127 ^ x807 ;
  assign n13563 = n13488 & n13562 ;
  assign n13564 = n13563 ^ x807 ;
  assign n13565 = x1101 ^ x808 ;
  assign n13566 = n13488 & n13565 ;
  assign n13567 = n13566 ^ x808 ;
  assign n13568 = x1103 ^ x809 ;
  assign n13569 = n13488 & ~n13568 ;
  assign n13570 = n13569 ^ x809 ;
  assign n13571 = x1108 ^ x810 ;
  assign n13572 = n13488 & n13571 ;
  assign n13573 = n13572 ^ x810 ;
  assign n13574 = x1102 ^ x811 ;
  assign n13575 = n13488 & n13574 ;
  assign n13576 = n13575 ^ x811 ;
  assign n13577 = x1104 ^ x812 ;
  assign n13578 = n13488 & ~n13577 ;
  assign n13579 = n13578 ^ x812 ;
  assign n13580 = x1131 ^ x813 ;
  assign n13581 = n13488 & n13580 ;
  assign n13582 = n13581 ^ x813 ;
  assign n13583 = x1105 ^ x814 ;
  assign n13584 = n13488 & ~n13583 ;
  assign n13585 = n13584 ^ x814 ;
  assign n13586 = x1110 ^ x815 ;
  assign n13587 = n13488 & n13586 ;
  assign n13588 = n13587 ^ x815 ;
  assign n13589 = x1129 ^ x816 ;
  assign n13590 = n13488 & n13589 ;
  assign n13591 = n13590 ^ x816 ;
  assign n13592 = n9340 ^ x269 ;
  assign n13593 = n9346 ^ x265 ;
  assign n13594 = ~x270 & n9343 ;
  assign n13595 = n13594 ^ x277 ;
  assign n13596 = ~x811 & ~x893 ;
  assign n13597 = n1564 & n1567 ;
  assign n13598 = n2991 & n13597 ;
  assign n13599 = n13598 ^ n1564 ;
  assign n13601 = ~x982 & ~n1569 ;
  assign n13602 = n13599 & n13601 ;
  assign n13603 = n13602 ^ n13598 ;
  assign n13604 = ~x222 & n9367 ;
  assign n13605 = x123 & n13604 ;
  assign n13610 = x1131 ^ x1130 ;
  assign n13609 = x1129 ^ x1128 ;
  assign n13611 = n13610 ^ n13609 ;
  assign n13607 = x1125 ^ x1124 ;
  assign n13606 = x1127 ^ x1126 ;
  assign n13608 = n13607 ^ n13606 ;
  assign n13612 = n13611 ^ n13608 ;
  assign n13613 = n13612 ^ x825 ;
  assign n13614 = ~n13605 & ~n13613 ;
  assign n13615 = n13614 ^ x825 ;
  assign n13620 = x1123 ^ x1122 ;
  assign n13619 = x1121 ^ x1120 ;
  assign n13621 = n13620 ^ n13619 ;
  assign n13617 = x1117 ^ x1116 ;
  assign n13616 = x1119 ^ x1118 ;
  assign n13618 = n13617 ^ n13616 ;
  assign n13622 = n13621 ^ n13618 ;
  assign n13623 = n13622 ^ x826 ;
  assign n13624 = ~n13605 & ~n13623 ;
  assign n13625 = n13624 ^ x826 ;
  assign n13630 = x1107 ^ x1106 ;
  assign n13629 = x1105 ^ x1104 ;
  assign n13631 = n13630 ^ n13629 ;
  assign n13627 = x1103 ^ x1102 ;
  assign n13626 = x1101 ^ x1100 ;
  assign n13628 = n13627 ^ n13626 ;
  assign n13632 = n13631 ^ n13628 ;
  assign n13633 = n13632 ^ x827 ;
  assign n13634 = ~n13605 & ~n13633 ;
  assign n13635 = n13634 ^ x827 ;
  assign n13640 = x1109 ^ x1108 ;
  assign n13639 = x1111 ^ x1110 ;
  assign n13641 = n13640 ^ n13639 ;
  assign n13637 = x1113 ^ x1112 ;
  assign n13636 = x1115 ^ x1114 ;
  assign n13638 = n13637 ^ n13636 ;
  assign n13642 = n13641 ^ n13638 ;
  assign n13643 = n13642 ^ x828 ;
  assign n13644 = ~n13605 & ~n13643 ;
  assign n13645 = n13644 ^ x828 ;
  assign n13646 = n2991 & n7783 ;
  assign n13647 = ~x951 & x1092 ;
  assign n13648 = ~n13646 & n13647 ;
  assign n13649 = n13648 ^ n13646 ;
  assign n13650 = n13538 ^ x281 ;
  assign n13651 = ~x832 & ~x1163 ;
  assign n13652 = n2989 & n13651 ;
  assign n13653 = n7783 & n13652 ;
  assign n13654 = x1091 ^ x833 ;
  assign n13655 = n2985 & n13654 ;
  assign n13656 = n13655 ^ x833 ;
  assign n13657 = x946 & n2985 ;
  assign n13658 = ~x281 & n9341 ;
  assign n13659 = n13658 ^ x282 ;
  assign n13660 = x1049 ^ x837 ;
  assign n13661 = ~x955 & n13660 ;
  assign n13662 = n13661 ^ x837 ;
  assign n13663 = x1047 ^ x838 ;
  assign n13664 = ~x955 & n13663 ;
  assign n13665 = n13664 ^ x838 ;
  assign n13666 = x1074 ^ x839 ;
  assign n13667 = ~x955 & n13666 ;
  assign n13668 = n13667 ^ x839 ;
  assign n13669 = x1196 ^ x840 ;
  assign n13670 = n2985 & n13669 ;
  assign n13671 = n13670 ^ x840 ;
  assign n13672 = n3494 & n5601 ;
  assign n13673 = x1035 ^ x842 ;
  assign n13674 = ~x955 & n13673 ;
  assign n13675 = n13674 ^ x842 ;
  assign n13676 = x1079 ^ x843 ;
  assign n13677 = ~x955 & n13676 ;
  assign n13678 = n13677 ^ x843 ;
  assign n13679 = x1078 ^ x844 ;
  assign n13680 = ~x955 & n13679 ;
  assign n13681 = n13680 ^ x844 ;
  assign n13682 = x1043 ^ x845 ;
  assign n13683 = ~x955 & n13682 ;
  assign n13684 = n13683 ^ x845 ;
  assign n13685 = x1134 ^ x846 ;
  assign n13686 = ~n7353 & n13685 ;
  assign n13687 = n13686 ^ x846 ;
  assign n13688 = x1055 ^ x847 ;
  assign n13689 = ~x955 & n13688 ;
  assign n13690 = n13689 ^ x847 ;
  assign n13691 = x1039 ^ x848 ;
  assign n13692 = ~x955 & n13691 ;
  assign n13693 = n13692 ^ x848 ;
  assign n13694 = x1198 ^ x849 ;
  assign n13695 = n2985 & n13694 ;
  assign n13696 = n13695 ^ x849 ;
  assign n13697 = x1048 ^ x850 ;
  assign n13698 = ~x955 & n13697 ;
  assign n13699 = n13698 ^ x850 ;
  assign n13700 = x1045 ^ x851 ;
  assign n13701 = ~x955 & n13700 ;
  assign n13702 = n13701 ^ x851 ;
  assign n13703 = x1062 ^ x852 ;
  assign n13704 = ~x955 & n13703 ;
  assign n13705 = n13704 ^ x852 ;
  assign n13706 = x1080 ^ x853 ;
  assign n13707 = ~x955 & n13706 ;
  assign n13708 = n13707 ^ x853 ;
  assign n13709 = x1051 ^ x854 ;
  assign n13710 = ~x955 & n13709 ;
  assign n13711 = n13710 ^ x854 ;
  assign n13712 = x1065 ^ x855 ;
  assign n13713 = ~x955 & n13712 ;
  assign n13714 = n13713 ^ x855 ;
  assign n13715 = x1067 ^ x856 ;
  assign n13716 = ~x955 & n13715 ;
  assign n13717 = n13716 ^ x856 ;
  assign n13718 = x1058 ^ x857 ;
  assign n13719 = ~x955 & n13718 ;
  assign n13720 = n13719 ^ x857 ;
  assign n13721 = x1087 ^ x858 ;
  assign n13722 = ~x955 & n13721 ;
  assign n13723 = n13722 ^ x858 ;
  assign n13724 = x1070 ^ x859 ;
  assign n13725 = ~x955 & n13724 ;
  assign n13726 = n13725 ^ x859 ;
  assign n13727 = x1076 ^ x860 ;
  assign n13728 = ~x955 & n13727 ;
  assign n13729 = n13728 ^ x860 ;
  assign n13730 = x1141 ^ x861 ;
  assign n13731 = ~n7353 & n13730 ;
  assign n13732 = n13731 ^ x861 ;
  assign n13733 = x1139 ^ x862 ;
  assign n13734 = ~n7353 & n13733 ;
  assign n13735 = n13734 ^ x862 ;
  assign n13736 = x1199 ^ x863 ;
  assign n13737 = n2985 & n13736 ;
  assign n13738 = n13737 ^ x863 ;
  assign n13739 = x1197 ^ x864 ;
  assign n13740 = n2985 & n13739 ;
  assign n13741 = n13740 ^ x864 ;
  assign n13742 = x1040 ^ x865 ;
  assign n13743 = ~x955 & n13742 ;
  assign n13744 = n13743 ^ x865 ;
  assign n13745 = x1053 ^ x866 ;
  assign n13746 = ~x955 & n13745 ;
  assign n13747 = n13746 ^ x866 ;
  assign n13748 = x1057 ^ x867 ;
  assign n13749 = ~x955 & n13748 ;
  assign n13750 = n13749 ^ x867 ;
  assign n13751 = x1063 ^ x868 ;
  assign n13752 = ~x955 & n13751 ;
  assign n13753 = n13752 ^ x868 ;
  assign n13754 = x1140 ^ x869 ;
  assign n13755 = ~n7353 & n13754 ;
  assign n13756 = n13755 ^ x869 ;
  assign n13757 = x1069 ^ x870 ;
  assign n13758 = ~x955 & n13757 ;
  assign n13759 = n13758 ^ x870 ;
  assign n13760 = x1072 ^ x871 ;
  assign n13761 = ~x955 & n13760 ;
  assign n13762 = n13761 ^ x871 ;
  assign n13763 = x1084 ^ x872 ;
  assign n13764 = ~x955 & n13763 ;
  assign n13765 = n13764 ^ x872 ;
  assign n13766 = x1044 ^ x873 ;
  assign n13767 = ~x955 & n13766 ;
  assign n13768 = n13767 ^ x873 ;
  assign n13769 = x1036 ^ x874 ;
  assign n13770 = ~x955 & n13769 ;
  assign n13771 = n13770 ^ x874 ;
  assign n13772 = x1136 ^ x875 ;
  assign n13773 = ~n7353 & n13772 ;
  assign n13774 = n13773 ^ x875 ;
  assign n13775 = x1037 ^ x876 ;
  assign n13776 = ~x955 & n13775 ;
  assign n13777 = n13776 ^ x876 ;
  assign n13778 = x1138 ^ x877 ;
  assign n13779 = ~n7353 & n13778 ;
  assign n13780 = n13779 ^ x877 ;
  assign n13781 = x1137 ^ x878 ;
  assign n13782 = ~n7353 & n13781 ;
  assign n13783 = n13782 ^ x878 ;
  assign n13784 = x1135 ^ x879 ;
  assign n13785 = ~n7353 & n13784 ;
  assign n13786 = n13785 ^ x879 ;
  assign n13787 = x1081 ^ x880 ;
  assign n13788 = ~x955 & n13787 ;
  assign n13789 = n13788 ^ x880 ;
  assign n13790 = x1059 ^ x881 ;
  assign n13791 = ~x955 & n13790 ;
  assign n13792 = n13791 ^ x881 ;
  assign n13793 = x1107 ^ x883 ;
  assign n13794 = ~n13605 & ~n13793 ;
  assign n13795 = n13794 ^ x883 ;
  assign n13796 = x1124 ^ x884 ;
  assign n13797 = ~n13605 & ~n13796 ;
  assign n13798 = n13797 ^ x884 ;
  assign n13799 = x1125 ^ x885 ;
  assign n13800 = ~n13605 & ~n13799 ;
  assign n13801 = n13800 ^ x885 ;
  assign n13802 = x1109 ^ x886 ;
  assign n13803 = ~n13605 & ~n13802 ;
  assign n13804 = n13803 ^ x886 ;
  assign n13805 = x1100 ^ x887 ;
  assign n13806 = ~n13605 & ~n13805 ;
  assign n13807 = n13806 ^ x887 ;
  assign n13808 = x1120 ^ x888 ;
  assign n13809 = ~n13605 & ~n13808 ;
  assign n13810 = n13809 ^ x888 ;
  assign n13811 = x1103 ^ x889 ;
  assign n13812 = ~n13605 & ~n13811 ;
  assign n13813 = n13812 ^ x889 ;
  assign n13814 = x1126 ^ x890 ;
  assign n13815 = ~n13605 & ~n13814 ;
  assign n13816 = n13815 ^ x890 ;
  assign n13817 = x1116 ^ x891 ;
  assign n13818 = ~n13605 & ~n13817 ;
  assign n13819 = n13818 ^ x891 ;
  assign n13820 = x1101 ^ x892 ;
  assign n13821 = ~n13605 & ~n13820 ;
  assign n13822 = n13821 ^ x892 ;
  assign n13823 = x1119 ^ x894 ;
  assign n13824 = ~n13605 & ~n13823 ;
  assign n13825 = n13824 ^ x894 ;
  assign n13826 = x1113 ^ x895 ;
  assign n13827 = ~n13605 & ~n13826 ;
  assign n13828 = n13827 ^ x895 ;
  assign n13829 = x1118 ^ x896 ;
  assign n13830 = ~n13605 & ~n13829 ;
  assign n13831 = n13830 ^ x896 ;
  assign n13832 = x1129 ^ x898 ;
  assign n13833 = ~n13605 & ~n13832 ;
  assign n13834 = n13833 ^ x898 ;
  assign n13835 = x1115 ^ x899 ;
  assign n13836 = ~n13605 & ~n13835 ;
  assign n13837 = n13836 ^ x899 ;
  assign n13838 = x1110 ^ x900 ;
  assign n13839 = ~n13605 & ~n13838 ;
  assign n13840 = n13839 ^ x900 ;
  assign n13841 = x1111 ^ x902 ;
  assign n13842 = ~n13605 & ~n13841 ;
  assign n13843 = n13842 ^ x902 ;
  assign n13844 = x1121 ^ x903 ;
  assign n13845 = ~n13605 & ~n13844 ;
  assign n13846 = n13845 ^ x903 ;
  assign n13847 = x1127 ^ x904 ;
  assign n13848 = ~n13605 & ~n13847 ;
  assign n13849 = n13848 ^ x904 ;
  assign n13850 = x1131 ^ x905 ;
  assign n13851 = ~n13605 & ~n13850 ;
  assign n13852 = n13851 ^ x905 ;
  assign n13853 = x1128 ^ x906 ;
  assign n13854 = ~n13605 & ~n13853 ;
  assign n13855 = n13854 ^ x906 ;
  assign n13858 = ~x598 & x979 ;
  assign n13859 = ~x615 & n13858 ;
  assign n13856 = ~x624 & ~x979 ;
  assign n13857 = x604 & n13856 ;
  assign n13860 = n13859 ^ n13857 ;
  assign n13861 = n13860 ^ x907 ;
  assign n13862 = x782 & n13861 ;
  assign n13863 = n13862 ^ x907 ;
  assign n13864 = x1122 ^ x908 ;
  assign n13865 = ~n13605 & ~n13864 ;
  assign n13866 = n13865 ^ x908 ;
  assign n13867 = x1105 ^ x909 ;
  assign n13868 = ~n13605 & ~n13867 ;
  assign n13869 = n13868 ^ x909 ;
  assign n13870 = x1117 ^ x910 ;
  assign n13871 = ~n13605 & ~n13870 ;
  assign n13872 = n13871 ^ x910 ;
  assign n13873 = x1130 ^ x911 ;
  assign n13874 = ~n13605 & ~n13873 ;
  assign n13875 = n13874 ^ x911 ;
  assign n13876 = x1114 ^ x912 ;
  assign n13877 = ~n13605 & ~n13876 ;
  assign n13878 = n13877 ^ x912 ;
  assign n13879 = x1106 ^ x913 ;
  assign n13880 = ~n13605 & ~n13879 ;
  assign n13881 = n13880 ^ x913 ;
  assign n13882 = n9339 ^ x280 ;
  assign n13883 = x1108 ^ x915 ;
  assign n13884 = ~n13605 & ~n13883 ;
  assign n13885 = n13884 ^ x915 ;
  assign n13886 = x1123 ^ x916 ;
  assign n13887 = ~n13605 & ~n13886 ;
  assign n13888 = n13887 ^ x916 ;
  assign n13889 = x1112 ^ x917 ;
  assign n13890 = ~n13605 & ~n13889 ;
  assign n13891 = n13890 ^ x917 ;
  assign n13892 = x1104 ^ x918 ;
  assign n13893 = ~n13605 & ~n13892 ;
  assign n13894 = n13893 ^ x918 ;
  assign n13895 = x1102 ^ x919 ;
  assign n13896 = ~n13605 & ~n13895 ;
  assign n13897 = n13896 ^ x919 ;
  assign n13898 = x1139 ^ x920 ;
  assign n13899 = x1093 & n13898 ;
  assign n13900 = n13899 ^ x920 ;
  assign n13901 = x1140 ^ x921 ;
  assign n13902 = x1093 & n13901 ;
  assign n13903 = n13902 ^ x921 ;
  assign n13904 = x1152 ^ x922 ;
  assign n13905 = x1093 & n13904 ;
  assign n13906 = n13905 ^ x922 ;
  assign n13907 = x1154 ^ x923 ;
  assign n13908 = x1093 & n13907 ;
  assign n13909 = n13908 ^ x923 ;
  assign n13910 = x311 & n7713 ;
  assign n13911 = x1155 ^ x925 ;
  assign n13912 = x1093 & n13911 ;
  assign n13913 = n13912 ^ x925 ;
  assign n13914 = x1157 ^ x926 ;
  assign n13915 = x1093 & n13914 ;
  assign n13916 = n13915 ^ x926 ;
  assign n13917 = x1145 ^ x927 ;
  assign n13918 = x1093 & n13917 ;
  assign n13919 = n13918 ^ x927 ;
  assign n13920 = x1136 ^ x928 ;
  assign n13921 = x1093 & n13920 ;
  assign n13922 = n13921 ^ x928 ;
  assign n13923 = x1144 ^ x929 ;
  assign n13924 = x1093 & n13923 ;
  assign n13925 = n13924 ^ x929 ;
  assign n13926 = x1134 ^ x930 ;
  assign n13927 = x1093 & n13926 ;
  assign n13928 = n13927 ^ x930 ;
  assign n13929 = x1150 ^ x931 ;
  assign n13930 = x1093 & n13929 ;
  assign n13931 = n13930 ^ x931 ;
  assign n13932 = x1093 & n2075 ;
  assign n13933 = n13932 ^ x932 ;
  assign n13934 = x1137 ^ x933 ;
  assign n13935 = x1093 & n13934 ;
  assign n13936 = n13935 ^ x933 ;
  assign n13937 = x1147 ^ x934 ;
  assign n13938 = x1093 & n13937 ;
  assign n13939 = n13938 ^ x934 ;
  assign n13940 = x1141 ^ x935 ;
  assign n13941 = x1093 & n13940 ;
  assign n13942 = n13941 ^ x935 ;
  assign n13943 = x1149 ^ x936 ;
  assign n13944 = x1093 & n13943 ;
  assign n13945 = n13944 ^ x936 ;
  assign n13946 = x1148 ^ x937 ;
  assign n13947 = x1093 & n13946 ;
  assign n13948 = n13947 ^ x937 ;
  assign n13949 = x1135 ^ x938 ;
  assign n13950 = x1093 & n13949 ;
  assign n13951 = n13950 ^ x938 ;
  assign n13952 = x1146 ^ x939 ;
  assign n13953 = x1093 & n13952 ;
  assign n13954 = n13953 ^ x939 ;
  assign n13955 = x1138 ^ x940 ;
  assign n13956 = x1093 & n13955 ;
  assign n13957 = n13956 ^ x940 ;
  assign n13958 = x1153 ^ x941 ;
  assign n13959 = x1093 & n13958 ;
  assign n13960 = n13959 ^ x941 ;
  assign n13961 = x1156 ^ x942 ;
  assign n13962 = x1093 & n13961 ;
  assign n13963 = n13962 ^ x942 ;
  assign n13964 = x1151 ^ x943 ;
  assign n13965 = x1093 & n13964 ;
  assign n13966 = n13965 ^ x943 ;
  assign n13967 = x1143 ^ x944 ;
  assign n13968 = x1093 & n13967 ;
  assign n13969 = n13968 ^ x944 ;
  assign n13970 = x230 & n2985 ;
  assign n13971 = n13858 ^ x947 ;
  assign n13972 = n13971 ^ n13856 ;
  assign n13973 = x782 & ~n13972 ;
  assign n13974 = n13973 ^ x947 ;
  assign n13975 = x992 ^ x266 ;
  assign n13976 = x949 ^ x313 ;
  assign n13977 = x954 & ~n13976 ;
  assign n13978 = n13977 ^ x313 ;
  assign n13979 = x1092 & n1569 ;
  assign n13980 = ~x31 & x957 ;
  assign n13981 = x1092 & n13980 ;
  assign n13982 = n13981 ^ x31 ;
  assign n13983 = ~x782 & x960 ;
  assign n13984 = ~x230 & x961 ;
  assign n13985 = ~x782 & x963 ;
  assign n13986 = ~x230 & x967 ;
  assign n13987 = ~x230 & x969 ;
  assign n13988 = ~x782 & x970 ;
  assign n13989 = ~x230 & x971 ;
  assign n13990 = ~x782 & x972 ;
  assign n13991 = ~x230 & x974 ;
  assign n13992 = ~x782 & x975 ;
  assign n13993 = ~x230 & x977 ;
  assign n13994 = ~x782 & x978 ;
  assign n13995 = ~x598 & x615 ;
  assign n13996 = x824 & x1092 ;
  assign n13997 = ~x604 & ~x624 ;
  assign y0 = x668 ;
  assign y1 = x672 ;
  assign y2 = x664 ;
  assign y3 = x667 ;
  assign y4 = x676 ;
  assign y5 = x673 ;
  assign y6 = x675 ;
  assign y7 = x666 ;
  assign y8 = x679 ;
  assign y9 = x674 ;
  assign y10 = x663 ;
  assign y11 = x670 ;
  assign y12 = x677 ;
  assign y13 = x682 ;
  assign y14 = x671 ;
  assign y15 = x678 ;
  assign y16 = x718 ;
  assign y17 = x707 ;
  assign y18 = x708 ;
  assign y19 = x713 ;
  assign y20 = x711 ;
  assign y21 = x716 ;
  assign y22 = x733 ;
  assign y23 = x712 ;
  assign y24 = x689 ;
  assign y25 = x717 ;
  assign y26 = x692 ;
  assign y27 = x719 ;
  assign y28 = x722 ;
  assign y29 = x714 ;
  assign y30 = x720 ;
  assign y31 = x685 ;
  assign y32 = x837 ;
  assign y33 = x850 ;
  assign y34 = x872 ;
  assign y35 = x871 ;
  assign y36 = x881 ;
  assign y37 = x866 ;
  assign y38 = x876 ;
  assign y39 = x873 ;
  assign y40 = x874 ;
  assign y41 = x859 ;
  assign y42 = x855 ;
  assign y43 = x852 ;
  assign y44 = x870 ;
  assign y45 = x848 ;
  assign y46 = x865 ;
  assign y47 = x856 ;
  assign y48 = x853 ;
  assign y49 = x847 ;
  assign y50 = x857 ;
  assign y51 = x854 ;
  assign y52 = x858 ;
  assign y53 = x845 ;
  assign y54 = x838 ;
  assign y55 = x842 ;
  assign y56 = x843 ;
  assign y57 = x839 ;
  assign y58 = x844 ;
  assign y59 = x868 ;
  assign y60 = x851 ;
  assign y61 = x867 ;
  assign y62 = x880 ;
  assign y63 = x860 ;
  assign y64 = x1030 ;
  assign y65 = x1034 ;
  assign y66 = x1015 ;
  assign y67 = x1020 ;
  assign y68 = x1025 ;
  assign y69 = x1005 ;
  assign y70 = x996 ;
  assign y71 = x1012 ;
  assign y72 = x993 ;
  assign y73 = x1016 ;
  assign y74 = x1021 ;
  assign y75 = x1010 ;
  assign y76 = x1027 ;
  assign y77 = x1018 ;
  assign y78 = x1017 ;
  assign y79 = x1024 ;
  assign y80 = x1009 ;
  assign y81 = x1032 ;
  assign y82 = x1003 ;
  assign y83 = x997 ;
  assign y84 = x1013 ;
  assign y85 = x1011 ;
  assign y86 = x1008 ;
  assign y87 = x1019 ;
  assign y88 = x1031 ;
  assign y89 = x1022 ;
  assign y90 = x1000 ;
  assign y91 = x1023 ;
  assign y92 = x1002 ;
  assign y93 = x1026 ;
  assign y94 = x1006 ;
  assign y95 = x998 ;
  assign y96 = x31 ;
  assign y97 = x80 ;
  assign y98 = x893 ;
  assign y99 = x467 ;
  assign y100 = x78 ;
  assign y101 = x112 ;
  assign y102 = x13 ;
  assign y103 = x25 ;
  assign y104 = x226 ;
  assign y105 = x127 ;
  assign y106 = x822 ;
  assign y107 = x808 ;
  assign y108 = x227 ;
  assign y109 = x477 ;
  assign y110 = x834 ;
  assign y111 = x229 ;
  assign y112 = x12 ;
  assign y113 = x11 ;
  assign y114 = x10 ;
  assign y115 = x9 ;
  assign y116 = x8 ;
  assign y117 = x7 ;
  assign y118 = x6 ;
  assign y119 = x5 ;
  assign y120 = x4 ;
  assign y121 = x3 ;
  assign y122 = x0 ;
  assign y123 = x2 ;
  assign y124 = x1 ;
  assign y125 = x310 ;
  assign y126 = x302 ;
  assign y127 = x475 ;
  assign y128 = x474 ;
  assign y129 = x466 ;
  assign y130 = x473 ;
  assign y131 = x471 ;
  assign y132 = x472 ;
  assign y133 = x470 ;
  assign y134 = x469 ;
  assign y135 = x465 ;
  assign y136 = x1028 ;
  assign y137 = x1033 ;
  assign y138 = x995 ;
  assign y139 = x994 ;
  assign y140 = x28 ;
  assign y141 = x27 ;
  assign y142 = x26 ;
  assign y143 = x29 ;
  assign y144 = x15 ;
  assign y145 = x14 ;
  assign y146 = x21 ;
  assign y147 = x20 ;
  assign y148 = x19 ;
  assign y149 = x18 ;
  assign y150 = x17 ;
  assign y151 = x16 ;
  assign y152 = x1096 ;
  assign y153 = ~n1930 ;
  assign y154 = n1984 ;
  assign y155 = n2006 ;
  assign y156 = n2074 ;
  assign y157 = ~n2163 ;
  assign y158 = ~n2224 ;
  assign y159 = n2266 ;
  assign y160 = n2332 ;
  assign y161 = n2386 ;
  assign y162 = n2444 ;
  assign y163 = n2499 ;
  assign y164 = n2554 ;
  assign y165 = ~n2606 ;
  assign y166 = ~1'b0 ;
  assign y167 = ~n2736 ;
  assign y168 = x228 ;
  assign y169 = x22 ;
  assign y170 = ~x1090 ;
  assign y171 = ~n2857 ;
  assign y172 = ~n2876 ;
  assign y173 = ~n2881 ;
  assign y174 = ~n2912 ;
  assign y175 = ~n2916 ;
  assign y176 = ~n2920 ;
  assign y177 = ~n2924 ;
  assign y178 = ~n2928 ;
  assign y179 = x1089 ;
  assign y180 = x23 ;
  assign y181 = ~n2736 ;
  assign y182 = ~n2964 ;
  assign y183 = n2972 ;
  assign y184 = ~n2978 ;
  assign y185 = ~n2980 ;
  assign y186 = ~n2982 ;
  assign y187 = ~n2984 ;
  assign y188 = x37 ;
  assign y189 = ~n3434 ;
  assign y190 = ~n3480 ;
  assign y191 = ~n3673 ;
  assign y192 = n3785 ;
  assign y193 = n3872 ;
  assign y194 = n3878 ;
  assign y195 = ~n2961 ;
  assign y196 = ~n3895 ;
  assign y197 = ~n3934 ;
  assign y198 = n3937 ;
  assign y199 = n4000 ;
  assign y200 = n4043 ;
  assign y201 = n4053 ;
  assign y202 = n4059 ;
  assign y203 = n4060 ;
  assign y204 = n4068 ;
  assign y205 = n4082 ;
  assign y206 = n4083 ;
  assign y207 = n4150 ;
  assign y208 = ~n4172 ;
  assign y209 = n4176 ;
  assign y210 = n4253 ;
  assign y211 = n4261 ;
  assign y212 = n4268 ;
  assign y213 = n4272 ;
  assign y214 = n4279 ;
  assign y215 = n4285 ;
  assign y216 = n4288 ;
  assign y217 = n4292 ;
  assign y218 = ~n4297 ;
  assign y219 = n4299 ;
  assign y220 = n4308 ;
  assign y221 = ~n4312 ;
  assign y222 = n4315 ;
  assign y223 = n4317 ;
  assign y224 = n4325 ;
  assign y225 = n4330 ;
  assign y226 = n4336 ;
  assign y227 = n4341 ;
  assign y228 = ~n4357 ;
  assign y229 = n4378 ;
  assign y230 = ~n4397 ;
  assign y231 = n4406 ;
  assign y232 = ~n4418 ;
  assign y233 = n4422 ;
  assign y234 = n4447 ;
  assign y235 = n4450 ;
  assign y236 = n4451 ;
  assign y237 = ~n4578 ;
  assign y238 = n4610 ;
  assign y239 = ~n4615 ;
  assign y240 = n4621 ;
  assign y241 = n4627 ;
  assign y242 = n4628 ;
  assign y243 = n4631 ;
  assign y244 = n4632 ;
  assign y245 = n4633 ;
  assign y246 = n4641 ;
  assign y247 = n4646 ;
  assign y248 = n4648 ;
  assign y249 = n4659 ;
  assign y250 = n4666 ;
  assign y251 = n4671 ;
  assign y252 = n4710 ;
  assign y253 = ~n4776 ;
  assign y254 = n4787 ;
  assign y255 = ~n4791 ;
  assign y256 = n4793 ;
  assign y257 = n4808 ;
  assign y258 = n4828 ;
  assign y259 = n4834 ;
  assign y260 = n4835 ;
  assign y261 = n4836 ;
  assign y262 = ~n4841 ;
  assign y263 = x117 ;
  assign y264 = n4842 ;
  assign y265 = n4310 ;
  assign y266 = n4849 ;
  assign y267 = n4850 ;
  assign y268 = ~n4854 ;
  assign y269 = n4858 ;
  assign y270 = ~n4859 ;
  assign y271 = n4866 ;
  assign y272 = n4868 ;
  assign y273 = n4875 ;
  assign y274 = n4877 ;
  assign y275 = ~n2969 ;
  assign y276 = n5007 ;
  assign y277 = n5025 ;
  assign y278 = n5038 ;
  assign y279 = ~n5176 ;
  assign y280 = n5037 ;
  assign y281 = n5190 ;
  assign y282 = n5298 ;
  assign y283 = ~n5369 ;
  assign y284 = n5377 ;
  assign y285 = x131 ;
  assign y286 = ~n5392 ;
  assign y287 = ~n5426 ;
  assign y288 = ~n5022 ;
  assign y289 = n5475 ;
  assign y290 = ~n5500 ;
  assign y291 = n5523 ;
  assign y292 = n5544 ;
  assign y293 = n5573 ;
  assign y294 = n5581 ;
  assign y295 = ~n5611 ;
  assign y296 = n5617 ;
  assign y297 = ~n5784 ;
  assign y298 = ~n5795 ;
  assign y299 = n5806 ;
  assign y300 = ~n5817 ;
  assign y301 = n5828 ;
  assign y302 = ~n5839 ;
  assign y303 = n5848 ;
  assign y304 = ~n5859 ;
  assign y305 = ~n5868 ;
  assign y306 = n5894 ;
  assign y307 = n5906 ;
  assign y308 = ~n5917 ;
  assign y309 = n5928 ;
  assign y310 = ~n5939 ;
  assign y311 = n5951 ;
  assign y312 = n5963 ;
  assign y313 = n5975 ;
  assign y314 = ~n5986 ;
  assign y315 = n5998 ;
  assign y316 = ~n6009 ;
  assign y317 = ~n6020 ;
  assign y318 = n6029 ;
  assign y319 = ~n6038 ;
  assign y320 = ~n6049 ;
  assign y321 = ~n6060 ;
  assign y322 = n6070 ;
  assign y323 = n6081 ;
  assign y324 = ~n6092 ;
  assign y325 = ~n6103 ;
  assign y326 = ~n6114 ;
  assign y327 = ~n6125 ;
  assign y328 = ~n6136 ;
  assign y329 = ~n6147 ;
  assign y330 = ~n6156 ;
  assign y331 = n6165 ;
  assign y332 = ~n6174 ;
  assign y333 = ~n6183 ;
  assign y334 = ~n6192 ;
  assign y335 = ~n6201 ;
  assign y336 = ~n6210 ;
  assign y337 = ~n6219 ;
  assign y338 = ~n6228 ;
  assign y339 = ~n6237 ;
  assign y340 = ~n6246 ;
  assign y341 = ~n6255 ;
  assign y342 = ~n6264 ;
  assign y343 = ~n6273 ;
  assign y344 = ~n6282 ;
  assign y345 = ~n6291 ;
  assign y346 = n6300 ;
  assign y347 = ~n6309 ;
  assign y348 = ~n6318 ;
  assign y349 = ~n6327 ;
  assign y350 = ~n6336 ;
  assign y351 = ~n6345 ;
  assign y352 = ~n6362 ;
  assign y353 = n6373 ;
  assign y354 = ~n6382 ;
  assign y355 = n6393 ;
  assign y356 = n6404 ;
  assign y357 = n6415 ;
  assign y358 = n6450 ;
  assign y359 = n6459 ;
  assign y360 = n6466 ;
  assign y361 = n6484 ;
  assign y362 = n6489 ;
  assign y363 = n6498 ;
  assign y364 = ~n6509 ;
  assign y365 = ~n6520 ;
  assign y366 = ~n6531 ;
  assign y367 = n6540 ;
  assign y368 = n6549 ;
  assign y369 = n6559 ;
  assign y370 = n6569 ;
  assign y371 = ~n6578 ;
  assign y372 = n6589 ;
  assign y373 = n6600 ;
  assign y374 = ~n6611 ;
  assign y375 = n6616 ;
  assign y376 = n6626 ;
  assign y377 = n6632 ;
  assign y378 = n6643 ;
  assign y379 = n6652 ;
  assign y380 = n6661 ;
  assign y381 = n6670 ;
  assign y382 = ~n6691 ;
  assign y383 = n6702 ;
  assign y384 = ~n6713 ;
  assign y385 = ~n6721 ;
  assign y386 = x232 ;
  assign y387 = n6725 ;
  assign y388 = x236 ;
  assign y389 = ~n6733 ;
  assign y390 = ~n6849 ;
  assign y391 = n6902 ;
  assign y392 = n6950 ;
  assign y393 = n6699 ;
  assign y394 = ~n7052 ;
  assign y395 = n7084 ;
  assign y396 = n7097 ;
  assign y397 = n7124 ;
  assign y398 = n7142 ;
  assign y399 = n7159 ;
  assign y400 = ~n7191 ;
  assign y401 = n7199 ;
  assign y402 = n7217 ;
  assign y403 = n7235 ;
  assign y404 = n7244 ;
  assign y405 = n7262 ;
  assign y406 = n7271 ;
  assign y407 = ~n7274 ;
  assign y408 = n7284 ;
  assign y409 = ~n7290 ;
  assign y410 = n7299 ;
  assign y411 = n7308 ;
  assign y412 = n7314 ;
  assign y413 = n7320 ;
  assign y414 = n7326 ;
  assign y415 = n7332 ;
  assign y416 = n7338 ;
  assign y417 = n7344 ;
  assign y418 = n7350 ;
  assign y419 = ~n7361 ;
  assign y420 = ~n7370 ;
  assign y421 = ~n7381 ;
  assign y422 = ~n7392 ;
  assign y423 = n7403 ;
  assign y424 = n7412 ;
  assign y425 = n7421 ;
  assign y426 = ~n7432 ;
  assign y427 = ~n7443 ;
  assign y428 = n7452 ;
  assign y429 = n7461 ;
  assign y430 = n7470 ;
  assign y431 = ~n7481 ;
  assign y432 = n7490 ;
  assign y433 = n7499 ;
  assign y434 = ~n7510 ;
  assign y435 = n7521 ;
  assign y436 = n7532 ;
  assign y437 = ~n7543 ;
  assign y438 = ~n7554 ;
  assign y439 = ~n7565 ;
  assign y440 = n7574 ;
  assign y441 = ~n7586 ;
  assign y442 = n7598 ;
  assign y443 = n7605 ;
  assign y444 = ~n7608 ;
  assign y445 = n7611 ;
  assign y446 = n7619 ;
  assign y447 = n7622 ;
  assign y448 = n7625 ;
  assign y449 = n7628 ;
  assign y450 = n7631 ;
  assign y451 = n7634 ;
  assign y452 = n7637 ;
  assign y453 = n7640 ;
  assign y454 = n7643 ;
  assign y455 = n7646 ;
  assign y456 = ~n7653 ;
  assign y457 = ~n7661 ;
  assign y458 = n7669 ;
  assign y459 = ~n7684 ;
  assign y460 = n7687 ;
  assign y461 = n7690 ;
  assign y462 = n7693 ;
  assign y463 = n7696 ;
  assign y464 = n7699 ;
  assign y465 = n7702 ;
  assign y466 = n7705 ;
  assign y467 = ~n7712 ;
  assign y468 = n7720 ;
  assign y469 = n7722 ;
  assign y470 = ~n7733 ;
  assign y471 = n7734 ;
  assign y472 = n7738 ;
  assign y473 = n7741 ;
  assign y474 = n7745 ;
  assign y475 = n7749 ;
  assign y476 = n7752 ;
  assign y477 = n7755 ;
  assign y478 = n7758 ;
  assign y479 = n7761 ;
  assign y480 = n7764 ;
  assign y481 = n7767 ;
  assign y482 = n7770 ;
  assign y483 = n7773 ;
  assign y484 = n7776 ;
  assign y485 = n7779 ;
  assign y486 = n7782 ;
  assign y487 = n7787 ;
  assign y488 = n7791 ;
  assign y489 = ~n7795 ;
  assign y490 = n7798 ;
  assign y491 = n7801 ;
  assign y492 = n7804 ;
  assign y493 = n7807 ;
  assign y494 = n7810 ;
  assign y495 = n7813 ;
  assign y496 = n7816 ;
  assign y497 = ~n7819 ;
  assign y498 = n7822 ;
  assign y499 = n7825 ;
  assign y500 = n7828 ;
  assign y501 = n7831 ;
  assign y502 = n7834 ;
  assign y503 = n7837 ;
  assign y504 = n7840 ;
  assign y505 = n7843 ;
  assign y506 = n7846 ;
  assign y507 = n7849 ;
  assign y508 = n7852 ;
  assign y509 = n7855 ;
  assign y510 = n7858 ;
  assign y511 = n7861 ;
  assign y512 = n7864 ;
  assign y513 = n7867 ;
  assign y514 = n7870 ;
  assign y515 = n7873 ;
  assign y516 = n7876 ;
  assign y517 = n7879 ;
  assign y518 = n7882 ;
  assign y519 = n7885 ;
  assign y520 = n7888 ;
  assign y521 = n7891 ;
  assign y522 = n7894 ;
  assign y523 = n7897 ;
  assign y524 = n7900 ;
  assign y525 = n7903 ;
  assign y526 = n7906 ;
  assign y527 = n7909 ;
  assign y528 = n7912 ;
  assign y529 = n7915 ;
  assign y530 = n7918 ;
  assign y531 = n7921 ;
  assign y532 = n7924 ;
  assign y533 = n7927 ;
  assign y534 = n7930 ;
  assign y535 = n7933 ;
  assign y536 = n7936 ;
  assign y537 = n7939 ;
  assign y538 = n7942 ;
  assign y539 = n7945 ;
  assign y540 = n7948 ;
  assign y541 = n7951 ;
  assign y542 = n7954 ;
  assign y543 = n7957 ;
  assign y544 = n7960 ;
  assign y545 = n7963 ;
  assign y546 = n7966 ;
  assign y547 = n7969 ;
  assign y548 = n7972 ;
  assign y549 = n7975 ;
  assign y550 = n7978 ;
  assign y551 = n7981 ;
  assign y552 = n7984 ;
  assign y553 = n7987 ;
  assign y554 = n7990 ;
  assign y555 = n7993 ;
  assign y556 = n7996 ;
  assign y557 = n7999 ;
  assign y558 = n8002 ;
  assign y559 = n8005 ;
  assign y560 = n8008 ;
  assign y561 = n8011 ;
  assign y562 = n8014 ;
  assign y563 = n8017 ;
  assign y564 = n8020 ;
  assign y565 = n8023 ;
  assign y566 = n8026 ;
  assign y567 = n8029 ;
  assign y568 = n8032 ;
  assign y569 = n8035 ;
  assign y570 = n8038 ;
  assign y571 = n8041 ;
  assign y572 = n8044 ;
  assign y573 = n8047 ;
  assign y574 = n8050 ;
  assign y575 = n8053 ;
  assign y576 = n8056 ;
  assign y577 = n8059 ;
  assign y578 = n8062 ;
  assign y579 = n8065 ;
  assign y580 = n8068 ;
  assign y581 = n8071 ;
  assign y582 = n8074 ;
  assign y583 = n8077 ;
  assign y584 = n8080 ;
  assign y585 = n8083 ;
  assign y586 = n8086 ;
  assign y587 = n8089 ;
  assign y588 = n8092 ;
  assign y589 = n8095 ;
  assign y590 = n8098 ;
  assign y591 = n8101 ;
  assign y592 = n8104 ;
  assign y593 = n8107 ;
  assign y594 = n8110 ;
  assign y595 = n8113 ;
  assign y596 = n8116 ;
  assign y597 = n8119 ;
  assign y598 = n8122 ;
  assign y599 = n8125 ;
  assign y600 = n8128 ;
  assign y601 = n8131 ;
  assign y602 = n8134 ;
  assign y603 = n8137 ;
  assign y604 = n8140 ;
  assign y605 = n8143 ;
  assign y606 = n8146 ;
  assign y607 = n8149 ;
  assign y608 = n8152 ;
  assign y609 = n8155 ;
  assign y610 = n8158 ;
  assign y611 = n8161 ;
  assign y612 = n8164 ;
  assign y613 = n8167 ;
  assign y614 = n8215 ;
  assign y615 = n8218 ;
  assign y616 = n8221 ;
  assign y617 = n8224 ;
  assign y618 = n8227 ;
  assign y619 = n8230 ;
  assign y620 = n8233 ;
  assign y621 = n8236 ;
  assign y622 = n8241 ;
  assign y623 = n8246 ;
  assign y624 = ~n8251 ;
  assign y625 = n8254 ;
  assign y626 = n8259 ;
  assign y627 = n8264 ;
  assign y628 = n8269 ;
  assign y629 = n8274 ;
  assign y630 = n8279 ;
  assign y631 = n8284 ;
  assign y632 = n8289 ;
  assign y633 = n8292 ;
  assign y634 = ~n7730 ;
  assign y635 = n8293 ;
  assign y636 = x583 ;
  assign y637 = n7587 ;
  assign y638 = n8296 ;
  assign y639 = n8299 ;
  assign y640 = n8302 ;
  assign y641 = n8305 ;
  assign y642 = n8308 ;
  assign y643 = n8311 ;
  assign y644 = n8314 ;
  assign y645 = n8317 ;
  assign y646 = n8320 ;
  assign y647 = n8323 ;
  assign y648 = n8326 ;
  assign y649 = n8329 ;
  assign y650 = n8332 ;
  assign y651 = n8335 ;
  assign y652 = n8338 ;
  assign y653 = n8341 ;
  assign y654 = n8344 ;
  assign y655 = n8347 ;
  assign y656 = n8350 ;
  assign y657 = n8353 ;
  assign y658 = n8356 ;
  assign y659 = n8359 ;
  assign y660 = n8362 ;
  assign y661 = n8365 ;
  assign y662 = n8368 ;
  assign y663 = n8371 ;
  assign y664 = n8374 ;
  assign y665 = n8377 ;
  assign y666 = n8380 ;
  assign y667 = n8383 ;
  assign y668 = n8386 ;
  assign y669 = n8389 ;
  assign y670 = n8392 ;
  assign y671 = n8395 ;
  assign y672 = n8398 ;
  assign y673 = n8401 ;
  assign y674 = n8404 ;
  assign y675 = n8407 ;
  assign y676 = n8410 ;
  assign y677 = n8413 ;
  assign y678 = n8416 ;
  assign y679 = n8419 ;
  assign y680 = n8422 ;
  assign y681 = n8425 ;
  assign y682 = n8428 ;
  assign y683 = n8431 ;
  assign y684 = n8434 ;
  assign y685 = n8437 ;
  assign y686 = n8440 ;
  assign y687 = n8443 ;
  assign y688 = n8446 ;
  assign y689 = n8449 ;
  assign y690 = n8452 ;
  assign y691 = n8455 ;
  assign y692 = n8458 ;
  assign y693 = n8461 ;
  assign y694 = n8464 ;
  assign y695 = n8467 ;
  assign y696 = n8470 ;
  assign y697 = n8473 ;
  assign y698 = n8476 ;
  assign y699 = n8479 ;
  assign y700 = n8482 ;
  assign y701 = n8485 ;
  assign y702 = n8488 ;
  assign y703 = n8491 ;
  assign y704 = n8494 ;
  assign y705 = n8497 ;
  assign y706 = n8500 ;
  assign y707 = n8503 ;
  assign y708 = n8506 ;
  assign y709 = n8509 ;
  assign y710 = n8512 ;
  assign y711 = n8515 ;
  assign y712 = n8518 ;
  assign y713 = n8521 ;
  assign y714 = n8524 ;
  assign y715 = n8527 ;
  assign y716 = n8530 ;
  assign y717 = n8533 ;
  assign y718 = n8536 ;
  assign y719 = n8539 ;
  assign y720 = n8542 ;
  assign y721 = n8545 ;
  assign y722 = n8548 ;
  assign y723 = n8551 ;
  assign y724 = n8560 ;
  assign y725 = n8563 ;
  assign y726 = n8566 ;
  assign y727 = n8569 ;
  assign y728 = n8572 ;
  assign y729 = n8575 ;
  assign y730 = n8578 ;
  assign y731 = n8581 ;
  assign y732 = n8584 ;
  assign y733 = n8587 ;
  assign y734 = n8590 ;
  assign y735 = n8593 ;
  assign y736 = n8596 ;
  assign y737 = n8599 ;
  assign y738 = n8602 ;
  assign y739 = n8605 ;
  assign y740 = ~n2640 ;
  assign y741 = n8608 ;
  assign y742 = n8611 ;
  assign y743 = n8614 ;
  assign y744 = n8617 ;
  assign y745 = n8625 ;
  assign y746 = n8653 ;
  assign y747 = ~n8659 ;
  assign y748 = n8665 ;
  assign y749 = n8671 ;
  assign y750 = ~n8797 ;
  assign y751 = n8805 ;
  assign y752 = n8816 ;
  assign y753 = n8821 ;
  assign y754 = n8823 ;
  assign y755 = ~n8895 ;
  assign y756 = n8902 ;
  assign y757 = n8904 ;
  assign y758 = n8908 ;
  assign y759 = n8911 ;
  assign y760 = n8928 ;
  assign y761 = n8938 ;
  assign y762 = n8940 ;
  assign y763 = n8949 ;
  assign y764 = n8955 ;
  assign y765 = n8961 ;
  assign y766 = n8967 ;
  assign y767 = n8973 ;
  assign y768 = n8979 ;
  assign y769 = n8985 ;
  assign y770 = n8991 ;
  assign y771 = n9000 ;
  assign y772 = ~n9065 ;
  assign y773 = n9074 ;
  assign y774 = n9083 ;
  assign y775 = n9089 ;
  assign y776 = n9095 ;
  assign y777 = n9101 ;
  assign y778 = n9107 ;
  assign y779 = n9113 ;
  assign y780 = n9119 ;
  assign y781 = n9128 ;
  assign y782 = n9140 ;
  assign y783 = n9146 ;
  assign y784 = n9152 ;
  assign y785 = n9158 ;
  assign y786 = n9164 ;
  assign y787 = n9170 ;
  assign y788 = n9176 ;
  assign y789 = n9182 ;
  assign y790 = n9188 ;
  assign y791 = n9194 ;
  assign y792 = n9200 ;
  assign y793 = n9206 ;
  assign y794 = n9212 ;
  assign y795 = n9218 ;
  assign y796 = n9224 ;
  assign y797 = n9230 ;
  assign y798 = n9236 ;
  assign y799 = n9242 ;
  assign y800 = n9248 ;
  assign y801 = n9254 ;
  assign y802 = n9260 ;
  assign y803 = n9266 ;
  assign y804 = n9272 ;
  assign y805 = n9278 ;
  assign y806 = n9284 ;
  assign y807 = n9290 ;
  assign y808 = n9296 ;
  assign y809 = n9302 ;
  assign y810 = n9308 ;
  assign y811 = n9314 ;
  assign y812 = n9320 ;
  assign y813 = n9326 ;
  assign y814 = n9332 ;
  assign y815 = n9338 ;
  assign y816 = ~n9348 ;
  assign y817 = n9354 ;
  assign y818 = n9360 ;
  assign y819 = n9366 ;
  assign y820 = n9500 ;
  assign y821 = n9624 ;
  assign y822 = n9630 ;
  assign y823 = n9754 ;
  assign y824 = n9878 ;
  assign y825 = n10002 ;
  assign y826 = n10008 ;
  assign y827 = ~n10071 ;
  assign y828 = ~n10184 ;
  assign y829 = n10308 ;
  assign y830 = n10432 ;
  assign y831 = n10556 ;
  assign y832 = n10680 ;
  assign y833 = n10804 ;
  assign y834 = ~n10921 ;
  assign y835 = ~n10977 ;
  assign y836 = ~n11098 ;
  assign y837 = n11104 ;
  assign y838 = n11110 ;
  assign y839 = ~n11223 ;
  assign y840 = n1571 ;
  assign y841 = n11229 ;
  assign y842 = ~n11347 ;
  assign y843 = n11353 ;
  assign y844 = n11359 ;
  assign y845 = n11365 ;
  assign y846 = n11485 ;
  assign y847 = n11491 ;
  assign y848 = n11497 ;
  assign y849 = ~n11614 ;
  assign y850 = n11620 ;
  assign y851 = n11626 ;
  assign y852 = n11632 ;
  assign y853 = n11638 ;
  assign y854 = n11644 ;
  assign y855 = n11650 ;
  assign y856 = n11656 ;
  assign y857 = n11662 ;
  assign y858 = n11668 ;
  assign y859 = n11674 ;
  assign y860 = n11680 ;
  assign y861 = n11686 ;
  assign y862 = n11692 ;
  assign y863 = n11698 ;
  assign y864 = ~n11815 ;
  assign y865 = ~n11934 ;
  assign y866 = n11940 ;
  assign y867 = n11946 ;
  assign y868 = ~n12063 ;
  assign y869 = ~n12180 ;
  assign y870 = ~n12297 ;
  assign y871 = n12418 ;
  assign y872 = n12424 ;
  assign y873 = ~n12488 ;
  assign y874 = n12608 ;
  assign y875 = ~n12659 ;
  assign y876 = n12779 ;
  assign y877 = n12900 ;
  assign y878 = n12927 ;
  assign y879 = ~n13045 ;
  assign y880 = n13051 ;
  assign y881 = n13057 ;
  assign y882 = n13063 ;
  assign y883 = n13069 ;
  assign y884 = n13075 ;
  assign y885 = n13081 ;
  assign y886 = n13087 ;
  assign y887 = n13093 ;
  assign y888 = n13101 ;
  assign y889 = n13107 ;
  assign y890 = ~n13226 ;
  assign y891 = n13232 ;
  assign y892 = n13238 ;
  assign y893 = n13244 ;
  assign y894 = n13250 ;
  assign y895 = n13256 ;
  assign y896 = ~n13262 ;
  assign y897 = n8918 ;
  assign y898 = ~n13268 ;
  assign y899 = ~n13274 ;
  assign y900 = ~n13280 ;
  assign y901 = ~n13286 ;
  assign y902 = ~n13292 ;
  assign y903 = ~n13298 ;
  assign y904 = n13305 ;
  assign y905 = ~n13311 ;
  assign y906 = ~n13317 ;
  assign y907 = ~n13323 ;
  assign y908 = ~n13329 ;
  assign y909 = ~n13335 ;
  assign y910 = ~n13341 ;
  assign y911 = ~n13347 ;
  assign y912 = ~n13353 ;
  assign y913 = ~n13359 ;
  assign y914 = ~n13365 ;
  assign y915 = ~n13371 ;
  assign y916 = ~n13377 ;
  assign y917 = ~n13383 ;
  assign y918 = ~n13389 ;
  assign y919 = ~n13395 ;
  assign y920 = ~n13401 ;
  assign y921 = ~n13407 ;
  assign y922 = n13419 ;
  assign y923 = ~n13425 ;
  assign y924 = ~n13431 ;
  assign y925 = ~n13437 ;
  assign y926 = n13439 ;
  assign y927 = ~n13445 ;
  assign y928 = n13449 ;
  assign y929 = ~n13455 ;
  assign y930 = n13457 ;
  assign y931 = ~n13463 ;
  assign y932 = n13470 ;
  assign y933 = ~n13476 ;
  assign y934 = ~n13482 ;
  assign y935 = n13491 ;
  assign y936 = ~n13492 ;
  assign y937 = ~n13493 ;
  assign y938 = n13496 ;
  assign y939 = ~n13498 ;
  assign y940 = n13501 ;
  assign y941 = n13504 ;
  assign y942 = n13507 ;
  assign y943 = ~n13510 ;
  assign y944 = n13513 ;
  assign y945 = n13516 ;
  assign y946 = n13519 ;
  assign y947 = n13522 ;
  assign y948 = n13525 ;
  assign y949 = n13528 ;
  assign y950 = n2647 ;
  assign y951 = n13531 ;
  assign y952 = n13534 ;
  assign y953 = ~n13541 ;
  assign y954 = n9135 ;
  assign y955 = n13544 ;
  assign y956 = ~n13547 ;
  assign y957 = n13550 ;
  assign y958 = n13553 ;
  assign y959 = n13554 ;
  assign y960 = ~n13557 ;
  assign y961 = n13560 ;
  assign y962 = ~n13561 ;
  assign y963 = n13417 ;
  assign y964 = n13564 ;
  assign y965 = n13567 ;
  assign y966 = ~n13570 ;
  assign y967 = n13573 ;
  assign y968 = n13576 ;
  assign y969 = ~n13579 ;
  assign y970 = n13582 ;
  assign y971 = ~n13585 ;
  assign y972 = n13588 ;
  assign y973 = n13591 ;
  assign y974 = ~n13592 ;
  assign y975 = ~n5031 ;
  assign y976 = ~n13593 ;
  assign y977 = ~n13595 ;
  assign y978 = n12915 ;
  assign y979 = n13596 ;
  assign y980 = n9134 ;
  assign y981 = n13603 ;
  assign y982 = ~n13615 ;
  assign y983 = ~n13625 ;
  assign y984 = ~n13635 ;
  assign y985 = ~n13645 ;
  assign y986 = n13649 ;
  assign y987 = ~n13650 ;
  assign y988 = n8917 ;
  assign y989 = n13653 ;
  assign y990 = n13656 ;
  assign y991 = n13657 ;
  assign y992 = ~n13659 ;
  assign y993 = n13662 ;
  assign y994 = n13665 ;
  assign y995 = n13668 ;
  assign y996 = n13671 ;
  assign y997 = n13672 ;
  assign y998 = n13675 ;
  assign y999 = n13678 ;
  assign y1000 = n13681 ;
  assign y1001 = n13684 ;
  assign y1002 = n13687 ;
  assign y1003 = n13690 ;
  assign y1004 = n13693 ;
  assign y1005 = n13696 ;
  assign y1006 = n13699 ;
  assign y1007 = n13702 ;
  assign y1008 = n13705 ;
  assign y1009 = n13708 ;
  assign y1010 = n13711 ;
  assign y1011 = n13714 ;
  assign y1012 = n13717 ;
  assign y1013 = n13720 ;
  assign y1014 = n13723 ;
  assign y1015 = n13726 ;
  assign y1016 = n13729 ;
  assign y1017 = n13732 ;
  assign y1018 = n13735 ;
  assign y1019 = n13738 ;
  assign y1020 = n13741 ;
  assign y1021 = n13744 ;
  assign y1022 = n13747 ;
  assign y1023 = n13750 ;
  assign y1024 = n13753 ;
  assign y1025 = n13756 ;
  assign y1026 = n13759 ;
  assign y1027 = n13762 ;
  assign y1028 = n13765 ;
  assign y1029 = n13768 ;
  assign y1030 = n13771 ;
  assign y1031 = n13774 ;
  assign y1032 = n13777 ;
  assign y1033 = n13780 ;
  assign y1034 = n13783 ;
  assign y1035 = n13786 ;
  assign y1036 = n13789 ;
  assign y1037 = n13792 ;
  assign y1038 = ~n1209 ;
  assign y1039 = ~n13795 ;
  assign y1040 = ~n13798 ;
  assign y1041 = ~n13801 ;
  assign y1042 = ~n13804 ;
  assign y1043 = ~n13807 ;
  assign y1044 = ~n13810 ;
  assign y1045 = ~n13813 ;
  assign y1046 = ~n13816 ;
  assign y1047 = ~n13819 ;
  assign y1048 = ~n13822 ;
  assign y1049 = ~n6726 ;
  assign y1050 = ~n13825 ;
  assign y1051 = ~n13828 ;
  assign y1052 = ~n13831 ;
  assign y1053 = x67 ;
  assign y1054 = ~n13834 ;
  assign y1055 = ~n13837 ;
  assign y1056 = ~n13840 ;
  assign y1057 = ~n2691 ;
  assign y1058 = ~n13843 ;
  assign y1059 = ~n13846 ;
  assign y1060 = ~n13849 ;
  assign y1061 = ~n13852 ;
  assign y1062 = ~n13855 ;
  assign y1063 = n13863 ;
  assign y1064 = ~n13866 ;
  assign y1065 = ~n13869 ;
  assign y1066 = ~n13872 ;
  assign y1067 = ~n13875 ;
  assign y1068 = ~n13878 ;
  assign y1069 = ~n13881 ;
  assign y1070 = ~n13882 ;
  assign y1071 = ~n13885 ;
  assign y1072 = ~n13888 ;
  assign y1073 = ~n13891 ;
  assign y1074 = ~n13894 ;
  assign y1075 = ~n13897 ;
  assign y1076 = n13900 ;
  assign y1077 = n13903 ;
  assign y1078 = n13906 ;
  assign y1079 = n13909 ;
  assign y1080 = n13910 ;
  assign y1081 = n13913 ;
  assign y1082 = n13916 ;
  assign y1083 = n13919 ;
  assign y1084 = n13922 ;
  assign y1085 = n13925 ;
  assign y1086 = n13928 ;
  assign y1087 = n13931 ;
  assign y1088 = n13933 ;
  assign y1089 = n13936 ;
  assign y1090 = n13939 ;
  assign y1091 = n13942 ;
  assign y1092 = n13945 ;
  assign y1093 = n13948 ;
  assign y1094 = n13951 ;
  assign y1095 = n13954 ;
  assign y1096 = n13957 ;
  assign y1097 = n13960 ;
  assign y1098 = n13963 ;
  assign y1099 = n13966 ;
  assign y1100 = n13969 ;
  assign y1101 = ~n2655 ;
  assign y1102 = n13970 ;
  assign y1103 = n13974 ;
  assign y1104 = n13975 ;
  assign y1105 = ~n13978 ;
  assign y1106 = n13979 ;
  assign y1107 = n2643 ;
  assign y1108 = x1134 ;
  assign y1109 = x964 ;
  assign y1110 = ~x954 ;
  assign y1111 = x965 ;
  assign y1112 = n13982 ;
  assign y1113 = x991 ;
  assign y1114 = x985 ;
  assign y1115 = n13983 ;
  assign y1116 = n13984 ;
  assign y1117 = x1014 ;
  assign y1118 = n13985 ;
  assign y1119 = x1029 ;
  assign y1120 = x1004 ;
  assign y1121 = x1007 ;
  assign y1122 = n13986 ;
  assign y1123 = x1135 ;
  assign y1124 = n13987 ;
  assign y1125 = n13988 ;
  assign y1126 = n13989 ;
  assign y1127 = n13990 ;
  assign y1128 = n13991 ;
  assign y1129 = n13992 ;
  assign y1130 = ~x278 ;
  assign y1131 = n13993 ;
  assign y1132 = n13994 ;
  assign y1133 = ~n13995 ;
  assign y1134 = x1064 ;
  assign y1135 = n13996 ;
  assign y1136 = x299 ;
  assign y1137 = ~n13997 ;
  assign y1138 = x1075 ;
  assign y1139 = x1052 ;
  assign y1140 = x771 ;
  assign y1141 = x765 ;
  assign y1142 = x605 ;
  assign y1143 = x601 ;
  assign y1144 = x278 ;
  assign y1145 = x279 ;
  assign y1146 = ~x915 ;
  assign y1147 = ~x825 ;
  assign y1148 = ~x826 ;
  assign y1149 = ~x913 ;
  assign y1150 = ~x894 ;
  assign y1151 = ~x905 ;
  assign y1152 = x1095 ;
  assign y1153 = ~x890 ;
  assign y1154 = x1094 ;
  assign y1155 = ~x906 ;
  assign y1156 = ~x896 ;
  assign y1157 = ~x909 ;
  assign y1158 = ~x911 ;
  assign y1159 = ~x908 ;
  assign y1160 = ~x891 ;
  assign y1161 = ~x902 ;
  assign y1162 = ~x903 ;
  assign y1163 = ~x883 ;
  assign y1164 = ~x888 ;
  assign y1165 = ~x919 ;
  assign y1166 = ~x886 ;
  assign y1167 = ~x912 ;
  assign y1168 = ~x895 ;
  assign y1169 = ~x916 ;
  assign y1170 = ~x889 ;
  assign y1171 = ~x900 ;
  assign y1172 = ~x885 ;
  assign y1173 = ~x904 ;
  assign y1174 = ~x899 ;
  assign y1175 = ~x918 ;
  assign y1176 = ~x898 ;
  assign y1177 = ~x917 ;
  assign y1178 = ~x827 ;
  assign y1179 = ~x887 ;
  assign y1180 = ~x884 ;
  assign y1181 = ~x910 ;
  assign y1182 = ~x828 ;
  assign y1183 = ~x892 ;
  assign y1184 = x1187 ;
  assign y1185 = x1172 ;
  assign y1186 = x1170 ;
  assign y1187 = x1138 ;
  assign y1188 = x1177 ;
  assign y1189 = x1178 ;
  assign y1190 = x863 ;
  assign y1191 = x1203 ;
  assign y1192 = x1185 ;
  assign y1193 = x1171 ;
  assign y1194 = x1192 ;
  assign y1195 = x1137 ;
  assign y1196 = x1186 ;
  assign y1197 = x1165 ;
  assign y1198 = x1164 ;
  assign y1199 = x1098 ;
  assign y1200 = x1183 ;
  assign y1201 = x230 ;
  assign y1202 = x1169 ;
  assign y1203 = x1136 ;
  assign y1204 = x1181 ;
  assign y1205 = x849 ;
  assign y1206 = x1193 ;
  assign y1207 = x1182 ;
  assign y1208 = x1168 ;
  assign y1209 = x1175 ;
  assign y1210 = x1191 ;
  assign y1211 = x1099 ;
  assign y1212 = x1174 ;
  assign y1213 = x1179 ;
  assign y1214 = x1202 ;
  assign y1215 = x1176 ;
  assign y1216 = x1173 ;
  assign y1217 = x1201 ;
  assign y1218 = x1167 ;
  assign y1219 = x840 ;
  assign y1220 = x1189 ;
  assign y1221 = x1195 ;
  assign y1222 = x864 ;
  assign y1223 = x1190 ;
  assign y1224 = x1188 ;
  assign y1225 = x1180 ;
  assign y1226 = x1194 ;
  assign y1227 = x1097 ;
  assign y1228 = x1166 ;
  assign y1229 = x1200 ;
  assign y1230 = x1184 ;
endmodule
