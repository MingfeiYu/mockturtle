module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n465 , n466 , n467 , n468 , n469 , n470 , n472 , n473 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n497 , n498 , n499 , n500 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n593 , n594 , n595 , n596 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n686 , n687 , n688 , n689 , n694 , n695 , n696 , n697 , n698 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n764 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n776 , n777 , n778 , n779 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n888 , n889 , n890 , n891 , n892 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1025 , n1026 , n1027 , n1028 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1141 , n1142 , n1143 , n1144 , n1147 , n1148 , n1149 , n1150 , n1153 , n1154 , n1155 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1233 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1282 , n1283 , n1284 , n1285 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1426 , n1427 , n1428 , n1429 , n1430 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1630 , n1631 , n1632 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1707 , n1708 , n1709 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1740 , n1741 , n1742 , n1744 , n1745 , n1746 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1788 , n1789 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2028 , n2029 , n2030 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2052 , n2053 , n2054 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2093 , n2094 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2120 , n2121 , n2122 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2519 , n2520 , n2521 , n2522 , n2525 , n2526 , n2527 , n2528 , n2533 , n2534 , n2535 , n2536 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2600 , n2601 , n2602 , n2603 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2961 , n2962 , n2963 , n2964 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3081 , n3082 , n3083 , n3084 , n3085 , n3087 , n3090 , n3091 , n3092 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3147 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3459 , n3460 , n3461 , n3462 , n3465 , n3466 , n3467 , n3468 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3492 , n3493 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4968 , n4969 , n4970 , n4971 , n4972 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5954 , n5955 , n5958 , n5959 , n5960 , n5961 , n5962 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6169 , n6170 , n6171 , n6172 , n6173 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7531 , n7532 , n7533 , n7534 , n7535 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8601 , n8602 , n8603 , n8604 , n8605 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8864 , n8865 , n8866 , n8867 , n8868 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9928 , n9929 , n9930 , n9931 , n9932 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11386 , n11387 , n11388 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11961 , n11962 , n11963 , n11964 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12517 , n12518 , n12519 , n12520 , n12521 , n12523 , n12524 , n12525 , n12526 , n12527 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15553 , n15554 , n15555 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15718 , n15719 , n15720 , n15721 , n15722 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16645 , n16646 , n16647 , n16648 , n16649 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16676 , n16677 , n16678 , n16679 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17760 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17817 , n17818 , n17819 , n17820 , n17821 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19756 , n19757 , n19758 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19772 , n19773 , n19774 , n19775 , n19776 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20749 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22320 , n22321 , n22322 , n22323 , n22324 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23767 , n23768 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23972 , n23973 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24813 , n24814 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24833 , n24834 , n24835 , n24836 , n24837 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 ;
  assign n803 = x89 ^ x50 ;
  assign n804 = x98 ^ x58 ;
  assign n805 = n803 & n804 ;
  assign n806 = x88 ^ x42 ;
  assign n807 = x107 ^ x34 ;
  assign n808 = ~n806 & n807 ;
  assign n824 = n808 ^ n806 ;
  assign n835 = n805 & ~n824 ;
  assign n809 = n808 ^ n807 ;
  assign n820 = n809 ^ n806 ;
  assign n827 = n805 & n820 ;
  assign n821 = n805 ^ n804 ;
  assign n826 = n809 & n821 ;
  assign n828 = n827 ^ n826 ;
  assign n836 = n835 ^ n828 ;
  assign n802 = x121 ^ x26 ;
  assign n812 = x66 ^ x0 ;
  assign n1352 = ~n802 & n812 ;
  assign n1822 = n836 & n1352 ;
  assign n1353 = n1352 ^ n802 ;
  assign n1354 = n1353 ^ n812 ;
  assign n1813 = n826 ^ n807 ;
  assign n813 = n805 ^ n803 ;
  assign n825 = n813 & ~n824 ;
  assign n1814 = n1813 ^ n825 ;
  assign n814 = n808 & n813 ;
  assign n810 = n805 & n809 ;
  assign n855 = n814 ^ n810 ;
  assign n854 = n806 ^ n804 ;
  assign n856 = n855 ^ n854 ;
  assign n829 = n828 ^ n825 ;
  assign n822 = n820 & n821 ;
  assign n815 = n813 ^ n804 ;
  assign n816 = n808 & ~n815 ;
  assign n823 = n822 ^ n816 ;
  assign n830 = n829 ^ n823 ;
  assign n857 = n856 ^ n830 ;
  assign n851 = n809 & n813 ;
  assign n852 = n851 ^ n809 ;
  assign n850 = n826 ^ n810 ;
  assign n853 = n852 ^ n850 ;
  assign n858 = n857 ^ n853 ;
  assign n849 = n816 ^ n815 ;
  assign n859 = n858 ^ n849 ;
  assign n839 = n826 ^ n821 ;
  assign n833 = n807 ^ n803 ;
  assign n834 = n804 & n833 ;
  assign n837 = n836 ^ n834 ;
  assign n838 = n837 ^ n822 ;
  assign n840 = n839 ^ n838 ;
  assign n1798 = n859 ^ n840 ;
  assign n1815 = n1814 ^ n1798 ;
  assign n1816 = n1354 & ~n1815 ;
  assign n819 = n812 ^ n802 ;
  assign n1807 = n815 ^ n814 ;
  assign n1808 = n1807 ^ n853 ;
  assign n1809 = ~n802 & ~n1808 ;
  assign n1804 = n1798 ^ n851 ;
  assign n832 = n813 & n820 ;
  assign n1797 = n853 ^ n832 ;
  assign n1799 = n1798 ^ n1797 ;
  assign n1800 = n1797 ^ n802 ;
  assign n1801 = n819 & n1800 ;
  assign n1802 = n1801 ^ n802 ;
  assign n1803 = n1799 & ~n1802 ;
  assign n1805 = n1804 ^ n1803 ;
  assign n1806 = n1805 ^ n825 ;
  assign n1810 = n1809 ^ n1806 ;
  assign n1811 = ~n819 & n1810 ;
  assign n1812 = n1811 ^ n1809 ;
  assign n1817 = n1816 ^ n1812 ;
  assign n868 = n837 ^ n808 ;
  assign n817 = n816 ^ n814 ;
  assign n869 = n868 ^ n817 ;
  assign n1795 = n869 ^ n838 ;
  assign n1796 = ~n819 & n1795 ;
  assign n1818 = n1817 ^ n1796 ;
  assign n1819 = n1818 ^ n810 ;
  assign n1820 = n1819 ^ x3 ;
  assign n1788 = n817 ^ n810 ;
  assign n1789 = n1788 ^ n850 ;
  assign n1792 = n802 & n1789 ;
  assign n1793 = n1792 ^ n850 ;
  assign n1794 = ~n812 & n1793 ;
  assign n1821 = n1820 ^ n1794 ;
  assign n1823 = n1822 ^ n1821 ;
  assign n1824 = n1823 ^ x77 ;
  assign n629 = x92 ^ x62 ;
  assign n630 = x110 ^ x36 ;
  assign n710 = n629 & ~n630 ;
  assign n632 = x68 ^ x20 ;
  assign n638 = x93 ^ x28 ;
  assign n639 = x116 ^ x12 ;
  assign n640 = n638 & n639 ;
  assign n641 = n640 ^ n638 ;
  assign n656 = n632 & ~n641 ;
  assign n657 = n656 ^ n632 ;
  assign n633 = x86 ^ x4 ;
  assign n634 = n632 & ~n633 ;
  assign n658 = n657 ^ n634 ;
  assign n635 = n634 ^ n633 ;
  assign n636 = n635 ^ n632 ;
  assign n650 = n636 & n640 ;
  assign n651 = n650 ^ n640 ;
  assign n648 = ~n635 & ~n638 ;
  assign n649 = n648 ^ n635 ;
  assign n652 = n651 ^ n649 ;
  assign n645 = n633 ^ n632 ;
  assign n646 = n645 ^ n638 ;
  assign n647 = ~n632 & n646 ;
  assign n653 = n652 ^ n647 ;
  assign n654 = n653 ^ n638 ;
  assign n655 = n654 ^ n645 ;
  assign n659 = n658 ^ n655 ;
  assign n660 = n659 ^ n650 ;
  assign n661 = n660 ^ n640 ;
  assign n662 = n661 ^ n652 ;
  assign n637 = n636 ^ n633 ;
  assign n643 = n637 & n638 ;
  assign n642 = n637 & n641 ;
  assign n644 = n643 ^ n642 ;
  assign n663 = n662 ^ n644 ;
  assign n664 = n663 ^ n651 ;
  assign n665 = n664 ^ n642 ;
  assign n697 = n665 ^ n662 ;
  assign n666 = n640 ^ n639 ;
  assign n673 = n637 & n666 ;
  assign n1732 = n697 ^ n673 ;
  assign n1733 = n710 & n1732 ;
  assign n674 = n673 ^ n637 ;
  assign n675 = n674 ^ n643 ;
  assign n1724 = n675 ^ n663 ;
  assign n1725 = n1724 ^ n660 ;
  assign n1721 = n666 ^ n658 ;
  assign n669 = n639 ^ n633 ;
  assign n670 = ~n639 & ~n669 ;
  assign n1722 = n1721 ^ n670 ;
  assign n1413 = n648 ^ n632 ;
  assign n1414 = n1413 ^ n647 ;
  assign n1415 = n1414 ^ n650 ;
  assign n1723 = n1722 ^ n1415 ;
  assign n1726 = n1725 ^ n1723 ;
  assign n1727 = n1726 ^ n1415 ;
  assign n1728 = n629 & ~n1727 ;
  assign n1729 = n1728 ^ n1723 ;
  assign n1730 = n630 & ~n1729 ;
  assign n667 = n634 & n666 ;
  assign n1717 = n1415 ^ n667 ;
  assign n631 = n630 ^ n629 ;
  assign n1435 = ~n630 & n663 ;
  assign n1429 = n658 ^ n650 ;
  assign n676 = n675 ^ n648 ;
  assign n677 = n676 ^ n669 ;
  assign n671 = n670 ^ n638 ;
  assign n672 = ~n632 & n671 ;
  assign n678 = n677 ^ n672 ;
  assign n1430 = n1429 ^ n678 ;
  assign n1436 = n1435 ^ n1430 ;
  assign n1437 = ~n631 & n1436 ;
  assign n1718 = n1717 ^ n1437 ;
  assign n679 = n678 ^ n650 ;
  assign n668 = n667 ^ n665 ;
  assign n680 = n679 ^ n668 ;
  assign n1449 = n680 ^ n636 ;
  assign n1450 = n1449 ^ n1414 ;
  assign n1451 = n1450 ^ n1430 ;
  assign n1714 = ~n629 & ~n1451 ;
  assign n1715 = n1714 ^ n1430 ;
  assign n1716 = ~n630 & n1715 ;
  assign n1719 = n1718 ^ n1716 ;
  assign n1720 = n1719 ^ x45 ;
  assign n1731 = n1730 ^ n1720 ;
  assign n1734 = n1733 ^ n1731 ;
  assign n1707 = ~n630 & n665 ;
  assign n1708 = n1707 ^ n667 ;
  assign n1709 = ~n629 & n1708 ;
  assign n1735 = n1734 ^ n1709 ;
  assign n1736 = n1735 ^ x109 ;
  assign n406 = x96 ^ x32 ;
  assign n399 = x72 ^ x8 ;
  assign n400 = x82 ^ x0 ;
  assign n401 = n399 & n400 ;
  assign n402 = n401 ^ n400 ;
  assign n421 = n402 ^ n399 ;
  assign n394 = x65 ^ x16 ;
  assign n395 = x120 ^ x24 ;
  assign n396 = ~n394 & ~n395 ;
  assign n397 = n396 ^ n394 ;
  assign n398 = n397 ^ n395 ;
  assign n479 = n398 ^ n394 ;
  assign n480 = ~n421 & ~n479 ;
  assign n420 = n396 & n402 ;
  assign n1744 = n480 ^ n420 ;
  assign n435 = n396 & n401 ;
  assign n413 = ~n398 & n401 ;
  assign n436 = n435 ^ n413 ;
  assign n404 = ~n397 & n401 ;
  assign n434 = n404 ^ n401 ;
  assign n437 = n436 ^ n434 ;
  assign n481 = n480 ^ n437 ;
  assign n422 = n421 ^ n400 ;
  assign n427 = ~n398 & n422 ;
  assign n403 = ~n398 & n402 ;
  assign n428 = n427 ^ n403 ;
  assign n429 = n428 ^ n422 ;
  assign n425 = n396 & n422 ;
  assign n423 = ~n397 & n422 ;
  assign n424 = n423 ^ n403 ;
  assign n426 = n425 ^ n424 ;
  assign n430 = n429 ^ n426 ;
  assign n482 = n481 ^ n430 ;
  assign n483 = n482 ^ n479 ;
  assign n446 = n396 & ~n421 ;
  assign n484 = n483 ^ n446 ;
  assign n1745 = n1744 ^ n484 ;
  assign n407 = x105 ^ x58 ;
  assign n1748 = n1745 ^ n407 ;
  assign n1749 = ~n406 & ~n1748 ;
  assign n1750 = n1749 ^ n407 ;
  assign n1315 = n427 ^ n404 ;
  assign n431 = n430 ^ n420 ;
  assign n1751 = n1315 ^ n431 ;
  assign n1746 = n1745 ^ n1315 ;
  assign n1752 = n1751 ^ n1746 ;
  assign n438 = n437 ^ n425 ;
  assign n1753 = n1752 ^ n438 ;
  assign n1754 = n1750 & ~n1753 ;
  assign n1755 = n1754 ^ n1746 ;
  assign n439 = ~n397 & n402 ;
  assign n1756 = n1755 ^ n439 ;
  assign n1765 = n1756 ^ n436 ;
  assign n1763 = n483 ^ n401 ;
  assign n1764 = n407 & ~n1763 ;
  assign n1766 = n1765 ^ n1764 ;
  assign n1767 = ~n406 & ~n1766 ;
  assign n408 = ~n406 & n407 ;
  assign n409 = n408 ^ n406 ;
  assign n410 = n409 ^ n407 ;
  assign n411 = n410 ^ n406 ;
  assign n468 = n413 ^ n398 ;
  assign n469 = n468 ^ n428 ;
  assign n492 = n411 & ~n469 ;
  assign n472 = n439 ^ n424 ;
  assign n441 = n472 ^ n397 ;
  assign n405 = n404 ^ n403 ;
  assign n442 = n441 ^ n405 ;
  assign n491 = n408 & ~n442 ;
  assign n493 = n492 ^ n491 ;
  assign n1757 = n1756 ^ n493 ;
  assign n500 = n469 ^ n423 ;
  assign n503 = n406 & ~n500 ;
  assign n504 = n503 ^ n469 ;
  assign n505 = ~n407 & ~n504 ;
  assign n1758 = n1757 ^ n505 ;
  assign n470 = n469 ^ n439 ;
  assign n1737 = n481 ^ n470 ;
  assign n1740 = n407 & ~n1737 ;
  assign n1741 = n1740 ^ n481 ;
  assign n1742 = ~n406 & n1741 ;
  assign n1759 = n1758 ^ n1742 ;
  assign n1282 = ~n407 & n429 ;
  assign n1283 = n1282 ^ n430 ;
  assign n1284 = ~n406 & n1283 ;
  assign n1760 = n1759 ^ n1284 ;
  assign n515 = n408 & n425 ;
  assign n1761 = n1760 ^ n515 ;
  assign n1762 = n1761 ^ x53 ;
  assign n1768 = n1767 ^ n1762 ;
  assign n1769 = n1768 ^ x94 ;
  assign n1770 = n1736 & ~n1769 ;
  assign n1771 = n1770 ^ n1769 ;
  assign n330 = x104 ^ x60 ;
  assign n329 = x122 ^ x34 ;
  assign n318 = x90 ^ x10 ;
  assign n321 = x81 ^ x2 ;
  assign n322 = x64 ^ x26 ;
  assign n323 = n321 & n322 ;
  assign n346 = ~n318 & n323 ;
  assign n317 = x99 ^ x18 ;
  assign n319 = n317 & ~n318 ;
  assign n320 = n319 ^ n317 ;
  assign n332 = n320 ^ n318 ;
  assign n335 = n323 ^ n321 ;
  assign n336 = n332 & n335 ;
  assign n337 = n336 ^ n323 ;
  assign n347 = n346 ^ n337 ;
  assign n340 = n318 & n321 ;
  assign n348 = n347 ^ n340 ;
  assign n343 = n317 & n322 ;
  assign n344 = n343 ^ n320 ;
  assign n349 = n348 ^ n344 ;
  assign n345 = ~n321 & n344 ;
  assign n350 = n349 ^ n345 ;
  assign n339 = n318 ^ n317 ;
  assign n341 = n340 ^ n335 ;
  assign n342 = ~n339 & n341 ;
  assign n351 = n350 ^ n342 ;
  assign n352 = n351 ^ n336 ;
  assign n333 = n332 ^ n317 ;
  assign n334 = n321 & ~n333 ;
  assign n338 = n337 ^ n334 ;
  assign n353 = n352 ^ n338 ;
  assign n1150 = n353 ^ n348 ;
  assign n1153 = n329 & n1150 ;
  assign n1154 = n1153 ^ n348 ;
  assign n1155 = n330 & n1154 ;
  assign n1133 = n322 ^ n317 ;
  assign n1131 = n343 ^ n321 ;
  assign n1132 = n339 & n1131 ;
  assign n1134 = n1133 ^ n1132 ;
  assign n1135 = ~n329 & n1134 ;
  assign n1157 = n1155 ^ n1135 ;
  assign n324 = n323 ^ n322 ;
  assign n326 = n324 ^ n321 ;
  assign n327 = n319 & ~n326 ;
  assign n359 = n347 ^ n327 ;
  assign n357 = n322 ^ n321 ;
  assign n358 = n357 ^ n317 ;
  assign n360 = n359 ^ n358 ;
  assign n325 = n320 & n324 ;
  assign n328 = n327 ^ n325 ;
  assign n384 = n360 ^ n328 ;
  assign n361 = n324 & ~n333 ;
  assign n362 = n361 ^ n333 ;
  assign n363 = n362 ^ n334 ;
  assign n364 = n363 ^ n360 ;
  assign n354 = n353 ^ n342 ;
  assign n355 = n354 ^ n341 ;
  assign n365 = n364 ^ n355 ;
  assign n385 = n384 ^ n365 ;
  assign n382 = n322 ^ n318 ;
  assign n383 = n382 ^ n354 ;
  assign n386 = n385 ^ n383 ;
  assign n1144 = n386 ^ n363 ;
  assign n1147 = ~n329 & ~n1144 ;
  assign n1148 = n1147 ^ n363 ;
  assign n1149 = n330 & ~n1148 ;
  assign n1158 = n1157 ^ n1149 ;
  assign n1159 = n1158 ^ x37 ;
  assign n1119 = n348 ^ n327 ;
  assign n1120 = n1119 ^ n361 ;
  assign n1129 = n1120 ^ n355 ;
  assign n1130 = n1129 ^ n325 ;
  assign n1141 = n329 & n1130 ;
  assign n379 = ~n326 & n332 ;
  assign n1136 = n1135 ^ n379 ;
  assign n1142 = n1141 ^ n1136 ;
  assign n1143 = n330 & n1142 ;
  assign n1160 = n1159 ^ n1143 ;
  assign n331 = n330 ^ n329 ;
  assign n1121 = n1120 ^ n345 ;
  assign n1122 = n1121 ^ n354 ;
  assign n1118 = n351 ^ n345 ;
  assign n1123 = n1122 ^ n1118 ;
  assign n1126 = ~n329 & ~n1123 ;
  assign n1127 = n1126 ^ n1122 ;
  assign n1128 = n331 & ~n1127 ;
  assign n1161 = n1160 ^ n1128 ;
  assign n1673 = n1161 ^ x92 ;
  assign n1037 = x73 ^ x6 ;
  assign n1001 = x114 ^ x56 ;
  assign n1002 = x123 ^ x40 ;
  assign n1003 = n1001 & n1002 ;
  assign n1008 = n1003 ^ n1001 ;
  assign n998 = x112 ^ x32 ;
  assign n999 = x97 ^ x48 ;
  assign n1007 = ~n998 & n999 ;
  assign n1013 = n1007 ^ n998 ;
  assign n1053 = n1008 & ~n1013 ;
  assign n1025 = n1001 ^ n999 ;
  assign n1026 = n1002 ^ n998 ;
  assign n1000 = n999 ^ n998 ;
  assign n1005 = n1000 & n1002 ;
  assign n1027 = n1026 ^ n1005 ;
  assign n1028 = ~n1025 & n1027 ;
  assign n1009 = n1008 ^ n1002 ;
  assign n1010 = n1009 ^ n1001 ;
  assign n1011 = n1007 & n1010 ;
  assign n1004 = n1000 & n1003 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1012 = n1011 ^ n1006 ;
  assign n1043 = n1028 ^ n1012 ;
  assign n1018 = n1002 ^ n999 ;
  assign n1019 = n998 & n1018 ;
  assign n1020 = n1019 ^ n999 ;
  assign n1021 = ~n1001 & n1020 ;
  assign n1016 = n1007 & ~n1009 ;
  assign n1017 = n1016 ^ n1010 ;
  assign n1022 = n1021 ^ n1017 ;
  assign n1014 = n1013 ^ n999 ;
  assign n1015 = ~n1009 & n1014 ;
  assign n1023 = n1022 ^ n1015 ;
  assign n1044 = n1043 ^ n1023 ;
  assign n1054 = n1053 ^ n1044 ;
  assign n1030 = n1003 & n1007 ;
  assign n1693 = n1054 ^ n1030 ;
  assign n997 = x80 ^ x24 ;
  assign n1032 = n1021 ^ n1020 ;
  assign n1689 = n1032 ^ n1030 ;
  assign n1690 = n1689 ^ n1044 ;
  assign n1079 = n1007 ^ n999 ;
  assign n1051 = n1008 & n1014 ;
  assign n1052 = n1051 ^ n1008 ;
  assign n1055 = n1054 ^ n1052 ;
  assign n1056 = n1055 ^ n1004 ;
  assign n1080 = n1079 ^ n1056 ;
  assign n1059 = n1010 ^ n1006 ;
  assign n1060 = n1059 ^ n1022 ;
  assign n1058 = n1056 ^ n1044 ;
  assign n1061 = n1060 ^ n1058 ;
  assign n1057 = n1056 ^ n1032 ;
  assign n1062 = n1061 ^ n1057 ;
  assign n1081 = n1080 ^ n1062 ;
  assign n1691 = n1690 ^ n1081 ;
  assign n1692 = n997 & n1691 ;
  assign n1694 = n1693 ^ n1692 ;
  assign n1695 = ~n1037 & n1694 ;
  assign n1069 = ~n997 & n1037 ;
  assign n1089 = n1069 ^ n997 ;
  assign n1678 = n1016 & n1089 ;
  assign n1677 = n1021 ^ n1015 ;
  assign n1679 = n1678 ^ n1677 ;
  assign n1680 = n1679 ^ n1069 ;
  assign n1685 = n1021 & ~n1089 ;
  assign n1386 = n1055 ^ n1003 ;
  assign n1387 = n1386 ^ n1032 ;
  assign n1682 = n1387 ^ n1055 ;
  assign n1683 = n1682 ^ n1057 ;
  assign n1681 = n1679 ^ n1044 ;
  assign n1684 = n1683 ^ n1681 ;
  assign n1686 = n1685 ^ n1684 ;
  assign n1687 = n1680 & ~n1686 ;
  assign n1688 = n1687 ^ n1069 ;
  assign n1696 = n1695 ^ n1688 ;
  assign n1929 = n1037 ^ n997 ;
  assign n1379 = n1051 & ~n1929 ;
  assign n1697 = n1696 ^ n1379 ;
  assign n1388 = n1387 ^ n1060 ;
  assign n1391 = ~n1037 & n1388 ;
  assign n1392 = n1391 ^ n1387 ;
  assign n1393 = n997 & n1392 ;
  assign n1698 = n1697 ^ n1393 ;
  assign n1033 = n1028 ^ n1025 ;
  assign n1034 = n1033 ^ n1032 ;
  assign n1031 = n1030 ^ n1004 ;
  assign n1035 = n1034 ^ n1031 ;
  assign n1036 = n1044 ^ n1035 ;
  assign n1040 = ~n1036 & n1037 ;
  assign n1041 = n1040 ^ n1035 ;
  assign n1042 = n997 & ~n1041 ;
  assign n1699 = n1698 ^ n1042 ;
  assign n1700 = n1699 ^ x61 ;
  assign n1088 = n1069 ^ n1037 ;
  assign n1674 = n1055 ^ n1006 ;
  assign n1366 = n1081 ^ n1022 ;
  assign n1675 = n1674 ^ n1366 ;
  assign n1676 = n1088 & n1675 ;
  assign n1701 = n1700 ^ n1676 ;
  assign n1702 = n1701 ^ x83 ;
  assign n1703 = n1673 & n1702 ;
  assign n1774 = n1703 ^ n1702 ;
  assign n1840 = n1774 ^ n1673 ;
  assign n1850 = ~n1771 & ~n1840 ;
  assign n1849 = n1770 & ~n1840 ;
  assign n1851 = n1850 ^ n1849 ;
  assign n1775 = n1770 ^ n1736 ;
  assign n1841 = n1775 & ~n1840 ;
  assign n1848 = n1841 ^ n1840 ;
  assign n1852 = n1851 ^ n1848 ;
  assign n1838 = n1703 ^ n1673 ;
  assign n1839 = n1770 & n1838 ;
  assign n1772 = n1771 ^ n1736 ;
  assign n1773 = n1703 & n1772 ;
  assign n1844 = n1839 ^ n1773 ;
  assign n1776 = n1774 & n1775 ;
  assign n1845 = n1844 ^ n1776 ;
  assign n1853 = n1852 ^ n1845 ;
  assign n3811 = n1853 ^ n1850 ;
  assign n1863 = n1852 ^ n1772 ;
  assign n1781 = n1770 & n1774 ;
  assign n1777 = n1703 & ~n1771 ;
  assign n1782 = n1781 ^ n1777 ;
  assign n1783 = n1782 ^ n1774 ;
  assign n1779 = ~n1771 & n1774 ;
  assign n1778 = n1777 ^ n1776 ;
  assign n1780 = n1779 ^ n1778 ;
  assign n1784 = n1783 ^ n1780 ;
  assign n1785 = n1784 ^ n1773 ;
  assign n1864 = n1863 ^ n1785 ;
  assign n1830 = n1703 & n1770 ;
  assign n1856 = n1830 ^ n1778 ;
  assign n1857 = n1856 ^ n1845 ;
  assign n1854 = n1839 ^ n1838 ;
  assign n1855 = n1854 ^ n1673 ;
  assign n1858 = n1857 ^ n1855 ;
  assign n1859 = n1858 ^ n1779 ;
  assign n1860 = n1859 ^ n1773 ;
  assign n1861 = n1860 ^ n1853 ;
  assign n1842 = n1841 ^ n1839 ;
  assign n1843 = n1842 ^ n1781 ;
  assign n1846 = n1845 ^ n1843 ;
  assign n1836 = n1702 ^ n1673 ;
  assign n1837 = n1836 ^ n1769 ;
  assign n1847 = n1846 ^ n1837 ;
  assign n1862 = n1861 ^ n1847 ;
  assign n1865 = n1864 ^ n1862 ;
  assign n1866 = n1865 ^ n1854 ;
  assign n3625 = n1866 ^ n1862 ;
  assign n3812 = n3811 ^ n3625 ;
  assign n3813 = n1824 & n3812 ;
  assign n129 = x94 ^ x56 ;
  assign n140 = x108 ^ x38 ;
  assign n146 = n129 & n140 ;
  assign n134 = x118 ^ x6 ;
  assign n130 = x125 ^ x14 ;
  assign n131 = x77 ^ x30 ;
  assign n133 = x76 ^ x22 ;
  assign n137 = ~n131 & n133 ;
  assign n138 = n130 & n137 ;
  assign n166 = n138 ^ n137 ;
  assign n167 = ~n134 & n166 ;
  assign n204 = n167 ^ n166 ;
  assign n154 = ~n133 & n134 ;
  assign n155 = n131 & n154 ;
  assign n156 = n155 ^ n154 ;
  assign n153 = n137 ^ n131 ;
  assign n157 = n156 ^ n153 ;
  assign n158 = n130 & ~n157 ;
  assign n159 = n158 ^ n157 ;
  assign n205 = n204 ^ n159 ;
  assign n955 = n146 & ~n205 ;
  assign n151 = ~n134 & n138 ;
  assign n947 = n155 ^ n151 ;
  assign n132 = n130 & n131 ;
  assign n181 = n132 & n133 ;
  assign n180 = n137 ^ n133 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = ~n134 & n182 ;
  assign n184 = n183 ^ n181 ;
  assign n168 = ~n130 & n156 ;
  assign n169 = n168 ^ n156 ;
  assign n170 = n169 ^ n167 ;
  assign n185 = n184 ^ n170 ;
  assign n174 = n138 ^ n130 ;
  assign n175 = n174 ^ n133 ;
  assign n176 = n175 ^ n138 ;
  assign n177 = ~n134 & n176 ;
  assign n178 = n177 ^ n174 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n132 & n135 ;
  assign n179 = n178 ^ n136 ;
  assign n186 = n185 ^ n179 ;
  assign n948 = n947 ^ n186 ;
  assign n943 = n182 ^ n138 ;
  assign n944 = n943 ^ n170 ;
  assign n187 = n155 ^ n136 ;
  assign n188 = n187 ^ n186 ;
  assign n945 = n944 ^ n188 ;
  assign n946 = ~n140 & n945 ;
  assign n949 = n948 ^ n946 ;
  assign n147 = n140 ^ n129 ;
  assign n148 = n147 ^ n146 ;
  assign n152 = n151 ^ n138 ;
  assign n171 = n170 ^ n152 ;
  assign n941 = n183 ^ n171 ;
  assign n942 = ~n148 & n941 ;
  assign n950 = n949 ^ n942 ;
  assign n149 = n136 ^ n132 ;
  assign n934 = n204 ^ n149 ;
  assign n935 = n934 ^ n136 ;
  assign n938 = n140 & n935 ;
  assign n939 = n938 ^ n136 ;
  assign n940 = ~n129 & n939 ;
  assign n951 = n950 ^ n940 ;
  assign n924 = n167 ^ n158 ;
  assign n952 = n951 ^ n924 ;
  assign n200 = n132 ^ n131 ;
  assign n201 = n200 ^ n182 ;
  assign n202 = n201 ^ n188 ;
  assign n932 = n202 ^ n136 ;
  assign n933 = ~n146 & n932 ;
  assign n953 = n952 ^ n933 ;
  assign n925 = n924 ^ n148 ;
  assign n926 = n156 ^ n146 ;
  assign n929 = ~n924 & ~n926 ;
  assign n930 = n929 ^ n146 ;
  assign n931 = ~n925 & ~n930 ;
  assign n954 = n953 ^ n931 ;
  assign n956 = n955 ^ n954 ;
  assign n957 = n956 ^ x29 ;
  assign n162 = n158 ^ n152 ;
  assign n163 = n162 ^ n149 ;
  assign n164 = n140 & n163 ;
  assign n165 = n164 ^ n149 ;
  assign n923 = n147 & n165 ;
  assign n958 = n957 ^ n923 ;
  assign n1672 = n958 ^ x126 ;
  assign n1831 = ~n1672 & n1824 ;
  assign n1832 = n1831 ^ n1672 ;
  assign n1833 = n1830 & ~n1832 ;
  assign n1827 = n1785 & ~n1824 ;
  assign n1828 = n1827 ^ n1784 ;
  assign n1829 = ~n1672 & n1828 ;
  assign n1834 = n1833 ^ n1829 ;
  assign n3817 = n3813 ^ n1834 ;
  assign n3462 = n1830 ^ n1782 ;
  assign n3465 = n1824 & n3462 ;
  assign n3466 = n3465 ^ n1782 ;
  assign n3467 = n1672 & n3466 ;
  assign n3818 = n3817 ^ n3467 ;
  assign n3819 = n3818 ^ x18 ;
  assign n1835 = n1824 ^ n1672 ;
  assign n3450 = n1849 ^ n1842 ;
  assign n3451 = n3450 ^ n1864 ;
  assign n3814 = n3813 ^ n3451 ;
  assign n1883 = n1865 ^ n1841 ;
  assign n1884 = n1883 ^ n1850 ;
  assign n3809 = n1884 ^ n1838 ;
  assign n3810 = ~n1824 & n3809 ;
  assign n3815 = n3814 ^ n3810 ;
  assign n3816 = n1835 & ~n3815 ;
  assign n3820 = n3819 ^ n3816 ;
  assign n3808 = n1780 & n1831 ;
  assign n3821 = n3820 ^ n3808 ;
  assign n3442 = n1858 ^ n1784 ;
  assign n3802 = n3442 ^ n1847 ;
  assign n3805 = n1672 & n3802 ;
  assign n3806 = n3805 ^ n1847 ;
  assign n3807 = ~n1824 & n3806 ;
  assign n3822 = n3821 ^ n3807 ;
  assign n3823 = n3822 ^ x104 ;
  assign n2057 = n482 ^ n435 ;
  assign n2058 = n2057 ^ n409 ;
  assign n2059 = ~n472 & n2058 ;
  assign n2060 = n2059 ^ n409 ;
  assign n494 = n442 ^ n427 ;
  assign n497 = n406 & ~n494 ;
  assign n498 = n497 ^ n427 ;
  assign n499 = ~n407 & n498 ;
  assign n2062 = n499 ^ n472 ;
  assign n2061 = n499 ^ n411 ;
  assign n2063 = n2062 ^ n2061 ;
  assign n2064 = ~n2060 & n2063 ;
  assign n2065 = n2064 ^ n2061 ;
  assign n433 = n407 ^ n406 ;
  assign n2048 = n438 ^ n404 ;
  assign n2047 = n435 ^ n423 ;
  assign n2049 = n2048 ^ n2047 ;
  assign n2052 = n406 & n2049 ;
  assign n2053 = n2052 ^ n2047 ;
  assign n2054 = n433 & n2053 ;
  assign n2066 = n2065 ^ n2054 ;
  assign n1292 = n410 & n428 ;
  assign n2067 = n2066 ^ n1292 ;
  assign n485 = n484 ^ n413 ;
  assign n488 = n406 & ~n485 ;
  assign n489 = n488 ^ n413 ;
  assign n490 = n433 & n489 ;
  assign n2068 = n2067 ^ n490 ;
  assign n1285 = n484 ^ n431 ;
  assign n1288 = ~n407 & ~n1285 ;
  assign n1289 = n1288 ^ n484 ;
  assign n1290 = ~n406 & ~n1289 ;
  assign n1291 = n1290 ^ n492 ;
  assign n2069 = n2068 ^ n1291 ;
  assign n2070 = n2069 ^ n1742 ;
  assign n2071 = n2070 ^ n515 ;
  assign n2072 = n2071 ^ x27 ;
  assign n2073 = n2072 ^ x113 ;
  assign n520 = x67 ^ x28 ;
  assign n521 = x85 ^ x2 ;
  assign n522 = ~n520 & n521 ;
  assign n523 = n522 ^ n520 ;
  assign n615 = n523 ^ n521 ;
  assign n616 = n615 ^ n520 ;
  assign n524 = x100 ^ x36 ;
  assign n526 = x117 ^ x44 ;
  assign n536 = ~n524 & n526 ;
  assign n525 = x102 ^ x52 ;
  assign n527 = ~n525 & n526 ;
  assign n528 = n524 & n527 ;
  assign n529 = n528 ^ n527 ;
  assign n558 = n536 ^ n529 ;
  assign n555 = n526 ^ n525 ;
  assign n556 = n526 ^ n524 ;
  assign n557 = ~n555 & n556 ;
  assign n559 = n558 ^ n557 ;
  assign n530 = x91 ^ x60 ;
  assign n543 = n524 & n530 ;
  assign n544 = ~n526 & n543 ;
  assign n545 = n525 & n544 ;
  assign n546 = n545 ^ n544 ;
  assign n564 = n559 ^ n546 ;
  assign n537 = n525 & ~n530 ;
  assign n540 = n524 & n537 ;
  assign n562 = n526 & n540 ;
  assign n563 = n562 ^ n540 ;
  assign n565 = n564 ^ n563 ;
  assign n554 = n527 ^ n525 ;
  assign n560 = n559 ^ n554 ;
  assign n552 = n536 ^ n524 ;
  assign n538 = n536 & n537 ;
  assign n539 = n538 ^ n537 ;
  assign n541 = n540 ^ n539 ;
  assign n553 = n552 ^ n541 ;
  assign n561 = n560 ^ n553 ;
  assign n566 = n565 ^ n561 ;
  assign n549 = n530 ^ n524 ;
  assign n550 = n549 ^ n526 ;
  assign n551 = ~n526 & n550 ;
  assign n567 = n566 ^ n551 ;
  assign n578 = n567 ^ n560 ;
  assign n2042 = n578 ^ n546 ;
  assign n576 = n562 ^ n561 ;
  assign n2043 = n2042 ^ n576 ;
  assign n2044 = n616 & ~n2043 ;
  assign n614 = n558 ^ n538 ;
  assign n568 = n567 ^ n563 ;
  assign n2019 = n614 ^ n568 ;
  assign n579 = n544 ^ n543 ;
  assign n535 = n528 & ~n530 ;
  assign n572 = n535 ^ n528 ;
  assign n580 = n579 ^ n572 ;
  assign n542 = n541 ^ n535 ;
  assign n2017 = n580 ^ n542 ;
  assign n531 = n529 & ~n530 ;
  assign n532 = n531 ^ n529 ;
  assign n587 = n568 ^ n532 ;
  assign n588 = n587 ^ n562 ;
  assign n2018 = n2017 ^ n588 ;
  assign n2020 = n2019 ^ n2018 ;
  assign n2021 = n521 & n2020 ;
  assign n2022 = n2021 ^ n2019 ;
  assign n1164 = n564 ^ n531 ;
  assign n1165 = n616 & n1164 ;
  assign n624 = n538 & n615 ;
  assign n1166 = n1165 ^ n624 ;
  assign n2036 = n2022 ^ n1166 ;
  assign n534 = n521 ^ n520 ;
  assign n2033 = n520 & n565 ;
  assign n2034 = n2033 ^ n564 ;
  assign n2035 = ~n534 & n2034 ;
  assign n2037 = n2036 ^ n2035 ;
  assign n610 = n521 & n546 ;
  assign n602 = n580 ^ n561 ;
  assign n603 = n602 ^ n572 ;
  assign n604 = ~n520 & n603 ;
  assign n605 = n604 ^ n572 ;
  assign n611 = n610 ^ n605 ;
  assign n612 = n534 & n611 ;
  assign n613 = n612 ^ n605 ;
  assign n2038 = n2037 ^ n613 ;
  assign n573 = n572 ^ n538 ;
  assign n596 = n573 ^ n564 ;
  assign n599 = ~n520 & n596 ;
  assign n600 = n599 ^ n564 ;
  assign n601 = ~n521 & n600 ;
  assign n2039 = n2038 ^ n601 ;
  assign n2040 = n2039 ^ x1 ;
  assign n1188 = n614 ^ n572 ;
  assign n1189 = n1188 ^ n532 ;
  assign n1190 = n1189 ^ n578 ;
  assign n2023 = n2022 ^ n1190 ;
  assign n570 = n545 ^ n535 ;
  assign n2024 = n2023 ^ n570 ;
  assign n2025 = n2024 ^ n2022 ;
  assign n2028 = ~n521 & ~n2025 ;
  assign n2029 = n2028 ^ n2022 ;
  assign n2030 = n520 & n2029 ;
  assign n2041 = n2040 ^ n2030 ;
  assign n2045 = n2044 ^ n2041 ;
  assign n2046 = n2045 ^ x123 ;
  assign n1919 = ~n329 & n385 ;
  assign n1920 = n1919 ^ n365 ;
  assign n1924 = n1920 ^ n1155 ;
  assign n1925 = n1924 ^ n1149 ;
  assign n1926 = n1925 ^ x51 ;
  assign n1918 = n352 ^ n328 ;
  assign n1921 = n1920 ^ n1918 ;
  assign n1915 = n379 ^ n352 ;
  assign n356 = n355 ^ n346 ;
  assign n1916 = n1915 ^ n356 ;
  assign n1917 = ~n329 & n1916 ;
  assign n1922 = n1921 ^ n1917 ;
  assign n1923 = n330 & ~n1922 ;
  assign n1927 = n1926 ^ n1923 ;
  assign n1928 = n1927 ^ x81 ;
  assign n1082 = n1081 ^ n1011 ;
  assign n1932 = n1082 ^ n1032 ;
  assign n1930 = n1366 ^ n1012 ;
  assign n1931 = n1930 ^ n1051 ;
  assign n1933 = n1932 ^ n1931 ;
  assign n1934 = n1037 & n1933 ;
  assign n1935 = n1934 ^ n1931 ;
  assign n1070 = n1035 ^ n1015 ;
  assign n1071 = n1069 & ~n1070 ;
  assign n1947 = n1935 ^ n1071 ;
  assign n1944 = n1053 ^ n1015 ;
  assign n1945 = n1944 ^ n1683 ;
  assign n1946 = ~n1089 & n1945 ;
  assign n1948 = n1947 ^ n1946 ;
  assign n1937 = n1935 ^ n1021 ;
  assign n1936 = n1935 ^ n1016 ;
  assign n1938 = n1937 ^ n1936 ;
  assign n1941 = ~n1037 & n1938 ;
  assign n1942 = n1941 ^ n1937 ;
  assign n1943 = ~n1929 & n1942 ;
  assign n1949 = n1948 ^ n1943 ;
  assign n1094 = n1053 & n1088 ;
  assign n1950 = n1949 ^ n1094 ;
  assign n1951 = n1950 ^ n1393 ;
  assign n1045 = n1044 ^ n1012 ;
  assign n1048 = n997 & n1045 ;
  assign n1049 = n1048 ^ n1012 ;
  assign n1050 = ~n1037 & n1049 ;
  assign n1952 = n1951 ^ n1050 ;
  assign n1953 = n1952 ^ n1042 ;
  assign n1954 = ~n1030 & ~n1953 ;
  assign n1955 = n1954 ^ x59 ;
  assign n1956 = n1955 ^ x90 ;
  assign n1957 = ~n1928 & n1956 ;
  assign n2007 = n1957 ^ n1928 ;
  assign n1408 = n666 ^ n638 ;
  assign n1438 = n1430 ^ n1408 ;
  assign n1439 = n1438 ^ n676 ;
  assign n1440 = n710 ^ n673 ;
  assign n1441 = n1440 ^ n630 ;
  assign n1442 = ~n1439 & n1441 ;
  assign n1443 = n1442 ^ n673 ;
  assign n1444 = n1439 ^ n710 ;
  assign n1445 = n1444 ^ n629 ;
  assign n1446 = n1443 & ~n1445 ;
  assign n1447 = n1446 ^ n1439 ;
  assign n1975 = n1447 ^ n667 ;
  assign n1976 = n1975 ^ n1716 ;
  assign n1452 = n1451 ^ n665 ;
  assign n1453 = n1452 ^ n1408 ;
  assign n1454 = n629 & n1453 ;
  assign n1455 = n1454 ^ n675 ;
  assign n1456 = ~n630 & n1455 ;
  assign n1977 = n1976 ^ n1456 ;
  assign n1978 = n1977 ^ x43 ;
  assign n701 = n657 ^ n642 ;
  assign n1416 = n1415 ^ n701 ;
  assign n1968 = n1416 ^ n680 ;
  assign n1966 = n663 ^ n642 ;
  assign n1967 = n1966 ^ n701 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n1972 = n630 & ~n1969 ;
  assign n1973 = n1972 ^ n1967 ;
  assign n1974 = ~n631 & n1973 ;
  assign n1979 = n1978 ^ n1974 ;
  assign n1965 = n629 & ~n660 ;
  assign n1980 = n1979 ^ n1965 ;
  assign n1960 = n643 ^ n639 ;
  assign n1961 = n1960 ^ n646 ;
  assign n1962 = ~n629 & n1961 ;
  assign n1963 = n1962 ^ n667 ;
  assign n1964 = n631 & n1963 ;
  assign n1981 = n1980 ^ n1964 ;
  assign n1982 = n1981 ^ x80 ;
  assign n221 = x78 ^ x38 ;
  assign n222 = x84 ^ x62 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = n223 ^ n222 ;
  assign n225 = x101 ^ x54 ;
  assign n226 = x126 ^ x46 ;
  assign n227 = ~n225 & n226 ;
  assign n228 = n227 ^ n225 ;
  assign n236 = n228 ^ n226 ;
  assign n252 = ~n224 & n236 ;
  assign n237 = n223 & n236 ;
  assign n231 = ~n224 & n227 ;
  assign n238 = n237 ^ n231 ;
  assign n234 = n227 ^ n226 ;
  assign n235 = n223 & n234 ;
  assign n239 = n238 ^ n235 ;
  assign n230 = n223 & n227 ;
  assign n232 = n231 ^ n230 ;
  assign n233 = n232 ^ n223 ;
  assign n240 = n239 ^ n233 ;
  assign n253 = n252 ^ n240 ;
  assign n266 = n253 ^ n230 ;
  assign n278 = n266 ^ n222 ;
  assign n243 = n224 ^ n221 ;
  assign n244 = n243 ^ n222 ;
  assign n256 = n234 & n244 ;
  assign n257 = n256 ^ n235 ;
  assign n258 = n257 ^ n234 ;
  assign n254 = n253 ^ n235 ;
  assign n229 = ~n224 & ~n228 ;
  assign n249 = n237 ^ n229 ;
  assign n250 = n249 ^ n232 ;
  assign n251 = n250 ^ n222 ;
  assign n255 = n254 ^ n251 ;
  assign n259 = n258 ^ n255 ;
  assign n277 = n259 ^ n233 ;
  assign n279 = n278 ^ n277 ;
  assign n275 = n226 ^ n222 ;
  assign n276 = n275 ^ n221 ;
  assign n280 = n279 ^ n276 ;
  assign n220 = x83 ^ x30 ;
  assign n269 = x124 ^ x4 ;
  assign n281 = n220 & n269 ;
  assign n282 = n281 ^ n269 ;
  assign n2001 = n280 & n282 ;
  assign n1989 = n277 ^ n238 ;
  assign n304 = n236 & n244 ;
  assign n1990 = n1989 ^ n304 ;
  assign n260 = n259 ^ n243 ;
  assign n247 = n236 & n243 ;
  assign n245 = n227 & n244 ;
  assign n242 = n232 ^ n227 ;
  assign n246 = n245 ^ n242 ;
  assign n248 = n247 ^ n246 ;
  assign n261 = n260 ^ n248 ;
  assign n987 = n261 ^ n256 ;
  assign n988 = n987 ^ n246 ;
  assign n1991 = n1990 ^ n988 ;
  assign n1992 = ~n220 & n1991 ;
  assign n1993 = n1992 ^ n277 ;
  assign n298 = n281 ^ n220 ;
  assign n262 = n261 ^ n228 ;
  assign n241 = n240 ^ n229 ;
  assign n263 = n262 ^ n241 ;
  assign n299 = n263 ^ n247 ;
  assign n300 = n298 & n299 ;
  assign n1996 = n1993 ^ n300 ;
  assign n285 = n255 ^ n252 ;
  assign n286 = n269 ^ n252 ;
  assign n287 = n286 ^ n252 ;
  assign n288 = ~n285 & ~n287 ;
  assign n289 = n288 ^ n252 ;
  assign n290 = n220 & n289 ;
  assign n1997 = n1996 ^ n290 ;
  assign n1998 = n1997 ^ x35 ;
  assign n1986 = n304 ^ n246 ;
  assign n1984 = n243 ^ n230 ;
  assign n1985 = n1984 ^ n248 ;
  assign n1987 = n1986 ^ n1985 ;
  assign n1988 = n220 & n1987 ;
  assign n1994 = n1993 ^ n1988 ;
  assign n1995 = n269 & ~n1994 ;
  assign n1999 = n1998 ^ n1995 ;
  assign n309 = n255 ^ n240 ;
  assign n977 = n269 ^ n220 ;
  assign n1983 = ~n309 & ~n977 ;
  assign n2000 = n1999 ^ n1983 ;
  assign n2002 = n2001 ^ n2000 ;
  assign n2003 = n2002 ^ x99 ;
  assign n2004 = n1982 & n2003 ;
  assign n2005 = n2004 ^ n2003 ;
  assign n2011 = n2005 ^ n1982 ;
  assign n2083 = n2011 ^ n2003 ;
  assign n2093 = ~n2007 & n2083 ;
  assign n2008 = n2004 & ~n2007 ;
  assign n2094 = n2093 ^ n2008 ;
  assign n2082 = ~n2007 & ~n2011 ;
  assign n2115 = n2094 ^ n2082 ;
  assign n2116 = n2115 ^ n2007 ;
  assign n1958 = n1957 ^ n1956 ;
  assign n1959 = n1958 ^ n1928 ;
  assign n2012 = n1959 & ~n2011 ;
  assign n2013 = n2012 ^ n2008 ;
  assign n2010 = n1959 & n2004 ;
  assign n2014 = n2013 ^ n2010 ;
  assign n2015 = n2014 ^ n1959 ;
  assign n2006 = n1959 & n2005 ;
  assign n2009 = n2008 ^ n2006 ;
  assign n2016 = n2015 ^ n2009 ;
  assign n2155 = n2116 ^ n2016 ;
  assign n2160 = ~n2046 & ~n2155 ;
  assign n2161 = n2160 ^ n2016 ;
  assign n2162 = n2073 & n2161 ;
  assign n2101 = n1957 & n2004 ;
  assign n2084 = n1958 & n2083 ;
  assign n2098 = n2084 ^ n2016 ;
  assign n2097 = n2093 ^ n2083 ;
  assign n2099 = n2098 ^ n2097 ;
  assign n2086 = n2082 ^ n2010 ;
  assign n2087 = n2086 ^ n2012 ;
  assign n2085 = n2084 ^ n2082 ;
  assign n2088 = n2087 ^ n2085 ;
  assign n2078 = n2003 ^ n1982 ;
  assign n2079 = n2078 ^ n1928 ;
  assign n2080 = n2079 ^ n1956 ;
  assign n2081 = n1928 & n2080 ;
  assign n2089 = n2088 ^ n2081 ;
  assign n2090 = n2089 ^ n2006 ;
  assign n2091 = n2090 ^ n2005 ;
  assign n2096 = n2116 ^ n2091 ;
  assign n2100 = n2099 ^ n2096 ;
  assign n2102 = n2101 ^ n2100 ;
  assign n3152 = n2046 & ~n2102 ;
  assign n3153 = n3152 ^ n2101 ;
  assign n3154 = n2073 & n3153 ;
  assign n2074 = n2046 & n2073 ;
  assign n2075 = n2074 ^ n2046 ;
  assign n3127 = n2075 & n2084 ;
  assign n2104 = n2101 ^ n2010 ;
  assign n2149 = n2046 & n2104 ;
  assign n2150 = n2149 ^ n2010 ;
  assign n2151 = ~n2073 & n2150 ;
  assign n3128 = n3127 ^ n2151 ;
  assign n3133 = n2014 ^ n2006 ;
  assign n2103 = n2102 ^ n1957 ;
  assign n3134 = n3133 ^ n2103 ;
  assign n3135 = n2046 & ~n3134 ;
  assign n3136 = n3135 ^ n2090 ;
  assign n3131 = n2096 ^ n2012 ;
  assign n2108 = n2100 ^ n2085 ;
  assign n2105 = n2008 ^ n2004 ;
  assign n2106 = n2105 ^ n2104 ;
  assign n2107 = n2106 ^ n2009 ;
  assign n2109 = n2108 ^ n2107 ;
  assign n2110 = n2109 ^ n2080 ;
  assign n2111 = n2110 ^ n2098 ;
  assign n2644 = n2111 ^ n2106 ;
  assign n3132 = n3131 ^ n2644 ;
  assign n3137 = n3136 ^ n3132 ;
  assign n2130 = n2099 ^ n2089 ;
  assign n3129 = n2130 ^ n2008 ;
  assign n3130 = n3129 ^ n2082 ;
  assign n3138 = n3137 ^ n3130 ;
  assign n3139 = n3138 ^ n3136 ;
  assign n3140 = ~n2046 & ~n3139 ;
  assign n3141 = n3140 ^ n3137 ;
  assign n3142 = ~n2073 & ~n3141 ;
  assign n3143 = n3142 ^ n3136 ;
  assign n3144 = ~n3128 & ~n3143 ;
  assign n3155 = n3154 ^ n3144 ;
  assign n2632 = n2074 ^ n2073 ;
  assign n2645 = n2632 & n2644 ;
  assign n2114 = n2073 ^ n2046 ;
  assign n2117 = n2116 ^ n2082 ;
  assign n2120 = n2046 & ~n2117 ;
  assign n2121 = n2120 ^ n2082 ;
  assign n2122 = n2114 & n2121 ;
  assign n3147 = n2645 ^ n2122 ;
  assign n3156 = n3155 ^ n3147 ;
  assign n2076 = n2075 ^ n2073 ;
  assign n2112 = n2111 ^ n2103 ;
  assign n2113 = ~n2076 & ~n2112 ;
  assign n3157 = n3156 ^ n2113 ;
  assign n2077 = n2016 & ~n2076 ;
  assign n3158 = n3157 ^ n2077 ;
  assign n3145 = n2093 & n2114 ;
  assign n3159 = n3158 ^ n3145 ;
  assign n3160 = ~n2162 & n3159 ;
  assign n3161 = n3160 ^ x2 ;
  assign n3801 = n3161 ^ x122 ;
  assign n1316 = n407 & n1315 ;
  assign n1311 = n481 ^ n446 ;
  assign n1308 = n446 ^ n425 ;
  assign n1309 = n1308 ^ n420 ;
  assign n1310 = n407 & n1309 ;
  assign n1312 = n1311 ^ n1310 ;
  assign n414 = n413 ^ n409 ;
  assign n1294 = n442 ^ n414 ;
  assign n1295 = n483 ^ n411 ;
  assign n1298 = n409 & n1295 ;
  assign n1299 = n1298 ^ n483 ;
  assign n1300 = n1294 & n1299 ;
  assign n1301 = n1300 ^ n408 ;
  assign n1302 = n1301 ^ n435 ;
  assign n1293 = n1292 ^ n1291 ;
  assign n1303 = n1302 ^ n1293 ;
  assign n1304 = n1303 ^ n1284 ;
  assign n473 = n472 ^ n470 ;
  assign n476 = ~n406 & ~n473 ;
  assign n477 = n476 ^ n470 ;
  assign n478 = n433 & ~n477 ;
  assign n1305 = n1304 ^ n478 ;
  assign n1306 = n1305 ^ x39 ;
  assign n1313 = n1312 ^ n1306 ;
  assign n1307 = n1306 ^ n435 ;
  assign n1314 = n1313 ^ n1307 ;
  assign n1317 = n1316 ^ n1314 ;
  assign n1318 = ~n406 & ~n1317 ;
  assign n1319 = n1318 ^ n1313 ;
  assign n1320 = n1319 ^ x100 ;
  assign n380 = n379 ^ n348 ;
  assign n381 = n380 ^ n363 ;
  assign n387 = n386 ^ n381 ;
  assign n388 = ~n329 & ~n387 ;
  assign n389 = n388 ^ n363 ;
  assign n390 = ~n330 & ~n389 ;
  assign n391 = n390 ^ x57 ;
  assign n366 = n365 ^ n356 ;
  assign n367 = ~n329 & n366 ;
  assign n368 = n367 ^ n365 ;
  assign n370 = n368 ^ n338 ;
  assign n369 = n368 ^ n360 ;
  assign n371 = n370 ^ n369 ;
  assign n374 = ~n329 & n371 ;
  assign n375 = n374 ^ n370 ;
  assign n376 = n331 & n375 ;
  assign n377 = n376 ^ n368 ;
  assign n378 = ~n328 & ~n377 ;
  assign n392 = n391 ^ n378 ;
  assign n1321 = n392 ^ x86 ;
  assign n1355 = ~n858 & n1354 ;
  assign n888 = n802 & ~n857 ;
  assign n880 = n822 ^ n810 ;
  assign n881 = n880 ^ n851 ;
  assign n882 = n802 & n881 ;
  assign n883 = n882 ^ n851 ;
  assign n889 = n888 ^ n883 ;
  assign n890 = n812 & n889 ;
  assign n891 = n890 ^ n883 ;
  assign n1356 = n1355 ^ n891 ;
  assign n1347 = ~n802 & ~n858 ;
  assign n1348 = n1347 ^ n859 ;
  assign n1349 = n819 & n1348 ;
  assign n1350 = n1349 ^ n859 ;
  assign n874 = n802 & n859 ;
  assign n875 = n874 ^ n869 ;
  assign n876 = n819 & n875 ;
  assign n877 = n876 ^ n869 ;
  assign n1340 = n877 ^ n814 ;
  assign n860 = n859 ^ n853 ;
  assign n863 = ~n802 & n860 ;
  assign n864 = n863 ^ n853 ;
  assign n865 = n812 & n864 ;
  assign n1341 = n1340 ^ n865 ;
  assign n897 = ~n802 & n851 ;
  assign n898 = n897 ^ n840 ;
  assign n899 = n819 & n898 ;
  assign n900 = n899 ^ n840 ;
  assign n1342 = n1341 ^ n900 ;
  assign n1351 = n1350 ^ n1342 ;
  assign n1357 = n1356 ^ n1351 ;
  assign n1358 = n1357 ^ x23 ;
  assign n902 = n837 ^ n835 ;
  assign n1334 = n902 ^ n826 ;
  assign n1335 = n1334 ^ n825 ;
  assign n1332 = n838 ^ n816 ;
  assign n1336 = n1335 ^ n1332 ;
  assign n1337 = n812 & n1336 ;
  assign n1333 = n1332 ^ n814 ;
  assign n1338 = n1337 ^ n1333 ;
  assign n1339 = ~n802 & n1338 ;
  assign n1359 = n1358 ^ n1339 ;
  assign n1331 = n810 & ~n819 ;
  assign n1360 = n1359 ^ n1331 ;
  assign n903 = n902 ^ n832 ;
  assign n1328 = ~n812 & n903 ;
  assign n1329 = n1328 ^ n832 ;
  assign n1330 = n802 & n1329 ;
  assign n1361 = n1360 ^ n1330 ;
  assign n1362 = n1361 ^ x68 ;
  assign n308 = n256 ^ n248 ;
  assign n310 = n309 ^ n308 ;
  assign n311 = n282 & ~n310 ;
  assign n305 = n304 ^ n249 ;
  assign n306 = n269 & n305 ;
  assign n267 = n266 ^ n246 ;
  assign n270 = n269 ^ n267 ;
  assign n271 = n270 ^ n267 ;
  assign n295 = n257 & ~n271 ;
  assign n296 = n295 ^ n235 ;
  assign n297 = n220 & n296 ;
  assign n301 = n300 ^ n297 ;
  assign n302 = n301 ^ n290 ;
  assign n303 = n302 ^ x7 ;
  assign n307 = n306 ^ n303 ;
  assign n312 = n311 ^ n307 ;
  assign n283 = n282 ^ n220 ;
  assign n284 = n280 & ~n283 ;
  assign n313 = n312 ^ n284 ;
  assign n264 = n263 ^ n259 ;
  assign n265 = n264 ^ n246 ;
  assign n268 = n267 ^ n265 ;
  assign n272 = ~n268 & n271 ;
  assign n273 = n272 ^ n267 ;
  assign n274 = n220 & n273 ;
  assign n314 = n313 ^ n274 ;
  assign n1363 = n314 ^ x110 ;
  assign n1364 = n1362 & ~n1363 ;
  assign n1400 = n1060 ^ n1011 ;
  assign n1401 = n1037 & n1400 ;
  assign n1381 = n1008 & ~n1089 ;
  assign n1380 = n1379 ^ n1057 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1394 = n1382 ^ n1094 ;
  assign n1395 = n1394 ^ n1393 ;
  assign n1396 = n1395 ^ n1050 ;
  assign n1397 = n1396 ^ x15 ;
  assign n1378 = n1023 ^ n1011 ;
  assign n1383 = n1382 ^ n1378 ;
  assign n1376 = n1034 ^ n998 ;
  assign n1377 = ~n997 & n1376 ;
  assign n1384 = n1383 ^ n1377 ;
  assign n1385 = n1384 & n1929 ;
  assign n1398 = n1397 ^ n1385 ;
  assign n1374 = n1081 ^ n1035 ;
  assign n1375 = n1088 & ~n1374 ;
  assign n1399 = n1398 ^ n1375 ;
  assign n1402 = n1401 ^ n1399 ;
  assign n1373 = ~n997 & n1011 ;
  assign n1403 = n1402 ^ n1373 ;
  assign n1367 = n1366 ^ n1056 ;
  assign n1370 = ~n997 & n1367 ;
  assign n1371 = n1370 ^ n1056 ;
  assign n1372 = ~n1037 & n1371 ;
  assign n1404 = n1403 ^ n1372 ;
  assign n1405 = n1404 ^ x117 ;
  assign n1409 = n1408 ^ n680 ;
  assign n1410 = n1409 ^ n676 ;
  assign n1411 = n1410 ^ n646 ;
  assign n1407 = n667 ^ n644 ;
  assign n1412 = n1411 ^ n1407 ;
  assign n1417 = n1416 ^ n1412 ;
  assign n1418 = ~n630 & ~n1417 ;
  assign n1419 = n1418 ^ n1411 ;
  assign n1448 = n1447 ^ n1419 ;
  assign n1457 = n1456 ^ n1448 ;
  assign n1458 = n1457 ^ n1437 ;
  assign n1459 = n1458 ^ x31 ;
  assign n1426 = n630 & n1732 ;
  assign n1406 = n673 ^ n659 ;
  assign n1420 = n1419 ^ n1406 ;
  assign n1427 = n1426 ^ n1420 ;
  assign n1428 = ~n631 & ~n1427 ;
  assign n1460 = n1459 ^ n1428 ;
  assign n1461 = n1460 ^ x69 ;
  assign n1462 = n1405 & n1461 ;
  assign n1463 = n1462 ^ n1461 ;
  assign n1491 = n1364 & n1463 ;
  assign n1509 = n1491 ^ n1463 ;
  assign n1365 = n1364 ^ n1363 ;
  assign n1471 = n1365 ^ n1362 ;
  assign n1479 = n1463 & n1471 ;
  assign n1478 = ~n1365 & n1463 ;
  assign n1480 = n1479 ^ n1478 ;
  assign n1510 = n1509 ^ n1480 ;
  assign n1464 = n1463 ^ n1405 ;
  assign n1472 = ~n1464 & n1471 ;
  assign n3078 = n1510 ^ n1472 ;
  assign n3081 = ~n1321 & n3078 ;
  assign n3082 = n3081 ^ n1472 ;
  assign n3083 = n1320 & n3082 ;
  assign n1468 = n1464 ^ n1461 ;
  assign n1490 = n1468 & n1471 ;
  assign n1470 = n1364 & ~n1464 ;
  assign n1501 = n1490 ^ n1470 ;
  assign n1465 = ~n1365 & ~n1464 ;
  assign n1502 = n1501 ^ n1465 ;
  assign n1503 = n1502 ^ n1472 ;
  assign n1481 = n1471 ^ n1363 ;
  assign n1482 = n1468 & n1481 ;
  assign n1469 = n1364 & n1468 ;
  assign n1483 = n1482 ^ n1469 ;
  assign n1504 = n1503 ^ n1483 ;
  assign n3838 = n1320 & n1504 ;
  assign n3839 = n3838 ^ n1483 ;
  assign n3073 = n1465 ^ n1461 ;
  assign n3074 = n3073 ^ n1504 ;
  assign n3075 = n1321 & ~n3074 ;
  assign n1475 = n1465 ^ n1464 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1476 = n1475 ^ n1473 ;
  assign n1514 = n1476 ^ n1461 ;
  assign n1515 = n1514 ^ n1504 ;
  assign n3076 = n3075 ^ n1515 ;
  assign n3077 = ~n1320 & n3076 ;
  assign n3847 = n3839 ^ n3077 ;
  assign n1467 = n1321 ^ n1320 ;
  assign n1487 = n1462 & n1471 ;
  assign n1523 = n1487 ^ n1462 ;
  assign n3841 = n1523 ^ n1478 ;
  assign n3842 = n3841 ^ n3839 ;
  assign n3837 = n1501 ^ n1476 ;
  assign n3840 = n3839 ^ n3837 ;
  assign n3843 = n3842 ^ n3840 ;
  assign n3844 = ~n1320 & ~n3843 ;
  assign n3845 = n3844 ^ n3842 ;
  assign n3846 = ~n1467 & n3845 ;
  assign n3848 = n3847 ^ n3846 ;
  assign n1322 = ~n1320 & n1321 ;
  assign n3835 = n1510 ^ n1487 ;
  assign n3836 = n1322 & n3835 ;
  assign n3849 = n3848 ^ n3836 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1324 = n1323 ^ n1321 ;
  assign n1325 = n1324 ^ n1320 ;
  assign n3399 = n1325 & n1501 ;
  assign n3850 = n3849 ^ n3399 ;
  assign n1484 = n1364 & n1462 ;
  assign n3827 = n1523 ^ n1484 ;
  assign n3828 = n3827 ^ n1478 ;
  assign n3829 = n3828 ^ n1523 ;
  assign n3832 = ~n1320 & n3829 ;
  assign n3833 = n3832 ^ n1523 ;
  assign n3834 = ~n1321 & n3833 ;
  assign n3851 = n3850 ^ n3834 ;
  assign n1466 = n1325 & n1465 ;
  assign n3852 = n3851 ^ n1466 ;
  assign n1521 = ~n1323 & n1491 ;
  assign n3853 = n3852 ^ n1521 ;
  assign n1493 = n1462 & n1481 ;
  assign n1524 = n1493 ^ n1484 ;
  assign n1525 = n1524 ^ n1523 ;
  assign n1526 = n1525 ^ n1479 ;
  assign n3826 = ~n1320 & n1526 ;
  assign n3854 = n3853 ^ n3826 ;
  assign n3855 = ~n3083 & ~n3854 ;
  assign n3856 = n3855 ^ x10 ;
  assign n3857 = n3856 ^ x66 ;
  assign n3868 = ~n3801 & ~n3857 ;
  assign n3869 = n3868 ^ n3801 ;
  assign n3895 = n3869 ^ n3857 ;
  assign n711 = n655 ^ n639 ;
  assign n712 = n711 ^ n638 ;
  assign n713 = n710 & ~n712 ;
  assign n698 = n697 ^ n650 ;
  assign n702 = n701 ^ n698 ;
  assign n703 = ~n656 & n702 ;
  assign n704 = n703 ^ n698 ;
  assign n705 = n630 & n704 ;
  assign n706 = n705 ^ n698 ;
  assign n707 = ~n631 & n706 ;
  assign n708 = n707 ^ x33 ;
  assign n694 = ~n629 & ~n678 ;
  assign n695 = n694 ^ n676 ;
  assign n696 = n630 & n695 ;
  assign n709 = n708 ^ n696 ;
  assign n714 = n713 ^ n709 ;
  assign n689 = ~n630 & ~n659 ;
  assign n715 = n714 ^ n689 ;
  assign n681 = n680 ^ n667 ;
  assign n682 = n681 ^ n675 ;
  assign n683 = n682 ^ n680 ;
  assign n686 = ~n630 & n683 ;
  assign n687 = n686 ^ n680 ;
  assign n688 = ~n631 & n687 ;
  assign n716 = n715 ^ n688 ;
  assign n2401 = n716 ^ x88 ;
  assign n2402 = n1955 ^ x97 ;
  assign n2403 = n2045 ^ x74 ;
  assign n911 = n802 & n825 ;
  assign n904 = n903 ^ n851 ;
  assign n905 = ~n802 & n904 ;
  assign n906 = n905 ^ n851 ;
  assign n912 = n911 ^ n906 ;
  assign n913 = ~n812 & n912 ;
  assign n914 = n913 ^ n906 ;
  assign n2422 = n914 ^ n869 ;
  assign n2413 = n1334 ^ n814 ;
  assign n2423 = n2422 ^ n2413 ;
  assign n2424 = n2423 ^ n1350 ;
  assign n2425 = n2424 ^ n1356 ;
  assign n2426 = n2425 ^ x17 ;
  assign n2414 = n2413 ^ n827 ;
  assign n2415 = n2414 ^ n816 ;
  assign n2416 = n2415 ^ n2413 ;
  assign n2419 = ~n812 & n2416 ;
  assign n2420 = n2419 ^ n2413 ;
  assign n2421 = n819 & n2420 ;
  assign n2427 = n2426 ^ n2421 ;
  assign n841 = n840 ^ n832 ;
  assign n2412 = n841 & ~n1353 ;
  assign n2428 = n2427 ^ n2412 ;
  assign n2404 = n869 ^ n840 ;
  assign n2405 = n2404 ^ n855 ;
  assign n2406 = n2405 ^ n869 ;
  assign n2409 = n812 & n2406 ;
  assign n2410 = n2409 ^ n869 ;
  assign n2411 = ~n802 & n2410 ;
  assign n2429 = n2428 ^ n2411 ;
  assign n2430 = n2429 ^ x122 ;
  assign n2431 = n2403 & ~n2430 ;
  assign n2453 = n304 ^ n255 ;
  assign n2454 = n282 & ~n2453 ;
  assign n2450 = n264 ^ x9 ;
  assign n2443 = n254 ^ n250 ;
  assign n2444 = n2443 ^ n261 ;
  assign n2442 = n231 & n281 ;
  assign n2445 = n2444 ^ n2442 ;
  assign n2446 = ~n977 & ~n2445 ;
  assign n2447 = n2446 ^ n250 ;
  assign n2440 = n1986 ^ n263 ;
  assign n2441 = n298 & n2440 ;
  assign n2448 = n2447 ^ n2441 ;
  assign n2449 = ~n290 & ~n2448 ;
  assign n2451 = n2450 ^ n2449 ;
  assign n2439 = n245 & ~n977 ;
  assign n2452 = n2451 ^ n2439 ;
  assign n2455 = n2454 ^ n2452 ;
  assign n2436 = ~n220 & n308 ;
  assign n2437 = n2436 ^ n264 ;
  assign n2438 = ~n269 & ~n2437 ;
  assign n2456 = n2455 ^ n2438 ;
  assign n2457 = n2456 ^ x64 ;
  assign n212 = n182 ^ n165 ;
  assign n190 = n183 ^ n169 ;
  assign n191 = n190 ^ n186 ;
  assign n192 = n191 ^ n159 ;
  assign n193 = n140 & ~n192 ;
  assign n189 = n188 ^ n183 ;
  assign n194 = n193 ^ n189 ;
  assign n195 = n194 ^ n182 ;
  assign n213 = n212 ^ n195 ;
  assign n199 = n184 ^ n180 ;
  assign n203 = n202 ^ n199 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = n205 ^ n140 ;
  assign n208 = n207 ^ n205 ;
  assign n209 = ~n206 & n208 ;
  assign n210 = n209 ^ n205 ;
  assign n211 = n147 & ~n210 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ x25 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ n165 ;
  assign n196 = n195 ^ n173 ;
  assign n160 = n159 ^ n152 ;
  assign n161 = n140 & ~n160 ;
  assign n197 = n196 ^ n161 ;
  assign n198 = ~n147 & n197 ;
  assign n216 = n215 ^ n198 ;
  assign n150 = ~n148 & n149 ;
  assign n217 = n216 ^ n150 ;
  assign n139 = n138 ^ n136 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = n139 & n142 ;
  assign n144 = n143 ^ n138 ;
  assign n145 = n129 & n144 ;
  assign n218 = n217 ^ n145 ;
  assign n2458 = n218 ^ x112 ;
  assign n2459 = n2457 & ~n2458 ;
  assign n2468 = n2459 ^ n2457 ;
  assign n2495 = n2431 & n2468 ;
  assign n2506 = n2495 ^ n2468 ;
  assign n2464 = n2431 ^ n2403 ;
  assign n2482 = n2464 & n2468 ;
  assign n2466 = n2431 ^ n2430 ;
  assign n2469 = ~n2466 & n2468 ;
  assign n2483 = n2482 ^ n2469 ;
  assign n2507 = n2506 ^ n2483 ;
  assign n2474 = n2464 ^ n2430 ;
  assign n2475 = n2459 & n2474 ;
  assign n2473 = n2431 & n2459 ;
  assign n2476 = n2475 ^ n2473 ;
  assign n2471 = n2459 & n2464 ;
  assign n2472 = n2471 ^ n2459 ;
  assign n2477 = n2476 ^ n2472 ;
  assign n2478 = n2477 ^ n2466 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2467 = ~n2460 & ~n2466 ;
  assign n2470 = n2469 ^ n2467 ;
  assign n2479 = n2478 ^ n2470 ;
  assign n2461 = n2460 ^ n2457 ;
  assign n2465 = n2461 & n2464 ;
  assign n2480 = n2479 ^ n2465 ;
  assign n2888 = n2507 ^ n2480 ;
  assign n2891 = n2402 & ~n2888 ;
  assign n2892 = n2891 ^ n2480 ;
  assign n2893 = ~n2401 & ~n2892 ;
  assign n2894 = n2893 ^ x26 ;
  assign n2462 = n2431 & n2461 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2481 = n2480 ^ n2463 ;
  assign n2496 = n2495 ^ n2481 ;
  assign n2553 = ~n2401 & ~n2402 ;
  assign n2558 = n2553 ^ n2401 ;
  assign n2566 = ~n2496 & ~n2558 ;
  assign n2560 = n2558 ^ n2402 ;
  assign n2565 = n2477 & ~n2560 ;
  assign n2567 = n2566 ^ n2565 ;
  assign n2528 = n2402 ^ n2401 ;
  assign n2877 = n2473 ^ n2469 ;
  assign n2878 = n2877 ^ n2471 ;
  assign n2508 = n2507 ^ n2481 ;
  assign n2505 = n2475 ^ n2474 ;
  assign n2509 = n2508 ^ n2505 ;
  assign n2487 = n2430 ^ n2403 ;
  assign n2488 = n2487 ^ n2458 ;
  assign n2489 = n2488 ^ n2457 ;
  assign n2485 = n2476 ^ n2462 ;
  assign n2484 = n2483 ^ n2467 ;
  assign n2486 = n2485 ^ n2484 ;
  assign n2490 = n2489 ^ n2486 ;
  assign n2491 = n2490 ^ n2481 ;
  assign n2510 = n2509 ^ n2491 ;
  assign n2504 = n2467 ^ n2460 ;
  assign n2511 = n2510 ^ n2504 ;
  assign n2512 = n2511 ^ n2509 ;
  assign n2503 = n2495 ^ n2479 ;
  assign n2513 = n2512 ^ n2503 ;
  assign n2879 = n2878 ^ n2513 ;
  assign n2880 = n2401 & n2879 ;
  assign n2881 = n2880 ^ n2473 ;
  assign n2882 = ~n2528 & n2881 ;
  assign n2536 = n2482 ^ n2462 ;
  assign n2867 = n2536 ^ n2508 ;
  assign n2866 = n2469 & n2553 ;
  assign n2868 = n2867 ^ n2866 ;
  assign n2561 = n2560 ^ n2401 ;
  assign n2869 = n2868 ^ n2561 ;
  assign n2872 = n2483 & n2553 ;
  assign n2554 = n2491 ^ n2475 ;
  assign n2870 = n2868 ^ n2554 ;
  assign n2864 = n2511 ^ n2477 ;
  assign n2871 = n2870 ^ n2864 ;
  assign n2873 = n2872 ^ n2871 ;
  assign n2874 = n2869 & n2873 ;
  assign n2875 = n2874 ^ n2561 ;
  assign n2865 = ~n2558 & n2864 ;
  assign n2876 = n2875 ^ n2865 ;
  assign n2883 = n2882 ^ n2876 ;
  assign n2559 = n2482 & ~n2558 ;
  assign n2884 = n2883 ^ n2559 ;
  assign n2858 = n2491 ^ n2467 ;
  assign n2861 = n2402 & n2858 ;
  assign n2862 = n2861 ^ n2467 ;
  assign n2863 = ~n2401 & n2862 ;
  assign n2885 = n2884 ^ n2863 ;
  assign n2555 = n2553 & n2554 ;
  assign n2547 = n2509 ^ n2465 ;
  assign n2550 = ~n2401 & ~n2547 ;
  assign n2551 = n2550 ^ n2465 ;
  assign n2552 = n2402 & n2551 ;
  assign n2556 = n2555 ^ n2552 ;
  assign n2886 = n2885 ^ n2556 ;
  assign n2887 = ~n2567 & n2886 ;
  assign n2895 = n2894 ^ n2887 ;
  assign n3825 = n2895 ^ x105 ;
  assign n3872 = n3801 & n3825 ;
  assign n3896 = n3895 ^ n3872 ;
  assign n3897 = n3823 & ~n3896 ;
  assign n3865 = n3823 & ~n3825 ;
  assign n3874 = n3865 ^ n3825 ;
  assign n3875 = n3874 ^ n3823 ;
  assign n617 = n614 & n616 ;
  assign n618 = n617 ^ n613 ;
  assign n581 = n580 ^ n578 ;
  assign n577 = n576 ^ n545 ;
  assign n582 = n581 ^ n577 ;
  assign n583 = ~n521 & ~n582 ;
  assign n584 = n583 ^ n581 ;
  assign n619 = n618 ^ n584 ;
  assign n620 = n619 ^ n601 ;
  assign n593 = ~n521 & n588 ;
  assign n594 = n593 ^ n562 ;
  assign n595 = n520 & n594 ;
  assign n621 = n620 ^ n595 ;
  assign n569 = n568 ^ n531 ;
  assign n571 = n570 ^ n569 ;
  assign n574 = n573 ^ n571 ;
  assign n575 = n521 & n574 ;
  assign n585 = n584 ^ n575 ;
  assign n586 = ~n520 & ~n585 ;
  assign n622 = n621 ^ n586 ;
  assign n547 = n546 ^ n542 ;
  assign n548 = ~n534 & n547 ;
  assign n623 = n622 ^ n548 ;
  assign n625 = n624 ^ n623 ;
  assign n626 = n625 ^ x41 ;
  assign n533 = ~n523 & n532 ;
  assign n627 = n626 ^ n533 ;
  assign n628 = n627 ^ x115 ;
  assign n717 = n716 ^ x104 ;
  assign n718 = ~n628 & ~n717 ;
  assign n393 = n392 ^ x106 ;
  assign n443 = n442 ^ n438 ;
  assign n447 = n446 ^ n431 ;
  assign n448 = n447 ^ n435 ;
  assign n444 = n438 ^ n420 ;
  assign n445 = n444 ^ n442 ;
  assign n449 = n448 ^ n445 ;
  assign n450 = n449 ^ n407 ;
  assign n451 = n450 ^ n445 ;
  assign n452 = ~n433 & n451 ;
  assign n453 = n452 ^ n433 ;
  assign n454 = n443 & ~n453 ;
  assign n455 = n454 ^ n445 ;
  assign n456 = n451 ^ n406 ;
  assign n457 = n456 ^ n452 ;
  assign n458 = ~n455 & n457 ;
  assign n459 = n458 ^ n445 ;
  assign n506 = n459 ^ n406 ;
  assign n507 = n506 ^ n505 ;
  assign n508 = n507 ^ n499 ;
  assign n509 = n508 ^ n493 ;
  assign n510 = n509 ^ n490 ;
  assign n511 = n510 ^ n478 ;
  assign n460 = n459 ^ n430 ;
  assign n461 = n460 ^ n437 ;
  assign n462 = n461 ^ n459 ;
  assign n465 = ~n407 & ~n462 ;
  assign n466 = n465 ^ n459 ;
  assign n467 = n433 & ~n466 ;
  assign n512 = n511 ^ n467 ;
  assign n432 = n408 & n431 ;
  assign n513 = n512 ^ n432 ;
  assign n412 = n411 ^ n405 ;
  assign n417 = ~n405 & n414 ;
  assign n418 = n417 ^ n409 ;
  assign n419 = n412 & ~n418 ;
  assign n514 = n513 ^ n419 ;
  assign n516 = n515 ^ n514 ;
  assign n517 = n516 ^ x49 ;
  assign n518 = n517 ^ x89 ;
  assign n519 = n393 & n518 ;
  assign n721 = n519 ^ n393 ;
  assign n758 = n718 & n721 ;
  assign n759 = n758 ^ n718 ;
  assign n726 = n721 ^ n518 ;
  assign n736 = n718 & ~n726 ;
  assign n727 = n726 ^ n393 ;
  assign n730 = n718 & n727 ;
  assign n739 = n736 ^ n730 ;
  assign n760 = n759 ^ n739 ;
  assign n719 = n718 ^ n717 ;
  assign n725 = n719 ^ n628 ;
  assign n741 = n721 & ~n725 ;
  assign n728 = ~n725 & n727 ;
  assign n742 = n741 ^ n728 ;
  assign n756 = n742 ^ n725 ;
  assign n731 = n725 ^ n717 ;
  assign n744 = ~n726 & ~n731 ;
  assign n745 = n744 ^ n726 ;
  assign n732 = n727 & ~n731 ;
  assign n733 = n732 ^ n730 ;
  assign n729 = n728 ^ n727 ;
  assign n734 = n733 ^ n729 ;
  assign n722 = ~n719 & n721 ;
  assign n720 = n519 & ~n719 ;
  assign n723 = n722 ^ n720 ;
  assign n724 = n723 ^ n719 ;
  assign n735 = n734 ^ n724 ;
  assign n737 = n736 ^ n735 ;
  assign n746 = n745 ^ n737 ;
  assign n757 = n756 ^ n746 ;
  assign n761 = n760 ^ n757 ;
  assign n219 = n218 ^ x72 ;
  assign n315 = n314 ^ x65 ;
  assign n316 = n219 & n315 ;
  assign n2574 = n316 ^ n315 ;
  assign n3278 = ~n761 & n2574 ;
  assign n785 = n316 ^ n219 ;
  assign n788 = n785 ^ n315 ;
  assign n2625 = n734 & ~n788 ;
  assign n3279 = n3278 ^ n2625 ;
  assign n786 = ~n735 & n785 ;
  assign n770 = n315 ^ n219 ;
  assign n747 = n746 ^ n734 ;
  assign n779 = n747 ^ n732 ;
  assign n782 = n315 & n779 ;
  assign n783 = n782 ^ n732 ;
  assign n784 = n770 & n783 ;
  assign n787 = n786 ^ n784 ;
  assign n3280 = n3279 ^ n787 ;
  assign n764 = n721 & ~n731 ;
  assign n789 = n764 ^ n732 ;
  assign n790 = ~n788 & n789 ;
  assign n3281 = n3280 ^ n790 ;
  assign n3282 = n3281 ^ x60 ;
  assign n796 = n720 ^ n519 ;
  assign n797 = n796 ^ n761 ;
  assign n2593 = n797 ^ n758 ;
  assign n2603 = n2593 ^ n732 ;
  assign n2606 = ~n219 & ~n2603 ;
  assign n2607 = n2606 ^ n732 ;
  assign n2608 = n315 & n2607 ;
  assign n750 = n742 ^ n730 ;
  assign n751 = n219 & n750 ;
  assign n752 = n751 ^ n730 ;
  assign n3267 = n739 ^ n723 ;
  assign n3268 = n219 & n3267 ;
  assign n771 = n744 ^ n736 ;
  assign n3261 = n771 ^ n760 ;
  assign n3260 = n764 ^ n720 ;
  assign n3262 = n3261 ^ n3260 ;
  assign n3263 = n219 & n3262 ;
  assign n3258 = n771 ^ n757 ;
  assign n3255 = n797 ^ n741 ;
  assign n3256 = n219 & ~n3255 ;
  assign n3257 = n3256 ^ n741 ;
  assign n3259 = n3258 ^ n3257 ;
  assign n3264 = n3263 ^ n3259 ;
  assign n3265 = n3264 ^ n723 ;
  assign n3266 = n3265 ^ n3257 ;
  assign n3269 = n3268 ^ n3266 ;
  assign n3272 = n3269 ^ n3265 ;
  assign n3273 = ~n752 & ~n3272 ;
  assign n3274 = n3273 ^ n3269 ;
  assign n3275 = n315 & n3274 ;
  assign n3276 = n3275 ^ n3269 ;
  assign n3277 = ~n2608 & n3276 ;
  assign n3283 = n3282 ^ n3277 ;
  assign n3799 = n3283 ^ x80 ;
  assign n1583 = n1460 ^ x75 ;
  assign n811 = ~n802 & n810 ;
  assign n818 = n812 & ~n817 ;
  assign n920 = n811 & n818 ;
  assign n866 = n817 ^ n812 ;
  assign n867 = n866 ^ n865 ;
  assign n878 = n877 ^ n867 ;
  assign n879 = n878 ^ n829 ;
  assign n892 = n891 ^ n879 ;
  assign n901 = n900 ^ n892 ;
  assign n915 = n914 ^ n901 ;
  assign n916 = n915 ^ x5 ;
  assign n842 = n841 ^ n829 ;
  assign n843 = n842 ^ n830 ;
  assign n846 = ~n812 & n843 ;
  assign n847 = n846 ^ n830 ;
  assign n848 = n819 & n847 ;
  assign n917 = n916 ^ n848 ;
  assign n918 = n917 ^ n818 ;
  assign n921 = n920 ^ n918 ;
  assign n1531 = n921 ^ x116 ;
  assign n1186 = n546 ^ n540 ;
  assign n1187 = n1186 ^ n531 ;
  assign n1191 = n1190 ^ n1187 ;
  assign n1192 = n521 & ~n1191 ;
  assign n1193 = n1192 ^ n546 ;
  assign n1194 = ~n520 & n1193 ;
  assign n1181 = n562 ^ n541 ;
  assign n1182 = n1181 ^ n532 ;
  assign n1183 = n616 & n1182 ;
  assign n1169 = n567 ^ n535 ;
  assign n1170 = n1169 ^ n1164 ;
  assign n1171 = ~n523 & n1170 ;
  assign n1172 = n1171 ^ n615 ;
  assign n1177 = ~n523 & n1164 ;
  assign n1173 = n567 ^ n544 ;
  assign n1174 = n1173 ^ n614 ;
  assign n1175 = n1174 ^ n562 ;
  assign n1176 = n1175 ^ n542 ;
  assign n1178 = n1177 ^ n1176 ;
  assign n1179 = n1172 & n1178 ;
  assign n1167 = n1166 ^ x63 ;
  assign n1168 = n1167 ^ n618 ;
  assign n1180 = n1179 ^ n1168 ;
  assign n1184 = n1183 ^ n1180 ;
  assign n1163 = ~n534 & n545 ;
  assign n1185 = n1184 ^ n1163 ;
  assign n1195 = n1194 ^ n1185 ;
  assign n1548 = n1195 ^ x76 ;
  assign n1564 = n168 ^ n151 ;
  assign n1555 = n178 ^ n131 ;
  assign n1556 = n1555 ^ n170 ;
  assign n1565 = n1564 ^ n1556 ;
  assign n1566 = n1565 ^ n211 ;
  assign n1557 = n1556 ^ n129 ;
  assign n1558 = n147 & n1557 ;
  assign n1559 = n1558 ^ n129 ;
  assign n1560 = n186 ^ n132 ;
  assign n1561 = n1560 ^ n1556 ;
  assign n1562 = n1561 ^ n183 ;
  assign n1563 = n1559 & n1562 ;
  assign n1567 = n1566 ^ n1563 ;
  assign n1570 = n1567 ^ n211 ;
  assign n1568 = n172 ^ n149 ;
  assign n1569 = ~n129 & n1568 ;
  assign n1571 = n1570 ^ n1569 ;
  assign n1572 = n147 & n1571 ;
  assign n1573 = n1572 ^ n1567 ;
  assign n1549 = n178 ^ n162 ;
  assign n1552 = n129 & n1549 ;
  assign n1553 = n1552 ^ n162 ;
  assign n1554 = ~n140 & n1553 ;
  assign n1574 = n1573 ^ n1554 ;
  assign n1575 = n1574 ^ n955 ;
  assign n1576 = n1575 ^ x47 ;
  assign n1577 = n1576 ^ x118 ;
  assign n1578 = ~n1548 & n1577 ;
  assign n1579 = n1578 ^ n1548 ;
  assign n1580 = n1579 ^ n1577 ;
  assign n1532 = n1319 ^ x70 ;
  assign n1543 = n390 ^ x55 ;
  assign n1537 = n1134 ^ n1118 ;
  assign n1538 = n330 & ~n1537 ;
  assign n1539 = n1538 ^ n1118 ;
  assign n1544 = n1543 ^ n1539 ;
  assign n1540 = n1539 ^ n1122 ;
  assign n1533 = n1122 ^ n353 ;
  assign n1534 = n1533 ^ n379 ;
  assign n1535 = n1534 ^ n1130 ;
  assign n1536 = ~n330 & n1535 ;
  assign n1541 = n1540 ^ n1536 ;
  assign n1542 = n329 & n1541 ;
  assign n1545 = n1544 ^ n1542 ;
  assign n1546 = n1545 ^ x93 ;
  assign n1547 = n1532 & ~n1546 ;
  assign n1589 = n1547 ^ n1532 ;
  assign n1594 = n1589 ^ n1546 ;
  assign n1601 = n1580 & n1594 ;
  assign n1590 = ~n1579 & n1589 ;
  assign n2727 = n1601 ^ n1590 ;
  assign n1587 = n1547 ^ n1546 ;
  assign n1592 = n1578 ^ n1577 ;
  assign n1597 = ~n1587 & n1592 ;
  assign n2728 = n2727 ^ n1597 ;
  assign n1602 = n1580 & ~n1587 ;
  assign n1585 = n1547 & n1578 ;
  assign n2725 = n1602 ^ n1585 ;
  assign n1609 = n1547 & ~n1579 ;
  assign n2726 = n2725 ^ n1609 ;
  assign n2729 = n2728 ^ n2726 ;
  assign n2973 = n1531 & n2729 ;
  assign n1603 = n1602 ^ n1601 ;
  assign n1581 = n1547 & n1580 ;
  assign n1600 = n1581 ^ n1580 ;
  assign n1604 = n1603 ^ n1600 ;
  assign n1598 = n1597 ^ n1592 ;
  assign n1595 = n1592 & n1594 ;
  assign n1593 = n1547 & n1592 ;
  assign n1596 = n1595 ^ n1593 ;
  assign n1599 = n1598 ^ n1596 ;
  assign n1605 = n1604 ^ n1599 ;
  assign n1591 = n1590 ^ n1589 ;
  assign n1606 = n1605 ^ n1591 ;
  assign n1588 = n1578 & ~n1587 ;
  assign n1607 = n1606 ^ n1588 ;
  assign n1586 = n1585 ^ n1578 ;
  assign n1608 = n1607 ^ n1586 ;
  assign n2717 = n1608 ^ n1597 ;
  assign n1622 = ~n1579 & ~n1587 ;
  assign n1623 = n1622 ^ n1590 ;
  assign n1661 = n1623 ^ n1579 ;
  assign n2716 = n1661 ^ n1604 ;
  assign n2718 = n2717 ^ n2716 ;
  assign n2969 = ~n1583 & ~n2718 ;
  assign n2970 = n2969 ^ n1595 ;
  assign n2971 = n1531 & n2970 ;
  assign n2972 = n2971 ^ n2726 ;
  assign n2974 = n2973 ^ n2972 ;
  assign n2730 = n1587 ^ n1579 ;
  assign n2731 = n2730 ^ n2729 ;
  assign n2723 = n1546 ^ n1532 ;
  assign n2724 = n2723 ^ n1548 ;
  assign n2732 = n2731 ^ n2724 ;
  assign n2733 = ~n1531 & ~n2732 ;
  assign n2980 = n2974 ^ n2733 ;
  assign n2981 = n2980 ^ n2971 ;
  assign n2982 = ~n1583 & n2981 ;
  assign n1650 = n1531 & ~n1583 ;
  assign n2976 = n1581 & n1650 ;
  assign n1613 = n1608 ^ n1590 ;
  assign n2738 = n1613 ^ n1607 ;
  assign n2741 = ~n1531 & n2738 ;
  assign n2742 = n2741 ^ n1607 ;
  assign n2743 = n1583 & n2742 ;
  assign n2977 = n2976 ^ n2743 ;
  assign n2961 = ~n1531 & n1604 ;
  assign n1640 = n1597 ^ n1581 ;
  assign n1641 = ~n1531 & n1640 ;
  assign n1642 = n1641 ^ n1581 ;
  assign n2962 = n2961 ^ n1642 ;
  assign n2963 = n1583 & n2962 ;
  assign n1651 = n1585 & n1650 ;
  assign n1647 = ~n1531 & n1605 ;
  assign n1648 = n1647 ^ n1604 ;
  assign n1649 = n1583 & n1648 ;
  assign n1652 = n1651 ^ n1649 ;
  assign n2964 = n2963 ^ n1652 ;
  assign n2975 = n2974 ^ n2964 ;
  assign n2978 = n2977 ^ n2975 ;
  assign n2979 = n2978 ^ x34 ;
  assign n2983 = n2982 ^ n2979 ;
  assign n3800 = n2983 ^ x98 ;
  assign n3917 = n3800 & ~n3857 ;
  assign n3918 = n3917 ^ n3868 ;
  assign n3919 = ~n3799 & n3918 ;
  assign n4482 = n3875 & n3919 ;
  assign n3906 = n3825 & ~n3869 ;
  assign n3858 = n3857 ^ n3801 ;
  assign n3891 = ~n3858 & ~n3874 ;
  assign n3877 = n3825 ^ n3823 ;
  assign n3888 = ~n3823 & n3868 ;
  assign n3889 = n3888 ^ n3801 ;
  assign n3890 = ~n3877 & ~n3889 ;
  assign n3892 = n3891 ^ n3890 ;
  assign n3879 = n3872 ^ n3801 ;
  assign n3880 = n3879 ^ n3865 ;
  assign n3876 = ~n3801 & ~n3875 ;
  assign n3878 = n3877 ^ n3876 ;
  assign n3881 = n3880 ^ n3878 ;
  assign n3885 = n3881 ^ n3877 ;
  assign n3893 = n3892 ^ n3885 ;
  assign n3866 = ~n3801 & n3865 ;
  assign n3903 = n3893 ^ n3866 ;
  assign n4470 = n3906 ^ n3903 ;
  assign n3882 = n3881 ^ n3801 ;
  assign n3883 = n3857 & n3882 ;
  assign n3884 = n3883 ^ n3876 ;
  assign n4469 = ~n3880 & ~n3884 ;
  assign n4471 = n4470 ^ n4469 ;
  assign n4472 = n3799 & n4471 ;
  assign n4473 = n4472 ^ n4470 ;
  assign n4483 = n4482 ^ n4473 ;
  assign n4475 = n4473 ^ n3892 ;
  assign n3894 = n3893 ^ n3884 ;
  assign n4474 = n4473 ^ n3894 ;
  assign n4476 = n4475 ^ n4474 ;
  assign n4479 = n3799 & n4476 ;
  assign n4480 = n4479 ^ n4475 ;
  assign n4481 = ~n3800 & n4480 ;
  assign n4484 = n4483 ^ n4481 ;
  assign n4485 = ~n3897 & ~n4484 ;
  assign n4486 = n4485 ^ n392 ;
  assign n5605 = n4486 ^ x117 ;
  assign n1873 = n1831 ^ n1824 ;
  assign n1909 = n1873 ^ n1672 ;
  assign n1910 = n1866 ^ n1852 ;
  assign n1911 = n1909 & ~n1910 ;
  assign n1912 = n1911 ^ x0 ;
  assign n1900 = ~n1672 & n1851 ;
  assign n1893 = n1850 ^ n1781 ;
  assign n1894 = ~n1672 & n1893 ;
  assign n1895 = n1894 ^ n1850 ;
  assign n1901 = n1900 ^ n1895 ;
  assign n1902 = n1824 & n1901 ;
  assign n1903 = n1902 ^ n1895 ;
  assign n1881 = n1856 ^ n1781 ;
  assign n1877 = n1845 ^ n1824 ;
  assign n1878 = ~n1835 & n1877 ;
  assign n1879 = n1878 ^ n1824 ;
  assign n1880 = n1857 & ~n1879 ;
  assign n1882 = n1881 ^ n1880 ;
  assign n1904 = n1903 ^ n1882 ;
  assign n1885 = n1884 ^ n1882 ;
  assign n1886 = n1885 ^ n1779 ;
  assign n1887 = n1886 ^ n1882 ;
  assign n1890 = ~n1824 & n1887 ;
  assign n1891 = n1890 ^ n1882 ;
  assign n1892 = ~n1835 & n1891 ;
  assign n1905 = n1904 ^ n1892 ;
  assign n1874 = n1849 ^ n1784 ;
  assign n1875 = n1874 ^ n1847 ;
  assign n1876 = n1873 & n1875 ;
  assign n1906 = n1905 ^ n1876 ;
  assign n1867 = n1866 ^ n1864 ;
  assign n1870 = n1824 & ~n1867 ;
  assign n1871 = n1870 ^ n1864 ;
  assign n1872 = n1835 & ~n1871 ;
  assign n1907 = n1906 ^ n1872 ;
  assign n1908 = ~n1834 & ~n1907 ;
  assign n1913 = n1912 ^ n1908 ;
  assign n1914 = n1913 ^ x123 ;
  assign n2138 = n2093 ^ n2006 ;
  assign n2136 = n2101 ^ n2096 ;
  assign n2131 = n2130 ^ n2106 ;
  assign n2132 = n2131 ^ n2013 ;
  assign n2135 = n2132 ^ n2109 ;
  assign n2137 = n2136 ^ n2135 ;
  assign n2139 = n2138 ^ n2137 ;
  assign n2140 = n2139 ^ n2132 ;
  assign n2141 = ~n2046 & n2140 ;
  assign n2142 = n2141 ^ n2135 ;
  assign n2143 = ~n2114 & ~n2142 ;
  assign n2127 = n2046 & n2098 ;
  assign n2128 = n2127 ^ n2084 ;
  assign n2129 = n2114 & n2128 ;
  assign n2133 = n2132 ^ n2129 ;
  assign n2134 = n2133 ^ n2122 ;
  assign n2144 = n2143 ^ n2134 ;
  assign n2152 = ~n2144 & ~n2151 ;
  assign n2153 = ~n2113 & n2152 ;
  assign n2154 = ~n2077 & n2153 ;
  assign n2163 = n2154 & ~n2162 ;
  assign n2164 = n2163 ^ x16 ;
  assign n2165 = n2164 ^ x106 ;
  assign n2166 = ~n1914 & n2165 ;
  assign n2167 = n2166 ^ n1914 ;
  assign n2168 = n2167 ^ n2165 ;
  assign n1527 = n1325 & n1526 ;
  assign n1516 = n1515 ^ n1476 ;
  assign n1492 = n1491 ^ n1490 ;
  assign n1494 = n1493 ^ n1492 ;
  assign n1488 = n1487 ^ n1484 ;
  assign n1486 = n1320 & n1462 ;
  assign n1489 = n1488 ^ n1486 ;
  assign n1495 = n1494 ^ n1489 ;
  assign n1485 = n1484 ^ n1483 ;
  assign n1496 = n1495 ^ n1485 ;
  assign n1497 = ~n1320 & n1496 ;
  assign n1498 = n1497 ^ n1495 ;
  assign n1513 = n1498 ^ n1489 ;
  assign n1517 = n1516 ^ n1513 ;
  assign n1511 = n1510 ^ n1478 ;
  assign n1512 = ~n1323 & n1511 ;
  assign n1518 = n1517 ^ n1512 ;
  assign n1506 = n1321 & ~n1516 ;
  assign n1499 = n1498 ^ n1480 ;
  assign n1474 = n1473 ^ n1469 ;
  assign n1477 = n1476 ^ n1474 ;
  assign n1500 = n1499 ^ n1477 ;
  assign n1507 = n1506 ^ n1500 ;
  assign n1508 = n1467 & ~n1507 ;
  assign n1519 = n1518 ^ n1508 ;
  assign n1520 = n1519 ^ n1466 ;
  assign n1522 = n1521 ^ n1520 ;
  assign n1528 = n1527 ^ n1522 ;
  assign n1529 = n1528 ^ x24 ;
  assign n1530 = n1529 ^ x96 ;
  assign n1662 = n1599 ^ n1597 ;
  assign n1663 = n1662 ^ n1661 ;
  assign n1664 = n1663 ^ n1603 ;
  assign n1660 = n1622 ^ n1606 ;
  assign n1665 = n1664 ^ n1660 ;
  assign n1666 = n1531 & ~n1665 ;
  assign n1659 = n1642 ^ n1602 ;
  assign n1667 = n1666 ^ n1659 ;
  assign n1668 = ~n1583 & n1667 ;
  assign n1653 = n1652 ^ n1642 ;
  assign n1612 = n1604 ^ n1588 ;
  assign n1614 = n1613 ^ n1612 ;
  assign n1620 = n1614 ^ n1596 ;
  assign n1610 = n1609 ^ n1588 ;
  assign n1611 = n1610 ^ n1608 ;
  assign n1615 = n1614 ^ n1611 ;
  assign n1584 = n1583 ^ n1531 ;
  assign n1616 = n1611 ^ n1531 ;
  assign n1617 = n1584 & ~n1616 ;
  assign n1618 = n1617 ^ n1531 ;
  assign n1619 = n1615 & n1618 ;
  assign n1621 = n1620 ^ n1619 ;
  assign n1654 = n1653 ^ n1621 ;
  assign n1637 = ~n1531 & n1603 ;
  assign n1638 = n1637 ^ n1602 ;
  assign n1639 = n1583 & n1638 ;
  assign n1655 = n1654 ^ n1639 ;
  assign n1656 = n1655 ^ x8 ;
  assign n1624 = n1623 ^ n1585 ;
  assign n1625 = n1624 ^ n1621 ;
  assign n1626 = n1625 ^ n1588 ;
  assign n1627 = n1626 ^ n1621 ;
  assign n1630 = ~n1531 & n1627 ;
  assign n1631 = n1630 ^ n1621 ;
  assign n1632 = n1584 & n1631 ;
  assign n1657 = n1656 ^ n1632 ;
  assign n1582 = ~n1531 & n1581 ;
  assign n1658 = n1657 ^ n1582 ;
  assign n1669 = n1668 ^ n1658 ;
  assign n1670 = n1669 ^ x113 ;
  assign n1671 = n1530 & n1670 ;
  assign n2179 = n1671 ^ n1530 ;
  assign n2180 = n2179 ^ n1670 ;
  assign n2183 = n2168 & ~n2180 ;
  assign n2181 = n2180 ^ n1530 ;
  assign n2182 = n2166 & n2181 ;
  assign n2184 = n2183 ^ n2182 ;
  assign n2170 = n1671 & n2166 ;
  assign n2185 = n2184 ^ n2170 ;
  assign n2175 = n1914 ^ n1670 ;
  assign n2176 = ~n1530 & n1914 ;
  assign n2177 = n2176 ^ n2165 ;
  assign n2178 = n2175 & n2177 ;
  assign n2186 = n2185 ^ n2178 ;
  assign n2173 = n1671 & ~n2167 ;
  assign n4970 = n2186 ^ n2173 ;
  assign n791 = n790 ^ n752 ;
  assign n792 = n791 ^ n787 ;
  assign n772 = n771 ^ n723 ;
  assign n773 = n772 ^ n758 ;
  assign n776 = n315 & n773 ;
  assign n777 = n776 ^ n758 ;
  assign n778 = n770 & n777 ;
  assign n793 = n792 ^ n778 ;
  assign n767 = n315 & n764 ;
  assign n768 = n767 ^ n761 ;
  assign n769 = n219 & ~n768 ;
  assign n794 = n793 ^ n769 ;
  assign n753 = n752 ^ n747 ;
  assign n740 = n739 ^ n720 ;
  assign n743 = n742 ^ n740 ;
  assign n748 = n747 ^ n743 ;
  assign n749 = ~n219 & n748 ;
  assign n754 = n753 ^ n749 ;
  assign n755 = ~n315 & n754 ;
  assign n795 = n794 ^ n755 ;
  assign n798 = n797 ^ n795 ;
  assign n799 = n798 ^ x58 ;
  assign n738 = n316 & ~n737 ;
  assign n800 = n799 ^ n738 ;
  assign n801 = n800 ^ x81 ;
  assign n1162 = n1161 ^ x102 ;
  assign n922 = n921 ^ x78 ;
  assign n959 = n958 ^ x85 ;
  assign n1220 = n922 & n959 ;
  assign n1221 = n1220 ^ n922 ;
  assign n1091 = n1023 & ~n1929 ;
  assign n1083 = n1082 ^ n1016 ;
  assign n1073 = n1022 ^ n1002 ;
  assign n1074 = n1073 ^ n1056 ;
  assign n1075 = n997 & n1074 ;
  assign n1084 = n1083 ^ n1075 ;
  assign n1077 = n1028 ^ n1026 ;
  assign n1078 = ~n997 & n1077 ;
  assign n1085 = n1084 ^ n1078 ;
  assign n1086 = n1037 & n1085 ;
  assign n1072 = n1071 ^ n1057 ;
  assign n1076 = n1075 ^ n1072 ;
  assign n1087 = n1086 ^ n1076 ;
  assign n1092 = n1091 ^ n1087 ;
  assign n1066 = ~n997 & n1061 ;
  assign n1067 = n1066 ^ n1057 ;
  assign n1068 = ~n1037 & n1067 ;
  assign n1093 = n1092 ^ n1068 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1096 = n1095 ^ n1050 ;
  assign n1097 = n1096 ^ n1042 ;
  assign n1098 = n1097 ^ x13 ;
  assign n1099 = n1098 ^ x108 ;
  assign n1103 = n959 & n1099 ;
  assign n1104 = n1103 ^ n1099 ;
  assign n1222 = n1221 ^ n1104 ;
  assign n1113 = ~n922 & ~n1099 ;
  assign n1114 = ~n959 & n1113 ;
  assign n989 = n988 ^ n263 ;
  assign n990 = n282 & ~n989 ;
  assign n980 = n304 ^ n245 ;
  assign n981 = n980 ^ n259 ;
  assign n971 = n235 ^ n232 ;
  assign n972 = n971 ^ n261 ;
  assign n973 = n220 & ~n972 ;
  assign n982 = n981 ^ n973 ;
  assign n983 = n982 ^ n247 ;
  assign n978 = n261 ^ n247 ;
  assign n979 = ~n220 & ~n978 ;
  assign n984 = n983 ^ n979 ;
  assign n985 = ~n977 & ~n984 ;
  assign n974 = n973 ^ n300 ;
  assign n975 = n974 ^ n297 ;
  assign n976 = n975 ^ x21 ;
  assign n986 = n985 ^ n976 ;
  assign n991 = n990 ^ n986 ;
  assign n969 = n253 ^ n232 ;
  assign n970 = ~n283 & n969 ;
  assign n992 = n991 ^ n970 ;
  assign n963 = n304 ^ n241 ;
  assign n966 = ~n269 & n963 ;
  assign n967 = n966 ^ n241 ;
  assign n968 = n220 & n967 ;
  assign n993 = n992 ^ n968 ;
  assign n961 = n255 ^ n239 ;
  assign n962 = n269 & ~n961 ;
  assign n994 = n993 ^ n962 ;
  assign n960 = n239 & n281 ;
  assign n995 = n994 ^ n960 ;
  assign n996 = n995 ^ x91 ;
  assign n1106 = ~n959 & n996 ;
  assign n1100 = ~n996 & n1099 ;
  assign n1101 = n959 & n1100 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1105 = n1104 ^ n1102 ;
  assign n1107 = n1106 ^ n1105 ;
  assign n1108 = ~n922 & n1107 ;
  assign n1115 = n1114 ^ n1108 ;
  assign n1111 = n1106 ^ n1102 ;
  assign n1112 = n1111 ^ n959 ;
  assign n1116 = n1115 ^ n1112 ;
  assign n1109 = n1108 ^ n1106 ;
  assign n1110 = n1109 ^ n1105 ;
  assign n1117 = n1116 ^ n1110 ;
  assign n1223 = n1222 ^ n1117 ;
  assign n1224 = n1223 ^ n1108 ;
  assign n1225 = n1224 ^ n1106 ;
  assign n1208 = n1099 ^ n922 ;
  assign n1209 = n1099 ^ n996 ;
  assign n1210 = n1208 & n1209 ;
  assign n1226 = n1225 ^ n1210 ;
  assign n1215 = n1103 ^ n959 ;
  assign n1204 = n1114 ^ n1113 ;
  assign n1216 = n1215 ^ n1204 ;
  assign n1217 = ~n996 & n1216 ;
  assign n1218 = n1217 ^ n1216 ;
  assign n1211 = n1210 ^ n1099 ;
  assign n1212 = n959 & n1211 ;
  assign n1205 = ~n996 & n1204 ;
  assign n1206 = n1205 ^ n1204 ;
  assign n1203 = n1106 ^ n996 ;
  assign n1207 = n1206 ^ n1203 ;
  assign n1213 = n1212 ^ n1207 ;
  assign n1214 = n1213 ^ n1101 ;
  assign n1219 = n1218 ^ n1214 ;
  assign n1227 = n1226 ^ n1219 ;
  assign n1270 = n1227 ^ n1116 ;
  assign n1271 = ~n1162 & n1270 ;
  assign n1196 = n1195 ^ x84 ;
  assign n1197 = ~n1162 & n1196 ;
  assign n1198 = n1197 ^ n1162 ;
  assign n1240 = n1220 ^ n1216 ;
  assign n1241 = n1240 ^ n1213 ;
  assign n1242 = n1241 ^ n1206 ;
  assign n1259 = n1242 ^ n1218 ;
  assign n1260 = n1259 ^ n1203 ;
  assign n1266 = n1260 ^ n1213 ;
  assign n1265 = n1217 ^ n1214 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1268 = ~n1198 & n1267 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1200 = n1199 ^ n1162 ;
  assign n1261 = n1260 ^ n1219 ;
  assign n1228 = n1227 ^ n1105 ;
  assign n1229 = n1228 ^ n1223 ;
  assign n1230 = n1229 ^ n1102 ;
  assign n1262 = n1261 ^ n1230 ;
  assign n1263 = n1200 & n1262 ;
  assign n1255 = n1108 & n1197 ;
  assign n1239 = n1200 & ~n1228 ;
  assign n1256 = n1255 ^ n1239 ;
  assign n1250 = n1217 ^ n1205 ;
  assign n1251 = n1250 ^ n1225 ;
  assign n1252 = n1199 & ~n1251 ;
  assign n1202 = n1196 ^ n1162 ;
  assign n1243 = n1242 ^ n1239 ;
  assign n1244 = n1243 ^ n1115 ;
  assign n1245 = n1244 ^ n1228 ;
  assign n1246 = n1245 ^ n1239 ;
  assign n1247 = ~n1202 & ~n1246 ;
  assign n1248 = n1247 ^ n1243 ;
  assign n1233 = n1229 ^ n1205 ;
  assign n1236 = n1196 & n1233 ;
  assign n1237 = n1236 ^ n1230 ;
  assign n1238 = n1202 & n1237 ;
  assign n1249 = n1248 ^ n1238 ;
  assign n1253 = n1252 ^ n1249 ;
  assign n1201 = ~n1117 & n1200 ;
  assign n1254 = n1253 ^ n1201 ;
  assign n1257 = n1256 ^ n1254 ;
  assign n1258 = n1257 ^ x32 ;
  assign n1264 = n1263 ^ n1258 ;
  assign n1269 = n1268 ^ n1264 ;
  assign n1272 = n1271 ^ n1269 ;
  assign n1273 = n1272 ^ x72 ;
  assign n1274 = ~n801 & n1273 ;
  assign n4971 = n4970 ^ n1274 ;
  assign n2196 = ~n2167 & n2181 ;
  assign n2197 = n2196 ^ n2186 ;
  assign n2198 = n2197 ^ n2170 ;
  assign n2193 = n2168 & n2179 ;
  assign n2194 = n2193 ^ n2184 ;
  assign n2195 = n2194 ^ n2173 ;
  assign n2199 = n2198 ^ n2195 ;
  assign n2200 = n2199 ^ n2175 ;
  assign n2204 = n2200 ^ n2182 ;
  assign n2203 = n2168 & n2181 ;
  assign n2205 = n2204 ^ n2203 ;
  assign n2201 = n2200 ^ n2196 ;
  assign n2202 = n2201 ^ n2181 ;
  assign n2206 = n2205 ^ n2202 ;
  assign n2191 = ~n2167 & ~n2180 ;
  assign n2223 = n2206 ^ n2191 ;
  assign n2253 = n2223 ^ n2203 ;
  assign n1275 = n1274 ^ n801 ;
  assign n1276 = n1275 ^ n1273 ;
  assign n4972 = n2253 ^ n1276 ;
  assign n4975 = ~n4970 & ~n4972 ;
  assign n4976 = n4975 ^ n1276 ;
  assign n4977 = n4971 & n4976 ;
  assign n2169 = n1671 & n2168 ;
  assign n4963 = n2184 ^ n2169 ;
  assign n2207 = n2206 ^ n2194 ;
  assign n2171 = n2170 ^ n2169 ;
  assign n2192 = n2191 ^ n2171 ;
  assign n2208 = n2207 ^ n2192 ;
  assign n2189 = n2165 ^ n1914 ;
  assign n2188 = n2180 ^ n2176 ;
  assign n2190 = n2189 ^ n2188 ;
  assign n2209 = n2208 ^ n2190 ;
  assign n2210 = n2209 ^ n2193 ;
  assign n4964 = n4963 ^ n2210 ;
  assign n4968 = ~n1275 & n4964 ;
  assign n1277 = n1276 ^ n1274 ;
  assign n2187 = n2186 ^ n2179 ;
  assign n2211 = n2210 ^ n2187 ;
  assign n2241 = n2211 ^ n2200 ;
  assign n2242 = n2200 ^ n801 ;
  assign n2243 = n2242 ^ n2200 ;
  assign n2244 = ~n2241 & ~n2243 ;
  assign n2245 = n2244 ^ n2200 ;
  assign n2246 = ~n1277 & n2245 ;
  assign n4965 = n2246 ^ n801 ;
  assign n4969 = n4968 ^ n4965 ;
  assign n4978 = n4977 ^ n4969 ;
  assign n4958 = n2192 ^ n1273 ;
  assign n4959 = n4958 ^ n2192 ;
  assign n4960 = n2208 & ~n4959 ;
  assign n4961 = n4960 ^ n2192 ;
  assign n4962 = n801 & n4961 ;
  assign n4979 = n4978 ^ n4962 ;
  assign n2239 = ~n1275 & n2201 ;
  assign n4980 = n4979 ^ n2239 ;
  assign n2172 = n2171 ^ n1671 ;
  assign n2174 = n2173 ^ n2172 ;
  assign n2212 = n2211 ^ n2174 ;
  assign n4489 = n2212 ^ n2209 ;
  assign n2254 = n2253 ^ n2188 ;
  assign n4490 = n4489 ^ n2254 ;
  assign n4491 = n2254 ^ n801 ;
  assign n4492 = n4491 ^ n2254 ;
  assign n4493 = ~n4490 & n4492 ;
  assign n4494 = n4493 ^ n2254 ;
  assign n4495 = n1273 & ~n4494 ;
  assign n4981 = n4980 ^ n4495 ;
  assign n2213 = n2212 ^ n2196 ;
  assign n2214 = n2196 ^ n801 ;
  assign n2215 = n2214 ^ n2196 ;
  assign n2216 = ~n2213 & ~n2215 ;
  assign n2217 = n2216 ^ n2196 ;
  assign n2218 = n1277 & n2217 ;
  assign n4982 = n4981 ^ n2218 ;
  assign n4488 = n1276 & ~n2254 ;
  assign n4983 = n4982 ^ n4488 ;
  assign n2237 = n1274 ^ n1273 ;
  assign n4533 = n2203 & n2237 ;
  assign n4984 = n4983 ^ n4533 ;
  assign n4985 = n4984 ^ n1319 ;
  assign n5606 = n4985 ^ x68 ;
  assign n5607 = ~n5605 & ~n5606 ;
  assign n5608 = n5607 ^ n5606 ;
  assign n5609 = n5608 ^ n5605 ;
  assign n2896 = n2895 ^ x97 ;
  assign n2857 = n1913 ^ x107 ;
  assign n3030 = n2896 ^ n2857 ;
  assign n2370 = n1701 ^ x96 ;
  assign n2359 = n2002 ^ x114 ;
  assign n2317 = n2072 ^ x121 ;
  assign n2342 = n2017 ^ n578 ;
  assign n2343 = n615 & ~n2342 ;
  assign n2340 = n2035 ^ n595 ;
  assign n2318 = n1174 ^ n535 ;
  assign n2327 = n2318 ^ n550 ;
  assign n2328 = n2327 ^ n537 ;
  assign n2329 = n2328 ^ n603 ;
  assign n2330 = n522 & ~n2329 ;
  assign n2331 = n2330 ^ n523 ;
  assign n2332 = n561 ^ n546 ;
  assign n2333 = n2332 ^ n1188 ;
  assign n2334 = n2333 ^ n546 ;
  assign n2337 = ~n522 & ~n2334 ;
  assign n2338 = n2337 ^ n546 ;
  assign n2339 = ~n2331 & ~n2338 ;
  assign n2341 = n2340 ^ n2339 ;
  assign n2344 = n2343 ^ n2341 ;
  assign n2326 = ~n523 & n1181 ;
  assign n2345 = n2344 ^ n2326 ;
  assign n2323 = n521 & n2318 ;
  assign n2324 = n2323 ^ n531 ;
  assign n2325 = ~n534 & n2324 ;
  assign n2346 = n2345 ^ n2325 ;
  assign n2347 = n2346 ^ n624 ;
  assign n2348 = n2347 ^ x19 ;
  assign n2349 = n2348 ^ x120 ;
  assign n2350 = n2317 & n2349 ;
  assign n2311 = ~n148 & n1560 ;
  assign n2306 = n955 ^ n202 ;
  assign n2292 = n133 ^ n131 ;
  assign n2293 = n2292 ^ n130 ;
  assign n2294 = n2293 ^ n155 ;
  assign n2283 = n1564 ^ n166 ;
  assign n2295 = n2294 ^ n2283 ;
  assign n2296 = n140 & ~n2295 ;
  assign n2297 = n2296 ^ n2283 ;
  assign n2307 = n2306 ^ n2297 ;
  assign n2308 = n2307 ^ x11 ;
  assign n2299 = n169 ^ n158 ;
  assign n2300 = n2299 ^ n2297 ;
  assign n2298 = n2297 ^ n1560 ;
  assign n2301 = n2300 ^ n2298 ;
  assign n2302 = n2301 ^ n199 ;
  assign n2303 = ~n140 & n2302 ;
  assign n2304 = n2303 ^ n2300 ;
  assign n2305 = n129 & n2304 ;
  assign n2309 = n2308 ^ n2305 ;
  assign n2291 = n146 & n184 ;
  assign n2310 = n2309 ^ n2291 ;
  assign n2312 = n2311 ^ n2310 ;
  assign n2288 = n129 & n2283 ;
  assign n2289 = n2288 ^ n202 ;
  assign n2290 = n147 & n2289 ;
  assign n2313 = n2312 ^ n2290 ;
  assign n2314 = n2313 ^ x82 ;
  assign n2315 = n1823 ^ x73 ;
  assign n2316 = ~n2314 & n2315 ;
  assign n2354 = n2316 ^ n2314 ;
  assign n2355 = n2354 ^ n2315 ;
  assign n2371 = n2350 & n2355 ;
  assign n2352 = n2349 ^ n2317 ;
  assign n2351 = ~n2316 & ~n2350 ;
  assign n2353 = n2352 ^ n2351 ;
  assign n2356 = ~n2317 & n2355 ;
  assign n2357 = ~n2353 & ~n2356 ;
  assign n2358 = n2357 ^ n2353 ;
  assign n2947 = n2371 ^ n2358 ;
  assign n2946 = n2356 ^ n2355 ;
  assign n2948 = n2947 ^ n2946 ;
  assign n2372 = n2371 ^ n2350 ;
  assign n2949 = n2948 ^ n2372 ;
  assign n2373 = n2315 & n2352 ;
  assign n2943 = n2373 ^ n2358 ;
  assign n2365 = n2352 ^ n2350 ;
  assign n2364 = ~n2317 & ~n2354 ;
  assign n2366 = n2365 ^ n2364 ;
  assign n2360 = ~n2315 & n2350 ;
  assign n2361 = n2360 ^ n2357 ;
  assign n2362 = n2361 ^ n2314 ;
  assign n2363 = n2362 ^ n2360 ;
  assign n2367 = n2366 ^ n2363 ;
  assign n2368 = n2359 & n2367 ;
  assign n2369 = n2368 ^ n2361 ;
  assign n2944 = n2943 ^ n2369 ;
  assign n2376 = n2316 & ~n2317 ;
  assign n2945 = n2944 ^ n2376 ;
  assign n2950 = n2949 ^ n2945 ;
  assign n2951 = n2950 ^ n2369 ;
  assign n2952 = ~n2359 & n2951 ;
  assign n2953 = n2952 ^ n2944 ;
  assign n2954 = ~n2370 & ~n2953 ;
  assign n3238 = n2355 ^ n2314 ;
  assign n2391 = ~n2349 & n3238 ;
  assign n2392 = n2391 ^ n2354 ;
  assign n2393 = ~n2317 & ~n2392 ;
  assign n2394 = n2393 ^ n2354 ;
  assign n2395 = n2359 & ~n2394 ;
  assign n2396 = n2370 & n2395 ;
  assign n2939 = n2396 ^ n2395 ;
  assign n2384 = n2355 & n2370 ;
  assign n2936 = n2384 ^ n2355 ;
  assign n2937 = ~n2359 & ~n2365 ;
  assign n2938 = n2936 & n2937 ;
  assign n2940 = n2939 ^ n2938 ;
  assign n2941 = n2940 ^ x50 ;
  assign n2942 = n2941 ^ n2369 ;
  assign n2955 = n2954 ^ n2942 ;
  assign n2956 = n2955 ^ x65 ;
  assign n2984 = n2983 ^ x112 ;
  assign n2985 = ~n2956 & n2984 ;
  assign n2897 = n800 ^ x74 ;
  assign n2669 = n1114 ^ n1112 ;
  assign n2670 = n2669 ^ n1213 ;
  assign n2673 = n1196 & ~n2670 ;
  assign n2674 = n2673 ^ n1213 ;
  assign n2675 = n1162 & n2674 ;
  assign n2928 = n1197 & n1229 ;
  assign n2915 = ~n1200 & ~n1206 ;
  assign n2920 = n1260 & ~n2915 ;
  assign n2916 = ~n1213 & n2915 ;
  assign n2918 = ~n1250 & n2916 ;
  assign n2917 = n2916 ^ n1250 ;
  assign n2919 = n2918 ^ n2917 ;
  assign n2921 = n2920 ^ n2919 ;
  assign n2667 = ~n1198 & n1206 ;
  assign n2914 = n2667 ^ n1218 ;
  assign n2922 = n2921 ^ n2914 ;
  assign n2923 = n2922 ^ n1227 ;
  assign n2909 = n1265 ^ n1110 ;
  assign n2910 = ~n1162 & n2909 ;
  assign n2924 = n2923 ^ n2910 ;
  assign n2925 = ~n1202 & ~n2924 ;
  assign n2905 = ~n1196 & n1214 ;
  assign n2906 = n2905 ^ n1230 ;
  assign n2907 = n1162 & n2906 ;
  assign n2908 = n2907 ^ n1230 ;
  assign n2911 = n2910 ^ n2908 ;
  assign n2695 = n1265 ^ n1242 ;
  assign n2698 = ~n1196 & n2695 ;
  assign n2699 = n2698 ^ n1242 ;
  assign n2700 = ~n1162 & n2699 ;
  assign n2912 = n2911 ^ n2700 ;
  assign n2900 = n1212 ^ n1208 ;
  assign n2901 = n2900 ^ n996 ;
  assign n2902 = n1199 & ~n2901 ;
  assign n2913 = n2912 ^ n2902 ;
  assign n2926 = n2925 ^ n2913 ;
  assign n2898 = n1229 ^ n1115 ;
  assign n2899 = ~n1162 & n2898 ;
  assign n2927 = n2926 ^ n2899 ;
  assign n2929 = n2928 ^ n2927 ;
  assign n2930 = ~n1256 & ~n2929 ;
  assign n2931 = ~n2675 & n2930 ;
  assign n2932 = n2931 ^ x42 ;
  assign n2933 = n2932 ^ x64 ;
  assign n2934 = ~n2897 & ~n2933 ;
  assign n2991 = n2934 ^ n2933 ;
  assign n3005 = n2991 ^ n2897 ;
  assign n3014 = n2985 & ~n3005 ;
  assign n2935 = n2934 ^ n2897 ;
  assign n3012 = ~n2935 & n2985 ;
  assign n3001 = n2984 ^ n2956 ;
  assign n3002 = n3001 ^ n2933 ;
  assign n3003 = n3002 ^ n2985 ;
  assign n3004 = n2897 & n3003 ;
  assign n3006 = n3005 ^ n3004 ;
  assign n2986 = n2985 ^ n2984 ;
  assign n2987 = n2986 ^ n2956 ;
  assign n2988 = ~n2935 & n2987 ;
  assign n3000 = n2988 ^ n2987 ;
  assign n3007 = n3006 ^ n3000 ;
  assign n2989 = n2934 & n2986 ;
  assign n3008 = n3007 ^ n2989 ;
  assign n2992 = n2987 ^ n2984 ;
  assign n2998 = n2934 & ~n2992 ;
  assign n2996 = ~n2935 & n2986 ;
  assign n2999 = n2998 ^ n2996 ;
  assign n3009 = n3008 ^ n2999 ;
  assign n2997 = n2996 ^ n2934 ;
  assign n3010 = n3009 ^ n2997 ;
  assign n3011 = n3010 ^ n2988 ;
  assign n3013 = n3012 ^ n3011 ;
  assign n3015 = n3014 ^ n3013 ;
  assign n5185 = n3014 ^ n2857 ;
  assign n5186 = n5185 ^ n3014 ;
  assign n5189 = ~n3015 & ~n5186 ;
  assign n5190 = n5189 ^ n3014 ;
  assign n5191 = n3030 & n5190 ;
  assign n2995 = n2988 ^ n2985 ;
  assign n3016 = n3015 ^ n2995 ;
  assign n3033 = n3016 ^ n2991 ;
  assign n3020 = n2986 & ~n2991 ;
  assign n2993 = ~n2991 & ~n2992 ;
  assign n3021 = n3020 ^ n2993 ;
  assign n3034 = n3033 ^ n3021 ;
  assign n3035 = n3034 ^ n3006 ;
  assign n4100 = n3035 ^ n3011 ;
  assign n4101 = n4100 ^ n3035 ;
  assign n4102 = n3035 ^ n2896 ;
  assign n4103 = n4102 ^ n3035 ;
  assign n4104 = ~n4101 & n4103 ;
  assign n4105 = n4104 ^ n3035 ;
  assign n4106 = ~n3030 & ~n4105 ;
  assign n4107 = n4106 ^ n3035 ;
  assign n3066 = ~n2857 & ~n2896 ;
  assign n3032 = ~n2992 & ~n3005 ;
  assign n3036 = n3035 ^ n3032 ;
  assign n3031 = n3014 ^ n3005 ;
  assign n3037 = n3036 ^ n3031 ;
  assign n5172 = n3037 ^ n2993 ;
  assign n5173 = n5172 ^ n3032 ;
  assign n5625 = n5173 ^ n3007 ;
  assign n5626 = n3066 & ~n5625 ;
  assign n3067 = n3066 ^ n2896 ;
  assign n3068 = n3067 ^ n2857 ;
  assign n4090 = n3068 ^ n2896 ;
  assign n5166 = n3014 ^ n2998 ;
  assign n5167 = n5166 ^ n2989 ;
  assign n5621 = n5167 ^ n3034 ;
  assign n5622 = ~n4090 & n5621 ;
  assign n3039 = n3012 ^ n2999 ;
  assign n4088 = ~n3039 & n3067 ;
  assign n3040 = n3011 ^ n3008 ;
  assign n3041 = n3040 ^ n2897 ;
  assign n3042 = n3041 ^ n3039 ;
  assign n4091 = n3042 ^ n3007 ;
  assign n5619 = n4091 ^ n3066 ;
  assign n5620 = ~n4088 & n5619 ;
  assign n5623 = n5622 ^ n5620 ;
  assign n5624 = n5623 ^ n3010 ;
  assign n5627 = n5626 ^ n5624 ;
  assign n4109 = n3034 ^ n3016 ;
  assign n4110 = n4109 ^ n3032 ;
  assign n5611 = n4110 ^ n3037 ;
  assign n5612 = n5611 ^ n2998 ;
  assign n5613 = n5612 ^ n4110 ;
  assign n5614 = n4110 ^ n2896 ;
  assign n5615 = n5614 ^ n4110 ;
  assign n5616 = n5613 & n5615 ;
  assign n5617 = n5616 ^ n4110 ;
  assign n5618 = n2857 & ~n5617 ;
  assign n5628 = n5627 ^ n5618 ;
  assign n5629 = n4107 & n5628 ;
  assign n5630 = ~n5191 & n5629 ;
  assign n3069 = n3012 & ~n3068 ;
  assign n5610 = n3069 ^ n1361 ;
  assign n5631 = n5630 ^ n5610 ;
  assign n5632 = n5631 ^ x67 ;
  assign n3239 = n3238 ^ n2354 ;
  assign n3236 = n2350 ^ n2317 ;
  assign n3237 = n3236 ^ n2946 ;
  assign n3240 = n3239 ^ n3237 ;
  assign n3245 = n3240 ^ n2370 ;
  assign n3226 = n2349 ^ n2314 ;
  assign n3227 = n2364 & ~n3226 ;
  assign n3241 = n3227 ^ n2949 ;
  assign n3242 = n3241 ^ n3240 ;
  assign n3243 = ~n2370 & n3242 ;
  assign n3244 = n3243 ^ n3241 ;
  assign n3246 = n3245 ^ n3244 ;
  assign n3247 = n3246 ^ n3241 ;
  assign n3225 = n2393 ^ n2366 ;
  assign n3228 = n3227 ^ n3225 ;
  assign n3222 = n2317 ^ n2314 ;
  assign n3223 = n3222 ^ n2376 ;
  assign n3224 = n3223 ^ n2946 ;
  assign n3229 = n3228 ^ n3224 ;
  assign n3230 = n3229 ^ n2360 ;
  assign n3248 = n3247 ^ n3230 ;
  assign n3232 = n3224 ^ n2373 ;
  assign n3233 = n3232 ^ n3227 ;
  assign n3231 = n3230 ^ n2946 ;
  assign n3234 = n3233 ^ n3231 ;
  assign n3235 = ~n2370 & ~n3234 ;
  assign n3249 = n3248 ^ n3235 ;
  assign n3250 = ~n2359 & ~n3249 ;
  assign n3251 = n3250 ^ n3247 ;
  assign n3252 = ~n2940 & n3251 ;
  assign n3253 = n3252 ^ x36 ;
  assign n4371 = n3253 ^ x86 ;
  assign n3483 = n1784 ^ n1778 ;
  assign n3484 = n1873 & n3483 ;
  assign n3479 = n1860 ^ n1841 ;
  assign n3480 = n1672 & n3479 ;
  assign n3474 = n1911 ^ n1860 ;
  assign n3468 = n1851 ^ n1784 ;
  assign n3471 = ~n1824 & n3468 ;
  assign n3472 = n3471 ^ n1851 ;
  assign n3473 = ~n1835 & n3472 ;
  assign n3475 = n3474 ^ n3473 ;
  assign n3476 = n3475 ^ n3467 ;
  assign n3477 = n3476 ^ x62 ;
  assign n3454 = n1883 ^ n1860 ;
  assign n3455 = n3454 ^ n1850 ;
  assign n3456 = n3455 ^ n1883 ;
  assign n3459 = ~n1672 & n3456 ;
  assign n3460 = n3459 ^ n1883 ;
  assign n3461 = n1824 & n3460 ;
  assign n3478 = n3477 ^ n3461 ;
  assign n3481 = n3480 ^ n3478 ;
  assign n3453 = n1849 & n1909 ;
  assign n3482 = n3481 ^ n3453 ;
  assign n3485 = n3484 ^ n3482 ;
  assign n3452 = ~n1832 & ~n3451 ;
  assign n3486 = n3485 ^ n3452 ;
  assign n3443 = n3442 ^ n1782 ;
  assign n3441 = n1839 ^ n1779 ;
  assign n3444 = n3443 ^ n3441 ;
  assign n3447 = n1824 & n3444 ;
  assign n3448 = n3447 ^ n3441 ;
  assign n3449 = n1835 & n3448 ;
  assign n3487 = n3486 ^ n3449 ;
  assign n4265 = n3487 ^ x68 ;
  assign n3114 = n1493 ^ n1478 ;
  assign n3115 = n3114 ^ n1515 ;
  assign n3112 = n1490 ^ n1465 ;
  assign n3113 = n3112 ^ n1482 ;
  assign n3116 = n3115 ^ n3113 ;
  assign n3117 = ~n1320 & n3116 ;
  assign n3118 = n3117 ^ n3115 ;
  assign n3119 = ~n1467 & n3118 ;
  assign n3105 = n1482 ^ n1472 ;
  assign n3106 = n3105 ^ n1492 ;
  assign n3107 = n1321 & ~n3106 ;
  assign n3108 = n3107 ^ n1488 ;
  assign n3109 = n1467 & n3108 ;
  assign n3087 = n3827 ^ n1467 ;
  assign n3090 = ~n1510 & n3087 ;
  assign n3091 = n3090 ^ n1467 ;
  assign n3097 = n1321 & n1483 ;
  assign n3098 = n3097 ^ n1482 ;
  assign n3099 = n1320 & n3098 ;
  assign n3101 = n3099 ^ n1320 ;
  assign n3092 = n1510 ^ n1322 ;
  assign n3100 = n3099 ^ n3092 ;
  assign n3102 = n3101 ^ n3100 ;
  assign n3103 = ~n3091 & ~n3102 ;
  assign n3104 = n3103 ^ n3101 ;
  assign n3110 = n3109 ^ n3104 ;
  assign n3084 = n1478 ^ n1474 ;
  assign n3085 = n1324 & n3084 ;
  assign n3111 = n3110 ^ n3085 ;
  assign n3120 = n3119 ^ n3111 ;
  assign n3121 = n3120 ^ n1521 ;
  assign n3122 = n3121 ^ n1527 ;
  assign n3123 = n3122 ^ n3083 ;
  assign n3124 = n3123 ^ n3077 ;
  assign n3125 = n3124 ^ x28 ;
  assign n4302 = n3125 ^ x69 ;
  assign n4323 = n1662 ^ n1602 ;
  assign n4324 = n4323 ^ n1624 ;
  assign n4325 = n1531 & n4324 ;
  assign n4315 = n1601 ^ n1585 ;
  assign n4326 = n4325 ^ n4315 ;
  assign n4327 = n1584 & n4326 ;
  assign n4303 = ~n1584 & ~n1661 ;
  assign n4314 = n4303 ^ n1608 ;
  assign n4316 = n4315 ^ n4314 ;
  assign n4317 = n4316 ^ n2963 ;
  assign n4318 = n4317 ^ n2977 ;
  assign n4319 = n4318 ^ n1639 ;
  assign n4320 = n4319 ^ x20 ;
  assign n4309 = n1660 ^ n1593 ;
  assign n4306 = n1595 ^ n1581 ;
  assign n4307 = n4306 ^ n1612 ;
  assign n4310 = n4309 ^ n4307 ;
  assign n4311 = n1583 & n4310 ;
  assign n4308 = n4307 ^ n1608 ;
  assign n4312 = n4311 ^ n4308 ;
  assign n4313 = ~n1531 & n4312 ;
  assign n4321 = n4320 ^ n4313 ;
  assign n4304 = n1583 & ~n1594 ;
  assign n4305 = n4303 & n4304 ;
  assign n4322 = n4321 ^ n4305 ;
  assign n4328 = n4327 ^ n4322 ;
  assign n4329 = n4328 ^ x75 ;
  assign n4330 = ~n4302 & ~n4329 ;
  assign n4331 = n4330 ^ n4302 ;
  assign n2633 = n2010 & n2632 ;
  assign n2634 = n2633 ^ n2129 ;
  assign n3549 = n2634 ^ x4 ;
  assign n3534 = n2103 ^ n2089 ;
  assign n3535 = n3534 ^ n2116 ;
  assign n3544 = n3535 ^ n3154 ;
  assign n3538 = n2097 ^ n2079 ;
  assign n3539 = n3538 ^ n2106 ;
  assign n3540 = n3539 ^ n2155 ;
  assign n3541 = ~n2046 & ~n3540 ;
  assign n3536 = n3535 ^ n2087 ;
  assign n2635 = n2116 ^ n2013 ;
  assign n2636 = n2046 & ~n2635 ;
  assign n2637 = n2636 ^ n2013 ;
  assign n3537 = n3536 ^ n2637 ;
  assign n3542 = n3541 ^ n3537 ;
  assign n3543 = ~n2114 & n3542 ;
  assign n3545 = n3544 ^ n3543 ;
  assign n3533 = n2075 & n2138 ;
  assign n3546 = n3545 ^ n3533 ;
  assign n3527 = n2644 ^ n2094 ;
  assign n3530 = n2046 & n3527 ;
  assign n3531 = n3530 ^ n2094 ;
  assign n3532 = n2073 & n3531 ;
  assign n3547 = n3546 ^ n3532 ;
  assign n3548 = ~n3128 & ~n3547 ;
  assign n3550 = n3549 ^ n3548 ;
  assign n4266 = n3550 ^ x125 ;
  assign n4298 = n219 & n720 ;
  assign n4295 = n732 & ~n788 ;
  assign n4284 = n746 ^ n736 ;
  assign n4293 = n2574 & n4284 ;
  assign n4282 = n728 ^ n722 ;
  assign n4283 = n4282 ^ n797 ;
  assign n4285 = n4284 ^ n4283 ;
  assign n4286 = n785 & ~n4285 ;
  assign n4275 = n744 ^ n735 ;
  assign n4278 = n4275 ^ n739 ;
  assign n4279 = n316 & ~n4278 ;
  assign n4280 = n4279 ^ n2625 ;
  assign n4276 = n4275 ^ n728 ;
  assign n4277 = ~n788 & ~n4276 ;
  assign n4281 = n4280 ^ n4277 ;
  assign n4287 = n4286 ^ n4281 ;
  assign n2594 = n2593 ^ n757 ;
  assign n4269 = n3260 ^ n2594 ;
  assign n4272 = ~n219 & n4269 ;
  assign n4273 = n4272 ^ n2594 ;
  assign n4274 = n315 & n4273 ;
  assign n4288 = n4287 ^ n4274 ;
  assign n4289 = n4288 ^ n3278 ;
  assign n4290 = n4289 ^ n786 ;
  assign n2617 = ~n315 & n741 ;
  assign n2610 = n764 ^ n733 ;
  assign n2611 = ~n219 & n2610 ;
  assign n2612 = n2611 ^ n764 ;
  assign n2618 = n2617 ^ n2612 ;
  assign n2619 = ~n770 & n2618 ;
  assign n2620 = n2619 ^ n2612 ;
  assign n4291 = n4290 ^ n2620 ;
  assign n4292 = n4291 ^ x12 ;
  assign n4294 = n4293 ^ n4292 ;
  assign n4296 = n4295 ^ n4294 ;
  assign n4267 = n760 ^ n720 ;
  assign n4268 = ~n315 & n4267 ;
  assign n4297 = n4296 ^ n4268 ;
  assign n4299 = n4298 ^ n4297 ;
  assign n4300 = n4299 ^ x92 ;
  assign n4301 = n4266 & ~n4300 ;
  assign n4352 = n4301 ^ n4300 ;
  assign n4373 = ~n4331 & ~n4352 ;
  assign n4334 = n4301 ^ n4266 ;
  assign n4335 = n4330 ^ n4329 ;
  assign n4336 = n4334 & ~n4335 ;
  assign n5061 = n4373 ^ n4336 ;
  assign n4364 = n4301 & n4330 ;
  assign n4395 = n4364 ^ n4330 ;
  assign n4359 = n4330 & ~n4352 ;
  assign n4358 = n4330 & n4334 ;
  assign n4360 = n4359 ^ n4358 ;
  assign n4396 = n4395 ^ n4360 ;
  assign n4760 = n4396 ^ n4364 ;
  assign n5062 = n5061 ^ n4760 ;
  assign n4353 = n4352 ^ n4266 ;
  assign n4357 = ~n4331 & n4353 ;
  assign n4361 = n4360 ^ n4357 ;
  assign n4339 = n4329 ^ n4302 ;
  assign n4341 = n4339 ^ n4266 ;
  assign n4342 = n4341 ^ n4300 ;
  assign n4343 = ~n4302 & ~n4342 ;
  assign n4362 = n4361 ^ n4343 ;
  assign n4346 = n4301 & ~n4335 ;
  assign n4347 = n4346 ^ n4301 ;
  assign n4338 = n4300 ^ n4266 ;
  assign n4340 = n4339 ^ n4300 ;
  assign n4344 = n4343 ^ n4340 ;
  assign n4345 = n4338 & ~n4344 ;
  assign n4348 = n4347 ^ n4345 ;
  assign n4349 = n4348 ^ n4346 ;
  assign n4337 = n4336 ^ n4335 ;
  assign n4350 = n4349 ^ n4337 ;
  assign n4332 = n4331 ^ n4329 ;
  assign n4333 = n4301 & ~n4332 ;
  assign n4351 = n4350 ^ n4333 ;
  assign n5060 = n4362 ^ n4351 ;
  assign n5063 = n5062 ^ n5060 ;
  assign n5064 = ~n4265 & ~n5063 ;
  assign n5065 = n5064 ^ n5060 ;
  assign n5066 = ~n4371 & ~n5065 ;
  assign n4372 = ~n4265 & ~n4371 ;
  assign n4381 = n4372 ^ n4371 ;
  assign n4382 = n4381 ^ n4265 ;
  assign n4388 = n4382 ^ n4371 ;
  assign n4374 = n4373 ^ n4359 ;
  assign n4375 = n4374 ^ n4352 ;
  assign n4376 = n4375 ^ n4350 ;
  assign n4354 = ~n4332 & n4353 ;
  assign n4402 = n4376 ^ n4354 ;
  assign n4401 = n4333 ^ n4332 ;
  assign n4403 = n4402 ^ n4401 ;
  assign n4404 = n4403 ^ n4350 ;
  assign n5056 = n4404 ^ n4376 ;
  assign n5057 = ~n4388 & n5056 ;
  assign n4363 = n4362 ^ n4357 ;
  assign n4397 = n4381 & ~n4396 ;
  assign n5037 = ~n4363 & n4397 ;
  assign n5039 = ~n4361 & n4382 ;
  assign n5040 = ~n5037 & n5039 ;
  assign n4390 = n4373 ^ n4331 ;
  assign n4391 = n4390 ^ n4363 ;
  assign n5038 = n5037 ^ n4391 ;
  assign n5041 = n5040 ^ n5038 ;
  assign n5053 = n5041 ^ n1460 ;
  assign n5050 = n4329 ^ n4266 ;
  assign n5051 = n4302 & ~n4382 ;
  assign n5052 = n5050 & n5051 ;
  assign n5054 = n5053 ^ n5052 ;
  assign n5043 = n5041 ^ n4343 ;
  assign n5042 = n5041 ^ n4332 ;
  assign n5044 = n5043 ^ n5042 ;
  assign n5045 = n5043 ^ n4371 ;
  assign n5046 = n5045 ^ n5043 ;
  assign n5047 = ~n5044 & ~n5046 ;
  assign n5048 = n5047 ^ n5043 ;
  assign n5049 = ~n4265 & n5048 ;
  assign n5055 = n5054 ^ n5049 ;
  assign n5058 = n5057 ^ n5055 ;
  assign n4387 = n4371 ^ n4265 ;
  assign n5036 = n4348 & n4387 ;
  assign n5059 = n5058 ^ n5036 ;
  assign n5067 = n5066 ^ n5059 ;
  assign n5633 = n5067 ^ x100 ;
  assign n5634 = ~n5632 & ~n5633 ;
  assign n5635 = n5634 ^ n5632 ;
  assign n3551 = n3550 ^ x100 ;
  assign n2562 = n2477 & ~n2561 ;
  assign n2563 = n2562 ^ n2559 ;
  assign n2541 = ~n2402 & n2536 ;
  assign n2542 = n2541 ^ n2462 ;
  assign n2543 = ~n2401 & n2542 ;
  assign n2497 = n2477 ^ n2469 ;
  assign n2498 = n2497 ^ n2496 ;
  assign n2499 = n2498 ^ n2488 ;
  assign n2492 = n2491 ^ n2476 ;
  assign n2493 = n2492 ^ n2479 ;
  assign n2494 = n2493 ^ n2465 ;
  assign n2500 = n2499 ^ n2494 ;
  assign n2501 = ~n2402 & ~n2500 ;
  assign n2502 = n2501 ^ n2493 ;
  assign n2544 = n2543 ^ n2502 ;
  assign n2533 = n2402 & ~n2508 ;
  assign n2534 = n2533 ^ n2481 ;
  assign n2535 = ~n2528 & ~n2534 ;
  assign n2545 = n2544 ^ n2535 ;
  assign n2522 = n2511 ^ n2471 ;
  assign n2525 = n2401 & n2522 ;
  assign n2526 = n2525 ^ n2471 ;
  assign n2527 = n2402 & n2526 ;
  assign n2546 = n2545 ^ n2527 ;
  assign n2557 = n2556 ^ n2546 ;
  assign n2564 = n2563 ^ n2557 ;
  assign n2568 = n2567 ^ n2564 ;
  assign n2569 = n2568 ^ x38 ;
  assign n2515 = n2502 ^ n2470 ;
  assign n2514 = n2513 ^ n2502 ;
  assign n2516 = n2515 ^ n2514 ;
  assign n2519 = ~n2402 & n2516 ;
  assign n2520 = n2519 ^ n2515 ;
  assign n2521 = ~n2401 & ~n2520 ;
  assign n2570 = n2569 ^ n2521 ;
  assign n3492 = n2570 ^ x117 ;
  assign n2385 = ~n2349 & ~n2359 ;
  assign n2386 = n2384 & n2385 ;
  assign n2397 = n2396 ^ n2386 ;
  assign n3428 = n3230 ^ n2371 ;
  assign n3429 = n3428 ^ n3233 ;
  assign n3430 = n2370 & n3429 ;
  assign n3431 = n3430 ^ n3230 ;
  assign n3432 = n3431 ^ n3244 ;
  assign n3435 = n2359 & n3432 ;
  assign n3436 = n3435 ^ n3431 ;
  assign n3437 = ~n2397 & n3436 ;
  assign n3438 = n3437 ^ x54 ;
  assign n3439 = n3438 ^ x77 ;
  assign n3559 = n3492 ^ n3439 ;
  assign n3488 = n3487 ^ x91 ;
  assign n3560 = n3559 ^ n3488 ;
  assign n3414 = n1484 ^ n1479 ;
  assign n3411 = n1487 ^ n1479 ;
  assign n3412 = n3411 ^ n1476 ;
  assign n3413 = n1320 & ~n3412 ;
  assign n3415 = n3414 ^ n3413 ;
  assign n3416 = n1321 & n3415 ;
  assign n3402 = n3827 ^ n3115 ;
  assign n3403 = n3402 ^ n1491 ;
  assign n3404 = n3827 ^ n3403 ;
  assign n3407 = ~n1321 & n3404 ;
  assign n3408 = n3827 ^ n3407 ;
  assign n3409 = n1320 & n3408 ;
  assign n3410 = n3827 ^ n3409 ;
  assign n3417 = n3416 ^ n3410 ;
  assign n3418 = n3417 ^ n1474 ;
  assign n3398 = n1501 ^ n1474 ;
  assign n3400 = n3399 ^ n3398 ;
  assign n3401 = n1323 & n3400 ;
  assign n3419 = n3418 ^ n3401 ;
  assign n3420 = n3419 ^ n1512 ;
  assign n3421 = n3420 ^ n3099 ;
  assign n3422 = n3421 ^ n1466 ;
  assign n3423 = n3422 ^ n1527 ;
  assign n3424 = n3423 ^ n3083 ;
  assign n3425 = n3424 ^ n3077 ;
  assign n3426 = n3425 ^ x46 ;
  assign n3427 = n3426 ^ x102 ;
  assign n3489 = n3488 ^ n3427 ;
  assign n3569 = n3439 & ~n3489 ;
  assign n3570 = ~n3560 & n3569 ;
  assign n3571 = n3570 ^ n3560 ;
  assign n3501 = ~n3427 & n3488 ;
  assign n3504 = n3439 & ~n3492 ;
  assign n3505 = n3504 ^ n3439 ;
  assign n3519 = n3501 & n3505 ;
  assign n3503 = n3501 ^ n3488 ;
  assign n3510 = n3503 ^ n3427 ;
  assign n3512 = n3510 ^ n3488 ;
  assign n3513 = n3504 & ~n3512 ;
  assign n3511 = n3504 & n3510 ;
  assign n3514 = n3513 ^ n3511 ;
  assign n3508 = n3503 & n3504 ;
  assign n3509 = n3508 ^ n3504 ;
  assign n3515 = n3514 ^ n3509 ;
  assign n3520 = n3519 ^ n3515 ;
  assign n3506 = n3505 ^ n3492 ;
  assign n3517 = n3501 & n3506 ;
  assign n3518 = n3517 ^ n3501 ;
  assign n3521 = n3520 ^ n3518 ;
  assign n3507 = n3503 & n3506 ;
  assign n3516 = n3515 ^ n3507 ;
  assign n3522 = n3521 ^ n3516 ;
  assign n3500 = n3488 & n3492 ;
  assign n3502 = n3501 ^ n3500 ;
  assign n3523 = n3522 ^ n3502 ;
  assign n3524 = n3523 ^ n3521 ;
  assign n3566 = n3524 ^ n3508 ;
  assign n3562 = n3492 ^ n3427 ;
  assign n3563 = n3562 ^ n3439 ;
  assign n3564 = n3563 ^ n3492 ;
  assign n3565 = n3564 ^ n3517 ;
  assign n3567 = n3566 ^ n3565 ;
  assign n3568 = n3567 ^ n3562 ;
  assign n3572 = n3571 ^ n3568 ;
  assign n3440 = n3439 ^ n3427 ;
  assign n3557 = n3500 ^ n3427 ;
  assign n3558 = ~n3440 & ~n3557 ;
  assign n3561 = n3560 ^ n3558 ;
  assign n3972 = n3572 ^ n3561 ;
  assign n3493 = n3492 ^ n3489 ;
  assign n3496 = ~n3427 & n3493 ;
  assign n3497 = n3496 ^ n3489 ;
  assign n3498 = ~n3440 & ~n3497 ;
  assign n3499 = n3498 ^ n3493 ;
  assign n3525 = n3524 ^ n3499 ;
  assign n3973 = n3972 ^ n3525 ;
  assign n3975 = n3973 ^ n3517 ;
  assign n2668 = ~n1202 & n1241 ;
  assign n2691 = n1197 & n1266 ;
  assign n2684 = n1230 ^ n1206 ;
  assign n2678 = n1225 ^ n1115 ;
  assign n2676 = n1107 ^ n959 ;
  assign n2677 = ~n1196 & ~n2676 ;
  assign n2679 = n2678 ^ n2677 ;
  assign n2685 = n2684 ^ n2679 ;
  assign n2681 = n1218 ^ n1106 ;
  assign n2682 = n2681 ^ n1233 ;
  assign n2683 = n2682 ^ n2679 ;
  assign n2686 = n2685 ^ n2683 ;
  assign n2687 = n1196 & n2686 ;
  assign n2688 = n2687 ^ n2683 ;
  assign n2689 = n1162 & ~n2688 ;
  assign n2680 = n2679 ^ n2675 ;
  assign n2690 = n2689 ^ n2680 ;
  assign n2692 = n2691 ^ n2690 ;
  assign n2693 = ~n2668 & n2692 ;
  assign n2694 = ~n2667 & n2693 ;
  assign n2701 = n2694 & ~n2700 ;
  assign n2704 = n2701 ^ x30 ;
  assign n2666 = n1265 ^ n1260 ;
  assign n2702 = n1200 & n2701 ;
  assign n2703 = n2666 & n2702 ;
  assign n2705 = n2704 ^ n2703 ;
  assign n3397 = n2705 ^ x126 ;
  assign n4552 = n3517 ^ n3397 ;
  assign n4553 = n4552 ^ n3517 ;
  assign n4554 = n3975 & ~n4553 ;
  assign n4555 = n4554 ^ n3517 ;
  assign n4556 = n3551 & n4555 ;
  assign n4557 = n4556 ^ n3397 ;
  assign n4558 = n4557 ^ n4556 ;
  assign n4027 = n3508 ^ n3507 ;
  assign n4028 = n4027 ^ n3503 ;
  assign n4559 = n4028 ^ n3523 ;
  assign n3979 = n3506 ^ n3439 ;
  assign n3980 = n3510 & ~n3979 ;
  assign n4565 = n3980 ^ n3512 ;
  assign n3976 = n3571 ^ n3562 ;
  assign n3977 = n3976 ^ n3975 ;
  assign n3978 = n3977 ^ n3513 ;
  assign n3981 = n3980 ^ n3978 ;
  assign n3974 = n3973 ^ n3524 ;
  assign n3982 = n3981 ^ n3974 ;
  assign n4562 = n3982 ^ n3513 ;
  assign n4566 = n4565 ^ n4562 ;
  assign n4010 = n3570 ^ n3508 ;
  assign n4567 = n4566 ^ n4010 ;
  assign n4568 = ~n3551 & ~n4567 ;
  assign n4014 = n3978 ^ n3512 ;
  assign n4560 = n4014 ^ n4010 ;
  assign n3997 = n3511 ^ n3510 ;
  assign n3983 = n3982 ^ n3980 ;
  assign n3998 = n3997 ^ n3983 ;
  assign n4561 = n4560 ^ n3998 ;
  assign n4563 = n4562 ^ n4561 ;
  assign n4564 = n4563 ^ n4559 ;
  assign n4569 = n4568 ^ n4564 ;
  assign n4570 = ~n4559 & n4569 ;
  assign n4571 = n4558 & n4570 ;
  assign n4572 = n4571 ^ n4557 ;
  assign n4573 = n4572 ^ n4556 ;
  assign n3992 = n3397 & ~n3551 ;
  assign n4574 = n3524 ^ n3519 ;
  assign n4575 = n3992 & n4574 ;
  assign n4576 = ~n4573 & n4575 ;
  assign n4577 = n4576 ^ n4572 ;
  assign n4578 = n4577 ^ n4027 ;
  assign n4579 = n4578 ^ n314 ;
  assign n4543 = n4027 ^ n3499 ;
  assign n4544 = n4543 ^ n4027 ;
  assign n4545 = n4027 ^ n3397 ;
  assign n4546 = n4545 ^ n4027 ;
  assign n4547 = n4544 & ~n4546 ;
  assign n4548 = n4547 ^ n4027 ;
  assign n4549 = ~n3551 & n4548 ;
  assign n4580 = n4579 ^ n4549 ;
  assign n5638 = n4580 ^ x78 ;
  assign n2744 = n2743 ^ n1649 ;
  assign n2711 = n1583 & n1610 ;
  assign n2712 = n2711 ^ n1596 ;
  assign n2713 = ~n1531 & n2712 ;
  assign n2714 = n2713 ^ n1663 ;
  assign n2715 = n2714 ^ n1606 ;
  assign n2719 = n2718 ^ n2715 ;
  assign n2720 = n2719 ^ n2713 ;
  assign n2721 = ~n1531 & n2720 ;
  assign n2722 = n2721 ^ n2714 ;
  assign n2745 = n2744 ^ n2722 ;
  assign n2746 = n2745 ^ n1639 ;
  assign n2747 = n2746 ^ x6 ;
  assign n2734 = n2733 ^ n2732 ;
  assign n2735 = n2734 ^ n2713 ;
  assign n2736 = n2735 ^ n2722 ;
  assign n2737 = n1584 & n2736 ;
  assign n2748 = n2747 ^ n2737 ;
  assign n3683 = n2748 ^ x114 ;
  assign n3684 = n1529 ^ x121 ;
  assign n3685 = ~n3683 & ~n3684 ;
  assign n3686 = n3685 ^ n3684 ;
  assign n2398 = n2397 ^ x56 ;
  assign n2374 = n2373 ^ n2369 ;
  assign n2375 = n2374 ^ n2372 ;
  assign n2377 = n2376 ^ n2375 ;
  assign n2378 = n2377 ^ n2369 ;
  assign n2379 = ~n2359 & n2378 ;
  assign n2380 = n2379 ^ n2374 ;
  assign n2381 = n2370 & ~n2380 ;
  assign n2382 = n2381 ^ n2369 ;
  assign n2383 = n2358 & n2382 ;
  assign n2399 = n2398 ^ n2383 ;
  assign n3613 = n2399 ^ x90 ;
  assign n3614 = n1272 ^ x88 ;
  assign n3615 = ~n3613 & n3614 ;
  assign n3616 = n3615 ^ n3613 ;
  assign n3638 = n1785 ^ n1772 ;
  assign n3639 = n3638 ^ n1830 ;
  assign n3640 = n3639 ^ n1842 ;
  assign n3641 = ~n1672 & n3640 ;
  assign n3642 = n3641 ^ n1842 ;
  assign n3643 = n1824 & n3642 ;
  assign n3633 = n1849 ^ n1773 ;
  assign n3634 = n3633 ^ n1862 ;
  assign n3635 = n1909 & ~n3634 ;
  assign n3626 = n3625 ^ n1842 ;
  assign n3629 = n3626 ^ n1859 ;
  assign n3624 = n1780 ^ n1773 ;
  assign n3627 = n3626 ^ n3624 ;
  assign n3628 = n1824 & ~n3627 ;
  assign n3630 = n3629 ^ n3628 ;
  assign n3631 = ~n1835 & ~n3630 ;
  assign n3619 = n1903 ^ n1859 ;
  assign n3620 = n3619 ^ n1829 ;
  assign n3621 = n3620 ^ n3473 ;
  assign n3622 = n3621 ^ n1911 ;
  assign n3623 = n3622 ^ x40 ;
  assign n3632 = n3631 ^ n3623 ;
  assign n3636 = n3635 ^ n3632 ;
  assign n3618 = n1776 & ~n1832 ;
  assign n3637 = n3636 ^ n3618 ;
  assign n3644 = n3643 ^ n3637 ;
  assign n3645 = n3644 ^ x99 ;
  assign n3669 = n2863 ^ n2565 ;
  assign n3652 = ~n2402 & n2507 ;
  assign n3653 = n3652 ^ n2509 ;
  assign n3654 = ~n2401 & ~n3653 ;
  assign n3655 = n3654 ^ n2486 ;
  assign n3656 = n3655 ^ n2503 ;
  assign n3657 = n3656 ^ n2473 ;
  assign n3658 = n3657 ^ n3654 ;
  assign n3659 = n2402 & ~n3658 ;
  assign n3660 = n3659 ^ n3655 ;
  assign n3670 = n3669 ^ n3660 ;
  assign n3671 = n3670 ^ n2543 ;
  assign n3672 = n3671 ^ n2527 ;
  assign n3173 = n2864 ^ n2510 ;
  assign n3176 = ~n2401 & ~n3173 ;
  assign n3177 = n3176 ^ n2510 ;
  assign n3178 = ~n2402 & ~n3177 ;
  assign n3673 = n3672 ^ n3178 ;
  assign n3674 = n3673 ^ n2893 ;
  assign n3675 = n3674 ^ x48 ;
  assign n3666 = n2402 & n2499 ;
  assign n3661 = n3660 ^ n3654 ;
  assign n3667 = n3666 ^ n3661 ;
  assign n3668 = ~n2528 & n3667 ;
  assign n3676 = n3675 ^ n3668 ;
  assign n3677 = n3676 ^ x73 ;
  assign n3678 = ~n3645 & ~n3677 ;
  assign n3679 = n3678 ^ n3645 ;
  assign n3680 = n3679 ^ n3677 ;
  assign n3713 = ~n3616 & ~n3680 ;
  assign n3696 = n3678 ^ n3677 ;
  assign n3697 = ~n3616 & ~n3696 ;
  assign n3714 = n3713 ^ n3697 ;
  assign n3702 = n3615 & ~n3679 ;
  assign n3688 = n3615 & n3678 ;
  assign n3703 = n3702 ^ n3688 ;
  assign n3704 = n3703 ^ n3615 ;
  assign n3701 = n3615 & ~n3680 ;
  assign n3705 = n3704 ^ n3701 ;
  assign n3617 = n3616 ^ n3614 ;
  assign n3692 = n3617 ^ n3613 ;
  assign n3694 = ~n3679 & n3692 ;
  assign n3681 = n3617 & ~n3680 ;
  assign n3646 = n3617 & ~n3645 ;
  assign n3647 = n3646 ^ n3617 ;
  assign n3682 = n3681 ^ n3647 ;
  assign n3700 = n3694 ^ n3682 ;
  assign n3706 = n3705 ^ n3700 ;
  assign n3698 = n3697 ^ n3694 ;
  assign n3699 = n3698 ^ n3696 ;
  assign n3707 = n3706 ^ n3699 ;
  assign n3708 = n3707 ^ n3692 ;
  assign n3693 = ~n3680 & n3692 ;
  assign n3695 = n3694 ^ n3693 ;
  assign n3709 = n3708 ^ n3695 ;
  assign n3690 = n3617 & ~n3679 ;
  assign n3691 = n3690 ^ n3646 ;
  assign n3710 = n3709 ^ n3691 ;
  assign n3689 = n3688 ^ n3678 ;
  assign n3711 = n3710 ^ n3689 ;
  assign n3712 = n3711 ^ n3616 ;
  assign n3715 = n3714 ^ n3712 ;
  assign n3716 = ~n3686 & n3715 ;
  assign n5658 = n3716 ^ n3698 ;
  assign n3754 = n3684 ^ n3683 ;
  assign n3755 = n3697 ^ n3693 ;
  assign n3722 = n3697 ^ n3684 ;
  assign n3756 = n3722 ^ n3697 ;
  assign n3757 = n3755 & ~n3756 ;
  assign n3758 = n3757 ^ n3697 ;
  assign n3759 = n3754 & n3758 ;
  assign n5659 = n5658 ^ n3759 ;
  assign n5660 = n5659 ^ n1404 ;
  assign n3719 = n3713 ^ n3705 ;
  assign n3750 = n3719 ^ n3710 ;
  assign n5653 = n3750 ^ n3700 ;
  assign n3744 = n3711 ^ n3701 ;
  assign n5654 = n5653 ^ n3744 ;
  assign n5655 = ~n3684 & n5654 ;
  assign n5656 = n5655 ^ n3698 ;
  assign n5657 = ~n3683 & ~n5656 ;
  assign n5661 = n5660 ^ n5657 ;
  assign n3729 = n3707 ^ n3681 ;
  assign n3730 = n3729 ^ n3709 ;
  assign n5646 = n3730 ^ n3688 ;
  assign n5647 = n5646 ^ n3691 ;
  assign n5648 = n5647 ^ n3730 ;
  assign n4048 = n3715 ^ n3701 ;
  assign n5649 = n5648 ^ n4048 ;
  assign n5650 = n3684 & ~n5649 ;
  assign n5651 = n5650 ^ n5646 ;
  assign n5652 = n3754 & ~n5651 ;
  assign n5662 = n5661 ^ n5652 ;
  assign n3734 = n3711 ^ n3702 ;
  assign n5639 = n3734 ^ n3690 ;
  assign n3727 = n3686 ^ n3683 ;
  assign n3728 = n3727 ^ n3684 ;
  assign n5640 = n5639 ^ n3728 ;
  assign n4063 = n3693 ^ n3682 ;
  assign n5641 = n5640 ^ n4063 ;
  assign n5642 = ~n3705 & ~n5641 ;
  assign n5643 = n5642 ^ n3728 ;
  assign n5644 = n3727 ^ n3705 ;
  assign n5645 = ~n5643 & ~n5644 ;
  assign n5663 = n5662 ^ n5645 ;
  assign n5664 = n5663 ^ x85 ;
  assign n5665 = ~n5638 & ~n5664 ;
  assign n5677 = n5665 ^ n5638 ;
  assign n5686 = n5677 ^ n5664 ;
  assign n5687 = ~n5635 & ~n5686 ;
  assign n5972 = ~n5609 & n5687 ;
  assign n5673 = n5638 ^ n5632 ;
  assign n5674 = n5638 ^ n5633 ;
  assign n5675 = n5673 & ~n5674 ;
  assign n5680 = n5675 ^ n5638 ;
  assign n5681 = n5673 ^ n5664 ;
  assign n5682 = ~n5680 & ~n5681 ;
  assign n5671 = n5634 & n5665 ;
  assign n5689 = n5682 ^ n5671 ;
  assign n5685 = ~n5635 & n5665 ;
  assign n5688 = n5687 ^ n5685 ;
  assign n5690 = n5689 ^ n5688 ;
  assign n5636 = n5635 ^ n5633 ;
  assign n5684 = ~n5636 & n5665 ;
  assign n5691 = n5690 ^ n5684 ;
  assign n5692 = n5691 ^ n5687 ;
  assign n5683 = n5682 ^ n5665 ;
  assign n5693 = n5692 ^ n5683 ;
  assign n5666 = n5665 ^ n5664 ;
  assign n5667 = ~n5633 & ~n5666 ;
  assign n5670 = n5632 & n5667 ;
  assign n5679 = n5670 ^ n5667 ;
  assign n5694 = n5693 ^ n5679 ;
  assign n5637 = n5636 ^ n5632 ;
  assign n5678 = ~n5637 & ~n5677 ;
  assign n5695 = n5694 ^ n5678 ;
  assign n5696 = n5695 ^ n5670 ;
  assign n5697 = n5696 ^ n5687 ;
  assign n5676 = n5675 ^ n5666 ;
  assign n5698 = n5697 ^ n5676 ;
  assign n5699 = n5698 ^ n5666 ;
  assign n5700 = n5699 ^ n5667 ;
  assign n5701 = n5700 ^ n5692 ;
  assign n5702 = n5701 ^ n5673 ;
  assign n5703 = n5702 ^ n5695 ;
  assign n5961 = n5703 ^ n5606 ;
  assign n5962 = n5961 ^ n5703 ;
  assign n5965 = n5690 & n5962 ;
  assign n5966 = n5965 ^ n5703 ;
  assign n5967 = n5605 & n5966 ;
  assign n5968 = n5967 ^ n5703 ;
  assign n5672 = n5671 ^ n5670 ;
  assign n5704 = n5703 ^ n5672 ;
  assign n5668 = n5667 ^ n5637 ;
  assign n5669 = n5668 ^ n5633 ;
  assign n5705 = n5704 ^ n5669 ;
  assign n5945 = n5705 ^ n5694 ;
  assign n5933 = n5678 ^ n5671 ;
  assign n5727 = n5700 ^ n5698 ;
  assign n5932 = n5727 ^ n5691 ;
  assign n5934 = n5933 ^ n5932 ;
  assign n5935 = n5934 ^ n5727 ;
  assign n5936 = n5727 ^ n5606 ;
  assign n5937 = n5936 ^ n5727 ;
  assign n5938 = n5935 & ~n5937 ;
  assign n5939 = n5938 ^ n5727 ;
  assign n5940 = ~n5605 & ~n5939 ;
  assign n5946 = n5945 ^ n5940 ;
  assign n5728 = n5700 ^ n5635 ;
  assign n5729 = n5728 ^ n5688 ;
  assign n5744 = n5729 ^ n5672 ;
  assign n5943 = n5744 ^ n5698 ;
  assign n5941 = n5633 ^ n5632 ;
  assign n5942 = n5664 & ~n5941 ;
  assign n5944 = n5943 ^ n5942 ;
  assign n5947 = n5946 ^ n5944 ;
  assign n5948 = n5947 ^ n5940 ;
  assign n5949 = ~n5606 & n5948 ;
  assign n5950 = n5949 ^ n5946 ;
  assign n5969 = n5968 ^ n5950 ;
  assign n5931 = n5606 ^ n5605 ;
  assign n5742 = n5695 ^ n5668 ;
  assign n5743 = n5742 ^ n5685 ;
  assign n5954 = n5743 ^ n5700 ;
  assign n5955 = n5954 ^ n5693 ;
  assign n5958 = n5606 & ~n5955 ;
  assign n5951 = n5950 ^ n5940 ;
  assign n5959 = n5958 ^ n5951 ;
  assign n5960 = ~n5931 & n5959 ;
  assign n5970 = n5969 ^ n5960 ;
  assign n5706 = n5705 ^ n5679 ;
  assign n5707 = ~n5609 & n5706 ;
  assign n5971 = n5970 ^ n5707 ;
  assign n5973 = n5972 ^ n5971 ;
  assign n5754 = n5698 ^ n5636 ;
  assign n5755 = n5754 ^ n5691 ;
  assign n5756 = n5755 ^ n5729 ;
  assign n5757 = n5756 ^ n5742 ;
  assign n5758 = n5742 ^ n5606 ;
  assign n5759 = n5758 ^ n5742 ;
  assign n5760 = n5757 & n5759 ;
  assign n5761 = n5760 ^ n5742 ;
  assign n5762 = ~n5605 & ~n5761 ;
  assign n5974 = n5973 ^ n5762 ;
  assign n5975 = n5974 ^ n1529 ;
  assign n5976 = n5975 ^ x89 ;
  assign n5068 = n5067 ^ x110 ;
  assign n4113 = n3032 ^ n2896 ;
  assign n4114 = n4113 ^ n3032 ;
  assign n4115 = ~n4110 & n4114 ;
  assign n4116 = n4115 ^ n3032 ;
  assign n4117 = ~n3030 & n4116 ;
  assign n3038 = n3037 ^ n3034 ;
  assign n3043 = n3042 ^ n3038 ;
  assign n3044 = n3042 ^ n2857 ;
  assign n3045 = n3044 ^ n3042 ;
  assign n3046 = ~n3043 & ~n3045 ;
  assign n3047 = n3046 ^ n3042 ;
  assign n3048 = ~n3030 & ~n3047 ;
  assign n4118 = n4117 ^ n3048 ;
  assign n4089 = n3007 & n4088 ;
  assign n4092 = n2996 ^ n2988 ;
  assign n4093 = n4092 ^ n4091 ;
  assign n4094 = n4090 & ~n4093 ;
  assign n4095 = ~n4089 & ~n4094 ;
  assign n4087 = n3021 ^ n3014 ;
  assign n4096 = n4095 ^ n4087 ;
  assign n4108 = n4107 ^ n4096 ;
  assign n4119 = n4118 ^ n4108 ;
  assign n4120 = n4119 ^ n921 ;
  assign n4085 = n3014 ^ n2996 ;
  assign n4086 = n4085 ^ n2989 ;
  assign n4097 = n4096 ^ n4086 ;
  assign n4083 = n3004 ^ n3002 ;
  assign n4084 = ~n2857 & n4083 ;
  assign n4098 = n4097 ^ n4084 ;
  assign n4099 = ~n3030 & n4098 ;
  assign n4121 = n4120 ^ n4099 ;
  assign n4920 = n4121 ^ x84 ;
  assign n3905 = n3857 ^ n3825 ;
  assign n3907 = n3906 ^ n3905 ;
  assign n3908 = n3823 & ~n3907 ;
  assign n3909 = n3908 ^ n3890 ;
  assign n3910 = n3909 ^ n3893 ;
  assign n3902 = n3895 ^ n3881 ;
  assign n3904 = n3903 ^ n3902 ;
  assign n3911 = n3910 ^ n3904 ;
  assign n3912 = ~n3800 & n3911 ;
  assign n3913 = n3912 ^ n3910 ;
  assign n4922 = n3913 ^ n3799 ;
  assign n3898 = n3897 ^ n3894 ;
  assign n3871 = n3857 ^ n3823 ;
  assign n3873 = n3872 ^ n3871 ;
  assign n3899 = n3898 ^ n3873 ;
  assign n3867 = n3866 ^ n3865 ;
  assign n3870 = n3869 ^ n3867 ;
  assign n3900 = n3899 ^ n3870 ;
  assign n3824 = n3823 ^ n3801 ;
  assign n3860 = n3825 & ~n3857 ;
  assign n3861 = n3860 ^ n3801 ;
  assign n3862 = n3824 & ~n3861 ;
  assign n3863 = n3862 ^ n3801 ;
  assign n3864 = n3800 & n3863 ;
  assign n3901 = n3900 ^ n3864 ;
  assign n3914 = n3913 ^ n3901 ;
  assign n3915 = ~n3799 & ~n3914 ;
  assign n3916 = n3915 ^ n3913 ;
  assign n4923 = n4922 ^ n3916 ;
  assign n4924 = n4923 ^ n3901 ;
  assign n4925 = n4924 ^ n4482 ;
  assign n4926 = n4925 ^ n1545 ;
  assign n4927 = n4926 ^ x124 ;
  assign n4986 = n4985 ^ x101 ;
  assign n4993 = n4927 & n4986 ;
  assign n4994 = n4993 ^ n4927 ;
  assign n4999 = n4994 ^ n4986 ;
  assign n3126 = n3125 ^ x110 ;
  assign n3162 = n3161 ^ x124 ;
  assign n3163 = ~n3126 & ~n3162 ;
  assign n3164 = n3163 ^ n3126 ;
  assign n3254 = n3253 ^ x76 ;
  assign n3284 = n3283 ^ x67 ;
  assign n3285 = n3254 & n3284 ;
  assign n3286 = n3285 ^ n3284 ;
  assign n3187 = ~n2401 & n2485 ;
  assign n3179 = n3178 ^ n2563 ;
  assign n3180 = n3179 ^ n2535 ;
  assign n3181 = n3180 ^ n2552 ;
  assign n3182 = n3181 ^ n2893 ;
  assign n3183 = n3182 ^ x52 ;
  assign n3170 = n2496 ^ n2471 ;
  assign n3171 = n3170 ^ n2483 ;
  assign n3172 = ~n2561 & ~n3171 ;
  assign n3184 = n3183 ^ n3172 ;
  assign n3167 = n2512 ^ n2484 ;
  assign n3168 = n3167 ^ n2473 ;
  assign n3169 = ~n2560 & ~n3168 ;
  assign n3185 = n3184 ^ n3169 ;
  assign n3165 = n2511 ^ n2469 ;
  assign n3166 = ~n2558 & n3165 ;
  assign n3186 = n3185 ^ n3166 ;
  assign n3188 = n3187 ^ n3186 ;
  assign n3189 = n3188 ^ x78 ;
  assign n3217 = n1201 ^ x44 ;
  assign n3198 = n1222 ^ n1214 ;
  assign n3199 = n3198 ^ n1233 ;
  assign n3200 = n1196 & n3199 ;
  assign n3201 = n3200 ^ n1222 ;
  assign n3210 = n3201 ^ n2668 ;
  assign n3203 = n3201 ^ n1261 ;
  assign n3202 = n3201 ^ n2918 ;
  assign n3204 = n3203 ^ n3202 ;
  assign n3207 = n1196 & ~n3204 ;
  assign n3208 = n3207 ^ n3203 ;
  assign n3209 = ~n1162 & n3208 ;
  assign n3211 = n3210 ^ n3209 ;
  assign n3197 = n1199 & n1259 ;
  assign n3212 = n3211 ^ n3197 ;
  assign n3196 = n1108 & ~n1202 ;
  assign n3213 = n3212 ^ n3196 ;
  assign n3190 = n1112 ^ n1109 ;
  assign n3193 = n1196 & ~n3190 ;
  assign n3194 = n3193 ^ n1112 ;
  assign n3195 = ~n1162 & ~n3194 ;
  assign n3214 = n3213 ^ n3195 ;
  assign n3215 = n3214 ^ n1239 ;
  assign n3216 = ~n2908 & ~n3215 ;
  assign n3218 = n3217 ^ n3216 ;
  assign n3219 = n3218 ^ x93 ;
  assign n3220 = ~n3189 & ~n3219 ;
  assign n3221 = n3220 ^ n3189 ;
  assign n3288 = n3221 ^ n3219 ;
  assign n3289 = n3288 ^ n3189 ;
  assign n3305 = n3286 & ~n3289 ;
  assign n3290 = n3285 & ~n3289 ;
  assign n3306 = n3305 ^ n3290 ;
  assign n3964 = n3306 ^ n3289 ;
  assign n3965 = ~n3164 & ~n3964 ;
  assign n3335 = n3163 ^ n3162 ;
  assign n3383 = n3335 ^ n3164 ;
  assign n3296 = n3286 ^ n3254 ;
  assign n3311 = ~n3288 & ~n3296 ;
  assign n3301 = n3219 ^ n3189 ;
  assign n3302 = n3284 ^ n3219 ;
  assign n3303 = n3301 & n3302 ;
  assign n3294 = n3285 ^ n3254 ;
  assign n3295 = ~n3221 & n3294 ;
  assign n3304 = n3303 ^ n3295 ;
  assign n3307 = n3306 ^ n3304 ;
  assign n3300 = n3220 & n3294 ;
  assign n3308 = n3307 ^ n3300 ;
  assign n3340 = n3311 ^ n3308 ;
  assign n3338 = n3219 & ~n3284 ;
  assign n3339 = n3338 ^ n3294 ;
  assign n3341 = n3340 ^ n3339 ;
  assign n3342 = n3341 ^ n3295 ;
  assign n3343 = n3342 ^ n3300 ;
  assign n3344 = n3343 ^ n3294 ;
  assign n3315 = n3220 & n3285 ;
  assign n3298 = n3254 ^ n3189 ;
  assign n3299 = ~n3284 & n3298 ;
  assign n3309 = n3308 ^ n3299 ;
  assign n3297 = n3296 ^ n3295 ;
  assign n3310 = n3309 ^ n3297 ;
  assign n3316 = n3315 ^ n3310 ;
  assign n3314 = n3300 ^ n3220 ;
  assign n3317 = n3316 ^ n3314 ;
  assign n3318 = n3317 ^ n3306 ;
  assign n3319 = n3318 ^ n3286 ;
  assign n3287 = ~n3221 & n3286 ;
  assign n3291 = n3290 ^ n3287 ;
  assign n3320 = n3319 ^ n3291 ;
  assign n3345 = n3344 ^ n3320 ;
  assign n3337 = n3311 ^ n3288 ;
  assign n3346 = n3345 ^ n3337 ;
  assign n3959 = n3346 ^ n3318 ;
  assign n3942 = n3335 & ~n3346 ;
  assign n3330 = n3315 ^ n3287 ;
  assign n3944 = n3942 ^ n3330 ;
  assign n3945 = ~n3164 & ~n3944 ;
  assign n3943 = n3306 & ~n3942 ;
  assign n3946 = n3945 ^ n3943 ;
  assign n3347 = n3346 ^ n3290 ;
  assign n3336 = n3315 ^ n3285 ;
  assign n3348 = n3347 ^ n3336 ;
  assign n3947 = n3946 ^ n3348 ;
  assign n3960 = n3959 ^ n3947 ;
  assign n3353 = n3341 ^ n3310 ;
  assign n3955 = n3353 ^ n3308 ;
  assign n3956 = n3955 ^ n3318 ;
  assign n3957 = n3956 ^ n3346 ;
  assign n3958 = n3126 & n3957 ;
  assign n3961 = n3960 ^ n3958 ;
  assign n3962 = ~n3383 & ~n3961 ;
  assign n3932 = n3335 ^ n3126 ;
  assign n3948 = n3348 ^ n3317 ;
  assign n3949 = ~n3932 & ~n3948 ;
  assign n3950 = n3949 ^ n3947 ;
  assign n3390 = ~n3317 & ~n3335 ;
  assign n3951 = n3950 ^ n3390 ;
  assign n3937 = n3344 ^ n3162 ;
  assign n3938 = n3937 ^ n3344 ;
  assign n3939 = ~n3345 & n3938 ;
  assign n3940 = n3939 ^ n3344 ;
  assign n3941 = n3383 & n3940 ;
  assign n3952 = n3951 ^ n3941 ;
  assign n3354 = n3353 ^ n3306 ;
  assign n3352 = n3310 ^ n3289 ;
  assign n3355 = n3354 ^ n3352 ;
  assign n3384 = n3355 ^ n3344 ;
  assign n3385 = n3355 ^ n3126 ;
  assign n3386 = n3385 ^ n3355 ;
  assign n3387 = ~n3384 & ~n3386 ;
  assign n3388 = n3387 ^ n3355 ;
  assign n3389 = n3383 & ~n3388 ;
  assign n3953 = n3952 ^ n3389 ;
  assign n3954 = n3953 ^ n1195 ;
  assign n3963 = n3962 ^ n3954 ;
  assign n3966 = n3965 ^ n3963 ;
  assign n3933 = n3346 ^ n3320 ;
  assign n3934 = ~n3932 & ~n3933 ;
  assign n3967 = n3966 ^ n3934 ;
  assign n3927 = n3308 ^ n3126 ;
  assign n3928 = n3927 ^ n3308 ;
  assign n3929 = n3309 & ~n3928 ;
  assign n3930 = n3929 ^ n3308 ;
  assign n3931 = ~n3162 & n3930 ;
  assign n3968 = n3967 ^ n3931 ;
  assign n4921 = n3968 ^ x75 ;
  assign n2571 = n2570 ^ x84 ;
  assign n2400 = n2399 ^ x70 ;
  assign n2706 = n2705 ^ x116 ;
  assign n2749 = n2748 ^ x94 ;
  assign n2750 = n2706 & ~n2749 ;
  assign n2591 = n760 ^ n722 ;
  assign n2589 = n219 & n393 ;
  assign n2590 = n628 & n2589 ;
  assign n2592 = n2591 ^ n2590 ;
  assign n2577 = n722 ^ n719 ;
  assign n2578 = n2577 ^ n736 ;
  assign n2579 = ~n219 & ~n2578 ;
  assign n2576 = n771 ^ n734 ;
  assign n2580 = n2579 ^ n2576 ;
  assign n2609 = n2592 ^ n2580 ;
  assign n2621 = n2620 ^ n2609 ;
  assign n2622 = n2621 ^ n2608 ;
  assign n2595 = n2594 ^ n2592 ;
  assign n2596 = n2595 ^ n742 ;
  assign n2597 = n2596 ^ n2592 ;
  assign n2600 = ~n315 & n2597 ;
  assign n2601 = n2600 ^ n2592 ;
  assign n2602 = n770 & n2601 ;
  assign n2623 = n2622 ^ n2602 ;
  assign n2586 = ~n219 & n746 ;
  assign n2581 = n2580 ^ n730 ;
  assign n2587 = n2586 ^ n2581 ;
  assign n2588 = ~n315 & n2587 ;
  assign n2624 = n2623 ^ n2588 ;
  assign n2626 = n2625 ^ n2624 ;
  assign n2627 = n2626 ^ n786 ;
  assign n2575 = ~n757 & n2574 ;
  assign n2628 = n2627 ^ n2575 ;
  assign n2629 = ~n790 & ~n2628 ;
  assign n2630 = n2629 ^ x14 ;
  assign n2631 = n2630 ^ x101 ;
  assign n2655 = n2009 & n2075 ;
  assign n2652 = n2644 ^ n2100 ;
  assign n2653 = ~n2076 & ~n2652 ;
  assign n2648 = n2075 & n2085 ;
  assign n2646 = n2645 ^ n2136 ;
  assign n2638 = n2637 ^ n2006 ;
  assign n2639 = n2638 ^ n2131 ;
  assign n2640 = n2639 ^ n2637 ;
  assign n2641 = n2046 & n2640 ;
  assign n2642 = n2641 ^ n2638 ;
  assign n2647 = n2646 ^ n2642 ;
  assign n2649 = n2648 ^ n2647 ;
  assign n2650 = n2114 & ~n2649 ;
  assign n2643 = n2642 ^ n2077 ;
  assign n2651 = n2650 ^ n2643 ;
  assign n2654 = n2653 ^ n2651 ;
  assign n2656 = n2655 ^ n2654 ;
  assign n2657 = ~n2634 & ~n2656 ;
  assign n2658 = ~n2162 & n2657 ;
  assign n2659 = ~n2012 & n2658 ;
  assign n2662 = n2659 ^ x22 ;
  assign n2660 = n2074 & n2659 ;
  assign n2661 = n2138 & n2660 ;
  assign n2663 = n2662 ^ n2661 ;
  assign n2664 = n2663 ^ x83 ;
  assign n2665 = ~n2631 & ~n2664 ;
  assign n2755 = n2665 ^ n2631 ;
  assign n2757 = n2755 ^ n2664 ;
  assign n2807 = n2750 & ~n2757 ;
  assign n2751 = n2750 ^ n2749 ;
  assign n2752 = n2665 & ~n2751 ;
  assign n4123 = n2807 ^ n2752 ;
  assign n4124 = n2400 & n4123 ;
  assign n4125 = n4124 ^ n2752 ;
  assign n2753 = n2750 ^ n2706 ;
  assign n2793 = n2753 & ~n2757 ;
  assign n4947 = n4125 ^ n2793 ;
  assign n2754 = n2753 ^ n2749 ;
  assign n2762 = n2665 ^ n2664 ;
  assign n2763 = n2754 & ~n2762 ;
  assign n2758 = ~n2751 & ~n2757 ;
  assign n2778 = n2763 ^ n2758 ;
  assign n2761 = ~n2751 & ~n2755 ;
  assign n2764 = n2763 ^ n2761 ;
  assign n2760 = n2664 & ~n2706 ;
  assign n2765 = n2764 ^ n2760 ;
  assign n2759 = n2758 ^ n2754 ;
  assign n2766 = n2765 ^ n2759 ;
  assign n2756 = n2754 & ~n2755 ;
  assign n2767 = n2766 ^ n2756 ;
  assign n2779 = n2778 ^ n2767 ;
  assign n2777 = n2706 ^ n2631 ;
  assign n2780 = n2779 ^ n2777 ;
  assign n2771 = n2749 ^ n2706 ;
  assign n2772 = n2771 ^ n2664 ;
  assign n2773 = n2631 & ~n2706 ;
  assign n2774 = n2773 ^ n2762 ;
  assign n2775 = n2774 ^ n2664 ;
  assign n2776 = n2772 & n2775 ;
  assign n2781 = n2780 ^ n2776 ;
  assign n2768 = n2767 ^ n2752 ;
  assign n2769 = n2768 ^ n2706 ;
  assign n2770 = n2769 ^ n2755 ;
  assign n2782 = n2781 ^ n2770 ;
  assign n4948 = n4947 ^ n2782 ;
  assign n2795 = n2782 ^ n2753 ;
  assign n2791 = n2779 ^ n2759 ;
  assign n2788 = n2750 & ~n2762 ;
  assign n2789 = n2788 ^ n2758 ;
  assign n2790 = n2789 ^ n2774 ;
  assign n2792 = n2791 ^ n2790 ;
  assign n2794 = n2793 ^ n2792 ;
  assign n2796 = n2795 ^ n2794 ;
  assign n2801 = n2796 ^ n2767 ;
  assign n2798 = n2772 ^ n2760 ;
  assign n2799 = ~n2631 & ~n2798 ;
  assign n2800 = n2799 ^ n2631 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2806 = n2802 ^ n2796 ;
  assign n2808 = n2807 ^ n2806 ;
  assign n4949 = n4948 ^ n2808 ;
  assign n4950 = n4949 ^ n4125 ;
  assign n4951 = n2400 & ~n4950 ;
  assign n4952 = n4951 ^ n4947 ;
  assign n4953 = n2571 & n4952 ;
  assign n4939 = n4125 ^ n2764 ;
  assign n4169 = n2758 ^ n2400 ;
  assign n4170 = n4169 ^ n2758 ;
  assign n4171 = n2789 & ~n4170 ;
  assign n4172 = n4171 ^ n2758 ;
  assign n4173 = ~n2571 & n4172 ;
  assign n4940 = n4939 ^ n4173 ;
  assign n2572 = ~n2400 & n2571 ;
  assign n4135 = n2572 & ~n2806 ;
  assign n4127 = n2793 ^ n2788 ;
  assign n4130 = n2793 ^ n2571 ;
  assign n4131 = n4130 ^ n2793 ;
  assign n4132 = n4127 & n4131 ;
  assign n4133 = n4132 ^ n2793 ;
  assign n4134 = ~n2400 & n4133 ;
  assign n4136 = n4135 ^ n4134 ;
  assign n4941 = n4940 ^ n4136 ;
  assign n2573 = n2572 ^ n2400 ;
  assign n4583 = ~n2573 & n2802 ;
  assign n4942 = n4941 ^ n4583 ;
  assign n2817 = n2573 ^ n2571 ;
  assign n2818 = n2817 ^ n2400 ;
  assign n2819 = n2791 ^ n2761 ;
  assign n2820 = n2819 ^ n2778 ;
  assign n2821 = n2820 ^ n2769 ;
  assign n2822 = n2821 ^ n2791 ;
  assign n2823 = n2818 & ~n2822 ;
  assign n4943 = n4942 ^ n2823 ;
  assign n4944 = n4943 ^ n1576 ;
  assign n4158 = n2571 ^ n2400 ;
  assign n4931 = n2779 ^ n2764 ;
  assign n4932 = n4931 ^ n2571 ;
  assign n4933 = n4932 ^ n4931 ;
  assign n4934 = n4931 ^ n2781 ;
  assign n4935 = n4934 ^ n4931 ;
  assign n4936 = ~n4933 & n4935 ;
  assign n4937 = n4936 ^ n4931 ;
  assign n4938 = n4158 & n4937 ;
  assign n4945 = n4944 ^ n4938 ;
  assign n4929 = n2792 ^ n2756 ;
  assign n4930 = ~n2573 & ~n4929 ;
  assign n4946 = n4945 ^ n4930 ;
  assign n4954 = n4953 ^ n4946 ;
  assign n4955 = n4954 ^ x86 ;
  assign n4995 = ~n4921 & n4955 ;
  assign n5006 = n4995 ^ n4955 ;
  assign n5008 = n5006 ^ n4921 ;
  assign n5009 = ~n4999 & n5008 ;
  assign n5007 = ~n4999 & n5006 ;
  assign n5010 = n5009 ^ n5007 ;
  assign n5000 = n4995 ^ n4921 ;
  assign n5001 = ~n4999 & ~n5000 ;
  assign n5005 = n5001 ^ n4999 ;
  assign n5011 = n5010 ^ n5005 ;
  assign n4997 = n4993 & n4995 ;
  assign n4996 = n4994 & n4995 ;
  assign n4998 = n4997 ^ n4996 ;
  assign n5014 = n5011 ^ n4998 ;
  assign n5015 = n5014 ^ n4995 ;
  assign n5013 = n4994 & ~n5000 ;
  assign n5016 = n5015 ^ n5013 ;
  assign n4991 = n4986 ^ n4927 ;
  assign n5017 = n5016 ^ n4991 ;
  assign n5004 = n4993 & ~n5000 ;
  assign n5012 = n5011 ^ n5004 ;
  assign n5018 = n5017 ^ n5012 ;
  assign n5002 = n5001 ^ n4998 ;
  assign n4992 = n4991 ^ n4921 ;
  assign n5003 = n5002 ^ n4992 ;
  assign n5019 = n5018 ^ n5003 ;
  assign n5109 = n5019 ^ n5016 ;
  assign n5110 = ~n4920 & n5109 ;
  assign n5111 = n5110 ^ n5016 ;
  assign n5112 = ~n5068 & ~n5111 ;
  assign n5069 = ~n4920 & n5068 ;
  assign n5070 = n5069 ^ n5068 ;
  assign n5071 = n5070 ^ n4920 ;
  assign n5103 = n5071 ^ n5068 ;
  assign n5104 = ~n5012 & ~n5103 ;
  assign n5029 = n4993 & n5006 ;
  assign n5024 = n5019 ^ n4996 ;
  assign n5025 = n5024 ^ n4994 ;
  assign n5022 = n5019 ^ n5013 ;
  assign n5021 = n4994 & n5006 ;
  assign n5023 = n5022 ^ n5021 ;
  assign n5026 = n5025 ^ n5023 ;
  assign n5079 = n5029 ^ n5026 ;
  assign n5096 = n5079 ^ n5009 ;
  assign n4987 = n4986 ^ n4955 ;
  assign n4988 = n4921 & ~n4987 ;
  assign n5097 = n5096 ^ n4988 ;
  assign n5100 = n5097 ^ n5009 ;
  assign n5027 = n5026 ^ n5015 ;
  assign n4928 = n4927 ^ n4921 ;
  assign n4989 = n4988 ^ n4986 ;
  assign n4990 = ~n4928 & n4989 ;
  assign n5020 = n5019 ^ n4990 ;
  assign n5028 = n5027 ^ n5020 ;
  assign n5095 = n5028 ^ n5008 ;
  assign n5098 = n5097 ^ n5095 ;
  assign n5099 = n4920 & n5098 ;
  assign n5101 = n5100 ^ n5099 ;
  assign n5102 = ~n5068 & n5101 ;
  assign n5105 = n5104 ^ n5102 ;
  assign n5082 = n4990 ^ n4955 ;
  assign n5080 = n5079 ^ n5001 ;
  assign n5030 = n5029 ^ n5007 ;
  assign n5072 = n5071 ^ n5030 ;
  assign n5073 = n5069 ^ n5024 ;
  assign n5074 = n5069 ^ n5030 ;
  assign n5075 = n5074 ^ n5069 ;
  assign n5076 = n5073 & ~n5075 ;
  assign n5077 = n5076 ^ n5069 ;
  assign n5078 = n5072 & n5077 ;
  assign n5081 = n5080 ^ n5078 ;
  assign n5083 = n5082 ^ n5081 ;
  assign n5084 = n5083 ^ n5078 ;
  assign n5085 = n5068 & ~n5084 ;
  assign n5086 = n5085 ^ n5081 ;
  assign n5106 = n5105 ^ n5086 ;
  assign n5107 = n5106 ^ n2748 ;
  assign n5087 = n5086 ^ n5078 ;
  assign n5033 = n5029 ^ n5011 ;
  assign n5031 = n5030 ^ n5026 ;
  assign n5032 = n5031 ^ n5028 ;
  assign n5034 = n5033 ^ n5032 ;
  assign n5035 = n5034 ^ n4992 ;
  assign n5088 = n5087 ^ n5035 ;
  assign n5089 = n5088 ^ n5087 ;
  assign n5092 = n5068 & ~n5089 ;
  assign n5093 = n5092 ^ n5087 ;
  assign n5094 = n4920 & ~n5093 ;
  assign n5108 = n5107 ^ n5094 ;
  assign n5113 = n5112 ^ n5108 ;
  assign n5977 = n5113 ^ x82 ;
  assign n5978 = n5976 & ~n5977 ;
  assign n5979 = n5978 ^ n5977 ;
  assign n4126 = ~n2571 & n4125 ;
  assign n2824 = n2806 ^ n2778 ;
  assign n2825 = n2778 ^ n2400 ;
  assign n2826 = n2825 ^ n2778 ;
  assign n2827 = ~n2824 & n2826 ;
  assign n2828 = n2827 ^ n2778 ;
  assign n2829 = ~n2571 & n2828 ;
  assign n2797 = n2796 ^ n2788 ;
  assign n2805 = n2797 ^ n2750 ;
  assign n2809 = n2808 ^ n2805 ;
  assign n4159 = n2809 ^ n2782 ;
  assign n4160 = ~n4158 & n4159 ;
  assign n4147 = n2752 ^ n2571 ;
  assign n4148 = n2758 ^ n2752 ;
  assign n4149 = n4148 ^ n2760 ;
  assign n4150 = n4149 ^ n4148 ;
  assign n4151 = n4148 ^ n2400 ;
  assign n4152 = n4151 ^ n4148 ;
  assign n4153 = n4150 & ~n4152 ;
  assign n4154 = n4153 ^ n4148 ;
  assign n4155 = n4147 & ~n4154 ;
  assign n4156 = n4155 ^ n2571 ;
  assign n4145 = n4127 ^ n2767 ;
  assign n4146 = n2817 & n4145 ;
  assign n4157 = n4156 ^ n4146 ;
  assign n4161 = n4160 ^ n4157 ;
  assign n4144 = ~n2573 & n2766 ;
  assign n4162 = n4161 ^ n4144 ;
  assign n4137 = n2792 ^ n2400 ;
  assign n4138 = n4137 ^ n2792 ;
  assign n4139 = n2792 ^ n2761 ;
  assign n4140 = n4139 ^ n2792 ;
  assign n4141 = n4138 & n4140 ;
  assign n4142 = n4141 ^ n2792 ;
  assign n4143 = n2571 & ~n4142 ;
  assign n4163 = n4162 ^ n4143 ;
  assign n4164 = ~n4136 & ~n4163 ;
  assign n4165 = ~n2829 & n4164 ;
  assign n4166 = ~n4126 & n4165 ;
  assign n4174 = n4166 & ~n4173 ;
  assign n4175 = ~n2823 & n4174 ;
  assign n4176 = n4175 ^ n958 ;
  assign n5395 = n4176 ^ x94 ;
  assign n3060 = n3036 ^ n3009 ;
  assign n3051 = n3042 ^ n3013 ;
  assign n3049 = n3037 ^ n3021 ;
  assign n3050 = n3049 ^ n3016 ;
  assign n3052 = n3051 ^ n3050 ;
  assign n3053 = ~n2857 & ~n3052 ;
  assign n3054 = n3053 ^ n3050 ;
  assign n3061 = n3060 ^ n3054 ;
  assign n3057 = n3014 ^ n2934 ;
  assign n3058 = n3057 ^ n3007 ;
  assign n3059 = ~n2857 & ~n3058 ;
  assign n3062 = n3061 ^ n3059 ;
  assign n3063 = n3030 & ~n3062 ;
  assign n2990 = n2989 ^ n2988 ;
  assign n2994 = n2993 ^ n2990 ;
  assign n3017 = n3016 ^ n2994 ;
  assign n3018 = ~n2896 & ~n3017 ;
  assign n3019 = n3018 ^ n2990 ;
  assign n3055 = n3054 ^ n3019 ;
  assign n3056 = n3055 ^ n3048 ;
  assign n3064 = n3063 ^ n3056 ;
  assign n3022 = n3021 ^ n3019 ;
  assign n3023 = n3022 ^ n2896 ;
  assign n3024 = n3023 ^ n3022 ;
  assign n3025 = n3022 ^ n2991 ;
  assign n3026 = n3025 ^ n3022 ;
  assign n3027 = n3024 & ~n3026 ;
  assign n3028 = n3027 ^ n3022 ;
  assign n3029 = ~n2857 & n3028 ;
  assign n3065 = n3064 ^ n3029 ;
  assign n3070 = n3069 ^ n3065 ;
  assign n3071 = n3070 ^ n1823 ;
  assign n5483 = n3071 ^ x108 ;
  assign n5533 = ~n5395 & n5483 ;
  assign n5539 = n5533 ^ n5483 ;
  assign n5534 = n5533 ^ n5395 ;
  assign n5980 = n5539 ^ n5534 ;
  assign n5418 = ~n801 & n2199 ;
  assign n5412 = n2206 ^ n2198 ;
  assign n4497 = n2203 ^ n2191 ;
  assign n4498 = n2203 ^ n801 ;
  assign n4499 = n4498 ^ n2203 ;
  assign n4500 = n4497 & ~n4499 ;
  assign n4501 = n4500 ^ n2203 ;
  assign n4502 = ~n1273 & n4501 ;
  assign n5413 = n5412 ^ n4502 ;
  assign n2247 = n2223 ^ n2210 ;
  assign n2248 = n2210 ^ n1273 ;
  assign n2249 = n2248 ^ n2210 ;
  assign n2250 = ~n2247 & n2249 ;
  assign n2251 = n2250 ^ n2210 ;
  assign n2252 = n801 & ~n2251 ;
  assign n5414 = n5413 ^ n2252 ;
  assign n2231 = n2210 ^ n2171 ;
  assign n2232 = n2171 ^ n801 ;
  assign n2233 = n2232 ^ n2171 ;
  assign n2234 = ~n2231 & n2233 ;
  assign n2235 = n2234 ^ n2171 ;
  assign n2236 = ~n1277 & n2235 ;
  assign n5415 = n5414 ^ n2236 ;
  assign n2219 = n1274 & n2196 ;
  assign n2220 = ~n2218 & n2219 ;
  assign n2221 = n2220 ^ n2218 ;
  assign n5416 = n5415 ^ n2221 ;
  assign n4518 = n1273 ^ n801 ;
  assign n5405 = n2178 ^ n2165 ;
  assign n5406 = n5405 ^ n2206 ;
  assign n5407 = n2206 ^ n1273 ;
  assign n5408 = n5407 ^ n2206 ;
  assign n5409 = n5406 & ~n5408 ;
  assign n5410 = n5409 ^ n2206 ;
  assign n5411 = ~n4518 & n5410 ;
  assign n5417 = n5416 ^ n5411 ;
  assign n5419 = n5418 ^ n5417 ;
  assign n5398 = n2198 ^ n2171 ;
  assign n5396 = n2199 ^ n2198 ;
  assign n5399 = n5398 ^ n5396 ;
  assign n5400 = n5396 ^ n801 ;
  assign n5401 = n5400 ^ n5396 ;
  assign n5402 = n5399 & n5401 ;
  assign n5403 = n5402 ^ n5396 ;
  assign n5404 = ~n1273 & n5403 ;
  assign n5420 = n5419 ^ n5404 ;
  assign n5421 = n5420 ^ n4488 ;
  assign n5422 = ~n4533 & ~n5421 ;
  assign n5423 = n5422 ^ n1768 ;
  assign n5424 = n5423 ^ x125 ;
  assign n4761 = n4358 ^ n4357 ;
  assign n5452 = n4387 & n4761 ;
  assign n5444 = n4364 ^ n4339 ;
  assign n5445 = n5444 ^ n4358 ;
  assign n5446 = n5445 ^ n4345 ;
  assign n5447 = n4265 & ~n5446 ;
  assign n5448 = n5447 ^ n4336 ;
  assign n5449 = n4371 & n5448 ;
  assign n4771 = n4376 ^ n4364 ;
  assign n4772 = n4364 ^ n4265 ;
  assign n4773 = n4772 ^ n4364 ;
  assign n4774 = n4771 & ~n4773 ;
  assign n4775 = n4774 ^ n4364 ;
  assign n4776 = ~n4371 & n4775 ;
  assign n5440 = n4776 ^ n4336 ;
  assign n5426 = n4351 ^ n4349 ;
  assign n5427 = n5426 ^ n4376 ;
  assign n5428 = n5427 ^ n4351 ;
  assign n5429 = n5428 ^ n4403 ;
  assign n5430 = n4265 & ~n5429 ;
  assign n5431 = n5430 ^ n5426 ;
  assign n5441 = n5440 ^ n5431 ;
  assign n5442 = n5441 ^ n1735 ;
  assign n5432 = n5431 ^ n4345 ;
  assign n5433 = n5432 ^ n4341 ;
  assign n5434 = n5433 ^ n5431 ;
  assign n5435 = n5431 ^ n4371 ;
  assign n5436 = n5435 ^ n5431 ;
  assign n5437 = n5434 & ~n5436 ;
  assign n5438 = n5437 ^ n5431 ;
  assign n5439 = ~n4387 & ~n5438 ;
  assign n5443 = n5442 ^ n5439 ;
  assign n5450 = n5449 ^ n5443 ;
  assign n4392 = n4391 ^ n4373 ;
  assign n5425 = ~n4388 & ~n4392 ;
  assign n5451 = n5450 ^ n5425 ;
  assign n5453 = n5452 ^ n5451 ;
  assign n5454 = n5453 ^ x77 ;
  assign n5455 = n5424 & n5454 ;
  assign n3687 = n3682 & ~n3686 ;
  assign n3717 = ~n3687 & ~n3716 ;
  assign n3751 = n3683 & ~n3750 ;
  assign n3745 = n3744 ^ n3690 ;
  assign n3746 = n3745 ^ n3693 ;
  assign n3747 = ~n3727 & ~n3746 ;
  assign n3737 = n3734 ^ n3694 ;
  assign n3733 = n3707 ^ n3646 ;
  assign n3735 = n3734 ^ n3733 ;
  assign n3736 = ~n3684 & n3735 ;
  assign n3738 = n3737 ^ n3736 ;
  assign n3740 = n3685 ^ n3683 ;
  assign n3739 = n3694 ^ n3685 ;
  assign n3741 = n3740 ^ n3739 ;
  assign n3742 = n3738 & ~n3741 ;
  assign n3743 = n3742 ^ n3740 ;
  assign n3748 = n3747 ^ n3743 ;
  assign n3731 = n3730 ^ n3682 ;
  assign n3732 = ~n3728 & n3731 ;
  assign n3749 = n3748 ^ n3732 ;
  assign n3752 = n3751 ^ n3749 ;
  assign n3718 = n3697 ^ n3685 ;
  assign n3720 = n3719 ^ n3688 ;
  assign n3721 = n3720 ^ n3684 ;
  assign n3724 = ~n3697 & n3721 ;
  assign n3725 = n3724 ^ n3684 ;
  assign n3726 = n3718 & ~n3725 ;
  assign n3753 = n3752 ^ n3726 ;
  assign n3760 = n3753 & ~n3759 ;
  assign n3761 = n3717 & n3760 ;
  assign n3762 = n3761 ^ n1701 ;
  assign n5456 = n3762 ^ x118 ;
  assign n3920 = n3919 ^ n3918 ;
  assign n3921 = n3875 & n3920 ;
  assign n3922 = n3921 ^ n3916 ;
  assign n3923 = n3922 ^ n1161 ;
  assign n5460 = n3923 ^ x91 ;
  assign n5461 = ~n5456 & n5460 ;
  assign n5487 = n5461 ^ n5460 ;
  assign n5501 = n5455 & n5487 ;
  assign n5491 = n5460 ^ n5424 ;
  assign n5492 = n5491 ^ n5454 ;
  assign n5493 = n5456 ^ n5454 ;
  assign n5471 = n5454 ^ n5424 ;
  assign n5494 = n5471 ^ n5454 ;
  assign n5495 = n5493 & n5494 ;
  assign n5496 = n5495 ^ n5454 ;
  assign n5497 = ~n5492 & ~n5496 ;
  assign n5462 = n5461 ^ n5456 ;
  assign n5476 = n5455 & ~n5462 ;
  assign n5498 = n5497 ^ n5476 ;
  assign n5459 = n5455 ^ n5424 ;
  assign n5464 = n5459 ^ n5454 ;
  assign n5465 = n5464 ^ n5424 ;
  assign n5468 = ~n5462 & n5465 ;
  assign n5466 = n5461 & n5465 ;
  assign n5475 = n5468 ^ n5466 ;
  assign n5477 = n5476 ^ n5475 ;
  assign n5478 = n5477 ^ n5462 ;
  assign n5463 = n5459 & ~n5462 ;
  assign n5467 = n5466 ^ n5463 ;
  assign n5479 = n5478 ^ n5467 ;
  assign n5472 = n5456 & n5471 ;
  assign n5473 = n5472 ^ n5471 ;
  assign n5469 = n5468 ^ n5467 ;
  assign n5474 = n5473 ^ n5469 ;
  assign n5480 = n5479 ^ n5474 ;
  assign n5499 = n5498 ^ n5480 ;
  assign n5488 = n5465 & n5487 ;
  assign n5489 = n5488 ^ n5465 ;
  assign n5490 = n5489 ^ n5475 ;
  assign n5500 = n5499 ^ n5490 ;
  assign n5502 = n5501 ^ n5500 ;
  assign n5457 = n5455 & ~n5456 ;
  assign n5485 = n5457 ^ n5455 ;
  assign n5484 = n5462 ^ n5460 ;
  assign n5486 = n5485 ^ n5484 ;
  assign n5503 = n5502 ^ n5486 ;
  assign n5504 = n5503 ^ n5501 ;
  assign n5505 = n5504 ^ n5488 ;
  assign n5506 = n5505 ^ n5499 ;
  assign n5507 = n5506 ^ n5472 ;
  assign n5508 = n5507 ^ n5502 ;
  assign n5519 = n5508 ^ n5488 ;
  assign n5518 = n5501 ^ n5487 ;
  assign n5520 = n5519 ^ n5518 ;
  assign n5985 = n5520 ^ n5508 ;
  assign n5981 = n5476 ^ n5457 ;
  assign n5982 = n5981 ^ n5480 ;
  assign n5983 = n5982 ^ n5485 ;
  assign n5984 = n5983 ^ n5981 ;
  assign n5986 = n5985 ^ n5984 ;
  assign n5987 = n5483 & ~n5986 ;
  assign n5988 = n5987 ^ n5982 ;
  assign n5989 = n5980 & ~n5988 ;
  assign n5990 = n5989 ^ n5981 ;
  assign n5992 = n5499 ^ n5485 ;
  assign n5458 = n5457 ^ n5456 ;
  assign n5470 = n5469 ^ n5458 ;
  assign n5481 = n5480 ^ n5470 ;
  assign n5993 = n5992 ^ n5481 ;
  assign n5994 = n5395 & ~n5993 ;
  assign n5995 = n5994 ^ n5506 ;
  assign n5996 = ~n5980 & n5995 ;
  assign n5991 = n5481 ^ n5466 ;
  assign n5997 = n5996 ^ n5991 ;
  assign n6008 = n5997 ^ n5458 ;
  assign n5998 = n5476 ^ n5395 ;
  assign n5999 = n5998 ^ n5476 ;
  assign n5547 = n5501 ^ n5485 ;
  assign n5548 = n5547 ^ n5488 ;
  assign n5509 = n5508 ^ n5490 ;
  assign n6000 = n5548 ^ n5509 ;
  assign n6001 = n6000 ^ n5476 ;
  assign n6002 = n5999 & ~n6001 ;
  assign n6003 = n6002 ^ n5476 ;
  assign n6004 = ~n5997 & ~n6003 ;
  assign n6009 = n6008 ^ n6004 ;
  assign n6005 = n5476 ^ n5462 ;
  assign n6006 = n6005 ^ n5474 ;
  assign n6007 = n5395 & ~n6006 ;
  assign n6010 = n6009 ^ n6007 ;
  assign n6011 = n5483 & n6010 ;
  assign n6012 = n6011 ^ n6004 ;
  assign n6013 = ~n5990 & n6012 ;
  assign n6015 = n5469 & n5539 ;
  assign n6016 = n6013 & n6015 ;
  assign n6014 = n6013 ^ n3644 ;
  assign n6017 = n6016 ^ n6014 ;
  assign n6018 = n6017 ^ x96 ;
  assign n2852 = n2817 & n2820 ;
  assign n2845 = n2766 ^ n2752 ;
  assign n2833 = n2793 ^ n2782 ;
  assign n2834 = n2833 ^ n2819 ;
  assign n2835 = n2400 & n2834 ;
  assign n2836 = n2835 ^ n2819 ;
  assign n2846 = n2845 ^ n2836 ;
  assign n2839 = n2572 & ~n2794 ;
  assign n2830 = n2572 & ~n2821 ;
  assign n2831 = n2830 ^ n2829 ;
  assign n2832 = n2831 ^ n2823 ;
  assign n2837 = n2836 ^ n2832 ;
  assign n2838 = n2837 ^ n2797 ;
  assign n2840 = n2839 ^ n2838 ;
  assign n2841 = n2840 ^ n2313 ;
  assign n2812 = n2807 ^ n2400 ;
  assign n2813 = n2812 ^ n2807 ;
  assign n2814 = n2809 & n2813 ;
  assign n2815 = n2814 ^ n2807 ;
  assign n2816 = n2571 & n2815 ;
  assign n2842 = n2841 ^ n2816 ;
  assign n2803 = n2802 ^ n2797 ;
  assign n2804 = ~n2400 & ~n2803 ;
  assign n2843 = n2842 ^ n2804 ;
  assign n2844 = n2843 ^ n2797 ;
  assign n2847 = n2846 ^ n2844 ;
  assign n2848 = n2847 ^ n2843 ;
  assign n2784 = n2760 ^ n2759 ;
  assign n2785 = n2784 ^ n2756 ;
  assign n2786 = n2785 ^ n2752 ;
  assign n2787 = ~n2400 & n2786 ;
  assign n2849 = n2848 ^ n2787 ;
  assign n2850 = n2571 & ~n2849 ;
  assign n2851 = n2850 ^ n2844 ;
  assign n2853 = n2852 ^ n2851 ;
  assign n2783 = ~n2573 & n2782 ;
  assign n2854 = n2853 ^ n2783 ;
  assign n2855 = n2854 ^ x115 ;
  assign n2276 = n2212 ^ n2203 ;
  assign n2277 = n1276 & ~n2276 ;
  assign n2260 = n2184 ^ n1274 ;
  assign n2255 = n2203 ^ n2183 ;
  assign n2256 = n2255 ^ n2254 ;
  assign n2258 = n1274 & n2256 ;
  assign n2259 = n2258 ^ n1277 ;
  assign n2261 = n2260 ^ n2259 ;
  assign n2262 = n2261 ^ n2260 ;
  assign n2264 = n2209 ^ n2169 ;
  assign n2265 = n1274 & n2264 ;
  assign n2271 = n2262 & ~n2265 ;
  assign n2263 = n2262 ^ n1274 ;
  assign n2266 = n2265 ^ n2263 ;
  assign n2267 = n2266 ^ n2252 ;
  assign n2272 = n2267 ^ n2184 ;
  assign n2273 = n2272 ^ n2252 ;
  assign n2274 = n2271 & n2273 ;
  assign n2268 = n2267 ^ n2246 ;
  assign n2238 = n2173 & n2237 ;
  assign n2240 = n2239 ^ n2238 ;
  assign n2269 = n2268 ^ n2240 ;
  assign n2270 = n2269 ^ n2236 ;
  assign n2275 = n2274 ^ n2270 ;
  assign n2278 = n2277 ^ n2275 ;
  assign n2224 = n2223 ^ n2186 ;
  assign n2222 = n2182 ^ n2174 ;
  assign n2225 = n2224 ^ n2222 ;
  assign n2226 = n2222 ^ n801 ;
  assign n2227 = n2226 ^ n2222 ;
  assign n2228 = n2225 & ~n2227 ;
  assign n2229 = n2228 ^ n2222 ;
  assign n2230 = ~n1277 & n2229 ;
  assign n2279 = n2278 ^ n2230 ;
  assign n2280 = ~n2221 & ~n2279 ;
  assign n2281 = n2280 ^ n2072 ;
  assign n2282 = n2281 ^ x89 ;
  assign n2856 = n2855 ^ n2282 ;
  assign n3072 = n3071 ^ x106 ;
  assign n3391 = n3390 ^ n2348 ;
  assign n3392 = n3391 ^ n3389 ;
  assign n3349 = n3348 ^ n3320 ;
  assign n3350 = ~n3335 & ~n3349 ;
  assign n3331 = n3330 ^ n3306 ;
  assign n3293 = n3162 ^ n3126 ;
  assign n3312 = n3311 ^ n3310 ;
  assign n3313 = n3312 ^ n3295 ;
  assign n3321 = n3320 ^ n3313 ;
  assign n3322 = n3321 ^ n3320 ;
  assign n3323 = n3316 ^ n3305 ;
  assign n3326 = n3322 & n3323 ;
  assign n3327 = n3326 ^ n3320 ;
  assign n3328 = ~n3293 & ~n3327 ;
  assign n3332 = ~n3162 & n3328 ;
  assign n3333 = n3331 & n3332 ;
  assign n3329 = n3328 ^ n3293 ;
  assign n3334 = n3333 ^ n3329 ;
  assign n3351 = n3350 ^ n3334 ;
  assign n3356 = n3355 ^ n3308 ;
  assign n3357 = n3356 ^ n3162 ;
  assign n3358 = ~n3293 & n3357 ;
  assign n3359 = n3358 ^ n3162 ;
  assign n3362 = n3356 ^ n3343 ;
  assign n3363 = n3359 & ~n3362 ;
  assign n3360 = n3346 ^ n3343 ;
  assign n3364 = n3363 ^ n3360 ;
  assign n3365 = n3364 ^ n3342 ;
  assign n3366 = n3365 ^ n3307 ;
  assign n3367 = n3366 ^ n3364 ;
  assign n3370 = n3162 & n3367 ;
  assign n3371 = n3370 ^ n3364 ;
  assign n3372 = ~n3293 & n3371 ;
  assign n3373 = n3372 ^ n3364 ;
  assign n3374 = n3351 & ~n3373 ;
  assign n3292 = ~n3164 & n3291 ;
  assign n3375 = n3374 ^ n3292 ;
  assign n3376 = n3317 ^ n3311 ;
  assign n3377 = n3311 ^ n3126 ;
  assign n3378 = n3377 ^ n3311 ;
  assign n3379 = ~n3376 & ~n3378 ;
  assign n3380 = n3379 ^ n3311 ;
  assign n3381 = n3162 & n3380 ;
  assign n3382 = n3375 & ~n3381 ;
  assign n3393 = n3392 ^ n3382 ;
  assign n3394 = n3393 ^ x88 ;
  assign n3395 = n3072 & ~n3394 ;
  assign n3396 = n2856 & n3395 ;
  assign n3582 = n3524 ^ n2002 ;
  assign n3573 = ~n3397 & ~n3572 ;
  assign n3574 = n3573 ^ n3571 ;
  assign n3583 = n3582 ^ n3574 ;
  assign n3575 = n3574 ^ n3561 ;
  assign n3576 = n3575 ^ n3574 ;
  assign n3579 = n3397 & n3576 ;
  assign n3580 = n3579 ^ n3574 ;
  assign n3581 = n3551 & ~n3580 ;
  assign n3584 = n3583 ^ n3581 ;
  assign n3526 = n3525 ^ n3524 ;
  assign n3554 = n3526 & n3551 ;
  assign n3555 = n3554 ^ n3524 ;
  assign n3556 = ~n3397 & n3555 ;
  assign n3585 = n3584 ^ n3556 ;
  assign n3586 = n3585 ^ x82 ;
  assign n3775 = n3395 ^ n3394 ;
  assign n3776 = n2282 & ~n3775 ;
  assign n3782 = n3776 ^ n3396 ;
  assign n3587 = n3072 ^ n2855 ;
  assign n3599 = n3394 ^ n2282 ;
  assign n3767 = n2855 & ~n3599 ;
  assign n3768 = n3767 ^ n2282 ;
  assign n3769 = ~n3587 & ~n3768 ;
  assign n3785 = n3782 ^ n3769 ;
  assign n3786 = n3785 ^ n2856 ;
  assign n3588 = n3587 ^ n3072 ;
  assign n3589 = n3072 ^ n2282 ;
  assign n3590 = n3589 ^ n3072 ;
  assign n3591 = n3588 & ~n3590 ;
  assign n3592 = n3591 ^ n3072 ;
  assign n3593 = n3394 & n3592 ;
  assign n3783 = n3782 ^ n3593 ;
  assign n3607 = n3394 ^ n2856 ;
  assign n3600 = n3599 ^ n3072 ;
  assign n3601 = n3600 ^ n3394 ;
  assign n3603 = n3395 ^ n3072 ;
  assign n3604 = n3603 ^ n2855 ;
  assign n3602 = n3072 & ~n3587 ;
  assign n3605 = n3604 ^ n3602 ;
  assign n3606 = ~n3601 & n3605 ;
  assign n3608 = n3607 ^ n3606 ;
  assign n3784 = n3783 ^ n3608 ;
  assign n3787 = n3786 ^ n3784 ;
  assign n3763 = n3762 ^ x64 ;
  assign n3770 = n3603 ^ n3394 ;
  assign n3594 = ~n2282 & ~n3394 ;
  assign n3595 = n3594 ^ n3072 ;
  assign n3771 = n3770 ^ n3595 ;
  assign n3772 = n3771 ^ n3072 ;
  assign n3773 = n2855 & n3772 ;
  assign n3774 = n3773 ^ n3600 ;
  assign n3777 = n3776 ^ n3774 ;
  assign n3778 = n3777 ^ n3769 ;
  assign n3779 = n3763 & ~n3778 ;
  assign n3780 = n3779 ^ n3774 ;
  assign n3788 = n3787 ^ n3780 ;
  assign n3596 = n3394 ^ n2855 ;
  assign n3597 = n3595 & ~n3596 ;
  assign n3598 = n3597 ^ n2856 ;
  assign n3609 = n3608 ^ n3598 ;
  assign n3610 = n3609 ^ n3602 ;
  assign n3611 = n3610 ^ n3593 ;
  assign n3612 = n3611 ^ n3607 ;
  assign n3781 = n3780 ^ n3612 ;
  assign n3789 = n3788 ^ n3781 ;
  assign n3790 = n3788 ^ n3763 ;
  assign n3791 = n3790 ^ n3788 ;
  assign n3792 = ~n3789 & ~n3791 ;
  assign n3793 = n3792 ^ n3788 ;
  assign n3794 = n3586 & ~n3793 ;
  assign n3795 = n3794 ^ n3780 ;
  assign n3796 = ~n3396 & n3795 ;
  assign n3797 = n3796 ^ n2399 ;
  assign n6019 = n3797 ^ x123 ;
  assign n6020 = ~n6018 & n6019 ;
  assign n3924 = n3923 ^ x70 ;
  assign n3969 = n3968 ^ x83 ;
  assign n3970 = n3924 & n3969 ;
  assign n4246 = n3970 ^ n3924 ;
  assign n4247 = n4246 ^ n3969 ;
  assign n4020 = n3983 ^ n3517 ;
  assign n3993 = n3992 ^ n3551 ;
  assign n4015 = n4014 ^ n3982 ;
  assign n4016 = n4015 ^ n3511 ;
  assign n4017 = ~n3993 & ~n4016 ;
  assign n4021 = n4020 ^ n4017 ;
  assign n4011 = ~n3993 & n4010 ;
  assign n4009 = n3517 ^ n3515 ;
  assign n4012 = n4011 ^ n4009 ;
  assign n4008 = n3519 ^ n3511 ;
  assign n4013 = n4012 ^ n4008 ;
  assign n4018 = n4017 ^ n4013 ;
  assign n4019 = n3992 & n4018 ;
  assign n4022 = n4021 ^ n4019 ;
  assign n4002 = n3551 ^ n3517 ;
  assign n3994 = n3993 ^ n3397 ;
  assign n4003 = n4002 ^ n3994 ;
  assign n3995 = n3994 ^ n3551 ;
  assign n4004 = n3566 ^ n3551 ;
  assign n4005 = n3995 & ~n4004 ;
  assign n4006 = n4005 ^ n3551 ;
  assign n4007 = n4003 & ~n4006 ;
  assign n4023 = n4022 ^ n4007 ;
  assign n4001 = n3522 & n3994 ;
  assign n4024 = n4023 ^ n4001 ;
  assign n3996 = n3995 ^ n3993 ;
  assign n3999 = n3998 ^ n3977 ;
  assign n4000 = n3996 & n3999 ;
  assign n4025 = n4024 ^ n4000 ;
  assign n3985 = n3983 ^ n3514 ;
  assign n3984 = n3983 ^ n3520 ;
  assign n3986 = n3985 ^ n3984 ;
  assign n3987 = n3985 ^ n3551 ;
  assign n3988 = n3987 ^ n3985 ;
  assign n3989 = n3986 & ~n3988 ;
  assign n3990 = n3989 ^ n3985 ;
  assign n3991 = ~n3397 & n3990 ;
  assign n4026 = n4025 ^ n3991 ;
  assign n4029 = n4028 ^ n4014 ;
  assign n4030 = n4014 ^ n3397 ;
  assign n4031 = n4030 ^ n4014 ;
  assign n4032 = ~n4029 & ~n4031 ;
  assign n4033 = n4032 ^ n4014 ;
  assign n4034 = ~n3996 & ~n4033 ;
  assign n4035 = ~n4026 & ~n4034 ;
  assign n4036 = n4035 ^ n995 ;
  assign n4037 = n4036 ^ x126 ;
  assign n4057 = n3713 ^ n3702 ;
  assign n4058 = n4057 ^ n3715 ;
  assign n4059 = n4058 ^ n3744 ;
  assign n4060 = n3684 & ~n4059 ;
  assign n4056 = n3713 ^ n3703 ;
  assign n4061 = n4060 ^ n4056 ;
  assign n4071 = n4061 ^ n3716 ;
  assign n4062 = n4061 ^ n3710 ;
  assign n4064 = n4063 ^ n4062 ;
  assign n4065 = n4064 ^ n4061 ;
  assign n4068 = n3684 & ~n4065 ;
  assign n4069 = n4068 ^ n4061 ;
  assign n4070 = ~n3683 & n4069 ;
  assign n4072 = n4071 ^ n4070 ;
  assign n4049 = n4048 ^ n3714 ;
  assign n4047 = n3707 ^ n3690 ;
  assign n4050 = n4049 ^ n4047 ;
  assign n4051 = n4047 ^ n3683 ;
  assign n4052 = n4051 ^ n4047 ;
  assign n4053 = ~n4050 & ~n4052 ;
  assign n4054 = n4053 ^ n4047 ;
  assign n4055 = ~n3684 & ~n4054 ;
  assign n4073 = n4072 ^ n4055 ;
  assign n4045 = n3719 ^ n3702 ;
  assign n4046 = ~n3728 & n4045 ;
  assign n4074 = n4073 ^ n4046 ;
  assign n4038 = n3706 ^ n3691 ;
  assign n4039 = n4038 ^ n3709 ;
  assign n4040 = n4039 ^ n3691 ;
  assign n4041 = n4040 ^ n3729 ;
  assign n4042 = ~n3684 & n4041 ;
  assign n4043 = n4042 ^ n4038 ;
  assign n4044 = ~n3754 & n4043 ;
  assign n4075 = n4074 ^ n4044 ;
  assign n4076 = n4075 ^ n3687 ;
  assign n4077 = n4076 ^ n3759 ;
  assign n4078 = n4077 ^ n1098 ;
  assign n4079 = n4078 ^ x76 ;
  assign n4080 = ~n4037 & ~n4079 ;
  assign n4081 = n4080 ^ n4079 ;
  assign n4122 = n4121 ^ x109 ;
  assign n4177 = n4176 ^ x116 ;
  assign n4178 = ~n4122 & n4177 ;
  assign n4184 = n4178 ^ n4122 ;
  assign n4204 = ~n4081 & ~n4184 ;
  assign n4179 = n4178 ^ n4177 ;
  assign n4180 = n4179 ^ n4122 ;
  assign n4194 = n4080 & n4180 ;
  assign n4205 = n4204 ^ n4194 ;
  assign n4082 = n4081 ^ n4037 ;
  assign n4188 = ~n4082 & n4178 ;
  assign n4187 = ~n4082 & n4179 ;
  assign n4189 = n4188 ^ n4187 ;
  assign n4182 = n4080 & ~n4177 ;
  assign n4185 = n4184 ^ n4182 ;
  assign n4186 = n4185 ^ n4082 ;
  assign n4190 = n4189 ^ n4186 ;
  assign n4191 = n4190 ^ n4184 ;
  assign n4181 = ~n4082 & n4180 ;
  assign n4183 = n4182 ^ n4181 ;
  assign n4192 = n4191 ^ n4183 ;
  assign n4206 = n4205 ^ n4192 ;
  assign n4209 = n4206 ^ n4185 ;
  assign n4196 = n4080 ^ n4037 ;
  assign n4229 = n4209 ^ n4196 ;
  assign n4215 = n4122 ^ n4037 ;
  assign n4216 = n4215 ^ n4079 ;
  assign n4217 = n4216 ^ n4190 ;
  assign n4211 = n4182 ^ n4080 ;
  assign n4202 = n4080 & n4178 ;
  assign n4212 = n4211 ^ n4202 ;
  assign n4210 = ~n4081 & n4178 ;
  assign n4213 = n4212 ^ n4210 ;
  assign n4214 = n4213 ^ n4187 ;
  assign n4218 = n4217 ^ n4214 ;
  assign n4197 = n4179 & ~n4196 ;
  assign n4219 = n4218 ^ n4197 ;
  assign n4230 = n4229 ^ n4219 ;
  assign n4228 = n4194 ^ n4182 ;
  assign n4231 = n4230 ^ n4228 ;
  assign n6022 = n4231 ^ n4181 ;
  assign n4233 = n4185 ^ n4177 ;
  assign n6026 = n6022 ^ n4233 ;
  assign n4259 = n4218 ^ n4212 ;
  assign n6027 = n6026 ^ n4259 ;
  assign n6028 = n6027 ^ n4188 ;
  assign n3971 = n3970 ^ n3969 ;
  assign n6024 = n4230 ^ n4205 ;
  assign n6025 = n3971 & ~n6024 ;
  assign n6029 = n6028 ^ n6025 ;
  assign n6030 = n6029 ^ n4183 ;
  assign n6031 = n6030 ^ n4183 ;
  assign n6032 = n4247 & ~n6031 ;
  assign n6033 = n6032 ^ n4183 ;
  assign n6034 = ~n3970 & n6033 ;
  assign n6035 = n6034 ^ n4183 ;
  assign n6023 = ~n4247 & ~n6022 ;
  assign n6036 = n6035 ^ n6023 ;
  assign n6056 = n4190 & n4246 ;
  assign n4200 = n3969 ^ n3924 ;
  assign n6044 = n4202 ^ n4197 ;
  assign n6045 = n6044 ^ n6026 ;
  assign n6046 = n6045 ^ n4187 ;
  assign n4251 = n4210 ^ n4187 ;
  assign n6047 = n6046 ^ n4251 ;
  assign n6048 = n6047 ^ n3924 ;
  assign n6049 = n6048 ^ n6047 ;
  assign n4201 = ~n4081 & n4179 ;
  assign n4203 = n4202 ^ n4201 ;
  assign n6050 = ~n4203 & ~n4251 ;
  assign n6051 = n6050 ^ n6047 ;
  assign n6052 = n6049 & n6051 ;
  assign n6053 = n6052 ^ n6047 ;
  assign n6054 = ~n4200 & ~n6053 ;
  assign n6055 = n6054 ^ n4192 ;
  assign n6057 = n6056 ^ n6055 ;
  assign n6039 = n4192 ^ n3969 ;
  assign n6040 = n6039 ^ n4192 ;
  assign n6041 = n4189 & n6040 ;
  assign n6042 = n6041 ^ n4192 ;
  assign n6043 = n4200 & ~n6042 ;
  assign n6058 = n6057 ^ n6043 ;
  assign n6059 = ~n6036 & n6058 ;
  assign n6060 = n6059 ^ n1272 ;
  assign n6061 = n6060 ^ x121 ;
  assign n6062 = n6020 & n6061 ;
  assign n4412 = n4265 & n4402 ;
  assign n4365 = n4364 ^ n4363 ;
  assign n4366 = n4365 ^ n4359 ;
  assign n4355 = n4354 ^ n4336 ;
  assign n4356 = n4355 ^ n4351 ;
  assign n4367 = n4366 ^ n4356 ;
  assign n4368 = ~n4265 & ~n4367 ;
  assign n4369 = n4368 ^ n4356 ;
  assign n4410 = n4369 ^ n4354 ;
  assign n4405 = n4404 ^ n4346 ;
  assign n4398 = ~n4360 & n4391 ;
  assign n4399 = n4397 & n4398 ;
  assign n4389 = n4358 ^ n4348 ;
  assign n4393 = n4392 ^ n4389 ;
  assign n4394 = n4388 & n4393 ;
  assign n4400 = n4399 ^ n4394 ;
  assign n4408 = n4405 ^ n4400 ;
  assign n4377 = n4376 ^ n4348 ;
  assign n4383 = ~n4355 & n4382 ;
  assign n4384 = ~n4377 & n4383 ;
  assign n4378 = n4377 ^ n4365 ;
  assign n4379 = n4378 ^ n4376 ;
  assign n4380 = ~n4372 & ~n4379 ;
  assign n4385 = n4384 ^ n4380 ;
  assign n4409 = n4408 ^ n4385 ;
  assign n4411 = n4410 ^ n4409 ;
  assign n4413 = n4412 ^ n4411 ;
  assign n4414 = n4387 & ~n4413 ;
  assign n4370 = n4369 ^ n716 ;
  assign n4386 = n4385 ^ n4370 ;
  assign n4415 = n4414 ^ n4386 ;
  assign n5126 = n4415 ^ x121 ;
  assign n4737 = n3734 ^ n3705 ;
  assign n4738 = ~n3686 & ~n4737 ;
  assign n4729 = n3730 ^ ~n3707 ;
  assign n4730 = n4729 ^ n3695 ;
  assign n4731 = n3695 ^ n3684 ;
  assign n4732 = n4731 ^ n3695 ;
  assign n4733 = n4730 & ~n4732 ;
  assign n4734 = n4733 ^ n3695 ;
  assign n4735 = n3683 & n4734 ;
  assign n4716 = n3714 ^ n3702 ;
  assign n4717 = n4716 ^ n3727 ;
  assign n4718 = n4717 ^ n3745 ;
  assign n4719 = ~n3691 & ~n4718 ;
  assign n4720 = n4719 ^ n3727 ;
  assign n4725 = ~n3707 ^ n3691 ;
  assign n4724 = n3728 ^ ~n3707 ;
  assign n4726 = n4725 ^ n4724 ;
  assign n4727 = n4720 & ~n4726 ;
  assign n4728 = n4727 ^ n4725 ;
  assign n4736 = n4735 ^ n4728 ;
  assign n4739 = n4738 ^ n4736 ;
  assign n4706 = n3713 ^ n3694 ;
  assign n4707 = n4706 ^ n3750 ;
  assign n4704 = n3614 ^ n3613 ;
  assign n4705 = n4704 ^ n3677 ;
  assign n4708 = n4707 ^ n4705 ;
  assign n4709 = n4708 ^ n3694 ;
  assign n4703 = n3720 ^ n3697 ;
  assign n4710 = n4709 ^ n4703 ;
  assign n4711 = n4709 ^ n3684 ;
  assign n4712 = n4711 ^ n4709 ;
  assign n4713 = ~n4710 & n4712 ;
  assign n4714 = n4713 ^ n4709 ;
  assign n4715 = ~n3754 & ~n4714 ;
  assign n4740 = n4739 ^ n4715 ;
  assign n4741 = n4740 ^ n3687 ;
  assign n4742 = n4741 ^ n3716 ;
  assign n4743 = n4742 ^ n1955 ;
  assign n5127 = n4743 ^ x65 ;
  assign n5128 = n5126 & ~n5127 ;
  assign n5204 = n5128 ^ n5127 ;
  assign n4837 = n3389 ^ n2045 ;
  assign n4417 = n3347 ^ n3344 ;
  assign n4418 = ~n3162 & n4417 ;
  assign n4419 = n4418 ^ n3344 ;
  assign n4421 = n4419 ^ n3291 ;
  assign n4420 = n4419 ^ n3933 ;
  assign n4422 = n4421 ^ n4420 ;
  assign n4425 = ~n3162 & ~n4422 ;
  assign n4426 = n4425 ^ n4421 ;
  assign n4427 = ~n3126 & n4426 ;
  assign n4428 = n4427 ^ n4419 ;
  assign n4830 = n3949 ^ n3295 ;
  assign n4818 = n3354 ^ n3339 ;
  assign n4819 = n4818 ^ n3323 ;
  assign n4820 = n4819 ^ n3313 ;
  assign n4821 = ~n3126 & ~n4820 ;
  assign n4822 = n4821 ^ n3354 ;
  assign n4831 = n4830 ^ n4822 ;
  assign n4832 = n4831 ^ n3941 ;
  assign n4833 = n4832 ^ n3381 ;
  assign n4823 = n4822 ^ n3316 ;
  assign n4824 = n4823 ^ n4822 ;
  assign n4825 = n4822 ^ n3162 ;
  assign n4826 = n4825 ^ n4822 ;
  assign n4827 = ~n4824 & n4826 ;
  assign n4828 = n4827 ^ n4822 ;
  assign n4829 = n3293 & ~n4828 ;
  assign n4834 = n4833 ^ n4829 ;
  assign n4811 = n3335 ^ n3295 ;
  assign n4431 = n3300 ^ n3287 ;
  assign n4432 = n4431 ^ n3311 ;
  assign n4812 = n4432 ^ n3164 ;
  assign n4815 = ~n3295 & n4812 ;
  assign n4816 = n4815 ^ n3164 ;
  assign n4817 = ~n4811 & n4816 ;
  assign n4835 = n4834 ^ n4817 ;
  assign n4836 = ~n4428 & n4835 ;
  assign n4838 = n4837 ^ n4836 ;
  assign n5129 = n4838 ^ x107 ;
  assign n5159 = n4034 ^ n2456 ;
  assign n5148 = n4011 ^ n3995 ;
  assign n5149 = n4028 ^ n4012 ;
  assign n5150 = n5148 & n5149 ;
  assign n5145 = n3516 ^ n3508 ;
  assign n5146 = n5145 ^ n3519 ;
  assign n5147 = n3996 & n5146 ;
  assign n5151 = n5150 ^ n5147 ;
  assign n5138 = n4561 ^ n3982 ;
  assign n5137 = n3981 ^ n3517 ;
  assign n5139 = n5138 ^ n5137 ;
  assign n5140 = n5138 ^ n3551 ;
  assign n5141 = n5140 ^ n5138 ;
  assign n5142 = ~n5139 & ~n5141 ;
  assign n5143 = n5142 ^ n5138 ;
  assign n5144 = ~n3397 & ~n5143 ;
  assign n5152 = n5151 ^ n5144 ;
  assign n5153 = n3521 ^ n3511 ;
  assign n5154 = n3996 ^ n3521 ;
  assign n5155 = n5154 ^ n3521 ;
  assign n5156 = n5153 & ~n5155 ;
  assign n5157 = n5156 ^ n3521 ;
  assign n5158 = ~n5152 & ~n5157 ;
  assign n5160 = n5159 ^ n5158 ;
  assign n5130 = n3998 ^ n3551 ;
  assign n5131 = n5130 ^ n3998 ;
  assign n5134 = n4562 & ~n5131 ;
  assign n5135 = n5134 ^ n3998 ;
  assign n5136 = n3397 & n5135 ;
  assign n5161 = n5160 ^ n5136 ;
  assign n5162 = n5161 ^ x97 ;
  assign n4602 = ~n2573 & ~n2801 ;
  assign n2810 = n2809 ^ n2807 ;
  assign n4599 = n2571 & n2810 ;
  assign n4591 = n2769 ^ n2766 ;
  assign n4592 = n4591 ^ n2834 ;
  assign n4593 = n4592 ^ n2807 ;
  assign n4589 = n2807 ^ n2772 ;
  assign n4590 = n4589 ^ n2799 ;
  assign n4594 = n4593 ^ n4590 ;
  assign n4595 = ~n2571 & n4594 ;
  assign n4596 = n4595 ^ n4593 ;
  assign n4597 = n2400 & ~n4596 ;
  assign n4584 = n2839 ^ n2807 ;
  assign n4585 = n4584 ^ n4134 ;
  assign n4586 = n4585 ^ n2831 ;
  assign n4587 = n4586 ^ n4583 ;
  assign n4588 = n4587 ^ n218 ;
  assign n4598 = n4597 ^ n4588 ;
  assign n4600 = n4599 ^ n4598 ;
  assign n4582 = n2572 & n2768 ;
  assign n4601 = n4600 ^ n4582 ;
  assign n4603 = n4602 ^ n4601 ;
  assign n5163 = n4603 ^ x80 ;
  assign n5175 = n3011 ^ n2989 ;
  assign n5176 = n5175 ^ n3035 ;
  assign n5177 = ~n2857 & n5176 ;
  assign n5174 = n5173 ^ n3040 ;
  assign n5178 = n5177 ^ n5174 ;
  assign n5192 = n5178 ^ n4118 ;
  assign n5193 = n5192 ^ n5191 ;
  assign n5170 = n3035 ^ n2999 ;
  assign n5171 = n5170 ^ n3020 ;
  assign n5179 = n5178 ^ n5171 ;
  assign n5180 = n5179 ^ n5178 ;
  assign n5168 = n3012 ^ n2988 ;
  assign n5169 = n5168 ^ n5167 ;
  assign n5181 = n5180 ^ n5169 ;
  assign n5182 = ~n2857 & ~n5181 ;
  assign n5183 = n5182 ^ n5179 ;
  assign n5184 = ~n3030 & ~n5183 ;
  assign n5194 = n5193 ^ n5184 ;
  assign n5195 = n5194 ^ n3069 ;
  assign n5196 = n5195 ^ n2429 ;
  assign n5197 = n5196 ^ x90 ;
  assign n5198 = n5163 & ~n5197 ;
  assign n5199 = n5162 & n5198 ;
  assign n5259 = n5129 & n5199 ;
  assign n5282 = n5259 ^ n5199 ;
  assign n5288 = ~n5204 & n5282 ;
  assign n5240 = n5199 ^ n5198 ;
  assign n5208 = n5198 ^ n5163 ;
  assign n5210 = ~n5129 & ~n5162 ;
  assign n5211 = n5208 & n5210 ;
  assign n5238 = n5211 ^ n5210 ;
  assign n5218 = ~n5163 & n5210 ;
  assign n5239 = n5238 ^ n5218 ;
  assign n5241 = n5240 ^ n5239 ;
  assign n6103 = n5241 ^ n5211 ;
  assign n6104 = ~n5204 & n6103 ;
  assign n5205 = n5204 ^ n5126 ;
  assign n5206 = n5205 ^ n5127 ;
  assign n5164 = n5162 & ~n5163 ;
  assign n5214 = ~n5129 & n5164 ;
  assign n5226 = n5197 & n5214 ;
  assign n5227 = n5226 ^ n5214 ;
  assign n5222 = n5164 ^ n5163 ;
  assign n5223 = n5222 ^ n5218 ;
  assign n5224 = ~n5197 & ~n5223 ;
  assign n5225 = n5224 ^ n5223 ;
  assign n5228 = n5227 ^ n5225 ;
  assign n5220 = ~n5197 & n5218 ;
  assign n5221 = n5220 ^ n5218 ;
  assign n5229 = n5228 ^ n5221 ;
  assign n5216 = n5197 ^ n5129 ;
  assign n5217 = ~n5163 & ~n5216 ;
  assign n5219 = n5218 ^ n5217 ;
  assign n5230 = n5229 ^ n5219 ;
  assign n5215 = n5214 ^ n5164 ;
  assign n5231 = n5230 ^ n5215 ;
  assign n5278 = n5231 ^ n5221 ;
  assign n5279 = n5206 & ~n5278 ;
  assign n6105 = n6104 ^ n5279 ;
  assign n5165 = n5164 ^ n5162 ;
  assign n5200 = n5199 ^ n5165 ;
  assign n6067 = n5128 & n5200 ;
  assign n5251 = n5226 ^ n5225 ;
  assign n6068 = n5251 ^ n5211 ;
  assign n6069 = n5127 & ~n6068 ;
  assign n6070 = n6069 ^ n5211 ;
  assign n5209 = n5208 ^ n5200 ;
  assign n5212 = n5211 ^ n5209 ;
  assign n6090 = n6070 ^ n5212 ;
  assign n6087 = n5227 ^ n5223 ;
  assign n5201 = ~n5129 & n5200 ;
  assign n5213 = n5212 ^ n5201 ;
  assign n6088 = n6087 ^ n5213 ;
  assign n6089 = ~n5127 & ~n6088 ;
  assign n6091 = n6090 ^ n6089 ;
  assign n6092 = ~n5126 & n6091 ;
  assign n5207 = n5206 ^ n5204 ;
  assign n6079 = n5259 ^ n5239 ;
  assign n5263 = n5227 ^ n5224 ;
  assign n6076 = n5263 ^ n5259 ;
  assign n6077 = ~n5128 & ~n6076 ;
  assign n6072 = n5259 ^ n5221 ;
  assign n6073 = n6072 ^ n5239 ;
  assign n6078 = n6077 ^ n6073 ;
  assign n6080 = n6079 ^ n6078 ;
  assign n6081 = n5217 ^ n5215 ;
  assign n6082 = ~n5205 & ~n6081 ;
  assign n6083 = ~n6080 & n6082 ;
  assign n6084 = n6083 ^ n6078 ;
  assign n6085 = n5207 & ~n6084 ;
  assign n6071 = n6070 ^ n5259 ;
  assign n6086 = n6085 ^ n6071 ;
  assign n6093 = n6092 ^ n6086 ;
  assign n5202 = n5201 ^ n5200 ;
  assign n5283 = n5282 ^ n5202 ;
  assign n5284 = n5206 & n5283 ;
  assign n6094 = n6093 ^ n5284 ;
  assign n6095 = ~n6067 & ~n6094 ;
  assign n6096 = n5241 ^ n5200 ;
  assign n6097 = n5200 ^ n5126 ;
  assign n6098 = n6097 ^ n5200 ;
  assign n6099 = n6096 & n6098 ;
  assign n6100 = n6099 ^ n5200 ;
  assign n6101 = n5127 & n6100 ;
  assign n6102 = n6095 & ~n6101 ;
  assign n6106 = n6105 ^ n6102 ;
  assign n6107 = ~n5288 & n6106 ;
  assign n6108 = n6107 ^ n3676 ;
  assign n6109 = n6108 ^ x106 ;
  assign n6120 = n6062 & n6109 ;
  assign n6142 = n6120 ^ n6062 ;
  assign n6110 = ~n6061 & n6109 ;
  assign n6123 = ~n6019 & n6110 ;
  assign n6021 = n6020 ^ n6019 ;
  assign n6116 = n6021 & n6110 ;
  assign n6117 = n6116 ^ n6110 ;
  assign n6132 = n6123 ^ n6117 ;
  assign n6143 = n6142 ^ n6132 ;
  assign n6139 = n6109 ^ n6061 ;
  assign n6140 = n6139 ^ n6019 ;
  assign n6141 = ~n6018 & ~n6140 ;
  assign n6144 = n6143 ^ n6141 ;
  assign n6136 = n6062 ^ n6020 ;
  assign n6137 = n6136 ^ n6132 ;
  assign n6111 = n6110 ^ n6061 ;
  assign n6112 = n6018 & ~n6111 ;
  assign n6113 = n6112 ^ n6111 ;
  assign n6138 = n6137 ^ n6113 ;
  assign n6145 = n6144 ^ n6138 ;
  assign n6064 = ~n6019 & n6061 ;
  assign n6128 = n6018 & n6064 ;
  assign n6135 = n6128 ^ n6064 ;
  assign n6146 = n6145 ^ n6135 ;
  assign n6194 = ~n5979 & ~n6146 ;
  assign n6192 = n5979 ^ n5976 ;
  assign n6193 = n6143 & n6192 ;
  assign n6195 = n6194 ^ n6193 ;
  assign n6196 = n6195 ^ n3762 ;
  assign n6063 = n6062 ^ n6061 ;
  assign n6065 = n6064 ^ n6063 ;
  assign n6126 = n6065 & ~n6109 ;
  assign n6154 = n6126 ^ n6065 ;
  assign n6186 = n6154 ^ n6138 ;
  assign n6187 = n6154 ^ n5976 ;
  assign n6188 = n6187 ^ n6154 ;
  assign n6189 = ~n6186 & ~n6188 ;
  assign n6190 = n6189 ^ n6154 ;
  assign n6191 = n5977 & n6190 ;
  assign n6197 = n6196 ^ n6191 ;
  assign n6066 = n6065 ^ n6021 ;
  assign n6114 = n6113 ^ n6066 ;
  assign n6115 = n6114 ^ n6061 ;
  assign n6118 = n6117 ^ n6115 ;
  assign n6119 = n6118 ^ n6112 ;
  assign n6121 = n6120 ^ n6119 ;
  assign n6122 = ~n5979 & n6121 ;
  assign n6129 = ~n6109 & n6128 ;
  assign n6149 = n6129 ^ n6119 ;
  assign n6150 = n6149 ^ n6142 ;
  assign n6124 = n6018 & n6123 ;
  assign n6125 = n6124 ^ n6123 ;
  assign n6147 = n6146 ^ n6125 ;
  assign n6148 = n6147 ^ n6138 ;
  assign n6151 = n6150 ^ n6148 ;
  assign n6130 = n6129 ^ n6020 ;
  assign n6131 = n6130 ^ n6126 ;
  assign n6133 = n6132 ^ n6131 ;
  assign n6134 = ~n5977 & n6133 ;
  assign n6152 = n6151 ^ n6134 ;
  assign n6181 = n6152 ^ n6116 ;
  assign n6172 = n6145 ^ n6112 ;
  assign n6173 = n6172 ^ n6126 ;
  assign n6176 = n6126 ^ n5977 ;
  assign n6177 = n6176 ^ n6126 ;
  assign n6178 = ~n6173 & ~n6177 ;
  assign n6179 = n6178 ^ n6126 ;
  assign n6180 = ~n5976 & n6179 ;
  assign n6182 = n6181 ^ n6180 ;
  assign n6164 = n5977 ^ n5976 ;
  assign n6165 = n6116 ^ n5977 ;
  assign n6166 = n6165 ^ n6116 ;
  assign n6169 = n6124 & ~n6166 ;
  assign n6170 = n6169 ^ n6116 ;
  assign n6171 = n6164 & n6170 ;
  assign n6183 = n6182 ^ n6171 ;
  assign n6156 = n6129 ^ n6128 ;
  assign n6157 = n6156 ^ n6118 ;
  assign n6155 = n6154 ^ n6137 ;
  assign n6158 = n6157 ^ n6155 ;
  assign n6159 = n6158 ^ n6152 ;
  assign n6127 = n6126 ^ n6125 ;
  assign n6153 = n6152 ^ n6127 ;
  assign n6160 = n6159 ^ n6153 ;
  assign n6161 = ~n5977 & n6160 ;
  assign n6162 = n6161 ^ n6159 ;
  assign n6163 = ~n5976 & n6162 ;
  assign n6184 = n6183 ^ n6163 ;
  assign n6185 = ~n6122 & ~n6184 ;
  assign n6198 = n6197 ^ n6185 ;
  assign n6911 = n6198 ^ x97 ;
  assign n5289 = n5288 ^ n2570 ;
  assign n5203 = n5128 & n5202 ;
  assign n5272 = n5223 ^ n5214 ;
  assign n5273 = n5205 & n5272 ;
  assign n5262 = n5228 ^ n5217 ;
  assign n5264 = n5263 ^ n5262 ;
  assign n5265 = n5264 ^ n5262 ;
  assign n5266 = n5262 ^ n5127 ;
  assign n5267 = n5266 ^ n5262 ;
  assign n5268 = ~n5265 & ~n5267 ;
  assign n5269 = n5268 ^ n5262 ;
  assign n5270 = n5126 & n5269 ;
  assign n5271 = n5270 ^ n5127 ;
  assign n5274 = n5273 ^ n5271 ;
  assign n5260 = n5259 ^ n5211 ;
  assign n5261 = n5207 & n5260 ;
  assign n5275 = n5274 ^ n5261 ;
  assign n5249 = n5239 ^ n5212 ;
  assign n5250 = n5249 ^ n5201 ;
  assign n5252 = n5251 ^ n5250 ;
  assign n5253 = n5252 ^ n5201 ;
  assign n5254 = n5201 ^ n5127 ;
  assign n5255 = n5254 ^ n5201 ;
  assign n5256 = ~n5253 & ~n5255 ;
  assign n5257 = n5256 ^ n5201 ;
  assign n5258 = ~n5126 & n5257 ;
  assign n5276 = n5275 ^ n5258 ;
  assign n5277 = n5276 ^ n5241 ;
  assign n5280 = n5279 ^ n5277 ;
  assign n5242 = n5241 ^ n5127 ;
  assign n5243 = n5242 ^ n5241 ;
  assign n5244 = n5241 ^ n5221 ;
  assign n5245 = n5244 ^ n5241 ;
  assign n5246 = ~n5243 & n5245 ;
  assign n5247 = n5246 ^ n5241 ;
  assign n5248 = n5126 & n5247 ;
  assign n5281 = n5280 ^ n5248 ;
  assign n5285 = n5284 ^ n5281 ;
  assign n5232 = n5231 ^ n5213 ;
  assign n5233 = n5231 ^ n5126 ;
  assign n5234 = n5233 ^ n5231 ;
  assign n5235 = ~n5232 & n5234 ;
  assign n5236 = n5235 ^ n5231 ;
  assign n5237 = ~n5207 & ~n5236 ;
  assign n5286 = n5285 ^ n5237 ;
  assign n5287 = ~n5203 & ~n5286 ;
  assign n5290 = n5289 ^ n5287 ;
  assign n6914 = n5290 ^ x85 ;
  assign n5708 = n5607 & n5695 ;
  assign n6930 = n5968 ^ n5708 ;
  assign n6919 = n5701 ^ n5680 ;
  assign n6377 = n5664 ^ n5633 ;
  assign n6920 = n6919 ^ n6377 ;
  assign n5730 = n5729 ^ n5727 ;
  assign n6918 = n5755 ^ n5730 ;
  assign n6921 = n6920 ^ n6918 ;
  assign n6922 = n5605 & n6921 ;
  assign n6923 = n6922 ^ n6918 ;
  assign n6931 = n6930 ^ n6923 ;
  assign n6924 = n6923 ^ n5943 ;
  assign n6916 = n5955 ^ n5684 ;
  assign n6915 = n5755 ^ n5678 ;
  assign n6917 = n6916 ^ n6915 ;
  assign n6925 = n6924 ^ n6917 ;
  assign n6926 = n6925 ^ n6923 ;
  assign n6927 = ~n5605 & ~n6926 ;
  assign n6928 = n6927 ^ n6924 ;
  assign n6929 = n5606 & n6928 ;
  assign n6932 = n6931 ^ n6929 ;
  assign n6933 = n6932 ^ n5707 ;
  assign n6934 = ~n5972 & ~n6933 ;
  assign n6935 = n6934 ^ n3426 ;
  assign n6936 = n6935 ^ x70 ;
  assign n6937 = n6914 & ~n6936 ;
  assign n6938 = n6937 ^ n6936 ;
  assign n5386 = n3598 ^ n3587 ;
  assign n5384 = n3602 ^ n3394 ;
  assign n5385 = n2282 & n5384 ;
  assign n5387 = n5386 ^ n5385 ;
  assign n5388 = n3586 & n5387 ;
  assign n5389 = n5388 ^ n3598 ;
  assign n5381 = n3586 & ~n3784 ;
  assign n5382 = n5381 ^ n3608 ;
  assign n5390 = n5389 ^ n5382 ;
  assign n5391 = n3763 & ~n5390 ;
  assign n6940 = n5391 ^ n5389 ;
  assign n6941 = n6940 ^ n3438 ;
  assign n6942 = n6941 ^ x108 ;
  assign n5549 = n5548 ^ n5504 ;
  assign n5544 = ~n5481 & ~n5539 ;
  assign n5545 = n5544 ^ n5480 ;
  assign n5546 = ~n5476 & ~n5545 ;
  assign n5550 = n5549 ^ n5546 ;
  assign n5551 = n5533 & ~n5550 ;
  assign n5532 = n5456 ^ n5424 ;
  assign n5535 = n5534 ^ n5532 ;
  assign n5536 = n5535 ^ n5497 ;
  assign n5537 = ~n5474 & n5536 ;
  assign n5538 = n5537 ^ n5534 ;
  assign n5540 = n5539 ^ n5474 ;
  assign n5541 = ~n5538 & n5540 ;
  assign n5542 = n5541 ^ n3487 ;
  assign n5512 = n5490 ^ n5395 ;
  assign n5513 = n5512 ^ n5490 ;
  assign n5514 = ~n5509 & n5513 ;
  assign n5515 = n5514 ^ n5490 ;
  assign n5516 = ~n5483 & n5515 ;
  assign n5517 = n5516 ^ n5504 ;
  assign n5521 = n5520 ^ n5517 ;
  assign n5529 = n5521 ^ n5477 ;
  assign n5526 = n5502 & n5508 ;
  assign n5527 = n5526 ^ n5521 ;
  assign n5528 = n5395 & ~n5527 ;
  assign n5530 = n5529 ^ n5528 ;
  assign n5531 = ~n5483 & ~n5530 ;
  assign n5543 = n5542 ^ n5531 ;
  assign n5552 = n5551 ^ n5543 ;
  assign n5482 = n5395 & n5481 ;
  assign n5553 = n5552 ^ n5482 ;
  assign n6943 = n5553 ^ x126 ;
  assign n6944 = ~n6942 & n6943 ;
  assign n6961 = ~n6938 & n6944 ;
  assign n4852 = n2281 ^ x81 ;
  assign n4702 = n3585 ^ x96 ;
  assign n4744 = n4743 ^ x123 ;
  assign n4745 = n4702 & ~n4744 ;
  assign n4781 = n4403 ^ n4349 ;
  assign n4782 = n4372 & ~n4781 ;
  assign n4762 = n4404 ^ n4354 ;
  assign n4763 = n4762 ^ n4333 ;
  assign n4764 = n4763 ^ n4761 ;
  assign n4765 = n4764 ^ n4760 ;
  assign n4766 = ~n4265 & n4765 ;
  assign n4767 = n4766 ^ n4763 ;
  assign n4777 = n4767 ^ n1981 ;
  assign n4778 = n4777 ^ n4776 ;
  assign n4768 = n4767 ^ n4349 ;
  assign n4757 = n4376 ^ n4333 ;
  assign n4758 = n4757 ^ n4388 ;
  assign n4759 = ~n4383 & ~n4758 ;
  assign n4769 = n4768 ^ n4759 ;
  assign n4770 = n4371 & n4769 ;
  assign n4779 = n4778 ^ n4770 ;
  assign n4756 = n4374 & n4387 ;
  assign n4780 = n4779 ^ n4756 ;
  assign n4783 = n4782 ^ n4780 ;
  assign n4755 = n4343 & ~n4382 ;
  assign n4784 = n4783 ^ n4755 ;
  assign n4748 = n4362 ^ n4358 ;
  assign n4749 = n4748 ^ n4391 ;
  assign n4750 = n4391 ^ n4265 ;
  assign n4751 = n4750 ^ n4391 ;
  assign n4752 = ~n4749 & ~n4751 ;
  assign n4753 = n4752 ^ n4391 ;
  assign n4754 = n4387 & ~n4753 ;
  assign n4785 = n4784 ^ n4754 ;
  assign n4786 = n4785 ^ x113 ;
  assign n4787 = n3799 & ~n3897 ;
  assign n4803 = n4787 ^ n1927 ;
  assign n4801 = n3921 ^ n3799 ;
  assign n4791 = n4469 ^ n3892 ;
  assign n4792 = ~n3799 & ~n4791 ;
  assign n4793 = n4792 ^ n3892 ;
  assign n4802 = n4801 ^ n4793 ;
  assign n4804 = n4803 ^ n4802 ;
  assign n4790 = n3800 ^ n3799 ;
  assign n4794 = n4793 ^ n3898 ;
  assign n4795 = n4794 ^ n4793 ;
  assign n4796 = n4793 ^ n3800 ;
  assign n4797 = n4796 ^ n4793 ;
  assign n4798 = ~n4795 & ~n4797 ;
  assign n4799 = n4798 ^ n4793 ;
  assign n4800 = ~n4790 & n4799 ;
  assign n4805 = n4804 ^ n4800 ;
  assign n4788 = n3800 & n4787 ;
  assign n4789 = n4470 & n4788 ;
  assign n4806 = n4805 ^ n4789 ;
  assign n4807 = n4806 ^ x114 ;
  assign n4808 = n4786 & n4807 ;
  assign n4845 = n4808 ^ n4786 ;
  assign n4860 = n4845 ^ n4807 ;
  assign n4886 = n4745 & ~n4860 ;
  assign n4746 = n4745 ^ n4744 ;
  assign n4809 = n4808 ^ n4807 ;
  assign n4885 = ~n4746 & n4809 ;
  assign n4887 = n4886 ^ n4885 ;
  assign n4747 = n4746 ^ n4702 ;
  assign n4840 = n4747 & n4808 ;
  assign n4910 = n4887 ^ n4840 ;
  assign n4839 = n4838 ^ x120 ;
  assign n4911 = n4840 ^ n4839 ;
  assign n4912 = n4911 ^ n4840 ;
  assign n4913 = n4910 & n4912 ;
  assign n4914 = n4913 ^ n4840 ;
  assign n4915 = ~n4852 & n4914 ;
  assign n4841 = n4747 ^ n4744 ;
  assign n4846 = n4841 & n4845 ;
  assign n4844 = n4809 & n4841 ;
  assign n4847 = n4846 ^ n4844 ;
  assign n4842 = n4808 & n4841 ;
  assign n4843 = n4842 ^ n4841 ;
  assign n4848 = n4847 ^ n4843 ;
  assign n4879 = n4839 & ~n4852 ;
  assign n4880 = n4879 ^ n4839 ;
  assign n4882 = n4880 ^ n4852 ;
  assign n4883 = n4882 ^ n4839 ;
  assign n5792 = n4848 & ~n4883 ;
  assign n4873 = n4852 ^ n4839 ;
  assign n4810 = n4747 & n4809 ;
  assign n5785 = n4846 ^ n4810 ;
  assign n5786 = n5785 ^ n4842 ;
  assign n4876 = n4842 ^ n4840 ;
  assign n4856 = n4745 & n4808 ;
  assign n4875 = n4856 ^ n4808 ;
  assign n4877 = n4876 ^ n4875 ;
  assign n4861 = n4747 & ~n4860 ;
  assign n4881 = n4877 ^ n4861 ;
  assign n4862 = n4861 ^ n4810 ;
  assign n4859 = n4840 ^ n4747 ;
  assign n4863 = n4862 ^ n4859 ;
  assign n5784 = n4881 ^ n4863 ;
  assign n5787 = n5786 ^ n5784 ;
  assign n5788 = ~n4852 & n5787 ;
  assign n4864 = n4863 ^ n4846 ;
  assign n4854 = n4745 & ~n4786 ;
  assign n4855 = n4854 ^ n4745 ;
  assign n4857 = n4856 ^ n4855 ;
  assign n4858 = n4857 ^ n4845 ;
  assign n4865 = n4864 ^ n4858 ;
  assign n4866 = n4865 ^ n4856 ;
  assign n5775 = n4887 ^ n4866 ;
  assign n5781 = n5775 ^ n4744 ;
  assign n5789 = n5788 ^ n5781 ;
  assign n5790 = n4873 & ~n5789 ;
  assign n5778 = n4844 ^ n4841 ;
  assign n5779 = n5778 ^ n4863 ;
  assign n5774 = n4859 ^ n4846 ;
  assign n5776 = n5775 ^ n5774 ;
  assign n5777 = n4882 & n5776 ;
  assign n5780 = n5779 ^ n5777 ;
  assign n5782 = n5781 ^ n5780 ;
  assign n4874 = n4863 ^ n4844 ;
  assign n5769 = n4841 ^ n4839 ;
  assign n5770 = n5769 ^ n4841 ;
  assign n5771 = n4874 & n5770 ;
  assign n5772 = n5771 ^ n4841 ;
  assign n5773 = ~n4852 & n5772 ;
  assign n5783 = n5782 ^ n5773 ;
  assign n5791 = n5790 ^ n5783 ;
  assign n5793 = n5792 ^ n5791 ;
  assign n5794 = ~n4915 & n5793 ;
  assign n5795 = n5794 ^ n3550 ;
  assign n6912 = n5795 ^ x68 ;
  assign n4248 = n4214 ^ n4202 ;
  assign n4249 = ~n4247 & n4248 ;
  assign n4235 = n4201 ^ n4188 ;
  assign n4236 = n3971 & n4235 ;
  assign n4234 = n4233 ^ n4218 ;
  assign n4237 = n4236 ^ n4234 ;
  assign n4220 = n4219 ^ n4209 ;
  assign n4221 = n4220 ^ n4196 ;
  assign n4222 = n4221 ^ n4209 ;
  assign n4223 = n4209 ^ n3924 ;
  assign n4224 = n4223 ^ n4209 ;
  assign n4225 = ~n4222 & n4224 ;
  assign n4226 = n4225 ^ n4209 ;
  assign n4227 = ~n3969 & n4226 ;
  assign n4238 = n4237 ^ n4227 ;
  assign n4232 = ~n3970 & ~n4231 ;
  assign n4239 = n4238 ^ n4232 ;
  assign n4240 = n4239 ^ n4236 ;
  assign n4241 = n4240 ^ n4227 ;
  assign n4207 = n4206 ^ n4203 ;
  assign n4208 = n3924 & ~n4207 ;
  assign n4242 = n4241 ^ n4208 ;
  assign n4243 = n4200 & n4242 ;
  assign n4244 = n4243 ^ n4239 ;
  assign n4193 = n4192 ^ n4184 ;
  assign n4195 = n4194 ^ n4193 ;
  assign n4198 = n4197 ^ n4195 ;
  assign n4199 = n3971 & n4198 ;
  assign n4245 = n4244 ^ n4199 ;
  assign n4250 = n4249 ^ n4245 ;
  assign n4252 = n4251 ^ n4230 ;
  assign n4253 = n4230 ^ n3924 ;
  assign n4254 = n4253 ^ n4230 ;
  assign n4255 = ~n4252 & n4254 ;
  assign n4256 = n4255 ^ n4230 ;
  assign n4257 = n3969 & ~n4256 ;
  assign n4258 = ~n4250 & ~n4257 ;
  assign n4262 = n4258 ^ n2705 ;
  assign n4260 = n3924 & n4259 ;
  assign n4261 = n4258 & n4260 ;
  assign n4263 = n4262 ^ n4261 ;
  assign n6913 = n4263 ^ x94 ;
  assign n7011 = n6912 & ~n6913 ;
  assign n7014 = n7011 ^ n6912 ;
  assign n7027 = n6961 & n7014 ;
  assign n6939 = n6938 ^ n6914 ;
  assign n6973 = n6939 & n6944 ;
  assign n6974 = n6973 ^ n6944 ;
  assign n6959 = n6939 ^ n6936 ;
  assign n6960 = n6944 & n6959 ;
  assign n6962 = n6961 ^ n6960 ;
  assign n6975 = n6974 ^ n6962 ;
  assign n6951 = n6943 ^ n6914 ;
  assign n6952 = ~n6936 & ~n6951 ;
  assign n6984 = n6975 ^ n6952 ;
  assign n6953 = n6952 ^ n6943 ;
  assign n6954 = n6942 ^ n6936 ;
  assign n6955 = ~n6953 & ~n6954 ;
  assign n6945 = n6944 ^ n6942 ;
  assign n6946 = n6945 ^ n6943 ;
  assign n6948 = ~n6938 & n6946 ;
  assign n6949 = n6948 ^ n6946 ;
  assign n6950 = n6949 ^ n6937 ;
  assign n6956 = n6955 ^ n6950 ;
  assign n6957 = n6956 ^ n6948 ;
  assign n6985 = n6984 ^ n6957 ;
  assign n6980 = ~n6945 & n6959 ;
  assign n7018 = n6985 ^ n6980 ;
  assign n6987 = n6937 & ~n6945 ;
  assign n7017 = n6987 ^ n6945 ;
  assign n7019 = n7018 ^ n7017 ;
  assign n6967 = n6937 & n6946 ;
  assign n6947 = n6939 & n6946 ;
  assign n6968 = n6967 ^ n6947 ;
  assign n6969 = n6968 ^ n6949 ;
  assign n7020 = n7019 ^ n6969 ;
  assign n7021 = n7020 ^ n7018 ;
  assign n7022 = n7018 ^ n6912 ;
  assign n7023 = n7022 ^ n7018 ;
  assign n7024 = ~n7021 & ~n7023 ;
  assign n7025 = n7024 ^ n7018 ;
  assign n7026 = n6913 & n7025 ;
  assign n7028 = n7027 ^ n7026 ;
  assign n7015 = n6973 & n7014 ;
  assign n7012 = n7011 ^ n6913 ;
  assign n7013 = n6947 & ~n7012 ;
  assign n7016 = n7015 ^ n7013 ;
  assign n7029 = n7028 ^ n7016 ;
  assign n6988 = n6987 ^ n6948 ;
  assign n6981 = n6980 ^ n6969 ;
  assign n6979 = n6960 ^ n6959 ;
  assign n6982 = n6981 ^ n6979 ;
  assign n6989 = n6988 ^ n6982 ;
  assign n6990 = n6989 ^ n6980 ;
  assign n6971 = n6946 ^ n6942 ;
  assign n6972 = n6939 & n6971 ;
  assign n6976 = n6975 ^ n6972 ;
  assign n6963 = n6943 ^ n6942 ;
  assign n6964 = n6963 ^ n6914 ;
  assign n6965 = n6959 ^ n6943 ;
  assign n6966 = ~n6964 & n6965 ;
  assign n6970 = n6969 ^ n6966 ;
  assign n6977 = n6976 ^ n6970 ;
  assign n6978 = n6977 ^ n6975 ;
  assign n6983 = n6982 ^ n6978 ;
  assign n6986 = n6985 ^ n6983 ;
  assign n6991 = n6990 ^ n6986 ;
  assign n6992 = n6990 ^ n6913 ;
  assign n6993 = n6992 ^ n6990 ;
  assign n6994 = n6991 & n6993 ;
  assign n6995 = n6994 ^ n6990 ;
  assign n6996 = ~n6962 & ~n6995 ;
  assign n7030 = n7029 ^ n6996 ;
  assign n7004 = n6913 ^ n6912 ;
  assign n7005 = n6982 ^ n6977 ;
  assign n7006 = n6982 ^ n6913 ;
  assign n7007 = n7006 ^ n6982 ;
  assign n7008 = n7005 & ~n7007 ;
  assign n7009 = n7008 ^ n6982 ;
  assign n7010 = ~n7004 & n7009 ;
  assign n7031 = n7030 ^ n7010 ;
  assign n7032 = n7031 ^ n3585 ;
  assign n6997 = n6964 ^ n6955 ;
  assign n6998 = n6997 ^ n6996 ;
  assign n6958 = n6957 ^ n6947 ;
  assign n6999 = n6998 ^ n6958 ;
  assign n7000 = n6999 ^ n6996 ;
  assign n7001 = n6913 & ~n7000 ;
  assign n7002 = n7001 ^ n6998 ;
  assign n7003 = n6912 & n7002 ;
  assign n7033 = n7032 ^ n7003 ;
  assign n7034 = n7033 ^ x115 ;
  assign n6304 = n5792 ^ n3161 ;
  assign n6293 = n4877 ^ n4810 ;
  assign n6294 = ~n4883 & n6293 ;
  assign n6283 = n4861 ^ n4846 ;
  assign n6273 = ~n4746 & ~n4860 ;
  assign n4894 = n4886 ^ n4854 ;
  assign n4895 = n4894 ^ n4865 ;
  assign n6274 = n6273 ^ n4895 ;
  assign n6284 = n6283 ^ n6274 ;
  assign n6285 = n6274 ^ n4852 ;
  assign n6286 = n6285 ^ n6274 ;
  assign n6287 = n6284 & ~n6286 ;
  assign n6288 = n6287 ^ n6274 ;
  assign n6289 = n4873 & n6288 ;
  assign n6277 = n4886 ^ n4876 ;
  assign n6278 = n4876 ^ n4852 ;
  assign n6279 = n6278 ^ n4876 ;
  assign n6280 = n6277 & n6279 ;
  assign n6281 = n6280 ^ n4876 ;
  assign n6282 = n4873 & n6281 ;
  assign n6290 = n6289 ^ n6282 ;
  assign n6275 = n6274 ^ n4885 ;
  assign n6276 = n4879 & n6275 ;
  assign n6291 = n6290 ^ n6276 ;
  assign n4888 = n4887 ^ n4855 ;
  assign n6266 = n4888 ^ n4854 ;
  assign n6267 = n6266 ^ n4888 ;
  assign n6268 = n4888 ^ n4852 ;
  assign n6269 = n6268 ^ n4888 ;
  assign n6270 = n6267 & n6269 ;
  assign n6271 = n6270 ^ n4888 ;
  assign n6272 = ~n4873 & n6271 ;
  assign n6292 = n6291 ^ n6272 ;
  assign n6295 = n6294 ^ n6292 ;
  assign n6258 = n4863 ^ n4861 ;
  assign n6259 = n6258 ^ n4844 ;
  assign n6260 = n6259 ^ n4863 ;
  assign n6261 = n4863 ^ n4852 ;
  assign n6262 = n6261 ^ n4863 ;
  assign n6263 = n6260 & n6262 ;
  assign n6264 = n6263 ^ n4863 ;
  assign n6265 = ~n4873 & n6264 ;
  assign n6296 = n6295 ^ n6265 ;
  assign n6305 = n6304 ^ n6296 ;
  assign n6299 = ~n4839 & ~n6296 ;
  assign n6300 = n5786 & n6299 ;
  assign n6301 = n6300 ^ n5786 ;
  assign n4849 = n4848 ^ n4840 ;
  assign n4850 = ~n4839 & n4849 ;
  assign n4851 = n4850 ^ n4848 ;
  assign n6254 = n5786 ^ n4851 ;
  assign n6302 = n6301 ^ n6254 ;
  assign n6303 = n4852 & n6302 ;
  assign n6306 = n6305 ^ n6303 ;
  assign n7199 = n6306 ^ x92 ;
  assign n5383 = n5382 ^ n3763 ;
  assign n5392 = n5391 ^ n5383 ;
  assign n5393 = n5392 ^ n3253 ;
  assign n7087 = n5393 ^ x75 ;
  assign n7097 = n6022 ^ n4204 ;
  assign n7111 = n7097 ^ n4188 ;
  assign n7110 = n6026 ^ n4182 ;
  assign n7112 = n7111 ^ n7110 ;
  assign n7113 = n7110 ^ n3924 ;
  assign n7114 = n7113 ^ n7110 ;
  assign n7115 = n7112 & ~n7114 ;
  assign n7116 = n7115 ^ n7110 ;
  assign n7117 = ~n3969 & ~n7116 ;
  assign n7095 = n4218 ^ n4189 ;
  assign n7096 = n7095 ^ n4201 ;
  assign n7098 = n7097 ^ n7096 ;
  assign n7099 = ~n3969 & ~n7098 ;
  assign n7100 = n7099 ^ n7097 ;
  assign n7101 = n7100 ^ n4209 ;
  assign n6729 = n6044 ^ n4181 ;
  assign n7102 = n7101 ^ n6729 ;
  assign n7103 = n7102 ^ n7100 ;
  assign n7104 = n7100 ^ n3969 ;
  assign n7105 = n7104 ^ n7100 ;
  assign n7106 = n7103 & n7105 ;
  assign n7107 = n7106 ^ n7100 ;
  assign n7108 = ~n4200 & ~n7107 ;
  assign n7109 = n7108 ^ n7100 ;
  assign n7118 = n7117 ^ n7109 ;
  assign n7119 = n7118 ^ n4213 ;
  assign n6708 = n4213 ^ n3924 ;
  assign n6709 = n6708 ^ n4213 ;
  assign n6700 = n6026 ^ n4192 ;
  assign n6710 = n6700 ^ n4213 ;
  assign n6711 = n6709 & n6710 ;
  assign n6712 = n6711 ^ n4213 ;
  assign n6713 = n3969 & n6712 ;
  assign n7120 = n7119 ^ n6713 ;
  assign n7121 = n7120 ^ n4227 ;
  assign n7122 = n7121 ^ n3218 ;
  assign n7088 = n4219 ^ n4213 ;
  assign n7089 = n7088 ^ n4213 ;
  assign n7090 = n4213 ^ n3969 ;
  assign n7091 = n7090 ^ n4213 ;
  assign n7092 = n7089 & n7091 ;
  assign n7093 = n7092 ^ n4213 ;
  assign n7094 = n4200 & n7093 ;
  assign n7123 = n7122 ^ n7094 ;
  assign n7124 = n7123 ^ x124 ;
  assign n7125 = ~n7087 & ~n7124 ;
  assign n7126 = n7125 ^ n7087 ;
  assign n7144 = n5205 & n6103 ;
  assign n7141 = n5282 ^ n5249 ;
  assign n7142 = n5126 & n7141 ;
  assign n7133 = ~n5126 & n5217 ;
  assign n7129 = n5229 ^ n5224 ;
  assign n7134 = n7133 ^ n7129 ;
  assign n6370 = ~n5204 & n5283 ;
  assign n7138 = n7134 ^ n6370 ;
  assign n7139 = n7138 ^ n6101 ;
  assign n7135 = n7134 ^ n5164 ;
  assign n7130 = n7129 ^ n5215 ;
  assign n7131 = n7130 ^ n6079 ;
  assign n7132 = ~n5126 & ~n7131 ;
  assign n7136 = n7135 ^ n7132 ;
  assign n7137 = ~n5207 & ~n7136 ;
  assign n7140 = n7139 ^ n7137 ;
  assign n7143 = n7142 ^ n7140 ;
  assign n7145 = n7144 ^ n7143 ;
  assign n7146 = ~n5203 & n7145 ;
  assign n7147 = n7146 ^ n3188 ;
  assign n7148 = n7147 ^ x109 ;
  assign n4416 = n4415 ^ x72 ;
  assign n4462 = n3390 ^ n627 ;
  assign n4437 = n3355 ^ n3342 ;
  assign n4438 = n4437 ^ n3310 ;
  assign n4439 = n3348 ^ n3290 ;
  assign n4440 = n3163 & ~n4439 ;
  assign n4441 = ~n4438 & n4440 ;
  assign n4442 = n4441 ^ n3163 ;
  assign n4448 = n4442 ^ n3305 ;
  assign n4443 = n3353 & n3942 ;
  assign n4444 = ~n3307 & n4443 ;
  assign n4445 = n4444 ^ n3383 ;
  assign n4446 = n3383 & n4445 ;
  assign n4447 = ~n4442 & n4446 ;
  assign n4449 = n4448 ^ n4447 ;
  assign n4450 = n4449 ^ n4442 ;
  assign n4451 = n4450 ^ n4447 ;
  assign n4452 = n4451 ^ n4450 ;
  assign n4453 = n4450 ^ n3339 ;
  assign n4454 = n4453 ^ n4450 ;
  assign n4455 = n4452 & n4454 ;
  assign n4456 = n4455 ^ n4450 ;
  assign n4457 = n3164 & n4456 ;
  assign n4458 = n4457 ^ n4449 ;
  assign n4459 = n4458 ^ n3315 ;
  assign n4429 = n3349 ^ n3305 ;
  assign n4430 = n4429 ^ n3313 ;
  assign n4433 = n4432 ^ n4430 ;
  assign n4434 = n3162 & n4433 ;
  assign n4435 = n4434 ^ n3315 ;
  assign n4436 = ~n3383 & n4435 ;
  assign n4460 = n4459 ^ n4436 ;
  assign n4461 = ~n4428 & ~n4460 ;
  assign n4463 = n4462 ^ n4461 ;
  assign n4464 = n4463 ^ x112 ;
  assign n4465 = ~n4416 & ~n4464 ;
  assign n4466 = n4465 ^ n4464 ;
  assign n4467 = n4466 ^ n4416 ;
  assign n4468 = n4467 ^ n4464 ;
  assign n4487 = n4486 ^ x74 ;
  assign n4504 = n801 & n2205 ;
  assign n4505 = n4504 ^ n2203 ;
  assign n4506 = n4505 ^ n2206 ;
  assign n4507 = n4506 ^ n2197 ;
  assign n4508 = n4507 ^ n4505 ;
  assign n4511 = ~n801 & n4508 ;
  assign n4512 = n4511 ^ n4505 ;
  assign n4513 = n1273 & n4512 ;
  assign n4514 = n4513 ^ n4505 ;
  assign n4516 = n2210 ^ n2174 ;
  assign n4523 = n4516 ^ n2186 ;
  assign n4515 = n2254 ^ n2206 ;
  assign n4517 = n4516 ^ n4515 ;
  assign n4519 = n4515 ^ n1273 ;
  assign n4520 = n4518 & n4519 ;
  assign n4521 = n4520 ^ n1273 ;
  assign n4522 = n4517 & n4521 ;
  assign n4524 = n4523 ^ n4522 ;
  assign n4534 = n4533 ^ n4524 ;
  assign n4530 = n1276 & n2173 ;
  assign n4528 = n1274 & n2169 ;
  assign n4525 = n2193 ^ n2170 ;
  assign n4526 = n4525 ^ n2211 ;
  assign n4527 = n4526 ^ n4524 ;
  assign n4529 = n4528 ^ n4527 ;
  assign n4531 = n4530 ^ n4529 ;
  assign n4532 = n1277 & n4531 ;
  assign n4535 = n4534 ^ n4532 ;
  assign n4536 = ~n4514 & n4535 ;
  assign n4496 = n4495 ^ n2240 ;
  assign n4503 = n4502 ^ n4496 ;
  assign n4537 = n4536 ^ n4503 ;
  assign n4538 = ~n4488 & n4537 ;
  assign n4539 = n4538 ^ n517 ;
  assign n4540 = n4539 ^ x122 ;
  assign n4541 = ~n4487 & n4540 ;
  assign n4542 = ~n4468 & n4541 ;
  assign n4581 = n4580 ^ x98 ;
  assign n4604 = n4603 ^ x105 ;
  assign n4605 = n4581 & n4604 ;
  assign n4606 = n4542 & n4605 ;
  assign n4619 = ~n4467 & n4541 ;
  assign n4678 = n4604 ^ n4581 ;
  assign n4679 = n4619 & n4678 ;
  assign n4607 = n4541 ^ n4487 ;
  assign n4613 = n4607 ^ n4540 ;
  assign n4641 = ~n4468 & n4613 ;
  assign n4672 = n4641 ^ n4542 ;
  assign n4675 = n4581 & n4672 ;
  assign n4676 = n4675 ^ n4542 ;
  assign n4677 = ~n4604 & n4676 ;
  assign n4680 = n4679 ^ n4677 ;
  assign n4609 = n4605 ^ n4581 ;
  assign n6224 = n4542 & n4609 ;
  assign n4608 = ~n4466 & ~n4607 ;
  assign n4610 = n4608 & n4609 ;
  assign n6225 = n6224 ^ n4610 ;
  assign n4620 = n4619 ^ n4542 ;
  assign n4614 = n4613 ^ n4487 ;
  assign n4618 = n4465 & n4614 ;
  assign n4621 = n4620 ^ n4618 ;
  assign n4616 = n4487 ^ n4464 ;
  assign n4617 = n4540 & n4616 ;
  assign n4622 = n4621 ^ n4617 ;
  assign n4615 = ~n4467 & n4614 ;
  assign n4623 = n4622 ^ n4615 ;
  assign n6217 = n4623 ^ n4618 ;
  assign n4611 = ~n4466 & n4541 ;
  assign n4645 = n4611 ^ n4541 ;
  assign n4646 = n4645 ^ n4620 ;
  assign n4647 = n4646 ^ n4608 ;
  assign n4648 = n4647 ^ n4542 ;
  assign n4643 = n4541 ^ n4466 ;
  assign n4634 = n4622 ^ n4619 ;
  assign n4644 = n4643 ^ n4634 ;
  assign n4649 = n4648 ^ n4644 ;
  assign n4642 = n4641 ^ n4615 ;
  assign n4650 = n4649 ^ n4642 ;
  assign n4662 = n4649 ^ n4641 ;
  assign n6210 = n4662 ^ n4604 ;
  assign n4690 = n4622 ^ n4604 ;
  assign n6211 = n6210 ^ n4690 ;
  assign n6212 = n6211 ^ n4604 ;
  assign n6213 = n4678 ^ n4604 ;
  assign n6214 = n6212 & ~n6213 ;
  assign n6215 = n6214 ^ n4604 ;
  assign n6216 = ~n4650 & n6215 ;
  assign n6218 = n6217 ^ n6216 ;
  assign n4627 = ~n4468 & ~n4607 ;
  assign n4632 = n4627 ^ n4608 ;
  assign n4631 = ~n4467 & n4613 ;
  assign n4633 = n4632 ^ n4631 ;
  assign n4635 = n4634 ^ n4633 ;
  assign n4624 = n4623 ^ n4608 ;
  assign n4636 = n4635 ^ n4624 ;
  assign n4630 = n4627 ^ n4467 ;
  assign n4637 = n4636 ^ n4630 ;
  assign n6219 = n6218 ^ n4637 ;
  assign n6226 = n6225 ^ n6219 ;
  assign n4657 = n4618 ^ n4614 ;
  assign n4658 = n4657 ^ n4623 ;
  assign n4628 = n4627 ^ n4611 ;
  assign n5810 = n4658 ^ n4628 ;
  assign n5811 = n4658 ^ n4604 ;
  assign n5812 = n5811 ^ n4658 ;
  assign n5813 = n5810 & n5812 ;
  assign n5814 = n5813 ^ n4658 ;
  assign n5815 = ~n4678 & n5814 ;
  assign n6227 = n6226 ^ n5815 ;
  assign n4661 = n4631 ^ n4613 ;
  assign n4663 = n4662 ^ n4661 ;
  assign n4659 = n4631 ^ n4618 ;
  assign n4660 = n4659 ^ n4658 ;
  assign n4664 = n4663 ^ n4660 ;
  assign n6220 = n6219 ^ n4664 ;
  assign n4638 = n4632 ^ n4607 ;
  assign n4639 = n4638 ^ n4637 ;
  assign n4640 = n4639 ^ n4611 ;
  assign n6207 = n4640 ^ n4615 ;
  assign n6221 = n6220 ^ n6207 ;
  assign n6204 = n4637 ^ n4634 ;
  assign n6205 = n6204 ^ n4646 ;
  assign n6203 = n4664 ^ n4649 ;
  assign n6206 = n6205 ^ n6203 ;
  assign n6208 = n6207 ^ n6206 ;
  assign n6209 = ~n4604 & ~n6208 ;
  assign n6222 = n6221 ^ n6209 ;
  assign n6223 = ~n4581 & n6222 ;
  assign n6228 = n6227 ^ n6223 ;
  assign n6229 = ~n4680 & n6228 ;
  assign n4669 = n4605 ^ n4604 ;
  assign n4670 = n4669 ^ n4581 ;
  assign n4671 = ~n4663 & ~n4670 ;
  assign n6230 = n6229 ^ n4671 ;
  assign n6231 = ~n4606 & n6230 ;
  assign n6232 = n6231 ^ n3283 ;
  assign n7149 = n6232 ^ x102 ;
  assign n7150 = ~n7148 & n7149 ;
  assign n7170 = n7150 ^ n7149 ;
  assign n7171 = n7170 ^ n7148 ;
  assign n7174 = ~n7126 & n7171 ;
  assign n7127 = n7126 ^ n7124 ;
  assign n7173 = ~n7127 & n7171 ;
  assign n7175 = n7174 ^ n7173 ;
  assign n7176 = n7175 ^ n7171 ;
  assign n7128 = n7127 ^ n7087 ;
  assign n7172 = ~n7128 & n7171 ;
  assign n7177 = n7176 ^ n7172 ;
  assign n7164 = n7125 & n7150 ;
  assign n7157 = ~n7127 & n7150 ;
  assign n7165 = n7164 ^ n7157 ;
  assign n7162 = ~n7128 & n7150 ;
  assign n7163 = n7162 ^ n7150 ;
  assign n7166 = n7165 ^ n7163 ;
  assign n7184 = n7177 ^ n7166 ;
  assign n7153 = n7124 & n7149 ;
  assign n7167 = n7166 ^ n7153 ;
  assign n7154 = n7148 ^ n7087 ;
  assign n7155 = n7154 ^ n7124 ;
  assign n7159 = ~n7087 & n7155 ;
  assign n7160 = n7159 ^ n7124 ;
  assign n7161 = n7149 & n7160 ;
  assign n7168 = n7167 ^ n7161 ;
  assign n7183 = n7168 ^ n7159 ;
  assign n7185 = n7184 ^ n7183 ;
  assign n7186 = n7185 ^ n7168 ;
  assign n7182 = n7166 ^ n7162 ;
  assign n7187 = n7186 ^ n7182 ;
  assign n7181 = n7175 ^ n7162 ;
  assign n7188 = n7187 ^ n7181 ;
  assign n7189 = n7188 ^ n7124 ;
  assign n7190 = n7189 ^ n7161 ;
  assign n7242 = n7190 ^ n7174 ;
  assign n7151 = n7150 ^ n7148 ;
  assign n7152 = ~n7128 & ~n7151 ;
  assign n7243 = n7242 ^ n7152 ;
  assign n5709 = ~n5605 & n5701 ;
  assign n5710 = n5709 ^ n5692 ;
  assign n5713 = n5710 ^ n5703 ;
  assign n5714 = n5713 ^ n5710 ;
  assign n5715 = n5605 & n5714 ;
  assign n5716 = n5715 ^ n5710 ;
  assign n5717 = n5606 & n5716 ;
  assign n5718 = n5717 ^ n5710 ;
  assign n5748 = ~n5609 & n5693 ;
  assign n5745 = n5744 ^ n5743 ;
  assign n5746 = ~n5608 & n5745 ;
  assign n5740 = n5607 & n5688 ;
  assign n5726 = n5678 ^ n5606 ;
  assign n5731 = n5730 ^ n5678 ;
  assign n5732 = n5731 ^ n5605 ;
  assign n5733 = n5732 ^ n5731 ;
  assign n5734 = n5704 ^ n5678 ;
  assign n5735 = n5734 ^ n5731 ;
  assign n5736 = ~n5733 & n5735 ;
  assign n5737 = n5736 ^ n5731 ;
  assign n5738 = n5726 & ~n5737 ;
  assign n5739 = n5738 ^ n5606 ;
  assign n5741 = n5740 ^ n5739 ;
  assign n5747 = n5746 ^ n5741 ;
  assign n5749 = n5748 ^ n5747 ;
  assign n5721 = n5684 ^ n5606 ;
  assign n5722 = n5721 ^ n5684 ;
  assign n5723 = ~n5698 & n5722 ;
  assign n5724 = n5723 ^ n5684 ;
  assign n5725 = ~n5605 & n5724 ;
  assign n5750 = n5749 ^ n5725 ;
  assign n5751 = ~n5718 & ~n5750 ;
  assign n5752 = ~n5708 & n5751 ;
  assign n5753 = ~n5707 & n5752 ;
  assign n5763 = n5753 & ~n5762 ;
  assign n5764 = n5763 ^ n3125 ;
  assign n7086 = n5764 ^ x78 ;
  assign n7244 = n7152 ^ n7086 ;
  assign n7245 = n7244 ^ n7152 ;
  assign n7246 = n7243 & n7245 ;
  assign n7247 = n7246 ^ n7152 ;
  assign n7248 = ~n7199 & n7247 ;
  assign n7249 = n7248 ^ n3393 ;
  assign n7212 = n7199 ^ n7086 ;
  assign n7216 = n7161 ^ n7155 ;
  assign n7156 = n7153 & ~n7155 ;
  assign n7158 = n7157 ^ n7156 ;
  assign n7214 = n7186 ^ n7158 ;
  assign n7213 = n7177 ^ n7157 ;
  assign n7215 = n7214 ^ n7213 ;
  assign n7217 = n7216 ^ n7215 ;
  assign n7218 = n7215 ^ n7086 ;
  assign n7219 = n7218 ^ n7215 ;
  assign n7220 = n7217 & n7219 ;
  assign n7221 = n7220 ^ n7215 ;
  assign n7222 = n7212 & n7221 ;
  assign n7223 = n7222 ^ n7215 ;
  assign n7205 = n7086 & ~n7199 ;
  assign n7206 = n7205 ^ n7199 ;
  assign n7208 = n7206 ^ n7086 ;
  assign n7178 = n7177 ^ n7125 ;
  assign n7169 = n7168 ^ n7164 ;
  assign n7179 = n7178 ^ n7169 ;
  assign n7191 = n7179 ^ n7173 ;
  assign n7192 = n7191 ^ n7190 ;
  assign n7193 = n7192 ^ n7157 ;
  assign n7180 = n7179 ^ n7127 ;
  assign n7194 = n7193 ^ n7180 ;
  assign n7209 = n7194 ^ n7155 ;
  assign n7210 = n7209 ^ n7156 ;
  assign n7211 = n7208 & n7210 ;
  assign n7224 = n7223 ^ n7211 ;
  assign n7207 = n7164 & ~n7206 ;
  assign n7225 = n7224 ^ n7207 ;
  assign n7228 = n7177 ^ n7086 ;
  assign n7229 = n7228 ^ n7177 ;
  assign n7230 = n7184 & ~n7229 ;
  assign n7231 = n7230 ^ n7177 ;
  assign n7232 = n7199 & n7231 ;
  assign n7233 = ~n7225 & ~n7232 ;
  assign n7196 = n7170 ^ n7168 ;
  assign n7195 = n7194 ^ n7158 ;
  assign n7197 = n7196 ^ n7195 ;
  assign n7198 = n7197 ^ n7152 ;
  assign n7202 = ~n7198 & n7199 ;
  assign n7203 = n7202 ^ n7197 ;
  assign n7204 = n7086 & ~n7203 ;
  assign n7234 = n7233 ^ n7204 ;
  assign n7235 = n7195 ^ n7191 ;
  assign n7236 = n7191 ^ n7086 ;
  assign n7237 = n7236 ^ n7191 ;
  assign n7238 = ~n7235 & ~n7237 ;
  assign n7239 = n7238 ^ n7191 ;
  assign n7240 = ~n7212 & n7239 ;
  assign n7241 = n7234 & ~n7240 ;
  assign n7250 = n7249 ^ n7241 ;
  assign n7251 = n7250 ^ x121 ;
  assign n5816 = n4605 & ~n4663 ;
  assign n5817 = n5816 ^ n4606 ;
  assign n6455 = n6225 ^ n5817 ;
  assign n6448 = n6207 ^ n4659 ;
  assign n6447 = n6205 ^ n4641 ;
  assign n6449 = n6448 ^ n6447 ;
  assign n6450 = ~n4604 & ~n6449 ;
  assign n6451 = n6450 ^ n6447 ;
  assign n6456 = n6455 ^ n6451 ;
  assign n6457 = n6456 ^ n4671 ;
  assign n4688 = n4637 ^ n4618 ;
  assign n4689 = n4688 ^ n4622 ;
  assign n4691 = n4690 ^ n4622 ;
  assign n4692 = ~n4689 & ~n4691 ;
  assign n4693 = n4692 ^ n4622 ;
  assign n4694 = ~n4581 & n4693 ;
  assign n6458 = n6457 ^ n4694 ;
  assign n6446 = n4647 ^ n4642 ;
  assign n6452 = n6451 ^ n6446 ;
  assign n6442 = n4647 ^ n4487 ;
  assign n6443 = n6442 ^ n4644 ;
  assign n6444 = n6443 ^ n4642 ;
  assign n6445 = n4604 & n6444 ;
  assign n6453 = n6452 ^ n6445 ;
  assign n6454 = ~n4581 & ~n6453 ;
  assign n6459 = n6458 ^ n6454 ;
  assign n6460 = ~n4658 & n6459 ;
  assign n6461 = n6460 ^ n800 ;
  assign n6462 = n6461 ^ x114 ;
  assign n5561 = n5011 ^ n4997 ;
  assign n6488 = n5561 ^ n5022 ;
  assign n6489 = ~n5103 & n6488 ;
  assign n6484 = n5096 ^ n5015 ;
  assign n6485 = n5071 & ~n6484 ;
  assign n6481 = n5028 ^ n5011 ;
  assign n6482 = n5070 & ~n6481 ;
  assign n6248 = n5028 & ~n5103 ;
  assign n6474 = n6248 ^ n5100 ;
  assign n6475 = n6474 ^ n5027 ;
  assign n5585 = n5028 ^ n5026 ;
  assign n6476 = n5585 ^ n5097 ;
  assign n6477 = ~n5103 & n6476 ;
  assign n6478 = n6477 ^ n5069 ;
  assign n6479 = ~n6475 & n6478 ;
  assign n5558 = n5068 ^ n4920 ;
  assign n5598 = ~n5023 & ~n5068 ;
  assign n5599 = n5598 ^ n5022 ;
  assign n5600 = ~n5558 & ~n5599 ;
  assign n6480 = n6479 ^ n5600 ;
  assign n6483 = n6482 ^ n6480 ;
  assign n6486 = n6485 ^ n6483 ;
  assign n6465 = n5004 ^ n5002 ;
  assign n6487 = n6486 ^ n6465 ;
  assign n6490 = n6489 ^ n6487 ;
  assign n5584 = n5009 ^ n5008 ;
  assign n5586 = n5585 ^ n5584 ;
  assign n6466 = n6465 ^ n5586 ;
  assign n6467 = n6466 ^ n5030 ;
  assign n6468 = n6467 ^ n6465 ;
  assign n6469 = n6465 ^ n4920 ;
  assign n6470 = n6469 ^ n6465 ;
  assign n6471 = n6468 & n6470 ;
  assign n6472 = n6471 ^ n6465 ;
  assign n6473 = ~n5558 & n6472 ;
  assign n6491 = n6490 ^ n6473 ;
  assign n5557 = n5021 & n5070 ;
  assign n6492 = n6491 ^ n5557 ;
  assign n6493 = n6492 ^ n1669 ;
  assign n6494 = n6493 ^ x81 ;
  assign n6311 = n5547 ^ n5479 ;
  assign n6525 = n6311 ^ n5505 ;
  assign n6526 = n5505 ^ n5483 ;
  assign n6527 = n6526 ^ n5505 ;
  assign n6528 = ~n6525 & n6527 ;
  assign n6529 = n6528 ^ n5505 ;
  assign n6530 = n5395 & n6529 ;
  assign n6510 = n5546 ^ n5476 ;
  assign n6511 = n6510 ^ n5545 ;
  assign n6508 = n5544 ^ n5501 ;
  assign n6509 = ~n5534 & ~n6508 ;
  assign n6512 = n6511 ^ n6509 ;
  assign n6513 = n6512 ^ n5467 ;
  assign n6507 = ~n5544 & n5981 ;
  assign n6514 = n6513 ^ n6507 ;
  assign n6504 = n5479 ^ n5468 ;
  assign n6505 = n6504 ^ n5985 ;
  assign n6506 = n6505 ^ n5492 ;
  assign n6515 = n6514 ^ n6506 ;
  assign n6310 = n5981 ^ n5468 ;
  assign n6502 = n6310 ^ n5481 ;
  assign n6503 = n6502 ^ n5479 ;
  assign n6516 = n6515 ^ n6503 ;
  assign n6517 = n6516 ^ n6514 ;
  assign n6518 = ~n5483 & ~n6517 ;
  assign n6519 = n6518 ^ n6515 ;
  assign n6521 = n6514 ^ n5395 ;
  assign n6520 = n6514 ^ n5483 ;
  assign n6522 = n6521 ^ n6520 ;
  assign n6523 = n6519 & n6522 ;
  assign n6524 = n6523 ^ n6521 ;
  assign n6531 = n6530 ^ n6524 ;
  assign n6495 = n5985 ^ n5534 ;
  assign n6496 = n5539 ^ n5499 ;
  assign n6499 = ~n5985 & n6496 ;
  assign n6500 = n6499 ^ n5539 ;
  assign n6501 = ~n6495 & n6500 ;
  assign n6532 = n6531 ^ n6501 ;
  assign n6533 = ~n5516 & ~n6532 ;
  assign n6534 = n6533 ^ n1913 ;
  assign n6535 = n6534 ^ x120 ;
  assign n6536 = n6494 & ~n6535 ;
  assign n6557 = n5792 ^ n2164 ;
  assign n6551 = n4895 ^ n4855 ;
  assign n6552 = ~n4883 & n6551 ;
  assign n6540 = n4866 ^ n4844 ;
  assign n6541 = n6540 ^ n4840 ;
  assign n6547 = n6541 ^ n4810 ;
  assign n6543 = n6273 ^ n4874 ;
  assign n6544 = n6543 ^ n4857 ;
  assign n6542 = n6541 ^ n4846 ;
  assign n6545 = n6544 ^ n6542 ;
  assign n6546 = ~n4852 & n6545 ;
  assign n6548 = n6547 ^ n6546 ;
  assign n6549 = n4873 & n6548 ;
  assign n6539 = n6282 ^ n5785 ;
  assign n6550 = n6549 ^ n6539 ;
  assign n6553 = n6552 ^ n6550 ;
  assign n6538 = n4852 & n4881 ;
  assign n6554 = n6553 ^ n6538 ;
  assign n4896 = n4895 ^ n4848 ;
  assign n4897 = n4896 ^ n4856 ;
  assign n6537 = n4880 & n4897 ;
  assign n6555 = n6554 ^ n6537 ;
  assign n6556 = ~n4915 & ~n6555 ;
  assign n6558 = n6557 ^ n6556 ;
  assign n6559 = n6558 ^ x74 ;
  assign n6560 = n5975 ^ x64 ;
  assign n6561 = n6559 & ~n6560 ;
  assign n6562 = n6561 ^ n6559 ;
  assign n6563 = n6562 ^ n6560 ;
  assign n6574 = n6563 ^ n6559 ;
  assign n6586 = n6536 & ~n6574 ;
  assign n6618 = n6586 ^ n6574 ;
  assign n6567 = n6536 ^ n6535 ;
  assign n6577 = ~n6567 & ~n6574 ;
  assign n6575 = n6536 ^ n6494 ;
  assign n6576 = ~n6574 & n6575 ;
  assign n6578 = n6577 ^ n6576 ;
  assign n6619 = n6618 ^ n6578 ;
  assign n6602 = n6562 & n6575 ;
  assign n6644 = n6619 ^ n6602 ;
  assign n6463 = n6060 ^ x105 ;
  assign n6645 = n6602 ^ n6463 ;
  assign n6646 = n6645 ^ n6602 ;
  assign n6647 = ~n6644 & n6646 ;
  assign n6648 = n6647 ^ n6602 ;
  assign n6649 = n6462 & n6648 ;
  assign n6464 = n6463 ^ n6462 ;
  assign n6568 = n6560 & ~n6567 ;
  assign n6579 = n6568 ^ n6567 ;
  assign n6580 = n6579 ^ n6577 ;
  assign n6597 = n6586 ^ n6580 ;
  assign n6583 = n6567 ^ n6494 ;
  assign n6584 = n6562 & n6583 ;
  assign n7076 = n6597 ^ n6584 ;
  assign n6625 = n6563 & ~n6567 ;
  assign n6626 = n6625 ^ n6568 ;
  assign n6622 = n6563 & n6583 ;
  assign n6627 = n6626 ^ n6622 ;
  assign n6628 = n6627 ^ n6563 ;
  assign n6564 = n6536 & n6563 ;
  assign n6569 = n6568 ^ n6564 ;
  assign n6629 = n6628 ^ n6569 ;
  assign n7074 = n6629 ^ n6625 ;
  assign n6588 = n6561 & n6575 ;
  assign n7075 = n7074 ^ n6588 ;
  assign n7077 = n7076 ^ n7075 ;
  assign n7078 = n6463 & ~n7077 ;
  assign n6585 = n6561 & n6583 ;
  assign n6587 = n6586 ^ n6585 ;
  assign n7056 = n6619 ^ n6587 ;
  assign n7079 = n7078 ^ n7056 ;
  assign n7080 = ~n6464 & ~n7079 ;
  assign n6582 = n6462 & n6463 ;
  assign n6616 = n6582 ^ n6462 ;
  assign n6617 = n6616 ^ n6463 ;
  assign n7071 = n6577 & ~n6617 ;
  assign n6589 = n6588 ^ n6587 ;
  assign n6596 = n6589 ^ n6561 ;
  assign n6598 = n6597 ^ n6596 ;
  assign n6599 = n6598 ^ n6564 ;
  assign n6595 = n6586 ^ n6536 ;
  assign n6600 = n6599 ^ n6595 ;
  assign n6642 = ~n6600 & n6616 ;
  assign n7072 = n7071 ^ n6642 ;
  assign n7067 = n6617 ^ n6462 ;
  assign n7068 = ~n6600 & n7067 ;
  assign n7060 = n6625 ^ n6602 ;
  assign n7061 = n7060 ^ n6580 ;
  assign n7062 = n6580 ^ n6462 ;
  assign n7063 = n7062 ^ n6580 ;
  assign n7064 = ~n7061 & ~n7063 ;
  assign n7065 = n7064 ^ n6580 ;
  assign n7066 = ~n6463 & ~n7065 ;
  assign n7069 = n7068 ^ n7066 ;
  assign n7051 = n6598 ^ n6462 ;
  assign n7052 = n7051 ^ n6598 ;
  assign n7053 = ~n6599 & n7052 ;
  assign n7054 = n7053 ^ n6598 ;
  assign n7055 = n6463 & ~n7054 ;
  assign n7057 = n7056 ^ n7055 ;
  assign n7042 = n6598 ^ n6585 ;
  assign n6630 = n6629 ^ n6626 ;
  assign n7043 = n7042 ^ n6630 ;
  assign n7044 = n6630 ^ n6462 ;
  assign n7045 = n7044 ^ n6630 ;
  assign n7046 = ~n7043 & ~n7045 ;
  assign n7047 = n7046 ^ n6630 ;
  assign n7048 = ~n6463 & n7047 ;
  assign n7058 = n7057 ^ n7048 ;
  assign n6651 = n6602 ^ n6584 ;
  assign n6652 = ~n6646 & n6651 ;
  assign n6653 = n6652 ^ n6602 ;
  assign n6654 = ~n6462 & n6653 ;
  assign n7059 = n7058 ^ n6654 ;
  assign n7070 = n7069 ^ n7059 ;
  assign n7073 = n7072 ^ n7070 ;
  assign n7081 = n7080 ^ n7073 ;
  assign n7035 = n6576 ^ n6564 ;
  assign n7036 = n7035 ^ n6627 ;
  assign n7037 = n6627 ^ n6463 ;
  assign n7038 = n7037 ^ n6627 ;
  assign n7039 = n7036 & ~n7038 ;
  assign n7040 = n7039 ^ n6627 ;
  assign n7041 = ~n6462 & n7040 ;
  assign n7082 = n7081 ^ n7041 ;
  assign n7083 = ~n6649 & n7082 ;
  assign n7084 = n7083 ^ n2281 ;
  assign n7085 = n7084 ^ x122 ;
  assign n7299 = n7251 ^ n7085 ;
  assign n6728 = n4189 ^ n4182 ;
  assign n6730 = n6729 ^ n6728 ;
  assign n6731 = ~n4247 & n6730 ;
  assign n6719 = n4219 ^ n4205 ;
  assign n6720 = n6719 ^ n4228 ;
  assign n6721 = n4228 ^ n3924 ;
  assign n6722 = n6721 ^ n4228 ;
  assign n6723 = n6720 & n6722 ;
  assign n6724 = n6723 ^ n4228 ;
  assign n6725 = n3969 & n6724 ;
  assign n6714 = n6713 ^ n4236 ;
  assign n6715 = n6714 ^ n4257 ;
  assign n6716 = n6715 ^ n4227 ;
  assign n6717 = n6716 ^ n2932 ;
  assign n6703 = n6700 ^ n3969 ;
  assign n6704 = n6703 ^ n6700 ;
  assign n6705 = n4209 & ~n6704 ;
  assign n6706 = n6705 ^ n6700 ;
  assign n6707 = n4200 & n6706 ;
  assign n6718 = n6717 ^ n6707 ;
  assign n6726 = n6725 ^ n6718 ;
  assign n6699 = n4217 & n4246 ;
  assign n6727 = n6726 ^ n6699 ;
  assign n6732 = n6731 ^ n6727 ;
  assign n6733 = n6732 ^ x97 ;
  assign n6734 = n3774 ^ n3612 ;
  assign n6735 = n3586 & n6734 ;
  assign n6736 = n6735 ^ n3774 ;
  assign n6744 = n6736 ^ n2955 ;
  assign n6737 = n6736 ^ n3785 ;
  assign n6738 = n6737 ^ n3396 ;
  assign n6739 = n6738 ^ n3787 ;
  assign n6740 = n6739 ^ n6736 ;
  assign n6741 = n3586 & n6740 ;
  assign n6742 = n6741 ^ n6737 ;
  assign n6743 = ~n3763 & n6742 ;
  assign n6745 = n6744 ^ n6743 ;
  assign n6746 = n6745 ^ x98 ;
  assign n6242 = n5035 ^ n5018 ;
  assign n6243 = ~n4920 & ~n6242 ;
  assign n6244 = n6243 ^ n5018 ;
  assign n6249 = n6248 ^ n6244 ;
  assign n6250 = n6249 ^ n5102 ;
  assign n6251 = n6250 ^ n2983 ;
  assign n5562 = n5561 ^ n5001 ;
  assign n6240 = n5562 ^ n5097 ;
  assign n6241 = n6240 ^ n5111 ;
  assign n6245 = n6244 ^ n6241 ;
  assign n6234 = n4955 ^ n4921 ;
  assign n6237 = n4986 & ~n6234 ;
  assign n6238 = n6237 ^ n4921 ;
  assign n6239 = ~n4920 & ~n6238 ;
  assign n6246 = n6245 ^ n6239 ;
  assign n6247 = ~n5068 & ~n6246 ;
  assign n6252 = n6251 ^ n6247 ;
  assign n6747 = n6252 ^ x80 ;
  assign n6748 = n6461 ^ x107 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6750 = n6746 & n6749 ;
  assign n6751 = n6750 ^ n6749 ;
  assign n6752 = ~n6733 & n6751 ;
  assign n6753 = n6752 ^ n6751 ;
  assign n6371 = n6370 ^ n6105 ;
  assign n6372 = n6371 ^ n5237 ;
  assign n6373 = n6372 ^ n2895 ;
  assign n6361 = n5225 ^ n5221 ;
  assign n6359 = n5128 & n5220 ;
  assign n6357 = n5282 ^ n5230 ;
  assign n6358 = n6357 ^ n5241 ;
  assign n6360 = n6359 ^ n6358 ;
  assign n6362 = n6361 ^ n6360 ;
  assign n6356 = n5205 & n5227 ;
  assign n6363 = n6362 ^ n6356 ;
  assign n6364 = n5127 ^ n5126 ;
  assign n6365 = ~n6363 & n6364 ;
  assign n6366 = n6365 ^ n5126 ;
  assign n6350 = n5220 ^ n5213 ;
  assign n6351 = n5220 ^ n5127 ;
  assign n6352 = n6351 ^ n5220 ;
  assign n6353 = ~n6350 & n6352 ;
  assign n6354 = n6353 ^ n5220 ;
  assign n6355 = ~n5126 & n6354 ;
  assign n6367 = n6366 ^ n6355 ;
  assign n6342 = n5226 ^ n5224 ;
  assign n6343 = n6342 ^ n5206 ;
  assign n6344 = n6079 ^ n5204 ;
  assign n6347 = ~n6342 & n6344 ;
  assign n6348 = n6347 ^ n5204 ;
  assign n6349 = n6343 & ~n6348 ;
  assign n6368 = n6367 ^ n6349 ;
  assign n6369 = ~n6067 & ~n6368 ;
  assign n6374 = n6373 ^ n6369 ;
  assign n6754 = n6374 ^ x65 ;
  assign n6755 = n6534 ^ x104 ;
  assign n6756 = ~n6754 & n6755 ;
  assign n6757 = n6756 ^ n6754 ;
  assign n6758 = n6757 ^ n6755 ;
  assign n6759 = n6753 & n6758 ;
  assign n6761 = ~n6746 & ~n6748 ;
  assign n6760 = n6748 ^ n6746 ;
  assign n6762 = n6761 ^ n6760 ;
  assign n6768 = n6733 & ~n6762 ;
  assign n6788 = ~n6747 & n6768 ;
  assign n6789 = n6756 ^ n6755 ;
  assign n6790 = n6788 & n6789 ;
  assign n6769 = ~n6733 & n6746 ;
  assign n6781 = n6749 & n6769 ;
  assign n6770 = n6769 ^ n6762 ;
  assign n6771 = n6770 ^ n6768 ;
  assign n6782 = n6781 ^ n6771 ;
  assign n6763 = n6762 ^ n6748 ;
  assign n6773 = n6733 & n6747 ;
  assign n6778 = ~n6763 & n6773 ;
  assign n6776 = n6746 & n6773 ;
  assign n6777 = n6776 ^ n6773 ;
  assign n6779 = n6778 ^ n6777 ;
  assign n6775 = n6761 ^ n6751 ;
  assign n6780 = n6779 ^ n6775 ;
  assign n6783 = n6782 ^ n6780 ;
  assign n6774 = n6773 ^ n6747 ;
  assign n6784 = n6783 ^ n6774 ;
  assign n6772 = n6771 ^ n6769 ;
  assign n6785 = n6784 ^ n6772 ;
  assign n6764 = n6733 & ~n6763 ;
  assign n6765 = n6764 ^ n6763 ;
  assign n6766 = ~n6747 & ~n6765 ;
  assign n6767 = n6766 ^ n6765 ;
  assign n6786 = n6785 ^ n6767 ;
  assign n6787 = n6756 & ~n6786 ;
  assign n6791 = n6790 ^ n6787 ;
  assign n6792 = ~n6759 & ~n6791 ;
  assign n6845 = n6754 ^ n6747 ;
  assign n6846 = n6845 ^ n6754 ;
  assign n6847 = n6756 & n6846 ;
  assign n6848 = n6847 ^ n6754 ;
  assign n6849 = ~n6765 & ~n6848 ;
  assign n6793 = n6755 ^ n6754 ;
  assign n6836 = n6778 ^ n6764 ;
  assign n6837 = n6836 ^ n6785 ;
  assign n6838 = n6837 ^ n6836 ;
  assign n6839 = n6836 ^ n6754 ;
  assign n6840 = n6839 ^ n6836 ;
  assign n6841 = n6838 & n6840 ;
  assign n6842 = n6841 ^ n6836 ;
  assign n6843 = ~n6793 & n6842 ;
  assign n6850 = n6849 ^ n6843 ;
  assign n6801 = n6781 ^ n6750 ;
  assign n6818 = n6801 ^ n6780 ;
  assign n6819 = n6818 ^ n6753 ;
  assign n6795 = n6776 ^ n6768 ;
  assign n6796 = n6795 ^ n6788 ;
  assign n6810 = n6796 ^ n6778 ;
  assign n6811 = n6810 ^ n6782 ;
  assign n6812 = n6811 ^ n6752 ;
  assign n6813 = n6812 ^ n6796 ;
  assign n6814 = ~n6754 & ~n6813 ;
  assign n6815 = n6814 ^ n6810 ;
  assign n6820 = n6819 ^ n6815 ;
  assign n6824 = n6820 ^ n6781 ;
  assign n6797 = n6796 ^ n6776 ;
  assign n6794 = n6786 ^ n6772 ;
  assign n6798 = n6797 ^ n6794 ;
  assign n6817 = n6798 ^ n6765 ;
  assign n6821 = n6820 ^ n6817 ;
  assign n6822 = n6821 ^ n6815 ;
  assign n6823 = n6754 & ~n6822 ;
  assign n6825 = n6824 ^ n6823 ;
  assign n6826 = n6793 & n6825 ;
  assign n6803 = n6780 ^ n6779 ;
  assign n6804 = n6779 ^ n6754 ;
  assign n6805 = n6804 ^ n6779 ;
  assign n6806 = n6803 & n6805 ;
  assign n6807 = n6806 ^ n6779 ;
  assign n6808 = n6755 & n6807 ;
  assign n6809 = n6808 ^ n6781 ;
  assign n6816 = n6815 ^ n6809 ;
  assign n6827 = n6826 ^ n6816 ;
  assign n6851 = n6850 ^ n6827 ;
  assign n6834 = n6758 & n6779 ;
  assign n6833 = ~n6757 & n6788 ;
  assign n6835 = n6834 ^ n6833 ;
  assign n6852 = n6851 ^ n6835 ;
  assign n6799 = n6798 ^ n6755 ;
  assign n6800 = n6799 ^ n6798 ;
  assign n6802 = n6801 ^ n6782 ;
  assign n6828 = ~n6802 & ~n6827 ;
  assign n6829 = n6828 ^ n6798 ;
  assign n6830 = ~n6800 & n6829 ;
  assign n6831 = n6830 ^ n6798 ;
  assign n6832 = n6793 & n6831 ;
  assign n6853 = n6852 ^ n6832 ;
  assign n6854 = n6792 & ~n6853 ;
  assign n6855 = n6854 ^ n3071 ;
  assign n7292 = n6855 ^ x74 ;
  assign n7321 = n7299 ^ n7292 ;
  assign n4264 = n4263 ^ x84 ;
  assign n4651 = n4646 ^ n4619 ;
  assign n4652 = n4651 ^ n4650 ;
  assign n4653 = n4652 ^ n4640 ;
  assign n4654 = n4604 & ~n4653 ;
  assign n4655 = n4654 ^ n4646 ;
  assign n4682 = n4663 ^ n4655 ;
  assign n4681 = n4680 ^ n4671 ;
  assign n4683 = n4682 ^ n4681 ;
  assign n4668 = ~n4604 & n4660 ;
  assign n4684 = n4683 ^ n4668 ;
  assign n4629 = n4628 ^ n4623 ;
  assign n4656 = n4655 ^ n4629 ;
  assign n4665 = n4664 ^ n4656 ;
  assign n4612 = n4611 ^ n4542 ;
  assign n4625 = n4624 ^ n4612 ;
  assign n4626 = n4604 & n4625 ;
  assign n4666 = n4665 ^ n4626 ;
  assign n4667 = ~n4581 & ~n4666 ;
  assign n4685 = n4684 ^ n4667 ;
  assign n4686 = n4685 ^ n4610 ;
  assign n4687 = ~n4606 & n4686 ;
  assign n4695 = n4687 & ~n4694 ;
  assign n4696 = n4695 ^ n2630 ;
  assign n4697 = n4696 ^ x69 ;
  assign n4698 = ~n4264 & n4697 ;
  assign n4699 = n4698 ^ n4697 ;
  assign n4700 = n4699 ^ n4264 ;
  assign n4701 = n4700 ^ n4697 ;
  assign n4867 = n4840 ^ n4810 ;
  assign n4868 = n4867 ^ n4866 ;
  assign n4869 = n4839 & n4868 ;
  assign n4853 = n4851 ^ n4847 ;
  assign n4870 = n4869 ^ n4853 ;
  assign n4871 = ~n4852 & n4870 ;
  assign n4872 = n4871 ^ n4851 ;
  assign n4906 = n4877 ^ n4842 ;
  assign n4907 = n4880 & n4906 ;
  assign n4878 = n4877 ^ n4807 ;
  assign n4884 = n4881 & ~n4883 ;
  assign n4889 = n4888 ^ n4884 ;
  assign n4890 = ~n4880 & n4889 ;
  assign n4891 = n4878 & n4890 ;
  assign n4892 = n4891 ^ n4889 ;
  assign n4893 = n4892 ^ n4874 ;
  assign n4898 = n4897 ^ n4893 ;
  assign n4899 = n4898 ^ n4892 ;
  assign n4900 = n4892 ^ n4852 ;
  assign n4901 = n4900 ^ n4892 ;
  assign n4902 = n4899 & n4901 ;
  assign n4903 = n4902 ^ n4892 ;
  assign n4904 = n4873 & n4903 ;
  assign n4905 = n4904 ^ n4892 ;
  assign n4908 = n4907 ^ n4905 ;
  assign n4909 = ~n4872 & ~n4908 ;
  assign n4916 = n4909 & ~n4915 ;
  assign n4917 = ~n4810 & n4916 ;
  assign n4918 = n4917 ^ n2663 ;
  assign n4919 = n4918 ^ x118 ;
  assign n5114 = n5113 ^ x125 ;
  assign n5115 = ~n4919 & n5114 ;
  assign n5116 = n5115 ^ n5114 ;
  assign n5117 = n5116 ^ n4919 ;
  assign n5118 = ~n4701 & n5117 ;
  assign n3798 = n3797 ^ x101 ;
  assign n5291 = n5290 ^ x83 ;
  assign n5297 = ~n3798 & n5291 ;
  assign n5298 = n5297 ^ n5291 ;
  assign n5299 = n5298 ^ n3798 ;
  assign n7287 = n5118 & n5299 ;
  assign n5322 = n4699 & n5116 ;
  assign n7284 = n5298 & n5322 ;
  assign n7275 = n4919 ^ n3798 ;
  assign n7276 = n7275 ^ n4919 ;
  assign n7277 = n5117 & n7276 ;
  assign n7278 = n7277 ^ n4919 ;
  assign n7279 = n5291 & n7278 ;
  assign n7280 = n4700 & n7279 ;
  assign n5121 = n5115 ^ n4919 ;
  assign n5123 = ~n4701 & ~n5121 ;
  assign n5119 = n4698 & n5116 ;
  assign n5311 = n5123 ^ n5119 ;
  assign n5312 = n5311 ^ n5118 ;
  assign n5310 = ~n4701 & n5116 ;
  assign n5313 = n5312 ^ n5310 ;
  assign n5309 = n5119 ^ n4701 ;
  assign n5314 = n5313 ^ n5309 ;
  assign n5315 = n5314 ^ n5115 ;
  assign n5304 = n4699 & ~n5121 ;
  assign n5305 = n5304 ^ n5121 ;
  assign n5122 = n4698 & ~n5121 ;
  assign n5124 = n5123 ^ n5122 ;
  assign n5306 = n5305 ^ n5124 ;
  assign n5302 = n4700 & n4919 ;
  assign n5303 = n5302 ^ n4700 ;
  assign n5307 = n5306 ^ n5303 ;
  assign n5301 = n4698 & n5115 ;
  assign n5308 = n5307 ^ n5301 ;
  assign n5316 = n5315 ^ n5308 ;
  assign n5324 = n5316 ^ n5304 ;
  assign n5323 = n5322 ^ n4699 ;
  assign n5325 = n5324 ^ n5323 ;
  assign n7262 = n5325 ^ n5304 ;
  assign n5350 = n5301 ^ n5122 ;
  assign n7263 = n7262 ^ n5350 ;
  assign n7264 = ~n5291 & n7263 ;
  assign n7265 = n7264 ^ n5350 ;
  assign n5372 = n5314 ^ n5118 ;
  assign n5373 = n5298 & ~n5372 ;
  assign n7271 = n7265 ^ n5373 ;
  assign n5300 = n5299 ^ n5297 ;
  assign n5351 = n5350 ^ n4264 ;
  assign n5352 = n5351 ^ n5309 ;
  assign n5353 = n5352 ^ n5291 ;
  assign n5354 = n5353 ^ n5352 ;
  assign n5333 = n4700 & n5116 ;
  assign n5334 = n5333 ^ n5302 ;
  assign n5355 = n5334 ^ n5316 ;
  assign n5356 = n5355 ^ n5352 ;
  assign n5357 = ~n5354 & n5356 ;
  assign n5358 = n5357 ^ n5352 ;
  assign n5359 = n5300 & n5358 ;
  assign n7272 = n7271 ^ n5359 ;
  assign n7281 = n7280 ^ n7272 ;
  assign n7267 = n5123 ^ n4701 ;
  assign n7268 = n5291 & ~n7267 ;
  assign n7266 = n7265 ^ n5313 ;
  assign n7269 = n7268 ^ n7266 ;
  assign n7270 = ~n3798 & n7269 ;
  assign n7282 = n7281 ^ n7270 ;
  assign n7260 = n5325 ^ n5307 ;
  assign n7261 = ~n5300 & ~n7260 ;
  assign n7283 = n7282 ^ n7261 ;
  assign n7285 = n7284 ^ n7283 ;
  assign n7254 = n5324 ^ n5311 ;
  assign n7255 = n5311 ^ n3798 ;
  assign n7256 = n7255 ^ n5311 ;
  assign n7257 = n7254 & ~n7256 ;
  assign n7258 = n7257 ^ n5311 ;
  assign n7259 = ~n5291 & n7258 ;
  assign n7286 = n7285 ^ n7259 ;
  assign n7288 = n7287 ^ n7286 ;
  assign n7289 = n7288 ^ n2854 ;
  assign n5317 = n5316 ^ n5306 ;
  assign n5318 = n5317 ^ n5310 ;
  assign n5319 = n5291 & ~n5318 ;
  assign n5320 = n5319 ^ n5310 ;
  assign n7253 = n5300 & n5320 ;
  assign n7290 = n7289 ^ n7253 ;
  assign n7291 = n7290 ^ x112 ;
  assign n7315 = n7299 ^ n7291 ;
  assign n7316 = n7291 ^ n7085 ;
  assign n7317 = n7315 & ~n7316 ;
  assign n7322 = n7317 ^ n7291 ;
  assign n7323 = n7321 & ~n7322 ;
  assign n7324 = n7323 ^ n7292 ;
  assign n7318 = n7317 ^ n7251 ;
  assign n7319 = ~n7292 & n7318 ;
  assign n7309 = n7292 ^ n7251 ;
  assign n7310 = ~n7299 & n7309 ;
  assign n7311 = n7309 ^ n7291 ;
  assign n7312 = ~n7310 & n7311 ;
  assign n7295 = ~n7085 & n7292 ;
  assign n7296 = n7291 & n7295 ;
  assign n7313 = n7312 ^ n7296 ;
  assign n7298 = n7291 ^ n7251 ;
  assign n7300 = ~n7291 & n7299 ;
  assign n7301 = n7300 ^ n7292 ;
  assign n7302 = n7298 & n7301 ;
  assign n7303 = n7302 ^ n7299 ;
  assign n7293 = n7292 ^ n7085 ;
  assign n7294 = ~n7291 & ~n7293 ;
  assign n7297 = n7296 ^ n7294 ;
  assign n7304 = n7303 ^ n7297 ;
  assign n7252 = n7085 & n7251 ;
  assign n7305 = n7304 ^ n7252 ;
  assign n7314 = n7313 ^ n7305 ;
  assign n7320 = n7319 ^ n7314 ;
  assign n7325 = n7324 ^ n7320 ;
  assign n7308 = n7297 ^ n7295 ;
  assign n7326 = n7325 ^ n7308 ;
  assign n7327 = n7326 ^ n7317 ;
  assign n7328 = n7327 ^ n7326 ;
  assign n7329 = n7326 ^ n7312 ;
  assign n7330 = n7329 ^ n7326 ;
  assign n7331 = ~n7328 & ~n7330 ;
  assign n7332 = n7331 ^ n7326 ;
  assign n7333 = ~n7034 & n7332 ;
  assign n7334 = n7333 ^ n7326 ;
  assign n7306 = n7034 & n7305 ;
  assign n7307 = n7306 ^ n7303 ;
  assign n7335 = n7334 ^ n7307 ;
  assign n7336 = ~n6911 & ~n7335 ;
  assign n7337 = n7336 ^ n7334 ;
  assign n9383 = n7337 ^ n6911 ;
  assign n9384 = n9383 ^ n7334 ;
  assign n9385 = n9384 ^ n7307 ;
  assign n9386 = n9385 ^ n5393 ;
  assign n10077 = n9386 ^ x85 ;
  assign n6199 = n6198 ^ x86 ;
  assign n5394 = n5393 ^ x117 ;
  assign n5554 = n5553 ^ x67 ;
  assign n5555 = n5394 & n5554 ;
  assign n5842 = n5555 ^ n5394 ;
  assign n5843 = n5842 ^ n5554 ;
  assign n5844 = n5843 ^ n5394 ;
  assign n5556 = n5032 & n5069 ;
  assign n5569 = n5028 ^ n4920 ;
  assign n5571 = n5028 ^ n5014 ;
  assign n5570 = n5100 ^ n5028 ;
  assign n5572 = n5571 ^ n5570 ;
  assign n5573 = n5571 ^ n5068 ;
  assign n5574 = n5573 ^ n5571 ;
  assign n5575 = ~n5572 & n5574 ;
  assign n5576 = n5575 ^ n5571 ;
  assign n5577 = n5569 & n5576 ;
  assign n5578 = n5577 ^ n4920 ;
  assign n5568 = ~n5016 & ~n5103 ;
  assign n5579 = n5578 ^ n5568 ;
  assign n5563 = n5562 ^ n5015 ;
  assign n5564 = n5563 ^ n5010 ;
  assign n5565 = n5068 & n5564 ;
  assign n5566 = n5565 ^ n5010 ;
  assign n5567 = n5558 & n5566 ;
  assign n5580 = n5579 ^ n5567 ;
  assign n5581 = ~n5557 & ~n5580 ;
  assign n5582 = ~n5104 & n5581 ;
  assign n5583 = ~n5556 & n5582 ;
  assign n5587 = n5586 ^ n4998 ;
  assign n5588 = n4998 ^ n4920 ;
  assign n5589 = n5588 ^ n4998 ;
  assign n5590 = n5587 & ~n5589 ;
  assign n5591 = n5590 ^ n4998 ;
  assign n5592 = ~n5558 & n5591 ;
  assign n5593 = n5583 & ~n5592 ;
  assign n5601 = n5593 & ~n5600 ;
  assign n5602 = ~n5102 & n5601 ;
  assign n5603 = n5602 ^ n4328 ;
  assign n5604 = n5603 ^ x110 ;
  assign n5765 = n5764 ^ x100 ;
  assign n5766 = n5604 & ~n5765 ;
  assign n5846 = n5766 ^ n5604 ;
  assign n5796 = n5795 ^ x93 ;
  assign n5828 = n4581 & n4646 ;
  assign n5804 = n4638 ^ n4620 ;
  assign n5805 = n5804 ^ n4650 ;
  assign n5806 = n5805 ^ n4638 ;
  assign n5807 = n5806 ^ n4658 ;
  assign n5808 = ~n4604 & ~n5807 ;
  assign n5809 = n5808 ^ n5804 ;
  assign n5822 = n4618 ^ n4605 ;
  assign n5823 = n5822 ^ n4642 ;
  assign n5824 = n4669 & n5823 ;
  assign n5819 = n5817 ^ n4678 ;
  assign n5820 = n5819 ^ n5815 ;
  assign n5818 = n5817 ^ n5815 ;
  assign n5821 = n5820 ^ n5818 ;
  assign n5825 = n5824 ^ n5821 ;
  assign n5826 = n5809 & n5825 ;
  assign n5827 = n5826 ^ n5820 ;
  assign n5829 = n5828 ^ n5827 ;
  assign n5797 = n4624 ^ n4604 ;
  assign n5798 = n5797 ^ n4624 ;
  assign n5801 = n4636 & ~n5798 ;
  assign n5802 = n5801 ^ n4624 ;
  assign n5803 = ~n4678 & n5802 ;
  assign n5830 = n5829 ^ n5803 ;
  assign n5831 = ~n4610 & ~n5830 ;
  assign n5832 = ~n4694 & n5831 ;
  assign n5833 = n5832 ^ n4299 ;
  assign n5834 = n5833 ^ x91 ;
  assign n5835 = n5796 & n5834 ;
  assign n5848 = n5835 ^ n5834 ;
  assign n5857 = n5848 ^ n5796 ;
  assign n5858 = n5846 & ~n5857 ;
  assign n5836 = n5835 ^ n5796 ;
  assign n5854 = n5836 & n5846 ;
  assign n5855 = n5854 ^ n5836 ;
  assign n5838 = n5766 ^ n5765 ;
  assign n5839 = n5836 & ~n5838 ;
  assign n5837 = n5766 & n5836 ;
  assign n5840 = n5839 ^ n5837 ;
  assign n5856 = n5855 ^ n5840 ;
  assign n5859 = n5858 ^ n5856 ;
  assign n5926 = n5844 & n5859 ;
  assign n5847 = n5846 ^ n5765 ;
  assign n5872 = n5835 & n5847 ;
  assign n5871 = n5847 & ~n5857 ;
  assign n5873 = n5872 ^ n5871 ;
  assign n5923 = n5844 & n5873 ;
  assign n5863 = n5846 & n5848 ;
  assign n5922 = n5555 & n5863 ;
  assign n5924 = n5923 ^ n5922 ;
  assign n5910 = n5554 ^ n5394 ;
  assign n5912 = ~n5838 & ~n5857 ;
  assign n5895 = n5766 & n5835 ;
  assign n5849 = n5847 & n5848 ;
  assign n5864 = n5863 ^ n5849 ;
  assign n5861 = n5766 & n5848 ;
  assign n5862 = n5861 ^ n5848 ;
  assign n5865 = n5864 ^ n5862 ;
  assign n5896 = n5895 ^ n5865 ;
  assign n5913 = n5912 ^ n5896 ;
  assign n5911 = n5896 ^ n5861 ;
  assign n5914 = n5913 ^ n5911 ;
  assign n5915 = n5913 ^ n5554 ;
  assign n5916 = n5915 ^ n5913 ;
  assign n5917 = n5914 & n5916 ;
  assign n5918 = n5917 ^ n5913 ;
  assign n5919 = ~n5910 & n5918 ;
  assign n5920 = n5919 ^ n5896 ;
  assign n5902 = n5766 & ~n5857 ;
  assign n5894 = n5873 ^ n5837 ;
  assign n5897 = n5896 ^ n5894 ;
  assign n5898 = ~n5554 & n5897 ;
  assign n5899 = n5898 ^ n5837 ;
  assign n5903 = n5902 ^ n5899 ;
  assign n5904 = n5903 ^ n5899 ;
  assign n5905 = n5554 & n5904 ;
  assign n5906 = n5905 ^ n5899 ;
  assign n5907 = n5394 & n5906 ;
  assign n5908 = n5907 ^ n5899 ;
  assign n5869 = n5835 & n5846 ;
  assign n5886 = n5869 ^ n5858 ;
  assign n5889 = n5858 ^ n5394 ;
  assign n5890 = n5889 ^ n5858 ;
  assign n5891 = n5886 & ~n5890 ;
  assign n5892 = n5891 ^ n5858 ;
  assign n5893 = ~n5554 & n5892 ;
  assign n5909 = n5908 ^ n5893 ;
  assign n5921 = n5920 ^ n5909 ;
  assign n5925 = n5924 ^ n5921 ;
  assign n5927 = n5926 ^ n5925 ;
  assign n5928 = n5927 ^ n5453 ;
  assign n5841 = n5555 & n5840 ;
  assign n5845 = n5844 ^ n5842 ;
  assign n5860 = n5859 ^ n5839 ;
  assign n5866 = n5865 ^ n5860 ;
  assign n5853 = n5765 ^ n5604 ;
  assign n5867 = n5866 ^ n5853 ;
  assign n5868 = ~n5554 & ~n5867 ;
  assign n5870 = n5869 ^ n5868 ;
  assign n5874 = n5873 ^ n5870 ;
  assign n5850 = n5849 ^ n5839 ;
  assign n5851 = ~n5554 & n5850 ;
  assign n5852 = n5851 ^ n5849 ;
  assign n5875 = n5874 ^ n5852 ;
  assign n5876 = n5875 ^ n5858 ;
  assign n5877 = n5876 ^ n5873 ;
  assign n5878 = n5877 ^ n5875 ;
  assign n5879 = n5875 ^ n5554 ;
  assign n5880 = n5879 ^ n5875 ;
  assign n5881 = n5878 & ~n5880 ;
  assign n5882 = n5881 ^ n5875 ;
  assign n5883 = ~n5845 & n5882 ;
  assign n5884 = n5883 ^ n5870 ;
  assign n5885 = ~n5841 & ~n5884 ;
  assign n5929 = n5928 ^ n5885 ;
  assign n5930 = n5929 ^ x108 ;
  assign n6673 = n6199 ^ n5930 ;
  assign n6233 = n6232 ^ x113 ;
  assign n6253 = n6252 ^ x66 ;
  assign n6375 = n6374 ^ x73 ;
  assign n6307 = n6306 ^ x90 ;
  assign n6404 = n6375 ^ n6307 ;
  assign n6387 = n5697 ^ n5693 ;
  assign n6388 = n6387 ^ n5942 ;
  assign n6389 = ~n5606 & n6388 ;
  assign n6385 = n5697 ^ n5685 ;
  assign n6379 = n5933 ^ n5698 ;
  assign n6380 = n6379 ^ n5706 ;
  assign n6378 = n6377 ^ n5682 ;
  assign n6381 = n6380 ^ n6378 ;
  assign n6382 = n5606 & n6381 ;
  assign n6383 = n6382 ^ n6380 ;
  assign n6386 = n6385 ^ n6383 ;
  assign n6390 = n6389 ^ n6386 ;
  assign n6391 = ~n5605 & ~n6390 ;
  assign n6376 = n5972 ^ n5718 ;
  assign n6384 = n6383 ^ n6376 ;
  assign n6392 = n6391 ^ n6384 ;
  assign n6393 = ~n5762 & n6392 ;
  assign n6394 = n6393 ^ n3856 ;
  assign n6395 = n6394 ^ x99 ;
  assign n6416 = n6395 ^ n6307 ;
  assign n6332 = n5481 ^ n5476 ;
  assign n6312 = n6311 ^ n6310 ;
  assign n6313 = n6312 ^ n5533 ;
  assign n6314 = n5503 ^ n5499 ;
  assign n6315 = n6314 ^ n6312 ;
  assign n6316 = ~n6313 & n6315 ;
  assign n6317 = n6316 ^ n5533 ;
  assign n6309 = n5539 ^ n5516 ;
  assign n6321 = n6317 ^ n6309 ;
  assign n6319 = ~n5490 & ~n5521 ;
  assign n6320 = n6309 & n6319 ;
  assign n6322 = n6321 ^ n6320 ;
  assign n6308 = ~n5395 & ~n5519 ;
  assign n6323 = n6322 ^ n6308 ;
  assign n6325 = n6312 ^ n5499 ;
  assign n6324 = n5501 ^ n5480 ;
  assign n6326 = n6325 ^ n6324 ;
  assign n6327 = n5395 & ~n6326 ;
  assign n6328 = n6327 ^ n6324 ;
  assign n6329 = ~n5483 & ~n6328 ;
  assign n6330 = ~n6323 & n6329 ;
  assign n6331 = n6330 ^ n6323 ;
  assign n6333 = ~n5980 & ~n6331 ;
  assign n6334 = n6332 & n6333 ;
  assign n6335 = n6334 ^ n6331 ;
  assign n6337 = n5395 & n5467 ;
  assign n6338 = ~n6335 & n6337 ;
  assign n6336 = n6335 ^ n3822 ;
  assign n6339 = n6338 ^ n6336 ;
  assign n6340 = n6339 ^ x72 ;
  assign n6417 = n6416 ^ n6340 ;
  assign n6418 = n6375 & n6417 ;
  assign n6419 = n6418 ^ n6340 ;
  assign n6420 = ~n6404 & ~n6419 ;
  assign n6428 = n6420 ^ n6419 ;
  assign n6401 = n6395 ^ n6340 ;
  assign n6405 = ~n6340 & ~n6404 ;
  assign n6406 = n6405 ^ n6375 ;
  assign n6402 = n6307 & n6340 ;
  assign n6403 = n6402 ^ n6340 ;
  assign n6407 = n6406 ^ n6403 ;
  assign n6408 = n6401 & ~n6407 ;
  assign n6427 = n6408 & ~n6416 ;
  assign n6429 = n6428 ^ n6427 ;
  assign n6425 = n6402 ^ n6307 ;
  assign n6412 = n6375 ^ n6340 ;
  assign n6413 = n6307 & ~n6412 ;
  assign n6426 = n6425 ^ n6413 ;
  assign n6430 = n6429 ^ n6426 ;
  assign n6431 = n6430 ^ n6340 ;
  assign n6432 = n6431 ^ n6395 ;
  assign n6433 = n6432 ^ n6427 ;
  assign n6423 = n6412 ^ n6307 ;
  assign n6414 = n6413 ^ n6375 ;
  assign n6415 = ~n6401 & ~n6414 ;
  assign n6421 = n6420 ^ n6415 ;
  assign n6409 = n6395 ^ n6375 ;
  assign n6410 = n6409 ^ n6408 ;
  assign n6422 = n6421 ^ n6410 ;
  assign n6424 = n6423 ^ n6422 ;
  assign n6434 = n6433 ^ n6424 ;
  assign n6435 = n6253 & n6434 ;
  assign n6436 = n6435 ^ n6424 ;
  assign n6341 = n6340 ^ n6307 ;
  assign n6396 = n6375 & n6395 ;
  assign n6397 = n6396 ^ n6340 ;
  assign n6398 = n6341 & ~n6397 ;
  assign n6399 = n6398 ^ n6340 ;
  assign n6400 = ~n6253 & n6399 ;
  assign n6411 = n6410 ^ n6400 ;
  assign n6437 = n6436 ^ n6411 ;
  assign n6438 = ~n6233 & n6437 ;
  assign n6439 = n6438 ^ n6436 ;
  assign n6440 = n6439 ^ n3923 ;
  assign n6441 = n6440 ^ x126 ;
  assign n6620 = ~n6617 & ~n6619 ;
  assign n6610 = n6598 ^ n6576 ;
  assign n6611 = n6610 ^ n6586 ;
  assign n6590 = n6589 ^ n6584 ;
  assign n6591 = n6462 & n6590 ;
  assign n6592 = n6591 ^ n6589 ;
  assign n6612 = n6611 ^ n6592 ;
  assign n6608 = n6578 ^ n6574 ;
  assign n6609 = n6462 & ~n6608 ;
  assign n6613 = n6612 ^ n6609 ;
  assign n6614 = ~n6463 & ~n6613 ;
  assign n6601 = n6600 ^ n6564 ;
  assign n6603 = n6602 ^ n6601 ;
  assign n6604 = n6463 & ~n6603 ;
  assign n6593 = n6592 ^ n6580 ;
  assign n6594 = n6593 ^ n6592 ;
  assign n6605 = n6604 ^ n6594 ;
  assign n6606 = ~n6464 & ~n6605 ;
  assign n6607 = n6606 ^ n6593 ;
  assign n6615 = n6614 ^ n6607 ;
  assign n6621 = n6620 ^ n6615 ;
  assign n6623 = n6622 ^ n6463 ;
  assign n6624 = n6623 ^ n6622 ;
  assign n6631 = ~n6462 & n6630 ;
  assign n6632 = n6631 ^ n6622 ;
  assign n6633 = n6624 & n6632 ;
  assign n6634 = n6633 ^ n6622 ;
  assign n6635 = n6621 & n6634 ;
  assign n6636 = n6635 ^ n6621 ;
  assign n6639 = n6636 ^ n6564 ;
  assign n6581 = n6580 ^ n6578 ;
  assign n6637 = n6582 & n6636 ;
  assign n6638 = ~n6581 & n6637 ;
  assign n6640 = n6639 ^ n6638 ;
  assign n6565 = n6564 ^ n6462 ;
  assign n6566 = n6565 ^ n6564 ;
  assign n6571 = ~n6566 & n6568 ;
  assign n6572 = n6571 ^ n6564 ;
  assign n6573 = ~n6464 & n6572 ;
  assign n6641 = n6640 ^ n6573 ;
  assign n6643 = n6642 ^ n6641 ;
  assign n6650 = n6643 & ~n6649 ;
  assign n6655 = n6650 & ~n6654 ;
  assign n6656 = n6655 ^ n5423 ;
  assign n6657 = n6656 ^ x93 ;
  assign n6674 = n6657 ^ n5930 ;
  assign n6675 = ~n6441 & ~n6674 ;
  assign n6676 = n6675 ^ n5930 ;
  assign n6677 = n6673 & ~n6676 ;
  assign n6678 = n6677 ^ n6199 ;
  assign n6200 = ~n5930 & ~n6199 ;
  assign n6201 = n6200 ^ n5930 ;
  assign n6658 = ~n6441 & n6657 ;
  assign n6664 = n6658 ^ n6441 ;
  assign n6665 = ~n6201 & ~n6664 ;
  assign n6202 = n6201 ^ n6199 ;
  assign n6672 = n6665 ^ n6202 ;
  assign n6679 = n6678 ^ n6672 ;
  assign n6667 = n6200 ^ n6199 ;
  assign n6659 = n6658 ^ n6657 ;
  assign n6670 = n6659 ^ n6441 ;
  assign n6671 = ~n6667 & n6670 ;
  assign n6680 = n6679 ^ n6671 ;
  assign n6668 = n6659 & ~n6667 ;
  assign n6669 = n6668 ^ n6667 ;
  assign n6681 = n6680 ^ n6669 ;
  assign n5376 = n5333 ^ n5325 ;
  assign n5377 = n5299 & n5376 ;
  assign n5337 = n5291 ^ n3798 ;
  assign n5360 = n5310 ^ n5301 ;
  assign n5361 = n5360 ^ n5291 ;
  assign n5362 = n5361 ^ n5360 ;
  assign n5363 = n5352 ^ n5310 ;
  assign n5364 = n5363 ^ n5360 ;
  assign n5365 = ~n5362 & n5364 ;
  assign n5366 = n5365 ^ n5360 ;
  assign n5367 = n5337 & n5366 ;
  assign n5368 = n5367 ^ n5310 ;
  assign n5342 = n5322 ^ n5304 ;
  assign n5335 = n5334 ^ n5307 ;
  assign n5343 = n5342 ^ n5335 ;
  assign n5332 = n5306 ^ n5119 ;
  assign n5336 = n5335 ^ n5332 ;
  assign n5338 = n5335 ^ n5291 ;
  assign n5339 = n5337 & ~n5338 ;
  assign n5340 = n5339 ^ n5291 ;
  assign n5341 = n5336 & n5340 ;
  assign n5344 = n5343 ^ n5341 ;
  assign n5345 = n5344 ^ n5301 ;
  assign n5326 = n5325 ^ n5122 ;
  assign n5329 = n5291 & n5326 ;
  assign n5330 = n5329 ^ n5122 ;
  assign n5331 = n5300 & n5330 ;
  assign n5346 = n5345 ^ n5331 ;
  assign n5369 = n5368 ^ n5346 ;
  assign n5370 = n5369 ^ n5359 ;
  assign n5321 = n5320 ^ n5307 ;
  assign n5347 = n5346 ^ n5321 ;
  assign n5348 = n5347 ^ n5331 ;
  assign n5349 = n5300 & n5348 ;
  assign n5371 = n5370 ^ n5349 ;
  assign n5374 = n5373 ^ n5371 ;
  assign n5120 = n5119 ^ n5118 ;
  assign n5125 = n5124 ^ n5120 ;
  assign n5294 = n5125 & n5291 ;
  assign n5295 = n5294 ^ n5124 ;
  assign n5296 = ~n3798 & n5295 ;
  assign n5375 = n5374 ^ n5296 ;
  assign n5378 = n5377 ^ n5375 ;
  assign n5379 = n5378 ^ n4176 ;
  assign n5380 = n5379 ^ x125 ;
  assign n6856 = n6855 ^ x76 ;
  assign n6869 = n5380 & ~n6856 ;
  assign n6907 = n6681 & n6869 ;
  assign n6908 = n6907 ^ n5553 ;
  assign n6862 = n6856 ^ n5380 ;
  assign n6863 = n6657 ^ n6441 ;
  assign n6864 = n6199 & n6863 ;
  assign n6865 = n6864 ^ n6199 ;
  assign n6684 = n6200 & ~n6664 ;
  assign n6690 = n6684 ^ n6681 ;
  assign n6691 = n6690 ^ n6668 ;
  assign n6661 = ~n6201 & n6658 ;
  assign n6692 = n6691 ^ n6661 ;
  assign n6686 = n6200 & n6658 ;
  assign n6687 = n6686 ^ n6200 ;
  assign n6683 = n6200 & n6670 ;
  assign n6685 = n6684 ^ n6683 ;
  assign n6688 = n6687 ^ n6685 ;
  assign n6689 = n6688 ^ n6684 ;
  assign n6693 = n6692 ^ n6689 ;
  assign n6682 = n6681 ^ n6659 ;
  assign n6694 = n6693 ^ n6682 ;
  assign n6660 = ~n6202 & n6659 ;
  assign n6662 = n6661 ^ n6660 ;
  assign n6695 = n6694 ^ n6662 ;
  assign n6666 = n6665 ^ n6660 ;
  assign n6696 = n6695 ^ n6666 ;
  assign n6866 = n6865 ^ n6696 ;
  assign n6867 = n6862 & n6866 ;
  assign n6663 = n6662 ^ n6201 ;
  assign n6697 = n6696 ^ n6663 ;
  assign n6698 = n6697 ^ n6695 ;
  assign n6859 = ~n6698 & n6856 ;
  assign n6860 = n6859 ^ n6695 ;
  assign n6861 = ~n5380 & n6860 ;
  assign n6868 = n6867 ^ n6861 ;
  assign n6893 = n6687 ^ n6679 ;
  assign n6892 = n6680 ^ n6662 ;
  assign n6894 = n6893 ^ n6892 ;
  assign n6895 = n6894 ^ n6680 ;
  assign n6896 = n6680 ^ n5380 ;
  assign n6897 = n6896 ^ n6680 ;
  assign n6898 = ~n6895 & ~n6897 ;
  assign n6899 = n6898 ^ n6680 ;
  assign n6900 = n6856 & n6899 ;
  assign n6901 = n6900 ^ n6680 ;
  assign n6885 = n6697 ^ n6665 ;
  assign n6886 = n6885 ^ n6864 ;
  assign n6887 = n6864 ^ n6856 ;
  assign n6888 = n6887 ^ n6864 ;
  assign n6889 = n6886 & ~n6888 ;
  assign n6890 = n6889 ^ n6864 ;
  assign n6891 = n5380 & n6890 ;
  assign n6902 = n6901 ^ n6891 ;
  assign n6876 = n6688 ^ n6681 ;
  assign n6872 = n6869 ^ n6856 ;
  assign n6877 = n6876 ^ n6872 ;
  assign n6878 = n6665 ^ n6662 ;
  assign n6873 = n6872 ^ n5380 ;
  assign n6874 = n6873 ^ n6856 ;
  assign n6879 = n6878 ^ n6874 ;
  assign n6880 = n6878 ^ n6872 ;
  assign n6881 = n6880 ^ n6878 ;
  assign n6882 = ~n6879 & n6881 ;
  assign n6883 = n6882 ^ n6878 ;
  assign n6884 = ~n6877 & ~n6883 ;
  assign n6903 = n6902 ^ n6884 ;
  assign n6875 = n6685 & n6874 ;
  assign n6904 = n6903 ^ n6875 ;
  assign n6870 = n6686 ^ n6668 ;
  assign n6871 = n6869 & n6870 ;
  assign n6905 = n6904 ^ n6871 ;
  assign n6906 = ~n6868 & ~n6905 ;
  assign n6909 = n6908 ^ n6906 ;
  assign n10078 = n6909 ^ x102 ;
  assign n10079 = n10077 & n10078 ;
  assign n10080 = n10079 ^ n10078 ;
  assign n10081 = n10080 ^ n10077 ;
  assign n7359 = n6600 ^ n6588 ;
  assign n7360 = n6588 ^ n6463 ;
  assign n7361 = n7360 ^ n6588 ;
  assign n7362 = ~n7359 & n7361 ;
  assign n7363 = n7362 ^ n6588 ;
  assign n7364 = n6462 & n7363 ;
  assign n7365 = n7364 ^ n6463 ;
  assign n7366 = n7365 ^ n7048 ;
  assign n7367 = n7366 ^ n7069 ;
  assign n7352 = n6630 ^ n6580 ;
  assign n7350 = n6610 ^ n6587 ;
  assign n7351 = n7350 ^ n6625 ;
  assign n7353 = n7352 ^ n7351 ;
  assign n7354 = n7351 ^ n6462 ;
  assign n7355 = n7354 ^ n7351 ;
  assign n7356 = ~n7353 & ~n7355 ;
  assign n7357 = n7356 ^ n7351 ;
  assign n7358 = ~n6464 & n7357 ;
  assign n7368 = n7367 ^ n7358 ;
  assign n7341 = n6622 ^ n6577 ;
  assign n7342 = n7341 ^ n6564 ;
  assign n7343 = n7342 ^ n7067 ;
  assign n7344 = n6616 ^ n6584 ;
  assign n7347 = n7067 & ~n7344 ;
  assign n7348 = n7347 ^ n6616 ;
  assign n7349 = n7343 & n7348 ;
  assign n7369 = n7368 ^ n7349 ;
  assign n7370 = n7369 ^ n6620 ;
  assign n7371 = n7370 ^ n6649 ;
  assign n7372 = n7371 ^ n4985 ;
  assign n7340 = n6463 & n6592 ;
  assign n7373 = n7372 ^ n7340 ;
  assign n7374 = n7373 ^ x67 ;
  assign n7480 = ~n5979 & n6154 ;
  assign n7491 = n6173 ^ n6147 ;
  assign n7492 = n5976 & ~n6164 ;
  assign n7493 = n7491 & n7492 ;
  assign n7494 = n7493 ^ n6164 ;
  assign n7496 = n6137 ^ n6120 ;
  assign n7497 = n7496 ^ n6116 ;
  assign n7498 = ~n7494 & n7497 ;
  assign n7503 = n5979 & ~n6137 ;
  assign n7504 = n7498 & n7503 ;
  assign n7499 = n6129 ^ n6124 ;
  assign n7500 = n5978 & n7499 ;
  assign n7501 = n7500 ^ n7498 ;
  assign n7502 = n7501 ^ n7493 ;
  assign n7505 = n7504 ^ n7502 ;
  assign n7488 = n6126 ^ n6124 ;
  assign n7489 = n7488 ^ n6135 ;
  assign n7490 = n6192 & n7489 ;
  assign n7506 = n7505 ^ n7490 ;
  assign n7481 = n6114 ^ n6019 ;
  assign n7482 = n7481 ^ n6157 ;
  assign n7483 = n6157 ^ n5976 ;
  assign n7484 = n7483 ^ n6157 ;
  assign n7485 = ~n7482 & n7484 ;
  assign n7486 = n7485 ^ n6157 ;
  assign n7487 = ~n5977 & n7486 ;
  assign n7507 = n7506 ^ n7487 ;
  assign n7508 = n6138 ^ n6119 ;
  assign n7509 = n6138 ^ n5977 ;
  assign n7510 = n7509 ^ n6138 ;
  assign n7511 = ~n7508 & n7510 ;
  assign n7512 = n7511 ^ n6138 ;
  assign n7513 = ~n5976 & ~n7512 ;
  assign n7514 = ~n7507 & ~n7513 ;
  assign n7515 = ~n6195 & n7514 ;
  assign n7516 = ~n7480 & n7515 ;
  assign n7517 = ~n6191 & n7516 ;
  assign n7518 = n7517 ^ n5663 ;
  assign n7519 = n7518 ^ x116 ;
  assign n7566 = n5856 ^ n5837 ;
  assign n7548 = n5835 & ~n5838 ;
  assign n7563 = n7548 ^ n5849 ;
  assign n7564 = n7563 ^ n5873 ;
  assign n7565 = n7564 ^ n5849 ;
  assign n7567 = n7566 ^ n7565 ;
  assign n7568 = ~n5554 & n7567 ;
  assign n7569 = n7568 ^ n7563 ;
  assign n7570 = ~n5845 & n7569 ;
  assign n7549 = n7548 ^ n5865 ;
  assign n7550 = n7548 ^ n5394 ;
  assign n7551 = n7550 ^ n7548 ;
  assign n7552 = n7549 & n7551 ;
  assign n7553 = n7552 ^ n7548 ;
  assign n7554 = n5554 & n7553 ;
  assign n7542 = n5861 ^ n5839 ;
  assign n7543 = n5861 ^ n5554 ;
  assign n7544 = n7543 ^ n5861 ;
  assign n7545 = n7542 & n7544 ;
  assign n7546 = n7545 ^ n5861 ;
  assign n7547 = ~n5910 & n7546 ;
  assign n7555 = n7554 ^ n7547 ;
  assign n7522 = n5871 ^ n5869 ;
  assign n7520 = n5873 ^ n5863 ;
  assign n7521 = n7520 ^ n5854 ;
  assign n7523 = n7522 ^ n7521 ;
  assign n7524 = n5554 & n7523 ;
  assign n7525 = n7524 ^ n7520 ;
  assign n7556 = n7555 ^ n7525 ;
  assign n7534 = n5902 ^ n5842 ;
  assign n7535 = n5844 ^ n5839 ;
  assign n7538 = ~n5902 & ~n7535 ;
  assign n7539 = n7538 ^ n5844 ;
  assign n7540 = n7534 & n7539 ;
  assign n7541 = n7540 ^ n5842 ;
  assign n7557 = n7556 ^ n7541 ;
  assign n7558 = n7557 ^ n5893 ;
  assign n7559 = n7558 ^ n5920 ;
  assign n7560 = n7559 ^ n5926 ;
  assign n7561 = n7560 ^ n5067 ;
  assign n7526 = n7525 ^ n5839 ;
  assign n7527 = n7526 ^ n5863 ;
  assign n7528 = n7527 ^ n7525 ;
  assign n7531 = n5554 & n7528 ;
  assign n7532 = n7531 ^ n7525 ;
  assign n7533 = ~n5394 & n7532 ;
  assign n7562 = n7561 ^ n7533 ;
  assign n7571 = n7570 ^ n7562 ;
  assign n7572 = n7571 ^ x68 ;
  assign n7573 = n7519 & ~n7572 ;
  assign n7574 = n7573 ^ n7572 ;
  assign n7575 = n7574 ^ n7519 ;
  assign n7577 = n7575 ^ n7572 ;
  assign n7399 = ~n6757 & n6778 ;
  assign n7400 = n7399 ^ n6808 ;
  assign n7407 = n6789 & n6801 ;
  assign n7401 = n6785 ^ n6779 ;
  assign n7402 = n6779 ^ n6755 ;
  assign n7403 = n7402 ^ n6779 ;
  assign n7404 = n7401 & ~n7403 ;
  assign n7405 = n7404 ^ n6779 ;
  assign n7406 = n6754 & n7405 ;
  assign n7408 = n7407 ^ n7406 ;
  assign n7431 = n6756 & n6781 ;
  assign n7432 = n7431 ^ n6790 ;
  assign n7433 = n7432 ^ n6835 ;
  assign n7416 = n6782 ^ n6778 ;
  assign n7417 = n7416 ^ n6786 ;
  assign n7418 = n7417 ^ n6837 ;
  assign n7419 = n6754 & n7418 ;
  assign n7420 = n7419 ^ n6837 ;
  assign n7434 = n7433 ^ n7420 ;
  assign n7421 = n7420 ^ n6752 ;
  assign n7409 = n6836 ^ n6797 ;
  assign n7413 = n7409 ^ n6818 ;
  assign n7414 = n6754 & n7413 ;
  assign n7415 = n7414 ^ n7409 ;
  assign n7422 = n7421 ^ n7415 ;
  assign n7423 = n7422 ^ n6766 ;
  assign n7424 = n7423 ^ n6752 ;
  assign n7425 = n7424 ^ n7422 ;
  assign n7426 = n7422 ^ n6755 ;
  assign n7427 = n7426 ^ n7422 ;
  assign n7428 = n7425 & n7427 ;
  assign n7429 = n7428 ^ n7422 ;
  assign n7430 = n6793 & n7429 ;
  assign n7435 = n7434 ^ n7430 ;
  assign n7411 = n6781 ^ n6753 ;
  assign n7412 = ~n6757 & n7411 ;
  assign n7436 = n7435 ^ n7412 ;
  assign n7410 = n6758 & n7409 ;
  assign n7437 = n7436 ^ n7410 ;
  assign n7438 = n6756 ^ n6752 ;
  assign n7439 = n7438 ^ n7437 ;
  assign n7440 = n6796 ^ n6755 ;
  assign n7441 = ~n6756 & ~n7440 ;
  assign n7442 = n7441 ^ n6796 ;
  assign n7443 = n7439 & ~n7442 ;
  assign n7444 = n7443 ^ n6756 ;
  assign n7445 = ~n7437 & ~n7444 ;
  assign n7446 = ~n7408 & n7445 ;
  assign n7447 = ~n7400 & n7446 ;
  assign n7448 = ~n6780 & n7447 ;
  assign n7449 = n7448 ^ n5631 ;
  assign n7450 = n7449 ^ x102 ;
  assign n7456 = n7019 ^ n6972 ;
  assign n7457 = n7456 ^ n6990 ;
  assign n7458 = n7457 ^ n6997 ;
  assign n7459 = n6912 & n7458 ;
  assign n7460 = n7459 ^ n6997 ;
  assign n7464 = n7460 ^ n7015 ;
  assign n7465 = n7464 ^ n7026 ;
  assign n7454 = n6969 ^ n6948 ;
  assign n7455 = n7454 ^ n6960 ;
  assign n7461 = n7460 ^ n7455 ;
  assign n7452 = n6966 ^ n6943 ;
  assign n7453 = ~n6912 & n7452 ;
  assign n7462 = n7461 ^ n7453 ;
  assign n7463 = n6913 & ~n7462 ;
  assign n7466 = n7465 ^ n7463 ;
  assign n7451 = n6976 & n7014 ;
  assign n7467 = n7466 ^ n7451 ;
  assign n7468 = n6987 ^ n6962 ;
  assign n7469 = n6962 ^ n6913 ;
  assign n7470 = n7469 ^ n6962 ;
  assign n7471 = n7468 & n7470 ;
  assign n7472 = n7471 ^ n6962 ;
  assign n7473 = n7004 & n7472 ;
  assign n7474 = n7467 & ~n7473 ;
  assign n7475 = n7474 ^ n4580 ;
  assign n7476 = n7475 ^ x109 ;
  assign n7477 = n7450 & n7476 ;
  assign n7478 = n7477 ^ n7450 ;
  assign n7479 = n7478 ^ n7476 ;
  assign n7592 = n7479 ^ n7450 ;
  assign n7599 = n7577 & n7592 ;
  assign n7576 = ~n7479 & n7575 ;
  assign n7600 = n7599 ^ n7576 ;
  assign n7579 = ~n7479 & n7577 ;
  assign n7578 = n7477 & n7577 ;
  assign n7580 = n7579 ^ n7578 ;
  assign n7604 = n7600 ^ n7580 ;
  assign n7603 = n7577 ^ n7576 ;
  assign n7605 = n7604 ^ n7603 ;
  assign n7606 = n7605 ^ n7599 ;
  assign n7583 = n7478 & n7575 ;
  assign n7584 = n7583 ^ n7579 ;
  assign n7582 = n7477 & n7575 ;
  assign n7585 = n7584 ^ n7582 ;
  assign n7581 = n7580 ^ n7576 ;
  assign n7586 = n7585 ^ n7581 ;
  assign n7587 = n7586 ^ n7575 ;
  assign n7588 = n7587 ^ n7578 ;
  assign n7650 = n7606 ^ n7588 ;
  assign n7593 = ~n7574 & n7592 ;
  assign n7591 = n7478 & ~n7574 ;
  assign n7594 = n7593 ^ n7591 ;
  assign n7595 = n7594 ^ n7574 ;
  assign n9261 = n7650 ^ n7595 ;
  assign n7377 = n6416 ^ n6415 ;
  assign n7375 = n6423 & n6431 ;
  assign n7376 = n7375 ^ n6412 ;
  assign n7378 = n7377 ^ n7376 ;
  assign n7379 = n7378 ^ n6409 ;
  assign n7380 = n7379 ^ n6434 ;
  assign n7387 = n6420 ^ n6417 ;
  assign n7381 = n6395 & n6406 ;
  assign n7382 = n7381 ^ n6423 ;
  assign n7383 = n7382 ^ n7377 ;
  assign n7384 = n6233 & n7383 ;
  assign n7385 = n7384 ^ n7377 ;
  assign n7388 = n7387 ^ n7385 ;
  assign n7386 = n7385 ^ n7376 ;
  assign n7389 = n7388 ^ n7386 ;
  assign n7390 = n7388 ^ n6233 ;
  assign n7391 = n7390 ^ n7388 ;
  assign n7392 = n7389 & ~n7391 ;
  assign n7393 = n7392 ^ n7388 ;
  assign n7394 = ~n6253 & n7393 ;
  assign n7395 = n7394 ^ n7385 ;
  assign n7396 = ~n7380 & n7395 ;
  assign n7397 = n7396 ^ n4486 ;
  assign n7398 = n7397 ^ x85 ;
  assign n9262 = n7595 ^ n7398 ;
  assign n9263 = n9262 ^ n7595 ;
  assign n9264 = ~n9261 & n9263 ;
  assign n9265 = n9264 ^ n7595 ;
  assign n9266 = ~n7374 & ~n9265 ;
  assign n9232 = n7398 ^ n7374 ;
  assign n7596 = ~n7479 & n7573 ;
  assign n7607 = n7596 ^ n7593 ;
  assign n7608 = n7607 ^ n7606 ;
  assign n7601 = n7600 ^ n7584 ;
  assign n7602 = n7601 ^ n7476 ;
  assign n7609 = n7608 ^ n7602 ;
  assign n9238 = n7609 ^ n7580 ;
  assign n7611 = n7477 & ~n7574 ;
  assign n7610 = n7609 ^ n7574 ;
  assign n7612 = n7611 ^ n7610 ;
  assign n7598 = n7573 & n7592 ;
  assign n7613 = n7612 ^ n7598 ;
  assign n7597 = n7596 ^ n7573 ;
  assign n7614 = n7613 ^ n7597 ;
  assign n8445 = n7614 ^ n7612 ;
  assign n9233 = n8445 ^ n7609 ;
  assign n9234 = n8445 ^ n7374 ;
  assign n9235 = n9232 & n9234 ;
  assign n9236 = n9235 ^ n7374 ;
  assign n9237 = ~n9233 & ~n9236 ;
  assign n9239 = n9238 ^ n9237 ;
  assign n9240 = n9239 ^ n7398 ;
  assign n9241 = n9240 ^ n9239 ;
  assign n9242 = n9239 ^ n7613 ;
  assign n9243 = n9242 ^ n7608 ;
  assign n9244 = n9243 ^ n9239 ;
  assign n9245 = ~n9241 & n9244 ;
  assign n9246 = n9245 ^ n9239 ;
  assign n9247 = n9232 & ~n9246 ;
  assign n9248 = n9247 ^ n9239 ;
  assign n7621 = ~n7398 & n7583 ;
  assign n7589 = n7588 ^ n7398 ;
  assign n7590 = n7589 ^ n7588 ;
  assign n7615 = n7614 ^ n7595 ;
  assign n7616 = n7615 ^ n7611 ;
  assign n7617 = n7616 ^ n7588 ;
  assign n7618 = n7590 & ~n7617 ;
  assign n7619 = n7618 ^ n7588 ;
  assign n7620 = ~n7374 & n7619 ;
  assign n7622 = n7621 ^ n7620 ;
  assign n9249 = n9248 ^ n7622 ;
  assign n9231 = n7374 & n7582 ;
  assign n9252 = n9249 ^ n9231 ;
  assign n9267 = n9266 ^ n9252 ;
  assign n9253 = n9252 ^ n7622 ;
  assign n9254 = n9248 ^ n7398 ;
  assign n9255 = n7596 ^ n7583 ;
  assign n8440 = n7598 ^ n7576 ;
  assign n9256 = n9255 ^ n8440 ;
  assign n9257 = ~n7374 & n9256 ;
  assign n9258 = n9257 ^ n7596 ;
  assign n9259 = ~n9254 & n9258 ;
  assign n9260 = n9253 & n9259 ;
  assign n9268 = n9267 ^ n9260 ;
  assign n9269 = n9268 ^ n5764 ;
  assign n10117 = n9269 ^ x68 ;
  assign n7847 = n5377 ^ n4603 ;
  assign n7838 = n5299 ^ n5122 ;
  assign n7839 = n7838 ^ n5306 ;
  assign n7840 = n7839 ^ n5322 ;
  assign n7841 = n5297 & n7840 ;
  assign n7842 = n7841 ^ n5299 ;
  assign n7843 = n5314 ^ n5297 ;
  assign n7844 = n7842 & ~n7843 ;
  assign n7830 = n5352 ^ n5335 ;
  assign n7831 = n7830 ^ n5352 ;
  assign n7832 = n5354 & ~n7831 ;
  assign n7833 = n7832 ^ n5352 ;
  assign n7834 = ~n3798 & n7833 ;
  assign n7835 = n7834 ^ n5368 ;
  assign n7816 = n5342 ^ n5314 ;
  assign n7817 = n7816 ^ n5302 ;
  assign n7818 = n5291 & ~n7817 ;
  assign n7819 = n7818 ^ n5124 ;
  assign n7828 = n7819 ^ n5291 ;
  assign n7829 = n3798 & n7828 ;
  assign n7836 = n7835 ^ n7829 ;
  assign n7822 = n5376 ^ n5119 ;
  assign n7823 = n7822 ^ n5355 ;
  assign n7824 = n7823 ^ n5317 ;
  assign n7825 = n3798 & ~n7824 ;
  assign n7820 = n7819 ^ n5376 ;
  assign n7821 = n7820 ^ n5355 ;
  assign n7826 = n7825 ^ n7821 ;
  assign n7827 = ~n5291 & ~n7826 ;
  assign n7837 = n7836 ^ n7827 ;
  assign n7845 = n7844 ^ n7837 ;
  assign n7846 = ~n7287 & n7845 ;
  assign n7848 = n7847 ^ n7846 ;
  assign n8851 = n7848 ^ x73 ;
  assign n8852 = n7475 ^ x66 ;
  assign n8853 = ~n8851 & n8852 ;
  assign n8854 = n8853 ^ n8851 ;
  assign n8855 = n8854 ^ n8852 ;
  assign n8856 = n7397 ^ x107 ;
  assign n7699 = n5858 ^ n5854 ;
  assign n7694 = n5902 ^ n5861 ;
  assign n7691 = n5912 ^ n5863 ;
  assign n7692 = n7691 ^ n5895 ;
  assign n7693 = n7692 ^ n7548 ;
  assign n7695 = n7694 ^ n7693 ;
  assign n7696 = n7695 ^ n5895 ;
  assign n7697 = ~n5554 & n7696 ;
  assign n7698 = n7697 ^ n7692 ;
  assign n7700 = n7699 ^ n7698 ;
  assign n7701 = n5845 & n7700 ;
  assign n7689 = n5872 ^ n5849 ;
  assign n7690 = n5842 & n7689 ;
  assign n7702 = n7701 ^ n7690 ;
  assign n7704 = n5871 ^ n5848 ;
  assign n7705 = n7704 ^ n5858 ;
  assign n7706 = n7705 ^ n7694 ;
  assign n7707 = ~n5554 & n7706 ;
  assign n7703 = n5886 ^ n5852 ;
  assign n7708 = n7707 ^ n7703 ;
  assign n7709 = ~n5845 & ~n7708 ;
  assign n7710 = ~n5852 & n7709 ;
  assign n7711 = n7710 ^ n5845 ;
  assign n7712 = ~n7702 & n7711 ;
  assign n7713 = n7712 ^ n5841 ;
  assign n7714 = ~n5924 & n7713 ;
  assign n7717 = n5837 ^ n5554 ;
  assign n7718 = n7717 ^ n5837 ;
  assign n7719 = n7566 & n7718 ;
  assign n7720 = n7719 ^ n5837 ;
  assign n7721 = ~n5845 & n7720 ;
  assign n7722 = ~n7554 & ~n7721 ;
  assign n7723 = n7714 & n7722 ;
  assign n7724 = n7723 ^ n4415 ;
  assign n8857 = n7724 ^ x105 ;
  assign n8858 = ~n8856 & n8857 ;
  assign n7729 = n7165 & n7208 ;
  assign n8887 = n7729 ^ n4463 ;
  assign n7771 = n7194 ^ n7185 ;
  assign n7772 = n7208 & ~n7771 ;
  assign n8888 = n8887 ^ n7772 ;
  assign n8874 = n7771 ^ n7175 ;
  assign n8875 = n8874 ^ n7152 ;
  assign n8876 = ~n7086 & ~n8875 ;
  assign n8877 = n8876 ^ n7158 ;
  assign n8878 = ~n7199 & n8877 ;
  assign n8879 = n8878 ^ n7158 ;
  assign n8867 = n7193 ^ n7166 ;
  assign n8868 = n8867 ^ n7169 ;
  assign n8871 = ~n7199 & n8868 ;
  assign n8872 = n8871 ^ n7169 ;
  assign n8873 = n7086 & n8872 ;
  assign n8880 = n8879 ^ n8873 ;
  assign n8881 = n8880 ^ n7162 ;
  assign n7979 = n7197 ^ n7190 ;
  assign n7980 = n7190 ^ n7086 ;
  assign n7981 = n7980 ^ n7190 ;
  assign n7982 = ~n7979 & ~n7981 ;
  assign n7983 = n7982 ^ n7190 ;
  assign n7984 = n7199 & n7983 ;
  assign n8882 = n8881 ^ n7984 ;
  assign n7731 = n7172 ^ n7168 ;
  assign n7732 = n7731 ^ n7185 ;
  assign n7733 = n7086 & n7732 ;
  assign n7734 = n7733 ^ n7168 ;
  assign n7735 = n7734 ^ n7177 ;
  assign n7736 = n7735 ^ n7734 ;
  assign n7739 = n7086 & n7736 ;
  assign n7740 = n7739 ^ n7734 ;
  assign n7741 = n7212 & n7740 ;
  assign n7742 = n7741 ^ n7734 ;
  assign n8883 = n8882 ^ n7742 ;
  assign n7765 = n7197 ^ n7194 ;
  assign n7766 = n7194 ^ n7086 ;
  assign n7767 = n7766 ^ n7194 ;
  assign n7768 = n7765 & ~n7767 ;
  assign n7769 = n7768 ^ n7194 ;
  assign n7770 = ~n7199 & ~n7769 ;
  assign n8884 = n8883 ^ n7770 ;
  assign n8860 = n7162 ^ n7086 ;
  assign n8861 = n8860 ^ n7162 ;
  assign n8864 = n7191 & ~n8861 ;
  assign n8865 = n8864 ^ n7162 ;
  assign n8866 = n7212 & n8865 ;
  assign n8885 = n8884 ^ n8866 ;
  assign n8886 = ~n7204 & ~n8885 ;
  assign n8889 = n8888 ^ n8886 ;
  assign n8890 = n8889 ^ x80 ;
  assign n8936 = n8858 & ~n8890 ;
  assign n8898 = n7342 ^ n6602 ;
  assign n8897 = n7074 ^ n6622 ;
  assign n8899 = n8898 ^ n8897 ;
  assign n8900 = n8897 ^ n6462 ;
  assign n8901 = ~n6464 & ~n8900 ;
  assign n8902 = n8901 ^ n6462 ;
  assign n8903 = n8899 & ~n8902 ;
  assign n8904 = n8903 ^ n8897 ;
  assign n8905 = n8904 ^ n6585 ;
  assign n8906 = n8905 ^ n6576 ;
  assign n8892 = n7076 ^ n6600 ;
  assign n8891 = n7341 ^ n6589 ;
  assign n8893 = n8892 ^ n8891 ;
  assign n8894 = n8893 ^ n6619 ;
  assign n8895 = n6463 & ~n8894 ;
  assign n8896 = n8895 ^ n8892 ;
  assign n8907 = n8906 ^ n8896 ;
  assign n8913 = n8907 ^ n6580 ;
  assign n8914 = n8913 ^ n8907 ;
  assign n8915 = n8907 ^ n6462 ;
  assign n8916 = n8915 ^ n8907 ;
  assign n8917 = ~n8914 & ~n8916 ;
  assign n8918 = ~n8906 & n8917 ;
  assign n8919 = n8918 ^ n8906 ;
  assign n8920 = n8919 ^ n8896 ;
  assign n8921 = n6464 & n8920 ;
  assign n8922 = n8921 ^ n8896 ;
  assign n8923 = ~n7364 & ~n8922 ;
  assign n8924 = ~n7055 & n8923 ;
  assign n8925 = ~n7066 & n8924 ;
  assign n8926 = ~n7072 & n8925 ;
  assign n8927 = n8926 ^ n6620 ;
  assign n8928 = n8927 ^ n4539 ;
  assign n8929 = n8928 ^ x90 ;
  assign n8930 = n8890 & n8929 ;
  assign n8933 = n8930 ^ n8929 ;
  assign n8934 = n8933 ^ n8890 ;
  assign n8935 = n8858 & ~n8934 ;
  assign n8937 = n8936 ^ n8935 ;
  assign n8859 = n8858 ^ n8856 ;
  assign n8931 = n8930 ^ n8890 ;
  assign n8932 = ~n8859 & n8931 ;
  assign n8938 = n8937 ^ n8932 ;
  assign n8939 = n8855 & n8938 ;
  assign n10144 = n8939 ^ n5833 ;
  assign n8962 = n8858 ^ n8857 ;
  assign n8968 = ~n8934 & n8962 ;
  assign n8969 = n8968 ^ n8934 ;
  assign n8945 = ~n8859 & ~n8934 ;
  assign n8946 = n8945 ^ n8935 ;
  assign n8970 = n8969 ^ n8946 ;
  assign n8963 = n8962 ^ n8856 ;
  assign n8964 = n8931 & n8963 ;
  assign n8971 = n8970 ^ n8964 ;
  assign n8966 = n8933 & n8963 ;
  assign n8967 = n8966 ^ n8963 ;
  assign n8972 = n8971 ^ n8967 ;
  assign n8949 = n8936 ^ n8858 ;
  assign n8947 = n8858 & n8930 ;
  assign n8950 = n8949 ^ n8947 ;
  assign n8951 = n8950 ^ n8937 ;
  assign n8940 = ~n8859 & n8930 ;
  assign n8952 = n8951 ^ n8940 ;
  assign n8948 = n8947 ^ n8946 ;
  assign n8953 = n8952 ^ n8948 ;
  assign n8944 = n8932 ^ n8856 ;
  assign n8954 = n8953 ^ n8944 ;
  assign n9371 = n8972 ^ n8954 ;
  assign n9372 = n8954 ^ n8852 ;
  assign n9373 = n9372 ^ n8954 ;
  assign n9374 = n9371 & ~n9373 ;
  assign n9375 = n9374 ^ n8954 ;
  assign n9376 = n8851 & ~n9375 ;
  assign n10145 = n10144 ^ n9376 ;
  assign n9005 = n8950 ^ n8932 ;
  assign n9006 = n8853 & n9005 ;
  assign n8988 = n8930 & n8962 ;
  assign n8985 = n8968 ^ n8966 ;
  assign n9744 = n8988 ^ n8985 ;
  assign n10139 = n9744 ^ n8972 ;
  assign n10140 = ~n8854 & ~n10139 ;
  assign n8996 = n8852 ^ n8851 ;
  assign n8942 = n8855 ^ n8851 ;
  assign n9736 = ~n8942 & ~n8946 ;
  assign n10126 = n8948 ^ n8940 ;
  assign n10127 = ~n9736 & n10126 ;
  assign n10128 = n10127 ^ n8951 ;
  assign n10125 = n8854 & n8936 ;
  assign n10129 = n10128 ^ n10125 ;
  assign n8941 = n8940 ^ n8935 ;
  assign n9350 = n8966 ^ n8941 ;
  assign n10130 = n10129 ^ n9350 ;
  assign n8955 = n8954 ^ n8937 ;
  assign n8974 = n8955 ^ n8933 ;
  assign n8975 = n8974 ^ n8966 ;
  assign n8989 = n8988 ^ n8975 ;
  assign n8990 = n8989 ^ n8964 ;
  assign n8991 = n8990 ^ n8856 ;
  assign n8986 = n8972 ^ n8970 ;
  assign n8987 = n8986 ^ n8985 ;
  assign n8992 = n8991 ^ n8987 ;
  assign n9358 = n8992 ^ n8970 ;
  assign n9750 = n9358 ^ n8975 ;
  assign n10131 = n10130 ^ n9750 ;
  assign n10132 = n10131 ^ n10129 ;
  assign n10133 = n10129 ^ n8852 ;
  assign n10134 = n10133 ^ n10129 ;
  assign n10135 = ~n10132 & n10134 ;
  assign n10136 = n10135 ^ n10129 ;
  assign n10137 = n8996 & n10136 ;
  assign n10138 = n10137 ^ n10129 ;
  assign n10141 = n10140 ^ n10138 ;
  assign n9355 = n8989 ^ n8954 ;
  assign n9356 = n9355 ^ n8935 ;
  assign n10118 = n9356 ^ n8970 ;
  assign n10119 = n10118 ^ n8990 ;
  assign n10120 = n8990 ^ n8852 ;
  assign n10121 = n10120 ^ n8990 ;
  assign n10122 = n10119 & ~n10121 ;
  assign n10123 = n10122 ^ n8990 ;
  assign n10124 = n8851 & ~n10123 ;
  assign n10142 = n10141 ^ n10124 ;
  assign n10143 = ~n9006 & ~n10142 ;
  assign n10146 = n10145 ^ n10143 ;
  assign n10147 = n10146 ^ x126 ;
  assign n10148 = ~n10117 & n10147 ;
  assign n10149 = n10148 ^ n10117 ;
  assign n8230 = n7380 ^ n6253 ;
  assign n8231 = n8230 ^ n7380 ;
  assign n8232 = n7382 & n8231 ;
  assign n8233 = n8232 ^ n7380 ;
  assign n8234 = ~n6233 & n8233 ;
  assign n8216 = ~n6253 & n7378 ;
  assign n8217 = n8216 ^ n7377 ;
  assign n8222 = n8217 ^ n7387 ;
  assign n8223 = n8222 ^ n8217 ;
  assign n8224 = ~n6253 & n8223 ;
  assign n8225 = n8224 ^ n8217 ;
  assign n8226 = ~n6233 & ~n8225 ;
  assign n8218 = n8217 ^ n7380 ;
  assign n8219 = n8218 ^ n4806 ;
  assign n8227 = n8226 ^ n8219 ;
  assign n8235 = n8234 ^ n8227 ;
  assign n8236 = n8235 ^ x82 ;
  assign n8247 = n5863 ^ n5854 ;
  assign n8240 = n7522 ^ n5864 ;
  assign n8241 = ~n5554 & n8240 ;
  assign n8242 = n8241 ^ n5871 ;
  assign n8246 = n8242 ^ n7689 ;
  assign n8248 = n8247 ^ n8246 ;
  assign n8249 = n8248 ^ n8242 ;
  assign n8250 = ~n5554 & n8249 ;
  assign n8251 = n8250 ^ n8246 ;
  assign n8252 = ~n5394 & n8251 ;
  assign n8244 = n5554 & n5912 ;
  assign n8237 = n5912 ^ n5854 ;
  assign n8238 = n8237 ^ n5895 ;
  assign n8239 = n5394 & n8238 ;
  assign n8243 = n8242 ^ n8239 ;
  assign n8245 = n8244 ^ n8243 ;
  assign n8253 = n8252 ^ n8245 ;
  assign n8254 = n8253 ^ n5922 ;
  assign n8255 = n8254 ^ n7721 ;
  assign n8256 = n8255 ^ n7555 ;
  assign n8257 = n8256 ^ n7541 ;
  assign n8258 = n8257 ^ n5908 ;
  assign n8259 = ~n5926 & ~n8258 ;
  assign n8260 = n8259 ^ n4785 ;
  assign n8261 = n8260 ^ x81 ;
  assign n8262 = n8236 & n8261 ;
  assign n8263 = n8262 ^ n8236 ;
  assign n7660 = ~n6142 & ~n6194 ;
  assign n7683 = n7480 ^ n6122 ;
  assign n7662 = n7488 ^ n5976 ;
  assign n7664 = n6132 ^ n6120 ;
  assign n7665 = n7664 ^ n6146 ;
  assign n7666 = n7665 ^ n6157 ;
  assign n7667 = ~n5977 & ~n7666 ;
  assign n7663 = n7496 ^ n5976 ;
  assign n7668 = n7667 ^ n7663 ;
  assign n7669 = n7662 & n7668 ;
  assign n7670 = n7669 ^ n5976 ;
  assign n7672 = n6172 ^ n6128 ;
  assign n7671 = n6129 ^ n6125 ;
  assign n7673 = n7672 ^ n7671 ;
  assign n7674 = n7671 ^ n5977 ;
  assign n7675 = n7674 ^ n7671 ;
  assign n7676 = ~n7673 & n7675 ;
  assign n7677 = n7676 ^ n7671 ;
  assign n7678 = n6164 & n7677 ;
  assign n7679 = n7678 ^ n7671 ;
  assign n7680 = ~n7670 & ~n7679 ;
  assign n7661 = n6116 & n6192 ;
  assign n7681 = n7680 ^ n7661 ;
  assign n7682 = ~n7513 & n7681 ;
  assign n7684 = n7683 ^ n7682 ;
  assign n7685 = ~n6191 & n7684 ;
  assign n7686 = n7660 & n7685 ;
  assign n7687 = n7686 ^ n4743 ;
  assign n8265 = n7687 ^ x120 ;
  assign n8266 = n7033 ^ x64 ;
  assign n8267 = n8265 & n8266 ;
  assign n8283 = n8263 & n8267 ;
  assign n8269 = n7084 ^ x114 ;
  assign n7730 = ~n7248 & ~n7729 ;
  assign n7773 = n7772 ^ n7770 ;
  assign n7756 = n7173 ^ n7152 ;
  assign n7753 = n7195 ^ n7182 ;
  assign n7757 = n7756 ^ n7753 ;
  assign n7751 = n7190 ^ n7179 ;
  assign n7752 = n7751 ^ n7156 ;
  assign n7754 = n7753 ^ n7752 ;
  assign n7755 = ~n7086 & ~n7754 ;
  assign n7758 = n7757 ^ n7755 ;
  assign n7759 = ~n7212 & ~n7758 ;
  assign n7760 = n7759 ^ n7152 ;
  assign n7749 = n7197 ^ n7164 ;
  assign n7750 = n7205 & ~n7749 ;
  assign n7761 = n7760 ^ n7750 ;
  assign n7762 = ~n7232 & ~n7761 ;
  assign n7743 = n7172 ^ n7086 ;
  assign n7744 = n7743 ^ n7172 ;
  assign n7745 = n7731 ^ n7172 ;
  assign n7746 = ~n7744 & n7745 ;
  assign n7747 = n7746 ^ n7172 ;
  assign n7748 = n7212 & n7747 ;
  assign n7763 = n7762 ^ n7748 ;
  assign n7764 = ~n7742 & n7763 ;
  assign n7774 = n7773 ^ n7764 ;
  assign n7775 = n7730 & n7774 ;
  assign n7776 = n7775 ^ n4838 ;
  assign n8275 = n7776 ^ x88 ;
  assign n8281 = ~n8269 & n8275 ;
  assign n8303 = n8281 ^ n8275 ;
  assign n8324 = n8303 ^ n8269 ;
  assign n8325 = n8283 & n8324 ;
  assign n8276 = n8275 ^ n8269 ;
  assign n8271 = n8267 ^ n8266 ;
  assign n8272 = n8271 ^ n8265 ;
  assign n8264 = n8263 ^ n8261 ;
  assign n8279 = n8264 ^ n8236 ;
  assign n8290 = ~n8272 & n8279 ;
  assign n8291 = n8290 ^ n8272 ;
  assign n8288 = n8263 & ~n8272 ;
  assign n8287 = n8262 & ~n8272 ;
  assign n8289 = n8288 ^ n8287 ;
  assign n8292 = n8291 ^ n8289 ;
  assign n8273 = n8272 ^ n8266 ;
  assign n8274 = n8263 & n8273 ;
  assign n8293 = n8292 ^ n8274 ;
  assign n8284 = n8273 & n8279 ;
  assign n8309 = n8293 ^ n8284 ;
  assign n8310 = n8309 ^ n8273 ;
  assign n8299 = n8262 & n8273 ;
  assign n8308 = n8299 ^ n8292 ;
  assign n8311 = n8310 ^ n8308 ;
  assign n8268 = ~n8264 & n8267 ;
  assign n8312 = n8311 ^ n8268 ;
  assign n8307 = n8292 ^ n8264 ;
  assign n8313 = n8312 ^ n8307 ;
  assign n8318 = n8313 ^ n8271 ;
  assign n8304 = n8262 & n8271 ;
  assign n8297 = n8271 & n8279 ;
  assign n8317 = n8304 ^ n8297 ;
  assign n8319 = n8318 ^ n8317 ;
  assign n8320 = n8276 & n8319 ;
  assign n8296 = n8292 ^ n8287 ;
  assign n8298 = n8297 ^ n8296 ;
  assign n8321 = n8320 ^ n8298 ;
  assign n8314 = n8313 ^ n8288 ;
  assign n8305 = n8304 ^ n8290 ;
  assign n8306 = n8305 ^ n8284 ;
  assign n8315 = n8314 ^ n8306 ;
  assign n8316 = n8303 & n8315 ;
  assign n8322 = n8321 ^ n8316 ;
  assign n8300 = n8299 ^ n8298 ;
  assign n8285 = n8284 ^ n8283 ;
  assign n8286 = n8285 ^ n8268 ;
  assign n8294 = n8293 ^ n8286 ;
  assign n8295 = ~n8275 & ~n8294 ;
  assign n8301 = n8300 ^ n8295 ;
  assign n8302 = ~n8276 & ~n8301 ;
  assign n8323 = n8322 ^ n8302 ;
  assign n8326 = n8325 ^ n8323 ;
  assign n8280 = n8267 & n8279 ;
  assign n8282 = n8280 & n8281 ;
  assign n8327 = n8326 ^ n8282 ;
  assign n8277 = n8274 & n8276 ;
  assign n8270 = n8268 & n8269 ;
  assign n8278 = n8277 ^ n8270 ;
  assign n8328 = n8327 ^ n8278 ;
  assign n8329 = n8262 & n8267 ;
  assign n8336 = n8303 & n8329 ;
  assign n8330 = n8329 ^ n8305 ;
  assign n8331 = n8305 ^ n8269 ;
  assign n8332 = n8331 ^ n8305 ;
  assign n8333 = n8330 & n8332 ;
  assign n8334 = n8333 ^ n8305 ;
  assign n8335 = ~n8275 & n8334 ;
  assign n8337 = n8336 ^ n8335 ;
  assign n8338 = n8329 ^ n8311 ;
  assign n8339 = n8281 & n8338 ;
  assign n8340 = ~n8337 & ~n8339 ;
  assign n8341 = n8328 & n8340 ;
  assign n8342 = n8341 ^ n5795 ;
  assign n10082 = n8342 ^ x124 ;
  assign n8480 = n5317 ^ n5301 ;
  assign n8481 = n8480 ^ n5335 ;
  assign n8479 = n5316 ^ n5124 ;
  assign n8482 = n8481 ^ n8479 ;
  assign n8483 = n8481 ^ n5291 ;
  assign n8484 = n8483 ^ n8481 ;
  assign n8485 = n8482 & n8484 ;
  assign n8486 = n8485 ^ n8481 ;
  assign n8487 = ~n3798 & n8486 ;
  assign n8471 = n5376 ^ n5311 ;
  assign n8472 = n8471 ^ n5324 ;
  assign n8473 = n8472 ^ n5311 ;
  assign n8474 = n5311 ^ n5291 ;
  assign n8475 = n8474 ^ n5311 ;
  assign n8476 = n8473 & n8475 ;
  assign n8477 = n8476 ^ n5311 ;
  assign n8478 = ~n5337 & n8477 ;
  assign n8488 = n8487 ^ n8478 ;
  assign n8489 = n8488 ^ n5310 ;
  assign n8490 = n8489 ^ n7834 ;
  assign n8491 = n8490 ^ n5331 ;
  assign n8463 = n7816 ^ n5337 ;
  assign n8464 = n7816 ^ n5310 ;
  assign n8465 = n8464 ^ n5310 ;
  assign n8466 = n5310 ^ n5291 ;
  assign n8467 = n8466 ^ n5310 ;
  assign n8468 = ~n8465 & ~n8467 ;
  assign n8469 = n8468 ^ n5310 ;
  assign n8470 = n8463 & n8469 ;
  assign n8492 = n8491 ^ n8470 ;
  assign n8493 = n8492 ^ n7287 ;
  assign n8494 = n8493 ^ n5373 ;
  assign n8495 = n8494 ^ n5377 ;
  assign n8496 = n8495 ^ n4954 ;
  assign n8497 = n8496 ^ x117 ;
  assign n8499 = n6436 ^ n6233 ;
  assign n8500 = n8499 ^ n6439 ;
  assign n8501 = n8500 ^ n6411 ;
  assign n8502 = n8501 ^ n4926 ;
  assign n8503 = n8502 ^ x92 ;
  assign n8504 = n8497 & n8503 ;
  assign n8512 = n8504 ^ n8503 ;
  assign n8462 = n7373 ^ x69 ;
  assign n7999 = ~n7197 & ~n7212 ;
  assign n7992 = n7753 ^ n7179 ;
  assign n7990 = n7242 ^ n7184 ;
  assign n7985 = n7086 & n7188 ;
  assign n7986 = n7985 ^ n7181 ;
  assign n7991 = n7990 ^ n7986 ;
  assign n7993 = n7992 ^ n7991 ;
  assign n7994 = n7993 ^ n7986 ;
  assign n7995 = n7086 & ~n7994 ;
  assign n7996 = n7995 ^ n7991 ;
  assign n7997 = ~n7199 & n7996 ;
  assign n7987 = n7986 ^ n7748 ;
  assign n7988 = n7987 ^ n7984 ;
  assign n7989 = n7988 ^ n7240 ;
  assign n7998 = n7997 ^ n7989 ;
  assign n8000 = n7999 ^ n7998 ;
  assign n8001 = n7730 & ~n8000 ;
  assign n8002 = n8001 ^ n3968 ;
  assign n8507 = n8002 ^ x110 ;
  assign n8510 = n8462 & ~n8507 ;
  assign n8514 = n8510 ^ n8462 ;
  assign n8515 = n8514 ^ n8507 ;
  assign n8516 = n8515 ^ n8462 ;
  assign n8540 = n8512 & ~n8516 ;
  assign n8518 = n8504 & n8510 ;
  assign n8541 = n8540 ^ n8518 ;
  assign n8505 = n8504 ^ n8497 ;
  assign n8517 = n8505 & ~n8516 ;
  assign n8519 = n8518 ^ n8517 ;
  assign n8513 = n8510 & n8512 ;
  assign n8520 = n8519 ^ n8513 ;
  assign n8506 = n8505 ^ n8503 ;
  assign n8511 = ~n8506 & n8510 ;
  assign n8521 = n8520 ^ n8511 ;
  assign n8524 = n8521 ^ n8510 ;
  assign n8525 = n8524 ^ n8517 ;
  assign n8498 = n8497 ^ n8462 ;
  assign n8523 = ~n8498 & ~n8507 ;
  assign n8526 = n8525 ^ n8523 ;
  assign n8542 = n8541 ^ n8526 ;
  assign n7872 = n6781 & ~n6793 ;
  assign n8109 = n7872 ^ n4121 ;
  assign n8098 = n6801 & ~n7415 ;
  assign n8096 = n6794 ^ n6766 ;
  assign n8094 = n7415 ^ n6796 ;
  assign n8095 = n8094 ^ n6778 ;
  assign n8097 = n8096 ^ n8095 ;
  assign n8099 = n8098 ^ n8097 ;
  assign n8100 = ~n6793 & n8099 ;
  assign n8101 = n8100 ^ n8094 ;
  assign n8087 = n6796 ^ n6785 ;
  assign n8088 = n8087 ^ n6795 ;
  assign n8089 = n8087 ^ n6755 ;
  assign n8090 = n8089 ^ n8087 ;
  assign n8091 = n8088 & ~n8090 ;
  assign n8092 = n8091 ^ n8087 ;
  assign n8093 = ~n6754 & n8092 ;
  assign n8102 = n8101 ^ n8093 ;
  assign n7852 = n6796 ^ n6752 ;
  assign n8080 = n7852 ^ n6783 ;
  assign n8081 = n6783 ^ n6754 ;
  assign n8082 = n8081 ^ n6783 ;
  assign n8083 = ~n8080 & n8082 ;
  assign n8084 = n8083 ^ n6783 ;
  assign n8085 = n6755 & ~n8084 ;
  assign n8103 = n8102 ^ n8085 ;
  assign n8104 = n8103 ^ n6753 ;
  assign n8105 = n8104 ^ n7406 ;
  assign n8077 = ~n6755 & ~n7416 ;
  assign n8078 = n8077 ^ n6753 ;
  assign n8079 = n6754 & n8078 ;
  assign n8106 = n8105 ^ n8079 ;
  assign n8107 = ~n7432 & ~n8106 ;
  assign n8108 = ~n6759 & n8107 ;
  assign n8110 = n8109 ^ n8108 ;
  assign n8461 = n8110 ^ x83 ;
  assign n8532 = n7571 ^ x78 ;
  assign n8559 = n8461 & ~n8532 ;
  assign n8560 = n8559 ^ n8532 ;
  assign n8585 = n8542 & ~n8560 ;
  assign n8552 = n8532 ^ n8461 ;
  assign n9608 = n8540 ^ n8526 ;
  assign n9068 = n8504 & n8515 ;
  assign n9609 = n9608 ^ n9068 ;
  assign n9610 = n9068 ^ n8461 ;
  assign n9611 = n9610 ^ n9068 ;
  assign n9612 = n9609 & ~n9611 ;
  assign n9613 = n9612 ^ n9068 ;
  assign n9614 = n8552 & n9613 ;
  assign n9055 = n8540 ^ n8511 ;
  assign n9053 = n8512 & n8514 ;
  assign n9054 = n9053 ^ n8540 ;
  assign n9056 = n9055 ^ n9054 ;
  assign n9057 = n9055 ^ n8461 ;
  assign n9058 = n9057 ^ n9055 ;
  assign n9059 = n9056 & n9058 ;
  assign n9060 = n9059 ^ n9055 ;
  assign n9061 = n8552 & n9060 ;
  assign n9062 = n9061 ^ n8540 ;
  assign n8566 = ~n8506 & n8515 ;
  assign n8554 = n8505 & n8514 ;
  assign n8567 = n8566 ^ n8554 ;
  assign n8562 = n8505 & n8515 ;
  assign n8538 = n8504 & n8514 ;
  assign n8565 = n8562 ^ n8538 ;
  assign n8568 = n8567 ^ n8565 ;
  assign n8569 = n8567 ^ n8461 ;
  assign n8570 = n8569 ^ n8567 ;
  assign n8571 = n8568 & n8570 ;
  assign n8572 = n8571 ^ n8567 ;
  assign n8573 = n8532 & n8572 ;
  assign n10108 = n8511 & ~n8552 ;
  assign n8527 = n8526 ^ n8516 ;
  assign n8528 = n8527 ^ n8519 ;
  assign n8529 = n8528 ^ n8525 ;
  assign n10101 = n8562 ^ n8529 ;
  assign n10102 = n10101 ^ n9053 ;
  assign n10103 = n8532 & ~n10102 ;
  assign n10100 = n8554 ^ n8525 ;
  assign n10104 = n10103 ^ n10100 ;
  assign n10105 = ~n8461 & n10104 ;
  assign n8508 = n8507 ^ n8506 ;
  assign n8509 = ~n8498 & ~n8508 ;
  assign n8522 = n8521 ^ n8509 ;
  assign n8555 = n8554 ^ n8522 ;
  assign n8543 = n8542 ^ n8520 ;
  assign n8539 = n8538 ^ n8511 ;
  assign n8544 = n8543 ^ n8539 ;
  assign n8556 = n8555 ^ n8544 ;
  assign n8553 = ~n8506 & n8514 ;
  assign n8557 = n8556 ^ n8553 ;
  assign n10085 = n8557 ^ n8538 ;
  assign n10086 = n10085 ^ n9068 ;
  assign n10084 = n8540 ^ n8520 ;
  assign n10087 = n10086 ^ n10084 ;
  assign n10088 = n8461 & n10087 ;
  assign n10089 = n10088 ^ n10086 ;
  assign n10098 = n10089 ^ n8554 ;
  assign n9592 = n9068 ^ n8513 ;
  assign n10090 = n10089 ^ n9592 ;
  assign n10091 = n10090 ^ n8553 ;
  assign n10092 = n10091 ^ n10089 ;
  assign n10095 = n8461 & n10092 ;
  assign n10096 = n10095 ^ n10089 ;
  assign n10097 = n8532 & n10096 ;
  assign n10099 = n10098 ^ n10097 ;
  assign n10106 = n10105 ^ n10099 ;
  assign n10083 = n8559 & n8566 ;
  assign n10107 = n10106 ^ n10083 ;
  assign n10109 = n10108 ^ n10107 ;
  assign n10110 = ~n8573 & ~n10109 ;
  assign n10111 = ~n9062 & n10110 ;
  assign n10112 = ~n9614 & n10111 ;
  assign n10113 = ~n8585 & n10112 ;
  assign n10114 = n10113 ^ n5603 ;
  assign n10115 = n10114 ^ x78 ;
  assign n10116 = n10082 & ~n10115 ;
  assign n10150 = n10116 ^ n10115 ;
  assign n10155 = ~n10149 & ~n10150 ;
  assign n10154 = n10116 & n10148 ;
  assign n10156 = n10155 ^ n10154 ;
  assign n10440 = ~n10081 & n10156 ;
  assign n10151 = n10150 ^ n10082 ;
  assign n10152 = n10151 ^ n10115 ;
  assign n10153 = ~n10149 & n10152 ;
  assign n10443 = n10153 ^ n10080 ;
  assign n10160 = n10149 ^ n10147 ;
  assign n10161 = n10160 ^ n10117 ;
  assign n10179 = n10151 & n10161 ;
  assign n10170 = n10147 ^ n10117 ;
  assign n10171 = n10117 ^ n10115 ;
  assign n10172 = ~n10170 & ~n10171 ;
  assign n10176 = n10172 ^ n10161 ;
  assign n10177 = n10176 ^ n10155 ;
  assign n10162 = n10116 & n10161 ;
  assign n10157 = n10156 ^ n10153 ;
  assign n10158 = n10157 ^ n10117 ;
  assign n10159 = n10116 & ~n10158 ;
  assign n10163 = n10162 ^ n10159 ;
  assign n10178 = n10177 ^ n10163 ;
  assign n10180 = n10179 ^ n10178 ;
  assign n10181 = n10180 ^ n10162 ;
  assign n10191 = n10181 ^ n10161 ;
  assign n10164 = n10163 ^ n10154 ;
  assign n10165 = n10164 ^ n10116 ;
  assign n10189 = n10165 ^ n10160 ;
  assign n10187 = n10152 & n10160 ;
  assign n10186 = ~n10150 & n10160 ;
  assign n10188 = n10187 ^ n10186 ;
  assign n10190 = n10189 ^ n10188 ;
  assign n10192 = n10191 ^ n10190 ;
  assign n10193 = n10192 ^ n10178 ;
  assign n10185 = n10148 & ~n10150 ;
  assign n10194 = n10193 ^ n10185 ;
  assign n10183 = n10159 ^ n10155 ;
  assign n10184 = n10183 ^ n10153 ;
  assign n10195 = n10194 ^ n10184 ;
  assign n10196 = n10195 ^ n10188 ;
  assign n10168 = n10117 ^ n10082 ;
  assign n10169 = n10168 ^ n10147 ;
  assign n10173 = n10172 ^ n10160 ;
  assign n10174 = ~n10169 & ~n10173 ;
  assign n10175 = n10174 ^ n10165 ;
  assign n10182 = n10181 ^ n10175 ;
  assign n10197 = n10196 ^ n10182 ;
  assign n10444 = n10197 ^ n10077 ;
  assign n10447 = ~n10153 & ~n10444 ;
  assign n10448 = n10447 ^ n10077 ;
  assign n10449 = n10443 & ~n10448 ;
  assign n10450 = n10449 ^ n10080 ;
  assign n10441 = n10148 & n10152 ;
  assign n10442 = n10079 & n10441 ;
  assign n10451 = n10450 ^ n10442 ;
  assign n10452 = ~n10440 & ~n10451 ;
  assign n10468 = n10185 ^ n10179 ;
  assign n10469 = n10468 ^ n10441 ;
  assign n10470 = n10080 & n10469 ;
  assign n10167 = n10079 ^ n10077 ;
  assign n10463 = n10179 ^ n10163 ;
  assign n10464 = n10463 ^ n10187 ;
  assign n10465 = n10167 & n10464 ;
  assign n10455 = n10188 ^ n10160 ;
  assign n10456 = n10081 & ~n10455 ;
  assign n10457 = n10456 ^ n10162 ;
  assign n10458 = n10193 ^ n10186 ;
  assign n10459 = ~n10081 & ~n10458 ;
  assign n10460 = n10459 ^ n10077 ;
  assign n10461 = ~n10457 & ~n10460 ;
  assign n10202 = n10078 ^ n10077 ;
  assign n10204 = n10184 ^ n10149 ;
  assign n10203 = n10197 ^ n10192 ;
  assign n10205 = n10204 ^ n10203 ;
  assign n10206 = n10205 ^ n10197 ;
  assign n10207 = n10197 ^ n10078 ;
  assign n10208 = n10207 ^ n10197 ;
  assign n10209 = ~n10206 & ~n10208 ;
  assign n10210 = n10209 ^ n10197 ;
  assign n10211 = n10202 & ~n10210 ;
  assign n10212 = n10211 ^ n10197 ;
  assign n10462 = n10461 ^ n10212 ;
  assign n10466 = n10465 ^ n10462 ;
  assign n10453 = n10178 ^ n10157 ;
  assign n10454 = n10079 & n10453 ;
  assign n10467 = n10466 ^ n10454 ;
  assign n10471 = n10470 ^ n10467 ;
  assign n10217 = n10188 ^ n10078 ;
  assign n10218 = n10217 ^ n10188 ;
  assign n10472 = n10188 ^ n10185 ;
  assign n10473 = ~n10218 & n10472 ;
  assign n10474 = n10473 ^ n10188 ;
  assign n10475 = n10077 & n10474 ;
  assign n10476 = n10471 & ~n10475 ;
  assign n10477 = n10452 & n10476 ;
  assign n10478 = n10477 ^ n7571 ;
  assign n11239 = n10478 ^ x109 ;
  assign n7725 = n7724 ^ x89 ;
  assign n7688 = n7687 ^ x98 ;
  assign n7945 = n7725 ^ n7688 ;
  assign n7849 = n7848 ^ x113 ;
  assign n7873 = n7872 ^ n5196 ;
  assign n7851 = ~n6834 & ~n7408 ;
  assign n7867 = ~n6757 & n6780 ;
  assign n7865 = n6789 & n7409 ;
  assign n7863 = n6766 & ~n6793 ;
  assign n7860 = n6778 ^ n6752 ;
  assign n7861 = n6756 & n7860 ;
  assign n7856 = n7409 ^ n6802 ;
  assign n7853 = n7852 ^ n6788 ;
  assign n7854 = n7853 ^ n6794 ;
  assign n7855 = ~n6755 & n7854 ;
  assign n7857 = n7856 ^ n7855 ;
  assign n7858 = ~n6754 & ~n7857 ;
  assign n7859 = n7858 ^ n7855 ;
  assign n7862 = n7861 ^ n7859 ;
  assign n7864 = n7863 ^ n7862 ;
  assign n7866 = n7865 ^ n7864 ;
  assign n7868 = n7867 ^ n7866 ;
  assign n7869 = n7851 & ~n7868 ;
  assign n7850 = n7400 ^ n6791 ;
  assign n7870 = n7869 ^ n7850 ;
  assign n7871 = ~n6759 & n7870 ;
  assign n7874 = n7873 ^ n7871 ;
  assign n7875 = n7874 ^ x123 ;
  assign n7876 = n7849 & ~n7875 ;
  assign n7777 = n7776 ^ x104 ;
  assign n7809 = n7011 & n7018 ;
  assign n7803 = n6986 ^ n6949 ;
  assign n7804 = n6913 & n7803 ;
  assign n7797 = n6971 ^ n6959 ;
  assign n7798 = n7797 ^ n6981 ;
  assign n7805 = n7804 ^ n7798 ;
  assign n7793 = n7019 ^ n6967 ;
  assign n7794 = n7793 ^ n6988 ;
  assign n7795 = n7794 ^ n6975 ;
  assign n7796 = ~n7012 & ~n7795 ;
  assign n7799 = n7798 ^ n7796 ;
  assign n7800 = n7799 ^ n6961 ;
  assign n7801 = n7800 ^ n7799 ;
  assign n7806 = n7805 ^ n7801 ;
  assign n7807 = ~n7004 & n7806 ;
  assign n7808 = n7807 ^ n7800 ;
  assign n7810 = n7809 ^ n7808 ;
  assign n7790 = n6913 & ~n6961 ;
  assign n7791 = ~n6912 & n7454 ;
  assign n7792 = n7790 & n7791 ;
  assign n7811 = n7810 ^ n7792 ;
  assign n7812 = ~n7016 & ~n7811 ;
  assign n7778 = ~n6913 & n6981 ;
  assign n7779 = n7778 ^ n6980 ;
  assign n7780 = n7779 ^ n6982 ;
  assign n7781 = n7780 ^ n6973 ;
  assign n7782 = n7781 ^ n7779 ;
  assign n7783 = n7779 ^ n6912 ;
  assign n7784 = n7783 ^ n7779 ;
  assign n7785 = n7782 & ~n7784 ;
  assign n7786 = n7785 ^ n7779 ;
  assign n7787 = ~n7004 & n7786 ;
  assign n7788 = n7787 ^ n7779 ;
  assign n7789 = n7788 ^ n5161 ;
  assign n7813 = n7812 ^ n7789 ;
  assign n7814 = n7813 ^ x65 ;
  assign n7815 = ~n7777 & n7814 ;
  assign n7883 = n7815 ^ n7777 ;
  assign n7906 = n7883 ^ n7814 ;
  assign n7907 = n7876 & n7906 ;
  assign n7877 = n7876 ^ n7875 ;
  assign n7878 = n7877 ^ n7849 ;
  assign n7879 = n7815 & n7878 ;
  assign n9528 = n7907 ^ n7879 ;
  assign n7881 = n7815 ^ n7814 ;
  assign n7912 = n7876 & n7881 ;
  assign n7913 = n7912 ^ n7876 ;
  assign n7910 = n7876 & ~n7883 ;
  assign n7911 = n7910 ^ n7907 ;
  assign n7914 = n7913 ^ n7911 ;
  assign n7904 = n7876 ^ n7849 ;
  assign n7909 = n7881 & n7904 ;
  assign n7915 = n7914 ^ n7909 ;
  assign n9529 = n9528 ^ n7915 ;
  assign n9530 = n7725 & n9529 ;
  assign n7726 = n7688 & ~n7725 ;
  assign n7727 = n7726 ^ n7688 ;
  assign n7937 = n7904 & n7906 ;
  assign n9398 = ~n7727 & ~n7937 ;
  assign n8666 = n7726 & n7914 ;
  assign n9521 = n9398 ^ n8666 ;
  assign n7905 = n7815 & n7904 ;
  assign n7908 = n7907 ^ n7905 ;
  assign n9522 = n9521 ^ n7908 ;
  assign n9531 = n9530 ^ n9522 ;
  assign n9532 = ~n7945 & ~n9531 ;
  assign n7919 = ~n7877 & n7881 ;
  assign n7890 = n7815 & ~n7877 ;
  assign n7926 = n7919 ^ n7890 ;
  assign n7884 = ~n7877 & ~n7883 ;
  assign n7927 = n7926 ^ n7884 ;
  assign n9523 = n9522 ^ n7927 ;
  assign n7888 = n7875 ^ n7777 ;
  assign n7889 = n7849 & n7888 ;
  assign n7891 = n7890 ^ n7889 ;
  assign n7886 = n7875 ^ n7849 ;
  assign n7887 = n7886 ^ n7777 ;
  assign n7892 = n7891 ^ n7887 ;
  assign n7882 = n7878 & n7881 ;
  assign n7885 = n7884 ^ n7882 ;
  assign n7893 = n7892 ^ n7885 ;
  assign n7920 = n7919 ^ n7893 ;
  assign n7921 = n7893 ^ n7725 ;
  assign n7922 = n7921 ^ n7893 ;
  assign n7923 = ~n7920 & n7922 ;
  assign n7924 = n7923 ^ n7893 ;
  assign n7925 = n7688 & ~n7924 ;
  assign n9524 = n9523 ^ n7925 ;
  assign n7960 = n7915 ^ n7906 ;
  assign n7956 = n7909 ^ n7893 ;
  assign n7916 = n7915 ^ n7908 ;
  assign n7957 = n7956 ^ n7916 ;
  assign n7958 = n7957 ^ n7886 ;
  assign n7959 = n7958 ^ n7927 ;
  assign n7961 = n7960 ^ n7959 ;
  assign n8675 = n7727 & n7961 ;
  assign n7928 = n7927 ^ n7877 ;
  assign n7901 = n7893 ^ n7879 ;
  assign n7900 = n7882 ^ n7878 ;
  assign n7902 = n7901 ^ n7900 ;
  assign n8668 = n7928 ^ n7902 ;
  assign n8669 = n8668 ^ n7937 ;
  assign n8670 = n7937 ^ n7725 ;
  assign n8671 = n8670 ^ n7937 ;
  assign n8672 = n8669 & n8671 ;
  assign n8673 = n8672 ^ n7937 ;
  assign n8674 = ~n7945 & n8673 ;
  assign n8676 = n8675 ^ n8674 ;
  assign n9525 = n9524 ^ n8676 ;
  assign n9516 = n7927 ^ n7725 ;
  assign n9517 = n9516 ^ n7927 ;
  assign n9518 = ~n7958 & ~n9517 ;
  assign n9519 = n9518 ^ n7927 ;
  assign n9520 = ~n7945 & n9519 ;
  assign n9526 = n9525 ^ n9520 ;
  assign n7728 = n7727 ^ n7725 ;
  assign n9513 = n7910 ^ n7882 ;
  assign n9514 = n7728 & n9513 ;
  assign n9527 = n9526 ^ n9514 ;
  assign n9533 = n9532 ^ n9527 ;
  assign n7917 = n7728 ^ n7688 ;
  assign n7952 = ~n7917 & ~n7928 ;
  assign n9534 = n9533 ^ n7952 ;
  assign n9535 = n9534 ^ n6374 ;
  assign n9536 = n9535 ^ x98 ;
  assign n9019 = n6676 ^ n6657 ;
  assign n9020 = n9019 ^ n6199 ;
  assign n9021 = n9020 ^ n6864 ;
  assign n9022 = n5380 & n9021 ;
  assign n9017 = n6893 ^ n6665 ;
  assign n8714 = n6885 ^ n6661 ;
  assign n8708 = ~n6202 & n6658 ;
  assign n8715 = n8714 ^ n8708 ;
  assign n8713 = n6864 ^ n6202 ;
  assign n8716 = n8715 ^ n8713 ;
  assign n8717 = n8716 ^ n6672 ;
  assign n9018 = n9017 ^ n8717 ;
  assign n9023 = n9022 ^ n9018 ;
  assign n8706 = n6866 & ~n6872 ;
  assign n8707 = n8706 ^ n6871 ;
  assign n9036 = n9023 ^ n8707 ;
  assign n9034 = n8717 ^ n8708 ;
  assign n9035 = n6873 & ~n9034 ;
  assign n9037 = n9036 ^ n9035 ;
  assign n8709 = n8708 ^ n6695 ;
  assign n9032 = n8709 ^ n6671 ;
  assign n9033 = n6869 & n9032 ;
  assign n9038 = n9037 ^ n9033 ;
  assign n9024 = n9023 ^ n6689 ;
  assign n9025 = n9024 ^ n6856 ;
  assign n9026 = n9025 ^ n9024 ;
  assign n9027 = n9024 ^ n6693 ;
  assign n9028 = n9027 ^ n9024 ;
  assign n9029 = n9026 & n9028 ;
  assign n9030 = n9029 ^ n9024 ;
  assign n9031 = n6862 & n9030 ;
  assign n9039 = n9038 ^ n9031 ;
  assign n9040 = ~n6868 & ~n9039 ;
  assign n9041 = n9040 ^ n6534 ;
  assign n9537 = n9041 ^ x72 ;
  assign n9662 = n9536 & n9537 ;
  assign n9683 = n9662 ^ n9536 ;
  assign n9684 = n9683 ^ n9537 ;
  assign n9007 = n9006 ^ n8966 ;
  assign n8998 = n8986 ^ n8975 ;
  assign n8997 = n8988 ^ n8971 ;
  assign n8999 = n8998 ^ n8997 ;
  assign n9000 = n8997 ^ n8852 ;
  assign n9001 = n9000 ^ n8997 ;
  assign n9002 = n8999 & ~n9001 ;
  assign n9003 = n9002 ^ n8997 ;
  assign n9004 = ~n8996 & ~n9003 ;
  assign n9008 = n9007 ^ n9004 ;
  assign n8993 = n8992 ^ n8988 ;
  assign n8994 = n8993 ^ n8948 ;
  assign n8995 = n8855 & n8994 ;
  assign n9009 = n9008 ^ n8995 ;
  assign n8976 = n8975 ^ n8947 ;
  assign n8977 = n8976 ^ n8954 ;
  assign n8973 = n8972 ^ n8968 ;
  assign n8978 = n8977 ^ n8973 ;
  assign n8965 = n8964 ^ n8950 ;
  assign n8979 = n8978 ^ n8965 ;
  assign n8980 = n8978 ^ n8852 ;
  assign n8981 = n8980 ^ n8978 ;
  assign n8982 = ~n8979 & ~n8981 ;
  assign n8983 = n8982 ^ n8978 ;
  assign n8984 = ~n8851 & n8983 ;
  assign n9010 = n9009 ^ n8984 ;
  assign n8943 = n8942 ^ n8941 ;
  assign n8956 = n8955 ^ n8854 ;
  assign n8957 = n8941 ^ n8854 ;
  assign n8958 = n8957 ^ n8854 ;
  assign n8959 = ~n8956 & ~n8958 ;
  assign n8960 = n8959 ^ n8854 ;
  assign n8961 = n8943 & ~n8960 ;
  assign n9011 = n9010 ^ n8961 ;
  assign n9012 = ~n8939 & n9011 ;
  assign n9013 = n9012 ^ n6461 ;
  assign n9587 = n9013 ^ x104 ;
  assign n8574 = n8559 ^ n8461 ;
  assign n9620 = n9592 ^ n8566 ;
  assign n9621 = ~n8574 & n9620 ;
  assign n8575 = n8574 ^ n8532 ;
  assign n8576 = n8556 & n8575 ;
  assign n8577 = n8576 ^ n8573 ;
  assign n9615 = n8577 ^ n8566 ;
  assign n9063 = n8557 & n8559 ;
  assign n8578 = n8517 & n8575 ;
  assign n9064 = n9063 ^ n8578 ;
  assign n9616 = n9615 ^ n9064 ;
  assign n9617 = n9616 ^ n9614 ;
  assign n9618 = n9617 ^ n6252 ;
  assign n9601 = n8523 ^ n8511 ;
  assign n9602 = n9601 ^ n8523 ;
  assign n9605 = n8532 & n9602 ;
  assign n9606 = n9605 ^ n8523 ;
  assign n9607 = n8461 & n9606 ;
  assign n9619 = n9618 ^ n9607 ;
  assign n9622 = n9621 ^ n9619 ;
  assign n9594 = n9592 ^ n8522 ;
  assign n9593 = n9592 ^ n8554 ;
  assign n9595 = n9594 ^ n9593 ;
  assign n9596 = n9594 ^ n8461 ;
  assign n9597 = n9596 ^ n9594 ;
  assign n9598 = ~n9595 & n9597 ;
  assign n9599 = n9598 ^ n9594 ;
  assign n9600 = ~n8532 & ~n9599 ;
  assign n9623 = n9622 ^ n9600 ;
  assign n9624 = n9623 ^ x113 ;
  assign n8685 = n7315 ^ n7310 ;
  assign n8686 = n8685 ^ n7300 ;
  assign n8684 = n7292 ^ n7291 ;
  assign n8687 = n8686 ^ n8684 ;
  assign n8689 = ~n7298 & n8687 ;
  assign n8690 = n8689 ^ n8684 ;
  assign n9577 = ~n7034 & n8690 ;
  assign n9576 = n7319 ^ n6911 ;
  assign n9578 = n9577 ^ n9576 ;
  assign n9583 = n9578 ^ n6745 ;
  assign n9579 = n6911 & n9578 ;
  assign n9580 = n7314 & n9579 ;
  assign n9581 = n7034 & n9580 ;
  assign n9582 = n9581 ^ n9579 ;
  assign n9584 = n9583 ^ n9582 ;
  assign n9569 = n7034 ^ n6911 ;
  assign n8683 = n7313 ^ n7294 ;
  assign n8688 = n8687 ^ n8683 ;
  assign n9570 = n8688 ^ n7324 ;
  assign n9571 = n8688 ^ n6911 ;
  assign n9572 = n9571 ^ n8688 ;
  assign n9573 = ~n9570 & ~n9572 ;
  assign n9574 = n9573 ^ n8688 ;
  assign n9575 = n9569 & ~n9574 ;
  assign n9585 = n9584 ^ n9575 ;
  assign n9586 = n9585 ^ x66 ;
  assign n9644 = n9624 ^ n9586 ;
  assign n8003 = n8002 ^ x118 ;
  assign n8037 = n7500 ^ n7480 ;
  assign n8038 = n8037 ^ n6194 ;
  assign n8039 = n8038 ^ n4078 ;
  assign n8034 = n5978 & n6156 ;
  assign n8024 = n6126 ^ n6119 ;
  assign n8025 = n8024 ^ n6120 ;
  assign n8026 = n8025 ^ n6113 ;
  assign n8027 = n8026 ^ n6119 ;
  assign n8028 = ~n5976 & ~n8027 ;
  assign n8029 = n8028 ^ n8024 ;
  assign n8030 = n5977 & n8029 ;
  assign n8010 = n6149 ^ n6137 ;
  assign n8011 = n8010 ^ n6141 ;
  assign n8012 = ~n5977 & n8011 ;
  assign n8013 = n8012 ^ n6141 ;
  assign n8031 = n8030 ^ n8013 ;
  assign n8021 = ~n5977 & n6018 ;
  assign n8022 = n8021 ^ n5976 ;
  assign n8023 = n6123 & n8022 ;
  assign n8032 = n8031 ^ n8023 ;
  assign n8014 = n8013 ^ n6142 ;
  assign n8006 = n6156 ^ n6142 ;
  assign n8007 = n8006 ^ n6147 ;
  assign n8015 = n8014 ^ n8007 ;
  assign n8008 = n8007 ^ n7497 ;
  assign n8009 = n5976 & ~n8008 ;
  assign n8016 = n8015 ^ n8009 ;
  assign n8017 = n6164 & ~n8016 ;
  assign n8033 = n8032 ^ n8017 ;
  assign n8035 = n8034 ^ n8033 ;
  assign n8036 = ~n6180 & ~n8035 ;
  assign n8040 = n8039 ^ n8036 ;
  assign n8041 = n8040 ^ x75 ;
  assign n8063 = n6988 & n7011 ;
  assign n8058 = n7028 ^ n6956 ;
  assign n8049 = n6978 ^ n6947 ;
  assign n8059 = n8058 ^ n8049 ;
  assign n8060 = n8059 ^ n7788 ;
  assign n8061 = n8060 ^ n7010 ;
  assign n8050 = n8049 ^ n6968 ;
  assign n8051 = n8050 ^ n7018 ;
  assign n8052 = n8051 ^ n8049 ;
  assign n8053 = n8049 ^ n6913 ;
  assign n8054 = n8053 ^ n8049 ;
  assign n8055 = n8052 & ~n8054 ;
  assign n8056 = n8055 ^ n8049 ;
  assign n8057 = ~n7004 & n8056 ;
  assign n8062 = n8061 ^ n8057 ;
  assign n8064 = n8063 ^ n8062 ;
  assign n8044 = n6956 ^ n6913 ;
  assign n8045 = n8044 ^ n6956 ;
  assign n8046 = ~n7793 & n8045 ;
  assign n8047 = n8046 ^ n6956 ;
  assign n8048 = n6912 & n8047 ;
  assign n8065 = n8064 ^ n8048 ;
  assign n8066 = n8065 ^ n7451 ;
  assign n8067 = ~n7473 & ~n8066 ;
  assign n8068 = n8067 ^ n4036 ;
  assign n8069 = n8068 ^ x94 ;
  assign n8070 = n8041 & n8069 ;
  assign n8071 = n8070 ^ n8041 ;
  assign n8111 = n8110 ^ x77 ;
  assign n8112 = n5379 ^ x84 ;
  assign n8113 = n8111 & n8112 ;
  assign n8151 = n8071 & n8113 ;
  assign n7978 = n6440 ^ x101 ;
  assign n9564 = n8151 ^ n7978 ;
  assign n9565 = ~n8003 & n9564 ;
  assign n8004 = n7978 & ~n8003 ;
  assign n8114 = n8113 ^ n8112 ;
  assign n8147 = n8071 & n8114 ;
  assign n8118 = n8113 ^ n8111 ;
  assign n8119 = n8071 & n8118 ;
  assign n8115 = n8114 ^ n8111 ;
  assign n8117 = n8070 & ~n8115 ;
  assign n8120 = n8119 ^ n8117 ;
  assign n9557 = n8147 ^ n8120 ;
  assign n8072 = n8071 ^ n8069 ;
  assign n8128 = ~n8072 & n8118 ;
  assign n8121 = n8071 & ~n8115 ;
  assign n8129 = n8128 ^ n8121 ;
  assign n8124 = ~n8041 & n8112 ;
  assign n8125 = n8124 ^ n8041 ;
  assign n8126 = n8125 ^ n8112 ;
  assign n8122 = n8121 ^ n8120 ;
  assign n8127 = n8126 ^ n8122 ;
  assign n8130 = n8129 ^ n8127 ;
  assign n8131 = n8130 ^ n8117 ;
  assign n8123 = n8122 ^ n8118 ;
  assign n8132 = n8131 ^ n8123 ;
  assign n8116 = ~n8072 & ~n8115 ;
  assign n8133 = n8132 ^ n8116 ;
  assign n8154 = n8133 ^ n8128 ;
  assign n8155 = n8154 ^ n8125 ;
  assign n8156 = n8155 ^ n8132 ;
  assign n9558 = n9557 ^ n8156 ;
  assign n9559 = n8004 & ~n9558 ;
  assign n9548 = n8131 ^ n8003 ;
  assign n9549 = n9548 ^ n8131 ;
  assign n9550 = ~n8121 & ~n8154 ;
  assign n9551 = n9550 ^ n8131 ;
  assign n9552 = n9549 & ~n9551 ;
  assign n9553 = n9552 ^ n8131 ;
  assign n9554 = ~n7978 & ~n9553 ;
  assign n9555 = n9554 ^ n7978 ;
  assign n8182 = n8126 ^ n8041 ;
  assign n8148 = ~n8072 & n8113 ;
  assign n8149 = n8148 ^ n8147 ;
  assign n8143 = n8072 ^ n8041 ;
  assign n8144 = n8113 & n8143 ;
  assign n8145 = n8144 ^ n8124 ;
  assign n8146 = n8145 ^ n8114 ;
  assign n8150 = n8149 ^ n8146 ;
  assign n8152 = n8151 ^ n8150 ;
  assign n8181 = n8152 ^ n8147 ;
  assign n8183 = n8182 ^ n8181 ;
  assign n8135 = n8004 ^ n7978 ;
  assign n8005 = n8004 ^ n8003 ;
  assign n8198 = n8135 ^ n8005 ;
  assign n9547 = n8183 & n8198 ;
  assign n9556 = n9555 ^ n9547 ;
  assign n9560 = n9559 ^ n9556 ;
  assign n8206 = ~n7978 & n8150 ;
  assign n8157 = n8144 ^ n8143 ;
  assign n8158 = n8157 ^ n8156 ;
  assign n8199 = n8158 ^ n8003 ;
  assign n8200 = n8199 ^ n8158 ;
  assign n8159 = n8158 ^ n8148 ;
  assign n8160 = n8159 ^ n8145 ;
  assign n8201 = n8160 ^ n8151 ;
  assign n8202 = n8201 ^ n8158 ;
  assign n8203 = n8200 & n8202 ;
  assign n8204 = n8203 ^ n8158 ;
  assign n8205 = n8198 & ~n8204 ;
  assign n8207 = n8206 ^ n8205 ;
  assign n9546 = n8207 ^ n7978 ;
  assign n9561 = n9560 ^ n9546 ;
  assign n8192 = n8135 & n8149 ;
  assign n8190 = n8155 ^ n8127 ;
  assign n8191 = n8135 & ~n8190 ;
  assign n8193 = n8192 ^ n8191 ;
  assign n9562 = n9561 ^ n8193 ;
  assign n9563 = n9562 ^ n6732 ;
  assign n9566 = n9565 ^ n9563 ;
  assign n8161 = n8160 ^ n8144 ;
  assign n9539 = n8161 ^ n8135 ;
  assign n9540 = n8129 ^ n8005 ;
  assign n9543 = n8161 & n9540 ;
  assign n9544 = n9543 ^ n8005 ;
  assign n9545 = ~n9539 & ~n9544 ;
  assign n9567 = n9566 ^ n9545 ;
  assign n9568 = n9567 ^ x65 ;
  assign n9645 = n9644 ^ n9568 ;
  assign n9646 = n9587 & ~n9645 ;
  assign n9647 = n9646 ^ n9645 ;
  assign n9625 = n9587 & ~n9624 ;
  assign n9631 = n9625 ^ n9587 ;
  assign n9632 = n9631 ^ n9624 ;
  assign n9590 = ~n9568 & ~n9586 ;
  assign n9639 = n9590 ^ n9586 ;
  assign n9640 = n9632 & ~n9639 ;
  assign n9634 = n9625 ^ n9624 ;
  assign n9635 = n9590 & ~n9634 ;
  assign n9641 = n9640 ^ n9635 ;
  assign n9633 = n9590 & n9632 ;
  assign n9636 = n9635 ^ n9633 ;
  assign n9637 = n9636 ^ n9632 ;
  assign n9627 = n9624 ^ n9568 ;
  assign n9588 = n9587 ^ n9586 ;
  assign n9589 = ~n9568 & n9588 ;
  assign n9628 = n9589 ^ n9587 ;
  assign n9629 = ~n9627 & ~n9628 ;
  assign n9626 = n9590 & n9625 ;
  assign n9630 = n9629 ^ n9626 ;
  assign n9638 = n9637 ^ n9630 ;
  assign n9642 = n9641 ^ n9638 ;
  assign n9648 = n9647 ^ n9642 ;
  assign n9643 = n9642 ^ n9637 ;
  assign n9649 = n9648 ^ n9643 ;
  assign n9650 = n9649 ^ n9640 ;
  assign n9651 = n9650 ^ n9587 ;
  assign n9591 = n9590 ^ n9589 ;
  assign n9652 = n9651 ^ n9591 ;
  assign n11258 = n9652 ^ n9648 ;
  assign n11259 = ~n9684 & ~n11258 ;
  assign n9538 = n9537 ^ n9536 ;
  assign n9670 = n9639 ^ n9568 ;
  assign n9671 = n9625 & ~n9670 ;
  assign n9672 = n9671 ^ n9670 ;
  assign n9673 = n9672 ^ n9649 ;
  assign n9665 = n9625 & ~n9639 ;
  assign n9674 = n9673 ^ n9665 ;
  assign n9687 = n9674 ^ n9646 ;
  assign n11249 = n9687 ^ n9629 ;
  assign n11250 = n11249 ^ n9587 ;
  assign n11251 = n11250 ^ n9687 ;
  assign n11252 = n9687 ^ n9537 ;
  assign n11253 = n11252 ^ n9687 ;
  assign n11254 = ~n11251 & n11253 ;
  assign n11255 = n11254 ^ n9687 ;
  assign n11256 = ~n9538 & n11255 ;
  assign n9699 = n9652 ^ n9638 ;
  assign n9700 = n9699 ^ n9635 ;
  assign n9701 = n9700 ^ n9633 ;
  assign n9702 = n9701 ^ n9651 ;
  assign n9703 = n9702 ^ n9683 ;
  assign n9704 = n9684 ^ n9536 ;
  assign n9705 = n9704 ^ n9643 ;
  assign n9708 = n9702 & ~n9705 ;
  assign n9709 = n9708 ^ n9643 ;
  assign n9710 = n9703 & ~n9709 ;
  assign n9711 = n9710 ^ n9683 ;
  assign n11247 = n9711 ^ n9646 ;
  assign n9715 = n9646 ^ n9587 ;
  assign n10427 = n9715 ^ n9674 ;
  assign n10428 = ~n9684 & n10427 ;
  assign n11248 = n11247 ^ n10428 ;
  assign n11257 = n11256 ^ n11248 ;
  assign n11260 = n11259 ^ n11257 ;
  assign n11242 = n9641 ^ n9536 ;
  assign n11243 = n11242 ^ n9641 ;
  assign n11244 = n9642 & ~n11243 ;
  assign n11245 = n11244 ^ n9641 ;
  assign n11246 = n9538 & n11245 ;
  assign n11261 = n11260 ^ n11246 ;
  assign n11262 = n11261 ^ n8110 ;
  assign n11240 = n9643 ^ n9633 ;
  assign n11241 = ~n9536 & n11240 ;
  assign n11263 = n11262 ^ n11241 ;
  assign n11264 = n11263 ^ x118 ;
  assign n11265 = ~n11239 & n11264 ;
  assign n7962 = n7961 ^ n7919 ;
  assign n7955 = n7912 ^ n7910 ;
  assign n7963 = n7962 ^ n7955 ;
  assign n7964 = n7728 & n7963 ;
  assign n7946 = n7937 ^ n7890 ;
  assign n7947 = n7890 ^ n7725 ;
  assign n7948 = n7947 ^ n7890 ;
  assign n7949 = n7946 & n7948 ;
  assign n7950 = n7949 ^ n7890 ;
  assign n7951 = ~n7945 & n7950 ;
  assign n7953 = n7952 ^ n7951 ;
  assign n7954 = n7953 ^ n7885 ;
  assign n7965 = n7964 ^ n7954 ;
  assign n7936 = n7902 ^ n7885 ;
  assign n7938 = n7937 ^ n7936 ;
  assign n7939 = n7938 ^ n7885 ;
  assign n7940 = n7885 ^ n7688 ;
  assign n7941 = n7940 ^ n7885 ;
  assign n7942 = ~n7939 & ~n7941 ;
  assign n7943 = n7942 ^ n7885 ;
  assign n7944 = ~n7725 & n7943 ;
  assign n7966 = n7965 ^ n7944 ;
  assign n7929 = n7928 ^ n7891 ;
  assign n7930 = n7929 ^ n7913 ;
  assign n7931 = n7913 ^ n7725 ;
  assign n7932 = n7931 ^ n7913 ;
  assign n7933 = ~n7930 & ~n7932 ;
  assign n7934 = n7933 ^ n7913 ;
  assign n7935 = n7688 & n7934 ;
  assign n7967 = n7966 ^ n7935 ;
  assign n7968 = n7967 ^ n7879 ;
  assign n7969 = n7968 ^ n7925 ;
  assign n7970 = n7969 ^ n5290 ;
  assign n7918 = n7916 & ~n7917 ;
  assign n7971 = n7970 ^ n7918 ;
  assign n7903 = n7727 & ~n7902 ;
  assign n7972 = n7971 ^ n7903 ;
  assign n7880 = n7879 ^ n7728 ;
  assign n7894 = n7893 ^ n7726 ;
  assign n7897 = n7728 & n7894 ;
  assign n7898 = n7897 ^ n7726 ;
  assign n7899 = n7880 & ~n7898 ;
  assign n7973 = n7972 ^ n7899 ;
  assign n9728 = n7973 ^ x118 ;
  assign n8691 = n8690 ^ n8688 ;
  assign n8692 = ~n6911 & n8691 ;
  assign n8693 = n8692 ^ n8690 ;
  assign n8694 = n8693 ^ n7324 ;
  assign n8695 = n8694 ^ n7325 ;
  assign n8696 = n8695 ^ n8694 ;
  assign n8699 = ~n6911 & ~n8696 ;
  assign n8700 = n8699 ^ n8694 ;
  assign n8701 = n7034 & n8700 ;
  assign n8702 = n8701 ^ n8693 ;
  assign n8703 = ~n7319 & ~n8702 ;
  assign n8704 = n8703 ^ n3797 ;
  assign n9727 = n8704 ^ x69 ;
  assign n8208 = n8207 ^ n8003 ;
  assign n8171 = ~n8005 & ~n8159 ;
  assign n8169 = n8144 ^ n8127 ;
  assign n8142 = n8003 ^ n7978 ;
  assign n8153 = n8152 ^ n8128 ;
  assign n8162 = n8161 ^ n8153 ;
  assign n8163 = n8162 ^ n8128 ;
  assign n8164 = n8128 ^ n8003 ;
  assign n8165 = n8164 ^ n8128 ;
  assign n8166 = ~n8163 & ~n8165 ;
  assign n8167 = n8166 ^ n8128 ;
  assign n8168 = n8142 & n8167 ;
  assign n8170 = n8169 ^ n8168 ;
  assign n8172 = n8171 ^ n8170 ;
  assign n8209 = n8208 ^ n8172 ;
  assign n8194 = n8005 ^ n7978 ;
  assign n8195 = n8155 ^ n8119 ;
  assign n8196 = n8194 & ~n8195 ;
  assign n8197 = n8196 ^ n8193 ;
  assign n8210 = n8209 ^ n8197 ;
  assign n8184 = n8183 ^ n8120 ;
  assign n8185 = n8120 ^ n8003 ;
  assign n8186 = n8185 ^ n8120 ;
  assign n8187 = n8184 & n8186 ;
  assign n8188 = n8187 ^ n8120 ;
  assign n8189 = n7978 & n8188 ;
  assign n8211 = n8210 ^ n8189 ;
  assign n8212 = n8211 ^ n4263 ;
  assign n8173 = n8172 ^ n8168 ;
  assign n8174 = n8173 ^ n8117 ;
  assign n8175 = n8174 ^ n8173 ;
  assign n8176 = n8173 ^ n8003 ;
  assign n8177 = n8176 ^ n8173 ;
  assign n8178 = ~n8175 & n8177 ;
  assign n8179 = n8178 ^ n8173 ;
  assign n8180 = n7978 & ~n8179 ;
  assign n8213 = n8212 ^ n8180 ;
  assign n8134 = n8133 ^ n8005 ;
  assign n8136 = n8135 ^ n8121 ;
  assign n8137 = n8121 ^ n8005 ;
  assign n8138 = n8137 ^ n8121 ;
  assign n8139 = ~n8136 & n8138 ;
  assign n8140 = n8139 ^ n8121 ;
  assign n8141 = ~n8134 & ~n8140 ;
  assign n8214 = n8213 ^ n8141 ;
  assign n9762 = n8214 ^ x83 ;
  assign n9785 = n8337 ^ n8324 ;
  assign n9781 = n8311 ^ n8280 ;
  assign n9782 = n9781 ^ n8285 ;
  assign n9783 = ~n8269 & n9782 ;
  assign n9772 = n8314 ^ n8304 ;
  assign n9773 = n9772 ^ n8297 ;
  assign n9774 = n9773 ^ n9772 ;
  assign n9775 = n9772 ^ n8275 ;
  assign n9776 = n9775 ^ n9772 ;
  assign n9777 = n9774 & n9776 ;
  assign n9778 = n9777 ^ n9772 ;
  assign n9779 = ~n8276 & n9778 ;
  assign n9780 = n9779 ^ n8304 ;
  assign n9784 = n9783 ^ n9780 ;
  assign n9786 = n9785 ^ n9784 ;
  assign n9277 = n8313 ^ n8290 ;
  assign n9099 = n8280 ^ n8274 ;
  assign n9764 = n9277 ^ n9099 ;
  assign n9765 = n9277 ^ n8324 ;
  assign n9766 = n9765 ^ n9277 ;
  assign n9767 = ~n9764 & ~n9766 ;
  assign n9768 = n9767 ^ n9277 ;
  assign n9769 = n8292 ^ n8269 ;
  assign n9770 = n9769 ^ n8268 ;
  assign n9771 = ~n9768 & ~n9770 ;
  assign n9787 = n9786 ^ n9771 ;
  assign n9115 = n8303 & n8311 ;
  assign n9788 = n9787 ^ n9115 ;
  assign n9789 = n9788 ^ n8320 ;
  assign n9763 = n8281 & ~n8308 ;
  assign n9790 = n9789 ^ n9763 ;
  assign n9791 = ~n8284 & ~n9790 ;
  assign n9792 = n9791 ^ n4918 ;
  assign n9793 = n9792 ^ x86 ;
  assign n9794 = n9762 & ~n9793 ;
  assign n9753 = n8951 ^ n8945 ;
  assign n9754 = n9753 ^ n8954 ;
  assign n9755 = ~n8852 & ~n9754 ;
  assign n9756 = n9755 ^ n8964 ;
  assign n9757 = n8996 & n9756 ;
  assign n9751 = n8942 & ~n9750 ;
  assign n9745 = n8855 & n9744 ;
  assign n9739 = n8938 & ~n9736 ;
  assign n9737 = n9736 ^ n8947 ;
  assign n9738 = ~n8996 & n9737 ;
  assign n9740 = n9739 ^ n9738 ;
  assign n9741 = n9740 ^ n9376 ;
  assign n9735 = ~n8854 & n8954 ;
  assign n9742 = n9741 ^ n9735 ;
  assign n9732 = n8963 ^ n8952 ;
  assign n9733 = n9732 ^ n8968 ;
  assign n9734 = n8853 & n9733 ;
  assign n9743 = n9742 ^ n9734 ;
  assign n9746 = n9745 ^ n9743 ;
  assign n9730 = n8989 ^ n8972 ;
  assign n9731 = ~n8854 & n9730 ;
  assign n9747 = n9746 ^ n9731 ;
  assign n9748 = n9747 ^ n8964 ;
  assign n9749 = n9748 ^ n4696 ;
  assign n9752 = n9751 ^ n9749 ;
  assign n9758 = n9757 ^ n9752 ;
  assign n9759 = n9758 ^ x100 ;
  assign n8579 = n8578 ^ n8577 ;
  assign n8580 = n8579 ^ n8529 ;
  assign n8561 = n8554 ^ n8518 ;
  assign n8563 = n8562 ^ n8561 ;
  assign n8564 = ~n8560 & n8563 ;
  assign n8581 = n8580 ^ n8564 ;
  assign n8558 = ~n8552 & n8557 ;
  assign n8582 = n8581 ^ n8558 ;
  assign n8547 = n8539 ^ n8461 ;
  assign n8548 = n8547 ^ n8539 ;
  assign n8549 = n8544 & n8548 ;
  assign n8550 = n8549 ^ n8539 ;
  assign n8551 = n8532 & n8550 ;
  assign n8583 = n8582 ^ n8551 ;
  assign n8530 = n8529 ^ n8522 ;
  assign n8531 = n8530 ^ n8529 ;
  assign n8535 = ~n8531 & ~n8532 ;
  assign n8536 = n8535 ^ n8529 ;
  assign n8537 = n8461 & ~n8536 ;
  assign n8584 = n8583 ^ n8537 ;
  assign n8586 = n8585 ^ n8584 ;
  assign n8587 = n8586 ^ n5113 ;
  assign n9760 = n8587 ^ x93 ;
  assign n9761 = n9759 & ~n9760 ;
  assign n9826 = n9761 ^ n9760 ;
  assign n9842 = n9794 & ~n9826 ;
  assign n9798 = n9794 ^ n9762 ;
  assign n9796 = n9761 ^ n9759 ;
  assign n9804 = n9796 ^ n9760 ;
  assign n9805 = n9798 & n9804 ;
  assign n9799 = n9761 & n9798 ;
  assign n9797 = n9794 & n9796 ;
  assign n9800 = n9799 ^ n9797 ;
  assign n9840 = n9805 ^ n9800 ;
  assign n9802 = n9796 & n9798 ;
  assign n9803 = n9802 ^ n9799 ;
  assign n9806 = n9805 ^ n9803 ;
  assign n9807 = n9806 ^ n9798 ;
  assign n9841 = n9840 ^ n9807 ;
  assign n9843 = n9842 ^ n9841 ;
  assign n9795 = n9761 & n9794 ;
  assign n9838 = n9802 ^ n9795 ;
  assign n9839 = n9838 ^ n9762 ;
  assign n9844 = n9843 ^ n9839 ;
  assign n10288 = n9844 ^ n9807 ;
  assign n9809 = n9798 ^ n9793 ;
  assign n9829 = n9761 & n9809 ;
  assign n9827 = n9809 & ~n9826 ;
  assign n9810 = n9796 & n9809 ;
  assign n9828 = n9827 ^ n9810 ;
  assign n9830 = n9829 ^ n9828 ;
  assign n9831 = n9830 ^ n9809 ;
  assign n9811 = n9794 ^ n9793 ;
  assign n9815 = n9761 & ~n9811 ;
  assign n10287 = n9831 ^ n9815 ;
  assign n10289 = n10288 ^ n10287 ;
  assign n10290 = n9727 & n10289 ;
  assign n10291 = n10290 ^ n10288 ;
  assign n10294 = n10291 ^ n9800 ;
  assign n10295 = n10294 ^ n10291 ;
  assign n10296 = ~n9727 & n10295 ;
  assign n10297 = n10296 ^ n10291 ;
  assign n10298 = ~n9728 & n10297 ;
  assign n10299 = n10298 ^ n10291 ;
  assign n9859 = n9829 ^ n9727 ;
  assign n9860 = n9859 ^ n9829 ;
  assign n9812 = n9804 & ~n9811 ;
  assign n9861 = n9827 ^ n9812 ;
  assign n9862 = n9861 ^ n9829 ;
  assign n9863 = n9860 & n9862 ;
  assign n9864 = n9863 ^ n9829 ;
  assign n9865 = ~n9728 & n9864 ;
  assign n11284 = n10299 ^ n9865 ;
  assign n9814 = n9796 & ~n9811 ;
  assign n10266 = n9829 ^ n9814 ;
  assign n9847 = n9842 ^ n9797 ;
  assign n11269 = n10266 ^ n9847 ;
  assign n11267 = n9840 ^ n9795 ;
  assign n9816 = n9815 ^ n9814 ;
  assign n9813 = n9812 ^ n9811 ;
  assign n9817 = n9816 ^ n9813 ;
  assign n9818 = n9817 ^ n9810 ;
  assign n11268 = n11267 ^ n9818 ;
  assign n11270 = n11269 ^ n11268 ;
  assign n11271 = n11270 ^ n9818 ;
  assign n11272 = n9728 & n11271 ;
  assign n11273 = n11272 ^ n11268 ;
  assign n11285 = n11284 ^ n11273 ;
  assign n11286 = n11285 ^ n8496 ;
  assign n9729 = n9728 ^ n9727 ;
  assign n11276 = n10288 ^ n9815 ;
  assign n9832 = n9831 ^ n9817 ;
  assign n11277 = n11276 ^ n9832 ;
  assign n11278 = n11277 ^ n11273 ;
  assign n11274 = n9861 ^ n9799 ;
  assign n11080 = n9838 ^ n9805 ;
  assign n11275 = n11274 ^ n11080 ;
  assign n11279 = n11278 ^ n11275 ;
  assign n11280 = n11279 ^ n11273 ;
  assign n11281 = n9728 & ~n11280 ;
  assign n11282 = n11281 ^ n11278 ;
  assign n11283 = ~n9729 & n11282 ;
  assign n11287 = n11286 ^ n11283 ;
  assign n11288 = n11287 ^ x85 ;
  assign n9014 = n9013 ^ x82 ;
  assign n8616 = n8161 ^ n8113 ;
  assign n8591 = ~n8069 & n8111 ;
  assign n8617 = n8616 ^ n8591 ;
  assign n8620 = n8617 ^ n8121 ;
  assign n8615 = n8120 ^ n8116 ;
  assign n8618 = n8617 ^ n8615 ;
  assign n8619 = ~n7978 & ~n8618 ;
  assign n8621 = n8620 ^ n8619 ;
  assign n8622 = ~n8003 & n8621 ;
  assign n8614 = n8205 ^ n8196 ;
  assign n8623 = n8622 ^ n8614 ;
  assign n8611 = n8132 ^ n8121 ;
  assign n8612 = n8611 ^ n8003 ;
  assign n8613 = ~n7978 & n8612 ;
  assign n8624 = n8623 ^ n8613 ;
  assign n8592 = n8591 ^ n8112 ;
  assign n8593 = n8111 ^ n8041 ;
  assign n8594 = ~n8135 & n8593 ;
  assign n8595 = n8592 & n8594 ;
  assign n8596 = n8595 ^ n8135 ;
  assign n8597 = n8127 ^ n8005 ;
  assign n8598 = n8597 ^ n8127 ;
  assign n8601 = ~n8154 & n8598 ;
  assign n8602 = n8601 ^ n8127 ;
  assign n8603 = n8596 & ~n8602 ;
  assign n8604 = n8603 ^ n8135 ;
  assign n8605 = n8181 ^ n8005 ;
  assign n8608 = ~n8603 & n8605 ;
  assign n8609 = n8608 ^ n8005 ;
  assign n8610 = n8604 & ~n8609 ;
  assign n8625 = n8624 ^ n8610 ;
  assign n8590 = ~n8159 & n8194 ;
  assign n8626 = n8625 ^ n8590 ;
  assign n8627 = n8190 ^ n8144 ;
  assign n8628 = n8144 ^ n8003 ;
  assign n8629 = n8628 ^ n8144 ;
  assign n8630 = ~n8627 & ~n8629 ;
  assign n8631 = n8630 ^ n8144 ;
  assign n8632 = n7978 & n8631 ;
  assign n8633 = n8626 & ~n8632 ;
  assign n8634 = n8633 ^ n6060 ;
  assign n8850 = n8634 ^ x73 ;
  assign n9015 = n9014 ^ n8850 ;
  assign n9042 = n9041 ^ x88 ;
  assign n8427 = n7588 ^ n7374 ;
  assign n8428 = n7588 ^ n7585 ;
  assign n8429 = n8428 ^ n7398 ;
  assign n8430 = n8429 ^ n8428 ;
  assign n8433 = n7586 & n8430 ;
  assign n8434 = n8433 ^ n8428 ;
  assign n8435 = n8427 & ~n8434 ;
  assign n8436 = n8435 ^ n7374 ;
  assign n7623 = ~n7374 & n7398 ;
  assign n7625 = n7623 ^ n7374 ;
  assign n8425 = n7650 ^ n7576 ;
  assign n8426 = ~n7625 & n8425 ;
  assign n8437 = n8436 ^ n8426 ;
  assign n8422 = n7598 ^ n7591 ;
  assign n8421 = n7608 ^ n7582 ;
  assign n8423 = n8422 ^ n8421 ;
  assign n8424 = n7623 & n8423 ;
  assign n8438 = n8437 ^ n8424 ;
  assign n7624 = n7623 ^ n7398 ;
  assign n7626 = n7625 ^ n7624 ;
  assign n8420 = ~n7615 & ~n7626 ;
  assign n8439 = n8438 ^ n8420 ;
  assign n8441 = ~n7398 & n8440 ;
  assign n8442 = n8441 ^ n7576 ;
  assign n8443 = n8442 ^ n7374 ;
  assign n8444 = n8443 ^ n8442 ;
  assign n8446 = ~n7398 & n8445 ;
  assign n8447 = n8446 ^ n8442 ;
  assign n8448 = n8444 & n8447 ;
  assign n8449 = n8448 ^ n8442 ;
  assign n8450 = ~n8439 & n8449 ;
  assign n8451 = n8450 ^ n8439 ;
  assign n8452 = n7591 ^ n7398 ;
  assign n8453 = n8452 ^ n7591 ;
  assign n8455 = n7598 & ~n8453 ;
  assign n8456 = n8455 ^ n7591 ;
  assign n8457 = n7374 & n8456 ;
  assign n8458 = ~n8451 & ~n8457 ;
  assign n8459 = n8458 ^ n5975 ;
  assign n9016 = n8459 ^ x97 ;
  assign n9080 = n8541 & n8575 ;
  assign n9074 = n8519 ^ n8511 ;
  assign n9075 = n9074 ^ n9068 ;
  assign n9076 = ~n8532 & n9075 ;
  assign n9069 = n9068 ^ n8554 ;
  assign n9070 = n9069 ^ n9053 ;
  assign n9071 = n8532 & n9070 ;
  assign n9066 = n8554 ^ n8538 ;
  assign n9067 = n9066 ^ n8566 ;
  assign n9072 = n9071 ^ n9067 ;
  assign n9077 = n9076 ^ n9072 ;
  assign n9078 = n8461 & n9077 ;
  assign n9065 = n9064 ^ n9062 ;
  assign n9073 = n9072 ^ n9065 ;
  assign n9079 = n9078 ^ n9073 ;
  assign n9081 = n9080 ^ n9079 ;
  assign n9052 = n8559 & n8562 ;
  assign n9082 = n9081 ^ n9052 ;
  assign n9044 = n8529 ^ n8513 ;
  assign n9045 = n9044 ^ n8509 ;
  assign n9046 = n9045 ^ n9044 ;
  assign n9047 = n9044 ^ n8461 ;
  assign n9048 = n9047 ^ n9044 ;
  assign n9049 = n9046 & n9048 ;
  assign n9050 = n9049 ^ n9044 ;
  assign n9051 = ~n8552 & ~n9050 ;
  assign n9083 = n9082 ^ n9051 ;
  assign n9084 = n9083 ^ n8585 ;
  assign n9085 = n9084 ^ n6493 ;
  assign n9086 = n9085 ^ x114 ;
  assign n9132 = n9016 & ~n9086 ;
  assign n9134 = n9132 ^ n9016 ;
  assign n9163 = ~n9042 & n9134 ;
  assign n9101 = n8297 ^ n8285 ;
  assign n9102 = n9101 ^ n8314 ;
  assign n9112 = n9102 ^ n8339 ;
  assign n9106 = n8312 ^ n8304 ;
  assign n9107 = n8304 ^ n8275 ;
  assign n9108 = n9107 ^ n8304 ;
  assign n9109 = n9106 & ~n9108 ;
  assign n9110 = n9109 ^ n8304 ;
  assign n9111 = ~n8276 & n9110 ;
  assign n9113 = n9112 ^ n9111 ;
  assign n9114 = n9113 ^ n8335 ;
  assign n9116 = n9115 ^ n9114 ;
  assign n9117 = n9116 ^ n6558 ;
  assign n9118 = n9117 ^ n8319 ;
  assign n9100 = n9099 ^ n8287 ;
  assign n9103 = n9102 ^ n9100 ;
  assign n9095 = n8312 ^ n8287 ;
  assign n9096 = n9095 ^ n8261 ;
  assign n9097 = n9096 ^ n8319 ;
  assign n9098 = n8275 & ~n9097 ;
  assign n9104 = n9103 ^ n9098 ;
  assign n9105 = ~n8276 & n9104 ;
  assign n9119 = n9118 ^ n9105 ;
  assign n9087 = n8319 ^ n8299 ;
  assign n9088 = n9087 ^ n8275 ;
  assign n9089 = n9088 ^ n9087 ;
  assign n9092 = ~n8292 & ~n9089 ;
  assign n9093 = n9092 ^ n9087 ;
  assign n9094 = n8269 & n9093 ;
  assign n9120 = n9119 ^ n9094 ;
  assign n9121 = n9120 ^ x107 ;
  assign n9126 = ~n9042 & ~n9121 ;
  assign n9135 = n9126 & n9134 ;
  assign n9164 = n9163 ^ n9135 ;
  assign n9127 = n9126 ^ n9121 ;
  assign n9145 = n9127 ^ n9042 ;
  assign n9146 = ~n9016 & ~n9145 ;
  assign n9147 = n9146 ^ n9016 ;
  assign n9128 = n9086 & ~n9127 ;
  assign n9129 = n9128 ^ n9127 ;
  assign n9130 = n9016 & ~n9129 ;
  assign n9143 = n9130 ^ n9129 ;
  assign n9043 = ~n9016 & ~n9042 ;
  assign n9144 = n9143 ^ n9043 ;
  assign n9148 = n9147 ^ n9144 ;
  assign n9153 = n9148 ^ n9128 ;
  assign n10050 = n9164 ^ n9153 ;
  assign n10051 = n9153 ^ n8850 ;
  assign n10052 = n10051 ^ n9153 ;
  assign n10053 = n10050 & ~n10052 ;
  assign n10054 = n10053 ^ n9153 ;
  assign n10055 = n9015 & n10054 ;
  assign n9122 = ~n9086 & n9121 ;
  assign n9124 = ~n9042 & n9122 ;
  assign n9168 = n9124 ^ n9122 ;
  assign n9136 = n9043 & n9121 ;
  assign n9137 = n9136 ^ n9043 ;
  assign n9138 = n9137 ^ n9126 ;
  assign n9139 = n9138 ^ n9135 ;
  assign n9123 = n9043 & n9122 ;
  assign n9125 = n9124 ^ n9123 ;
  assign n9131 = n9130 ^ n9125 ;
  assign n9133 = n9132 ^ n9131 ;
  assign n9140 = n9139 ^ n9133 ;
  assign n9169 = n9168 ^ n9140 ;
  assign n9225 = n9169 ^ n9123 ;
  assign n9226 = n9014 & n9225 ;
  assign n9227 = n9226 ^ n9123 ;
  assign n9149 = n9148 ^ n9123 ;
  assign n10664 = n9227 ^ n9149 ;
  assign n10665 = ~n8850 & n10664 ;
  assign n9156 = n9131 ^ n8850 ;
  assign n9157 = n9156 ^ n9131 ;
  assign n9209 = n9169 ^ n9146 ;
  assign n9210 = n9209 ^ n9131 ;
  assign n9211 = ~n9157 & n9210 ;
  assign n9212 = n9211 ^ n9131 ;
  assign n9213 = ~n9015 & n9212 ;
  assign n10660 = n9213 ^ n9149 ;
  assign n9152 = n8850 & n9014 ;
  assign n9179 = n9152 ^ n9014 ;
  assign n9180 = n9179 ^ n8850 ;
  assign n10643 = n9132 ^ n9043 ;
  assign n10644 = n10643 ^ n9042 ;
  assign n10645 = ~n9180 & ~n10644 ;
  assign n9158 = n9136 ^ n9123 ;
  assign n10641 = n9158 ^ n9143 ;
  assign n9187 = n9153 ^ n9134 ;
  assign n9188 = n9187 ^ n9163 ;
  assign n9189 = n9188 ^ n9139 ;
  assign n9190 = ~n9179 & ~n9189 ;
  assign n10634 = n9190 ^ n9125 ;
  assign n10642 = n10641 ^ n10634 ;
  assign n10646 = n10645 ^ n10642 ;
  assign n9185 = n9152 ^ n8850 ;
  assign n10032 = n9153 ^ n9139 ;
  assign n10031 = n9140 ^ n9135 ;
  assign n10033 = n10032 ^ n10031 ;
  assign n10638 = ~n9190 & ~n10033 ;
  assign n10639 = n10638 ^ n9125 ;
  assign n10640 = ~n9185 & n10639 ;
  assign n10647 = n10646 ^ n10640 ;
  assign n10661 = n10660 ^ n10647 ;
  assign n9204 = n9188 ^ n8850 ;
  assign n9205 = n9204 ^ n9188 ;
  assign n9141 = n9086 & n9137 ;
  assign n9142 = n9141 ^ n9137 ;
  assign n9170 = n9169 ^ n9142 ;
  assign n10656 = n9188 ^ n9170 ;
  assign n10657 = ~n9205 & n10656 ;
  assign n10658 = n10657 ^ n9188 ;
  assign n10659 = ~n9015 & n10658 ;
  assign n10662 = n10661 ^ n10659 ;
  assign n10648 = n10647 ^ n10645 ;
  assign n10047 = n9209 ^ n9137 ;
  assign n10649 = n10648 ^ n10047 ;
  assign n10650 = n10649 ^ n10648 ;
  assign n10653 = n8850 & n10650 ;
  assign n10654 = n10653 ^ n10648 ;
  assign n10655 = ~n9015 & n10654 ;
  assign n10663 = n10662 ^ n10655 ;
  assign n10666 = n10665 ^ n10663 ;
  assign n10667 = ~n10055 & ~n10666 ;
  assign n10668 = n10667 ^ n7373 ;
  assign n11289 = n10668 ^ x100 ;
  assign n11290 = ~n11288 & n11289 ;
  assign n9359 = n9358 ^ n8972 ;
  assign n9360 = n9359 ^ n8988 ;
  assign n9349 = n8964 ^ n8955 ;
  assign n9351 = n9350 ^ n9349 ;
  assign n9352 = n9351 ^ n8993 ;
  assign n9353 = ~n8851 & n9352 ;
  assign n9361 = n9360 ^ n9353 ;
  assign n9354 = n8986 ^ n8951 ;
  assign n9357 = n9356 ^ n9354 ;
  assign n9362 = n9361 ^ n9357 ;
  assign n9363 = n9362 ^ n9353 ;
  assign n9364 = ~n8851 & ~n9363 ;
  assign n9365 = n9364 ^ n9361 ;
  assign n9366 = n8852 & ~n9365 ;
  assign n9367 = n9366 ^ n9353 ;
  assign n9346 = n8985 ^ n8964 ;
  assign n9347 = n9346 ^ n8976 ;
  assign n9348 = n8855 & ~n9347 ;
  assign n9368 = n9367 ^ n9348 ;
  assign n9369 = n9368 ^ n8939 ;
  assign n9345 = n8942 & n8948 ;
  assign n9370 = n9369 ^ n9345 ;
  assign n9377 = ~n9370 & ~n9376 ;
  assign n9378 = n9377 ^ n6232 ;
  assign n10004 = n9378 ^ x81 ;
  assign n9922 = n9623 ^ x99 ;
  assign n9956 = n9535 ^ x106 ;
  assign n9290 = n8275 & n8286 ;
  assign n9281 = n8297 ^ n8275 ;
  assign n9282 = n9281 ^ n8297 ;
  assign n9284 = n8304 & n9282 ;
  assign n9285 = n9284 ^ n8297 ;
  assign n9286 = ~n8269 & n9285 ;
  assign n9287 = n9286 ^ n9111 ;
  assign n9271 = n8267 ^ n8261 ;
  assign n9272 = n8265 ^ n8236 ;
  assign n9273 = ~n8275 & ~n9272 ;
  assign n9274 = n9271 & n9273 ;
  assign n9280 = n9274 ^ n8297 ;
  assign n9288 = n9287 ^ n9280 ;
  assign n9289 = n9288 ^ n8289 ;
  assign n9291 = n9290 ^ n9289 ;
  assign n9299 = n9291 ^ n9115 ;
  assign n9294 = n8309 ^ n8299 ;
  assign n9295 = n9294 ^ n9099 ;
  assign n9296 = ~n8269 & ~n9295 ;
  assign n9276 = n9099 ^ n8299 ;
  assign n9278 = n9277 ^ n9276 ;
  assign n9275 = n9274 ^ n8329 ;
  assign n9279 = n9278 ^ n9275 ;
  assign n9292 = n9291 ^ n9279 ;
  assign n9293 = n9292 ^ n9288 ;
  assign n9297 = n9296 ^ n9293 ;
  assign n9298 = n8276 & n9297 ;
  assign n9300 = n9299 ^ n9298 ;
  assign n9301 = ~n8320 & ~n9300 ;
  assign n9302 = n9301 ^ n6306 ;
  assign n9923 = n9302 ^ x123 ;
  assign n10016 = n9956 ^ n9923 ;
  assign n9947 = n6876 ^ n6680 ;
  assign n9948 = n6873 & ~n9947 ;
  assign n9930 = ~n6856 & ~n8716 ;
  assign n9931 = n9930 ^ n8715 ;
  assign n9925 = n6863 ^ n6677 ;
  assign n9926 = n9925 ^ n6856 ;
  assign n9928 = n6666 & ~n9926 ;
  assign n9929 = n9928 ^ n9926 ;
  assign n9932 = n9931 ^ n9929 ;
  assign n9940 = n9931 ^ n5380 ;
  assign n9937 = n6689 & ~n6856 ;
  assign n9938 = n9937 ^ n6668 ;
  assign n9939 = n5380 & n9938 ;
  assign n9941 = n9940 ^ n9939 ;
  assign n9942 = n9941 ^ n6856 ;
  assign n9943 = n9942 ^ n9929 ;
  assign n9944 = n9943 ^ n9939 ;
  assign n9945 = ~n9932 & ~n9944 ;
  assign n9946 = n9945 ^ n9941 ;
  assign n9951 = n9948 ^ n9946 ;
  assign n9952 = ~n6875 & n9951 ;
  assign n9924 = n6907 ^ n6339 ;
  assign n9953 = n9952 ^ n9924 ;
  assign n9954 = n9953 ^ x105 ;
  assign n10005 = n9956 ^ n9954 ;
  assign n9961 = n7607 ^ n7595 ;
  assign n9972 = n9961 ^ n7479 ;
  assign n9973 = n9972 ^ n7610 ;
  assign n9971 = n7519 ^ n7476 ;
  assign n9974 = n9973 ^ n9971 ;
  assign n9975 = n9974 ^ n8445 ;
  assign n9976 = ~n7398 & n9975 ;
  assign n9977 = n9976 ^ n8445 ;
  assign n9978 = n7374 & n9977 ;
  assign n9957 = n7596 ^ n7578 ;
  assign n9958 = n9957 ^ n7606 ;
  assign n9959 = n9958 ^ n7583 ;
  assign n9960 = ~n7374 & n9959 ;
  assign n9963 = n9960 ^ n7601 ;
  assign n9962 = n9961 ^ n9960 ;
  assign n9964 = n9963 ^ n9962 ;
  assign n9967 = ~n7374 & ~n9964 ;
  assign n9968 = n9967 ^ n9963 ;
  assign n9969 = n7398 & n9968 ;
  assign n9970 = n9969 ^ n9960 ;
  assign n9979 = n9978 ^ n9970 ;
  assign n9982 = n7398 & n7578 ;
  assign n9983 = n9982 ^ n7593 ;
  assign n9984 = n9232 & n9983 ;
  assign n9985 = n9984 ^ n7593 ;
  assign n9986 = ~n9979 & n9985 ;
  assign n9987 = n9986 ^ n9979 ;
  assign n9988 = ~n9266 & ~n9987 ;
  assign n9989 = ~n8457 & n9988 ;
  assign n9990 = n9989 ^ n6394 ;
  assign n9991 = n9990 ^ x96 ;
  assign n10014 = n10005 ^ n9991 ;
  assign n10017 = ~n9923 & n10014 ;
  assign n10001 = n9991 ^ n9956 ;
  assign n10018 = n10017 ^ n10001 ;
  assign n10019 = ~n10016 & n10018 ;
  assign n10006 = n10005 ^ n9923 ;
  assign n10010 = n9954 & n10006 ;
  assign n10011 = n10010 ^ n9923 ;
  assign n10012 = n9991 & ~n10011 ;
  assign n10013 = n10012 ^ n10006 ;
  assign n10015 = n10014 ^ n10013 ;
  assign n10020 = n10019 ^ n10015 ;
  assign n10021 = ~n9922 & ~n10020 ;
  assign n10022 = n10021 ^ n10013 ;
  assign n9997 = n9991 ^ n9954 ;
  assign n9998 = ~n9954 & n9956 ;
  assign n9999 = n9998 ^ n9923 ;
  assign n10000 = n9997 & ~n9999 ;
  assign n10002 = n10001 ^ n10000 ;
  assign n9955 = n9954 ^ n9923 ;
  assign n9992 = n9956 & ~n9991 ;
  assign n9993 = n9992 ^ n9954 ;
  assign n9994 = n9955 & n9993 ;
  assign n9995 = n9994 ^ n9954 ;
  assign n9996 = n9922 & ~n9995 ;
  assign n10003 = n10002 ^ n9996 ;
  assign n10023 = n10022 ^ n10003 ;
  assign n10024 = n10004 & n10023 ;
  assign n10025 = n10024 ^ n10022 ;
  assign n11293 = n10025 ^ n8502 ;
  assign n11294 = n11293 ^ x91 ;
  assign n9303 = n9302 ^ x91 ;
  assign n9270 = n9269 ^ x109 ;
  assign n9304 = n9303 ^ n9270 ;
  assign n9313 = n8119 ^ n8116 ;
  assign n9312 = n8152 ^ n8149 ;
  assign n9314 = n9313 ^ n9312 ;
  assign n9315 = ~n8003 & n9314 ;
  assign n9316 = n9315 ^ n9313 ;
  assign n9328 = n9316 ^ n8191 ;
  assign n9321 = n8160 ^ n8150 ;
  assign n9320 = n8156 ^ n8127 ;
  assign n9322 = n9321 ^ n9320 ;
  assign n9323 = n9320 ^ n8003 ;
  assign n9324 = n9323 ^ n9320 ;
  assign n9325 = n9322 & n9324 ;
  assign n9326 = n9325 ^ n9320 ;
  assign n9327 = ~n8198 & ~n9326 ;
  assign n9329 = n9328 ^ n9327 ;
  assign n9310 = n8183 ^ n8158 ;
  assign n9311 = n9310 ^ n8161 ;
  assign n9317 = n9316 ^ n9311 ;
  assign n9306 = n8147 ^ n8116 ;
  assign n9307 = n9306 ^ n8158 ;
  assign n9308 = n9307 ^ n8183 ;
  assign n9309 = ~n8003 & ~n9308 ;
  assign n9318 = n9317 ^ n9309 ;
  assign n9319 = n8198 & n9318 ;
  assign n9330 = n9329 ^ n9319 ;
  assign n9305 = n8122 & n8194 ;
  assign n9331 = n9330 ^ n9305 ;
  assign n9332 = n9331 ^ n9327 ;
  assign n9333 = n9331 ^ n8128 ;
  assign n9334 = n9333 ^ n9331 ;
  assign n9335 = n9331 ^ n7978 ;
  assign n9336 = n9335 ^ n9331 ;
  assign n9337 = n9334 & ~n9336 ;
  assign n9338 = ~n9332 & n9337 ;
  assign n9339 = n9338 ^ n9332 ;
  assign n9340 = n9339 ^ n9327 ;
  assign n9341 = ~n8189 & ~n8632 ;
  assign n9342 = ~n9340 & n9341 ;
  assign n9343 = n9342 ^ n7123 ;
  assign n9344 = n9343 ^ x92 ;
  assign n9379 = n9378 ^ x70 ;
  assign n9380 = n9344 & n9379 ;
  assign n9381 = n9380 ^ n9379 ;
  assign n9382 = n9381 ^ n9344 ;
  assign n9387 = n9386 ^ x110 ;
  assign n9391 = n7955 ^ n7908 ;
  assign n9390 = n7926 ^ n7879 ;
  assign n9392 = n9391 ^ n9390 ;
  assign n9393 = n9391 ^ n7725 ;
  assign n9394 = n9393 ^ n9391 ;
  assign n9395 = n9392 & n9394 ;
  assign n9396 = n9395 ^ n9391 ;
  assign n9397 = n7945 & n9396 ;
  assign n9402 = n9397 ^ n7915 ;
  assign n9400 = n9398 ^ n7910 ;
  assign n9401 = n7728 & ~n9400 ;
  assign n9403 = n9402 ^ n9401 ;
  assign n9399 = n7905 & ~n9398 ;
  assign n9404 = n9403 ^ n9399 ;
  assign n9413 = n9404 ^ n7953 ;
  assign n9405 = n9404 ^ n9397 ;
  assign n8646 = n7919 ^ n7879 ;
  assign n9406 = n9405 ^ n8646 ;
  assign n9407 = n9406 ^ n9405 ;
  assign n9408 = n9405 ^ n7688 ;
  assign n9409 = n9408 ^ n9405 ;
  assign n9410 = n9407 & ~n9409 ;
  assign n9411 = n9410 ^ n9405 ;
  assign n9412 = ~n7725 & n9411 ;
  assign n9414 = n9413 ^ n9412 ;
  assign n9388 = n8646 ^ n7885 ;
  assign n9389 = n7726 & n9388 ;
  assign n9415 = n9414 ^ n9389 ;
  assign n9416 = n7725 & ~n9415 ;
  assign n9417 = ~n7893 & n9416 ;
  assign n9419 = n9417 ^ n9415 ;
  assign n9420 = ~n8674 & ~n9419 ;
  assign n9429 = n9420 ^ n7147 ;
  assign n9418 = n9417 ^ n7945 ;
  assign n8648 = n7910 ^ n7909 ;
  assign n9421 = n8648 ^ n7961 ;
  assign n9422 = n9421 ^ n7884 ;
  assign n9423 = n7884 ^ n7725 ;
  assign n9424 = n9423 ^ n7884 ;
  assign n9425 = n9422 & ~n9424 ;
  assign n9426 = n9425 ^ n7884 ;
  assign n9427 = n9420 & n9426 ;
  assign n9428 = ~n9418 & n9427 ;
  assign n9430 = n9429 ^ n9428 ;
  assign n9431 = n9430 ^ x77 ;
  assign n9432 = ~n9387 & ~n9431 ;
  assign n9447 = ~n9382 & n9432 ;
  assign n9453 = n9447 ^ n9382 ;
  assign n9438 = n9432 ^ n9431 ;
  assign n9439 = n9438 ^ n9387 ;
  assign n9440 = ~n9382 & ~n9439 ;
  assign n9433 = n9432 ^ n9387 ;
  assign n9434 = ~n9382 & ~n9433 ;
  assign n9452 = n9440 ^ n9434 ;
  assign n9454 = n9453 ^ n9452 ;
  assign n9450 = n9380 & ~n9433 ;
  assign n11135 = n9454 ^ n9450 ;
  assign n11136 = n9450 ^ n9303 ;
  assign n11137 = n11136 ^ n9450 ;
  assign n11138 = ~n11135 & ~n11137 ;
  assign n11139 = n11138 ^ n9450 ;
  assign n11140 = n9304 & n11139 ;
  assign n9460 = n9381 & n9432 ;
  assign n9461 = n9460 ^ n9381 ;
  assign n9462 = n9461 ^ n9379 ;
  assign n9463 = n9439 & n9462 ;
  assign n9464 = n9463 ^ n9462 ;
  assign n11309 = n9464 ^ n9452 ;
  assign n11313 = n11309 ^ n9461 ;
  assign n9435 = n9382 ^ n9379 ;
  assign n9442 = n9435 & ~n9438 ;
  assign n9472 = n9442 ^ n9434 ;
  assign n10772 = n9472 ^ n9447 ;
  assign n11112 = n10772 ^ n9450 ;
  assign n11308 = n11112 ^ n9442 ;
  assign n11310 = n11309 ^ n11308 ;
  assign n9485 = n9380 & n9432 ;
  assign n9486 = n9485 ^ n9464 ;
  assign n9473 = n9472 ^ n9450 ;
  assign n9441 = ~n9433 & n9435 ;
  assign n9443 = n9442 ^ n9441 ;
  assign n9471 = n9443 ^ n9433 ;
  assign n9474 = n9473 ^ n9471 ;
  assign n9436 = n9432 & n9435 ;
  assign n9455 = n9436 ^ n9435 ;
  assign n9456 = n9455 ^ n9443 ;
  assign n9458 = n9456 ^ n9440 ;
  assign n9459 = n9458 ^ n9439 ;
  assign n9465 = n9464 ^ n9459 ;
  assign n9475 = n9474 ^ n9465 ;
  assign n9476 = n9475 ^ n9461 ;
  assign n9489 = n9486 ^ n9476 ;
  assign n11311 = n11310 ^ n9489 ;
  assign n11312 = n9270 & n11311 ;
  assign n11314 = n11313 ^ n11312 ;
  assign n11315 = ~n9303 & n11314 ;
  assign n11306 = n9270 & n9442 ;
  assign n11299 = n9485 ^ n9463 ;
  assign n11300 = n9463 ^ n9270 ;
  assign n11301 = n11300 ^ n9463 ;
  assign n11302 = n11299 & n11301 ;
  assign n11303 = n11302 ^ n9463 ;
  assign n11304 = ~n9304 & n11303 ;
  assign n11305 = n11304 ^ n9461 ;
  assign n11307 = n11306 ^ n11305 ;
  assign n11316 = n11315 ^ n11307 ;
  assign n9497 = ~n9270 & n9303 ;
  assign n11298 = n9458 & n9497 ;
  assign n11317 = n11316 ^ n11298 ;
  assign n11297 = n9303 & n9447 ;
  assign n11318 = n11317 ^ n11297 ;
  assign n11319 = ~n11140 & ~n11318 ;
  assign n9498 = n9436 & n9497 ;
  assign n11295 = n9498 ^ n8002 ;
  assign n10740 = n9497 ^ n9270 ;
  assign n10741 = n10740 ^ n9303 ;
  assign n10742 = n10741 ^ n9270 ;
  assign n10782 = n10742 ^ n9441 ;
  assign n10783 = n10740 ^ n9440 ;
  assign n10784 = n10740 ^ n9441 ;
  assign n10785 = n10784 ^ n10740 ;
  assign n10786 = n10783 & ~n10785 ;
  assign n10787 = n10786 ^ n10740 ;
  assign n10788 = n10782 & ~n10787 ;
  assign n10789 = n10788 ^ n10742 ;
  assign n11296 = n11295 ^ n10789 ;
  assign n11320 = n11319 ^ n11296 ;
  assign n11321 = n11320 ^ x78 ;
  assign n11322 = ~n11294 & ~n11321 ;
  assign n11343 = n11290 & n11322 ;
  assign n11291 = n11290 ^ n11289 ;
  assign n11292 = n11291 ^ n11288 ;
  assign n11342 = n11292 & n11322 ;
  assign n11344 = n11343 ^ n11342 ;
  assign n11323 = n11322 ^ n11321 ;
  assign n11327 = n11291 & ~n11323 ;
  assign n11328 = n11327 ^ n11323 ;
  assign n11345 = n11344 ^ n11328 ;
  assign n11330 = n11290 ^ n11288 ;
  assign n11331 = n11322 & ~n11330 ;
  assign n11332 = n11331 ^ n11327 ;
  assign n11341 = n11332 ^ n11321 ;
  assign n11346 = n11345 ^ n11341 ;
  assign n11347 = n11346 ^ n11331 ;
  assign n11414 = n11265 & n11347 ;
  assign n11578 = n11414 ^ n8587 ;
  assign n11348 = n11322 ^ n11294 ;
  assign n11349 = n11290 & ~n11348 ;
  assign n11350 = n11349 ^ n11347 ;
  assign n11337 = ~n11288 & ~n11321 ;
  assign n11338 = n11337 ^ n11289 ;
  assign n11339 = n11294 & n11338 ;
  assign n11340 = n11339 ^ n11338 ;
  assign n11351 = n11350 ^ n11340 ;
  assign n11376 = n11351 ^ n11348 ;
  assign n11361 = n11292 & ~n11348 ;
  assign n11362 = n11361 ^ n11349 ;
  assign n11377 = n11376 ^ n11362 ;
  assign n11359 = n11339 ^ n11331 ;
  assign n11335 = n11323 ^ n11294 ;
  assign n11336 = ~n11330 & ~n11335 ;
  assign n11352 = n11351 ^ n11336 ;
  assign n11325 = n11290 & ~n11323 ;
  assign n11354 = n11352 ^ n11325 ;
  assign n11355 = n11354 ^ n11342 ;
  assign n11353 = n11352 ^ n11350 ;
  assign n11356 = n11355 ^ n11353 ;
  assign n11334 = n11322 ^ n11290 ;
  assign n11357 = n11356 ^ n11334 ;
  assign n11324 = n11292 & ~n11323 ;
  assign n11326 = n11325 ^ n11324 ;
  assign n11329 = n11328 ^ n11326 ;
  assign n11333 = n11332 ^ n11329 ;
  assign n11358 = n11357 ^ n11333 ;
  assign n11360 = n11359 ^ n11358 ;
  assign n11572 = n11377 ^ n11360 ;
  assign n11573 = n11377 ^ n11264 ;
  assign n11574 = n11573 ^ n11377 ;
  assign n11575 = n11572 & ~n11574 ;
  assign n11576 = n11575 ^ n11377 ;
  assign n11577 = n11239 & ~n11576 ;
  assign n11579 = n11578 ^ n11577 ;
  assign n11391 = n11325 ^ n11264 ;
  assign n11392 = n11391 ^ n11325 ;
  assign n11393 = n11326 & n11392 ;
  assign n11394 = n11393 ^ n11325 ;
  assign n11395 = n11239 & n11394 ;
  assign n11372 = n11265 ^ n11264 ;
  assign n11266 = n11265 ^ n11239 ;
  assign n11373 = n11372 ^ n11266 ;
  assign n11568 = n11362 & n11373 ;
  assign n11564 = n11327 ^ n11324 ;
  assign n11565 = n11564 ^ n11352 ;
  assign n11566 = n11265 & n11565 ;
  assign n11550 = n11342 ^ n11332 ;
  assign n11551 = n11550 ^ n11336 ;
  assign n11547 = n11360 ^ n11344 ;
  assign n11548 = n11547 ^ n11352 ;
  assign n11549 = n11548 ^ n11346 ;
  assign n11552 = n11551 ^ n11549 ;
  assign n11553 = n11264 & ~n11552 ;
  assign n11554 = n11553 ^ n11551 ;
  assign n11567 = n11566 ^ n11554 ;
  assign n11569 = n11568 ^ n11567 ;
  assign n11555 = n11554 ^ n11264 ;
  assign n11556 = n11555 ^ n11554 ;
  assign n11557 = n11548 ^ n11325 ;
  assign n11558 = n11557 ^ n11332 ;
  assign n11561 = ~n11556 & n11558 ;
  assign n11562 = n11561 ^ n11554 ;
  assign n11563 = ~n11239 & n11562 ;
  assign n11570 = n11569 ^ n11563 ;
  assign n11571 = ~n11395 & ~n11570 ;
  assign n11580 = n11579 ^ n11571 ;
  assign n13147 = n11580 ^ x69 ;
  assign n10743 = n9456 & n10742 ;
  assign n10744 = n10743 ^ n9498 ;
  assign n10745 = n9485 ^ n9461 ;
  assign n10746 = n10741 & n10745 ;
  assign n10747 = n9464 ^ n9454 ;
  assign n10748 = ~n10740 & ~n10747 ;
  assign n10753 = n9303 & ~n9450 ;
  assign n10754 = n9474 ^ n9447 ;
  assign n9484 = n9450 ^ n9380 ;
  assign n9487 = n9486 ^ n9484 ;
  assign n10755 = n10754 ^ n9487 ;
  assign n9466 = n9465 ^ n9460 ;
  assign n9467 = n9466 ^ n9464 ;
  assign n10756 = n10755 ^ n9467 ;
  assign n10757 = n9270 & n10756 ;
  assign n10758 = n10757 ^ n9467 ;
  assign n10759 = n10753 & n10758 ;
  assign n10760 = n10759 ^ n9303 ;
  assign n10751 = n9465 ^ n9381 ;
  assign n10752 = ~n10740 & ~n10751 ;
  assign n10761 = n10760 ^ n10752 ;
  assign n9457 = n9456 ^ n9454 ;
  assign n10749 = n9457 ^ n9434 ;
  assign n10750 = n10741 & ~n10749 ;
  assign n10762 = n10761 ^ n10750 ;
  assign n10763 = n9487 ^ n9441 ;
  assign n10764 = n9441 ^ n9270 ;
  assign n10765 = n10764 ^ n9441 ;
  assign n10766 = n10763 & ~n10765 ;
  assign n10767 = n10766 ^ n9441 ;
  assign n10768 = ~n9303 & n10767 ;
  assign n10769 = ~n10762 & ~n10768 ;
  assign n10770 = ~n10748 & n10769 ;
  assign n10771 = ~n10746 & n10770 ;
  assign n10775 = n9436 ^ n9270 ;
  assign n10776 = n10775 ^ n9436 ;
  assign n10777 = n10772 & ~n10776 ;
  assign n10778 = n10777 ^ n9436 ;
  assign n10779 = n9304 & n10778 ;
  assign n10780 = n10779 ^ n9436 ;
  assign n10781 = n10771 & ~n10780 ;
  assign n10790 = n10781 & ~n10789 ;
  assign n10791 = ~n10744 & n10790 ;
  assign n10792 = n10791 ^ n7776 ;
  assign n10793 = n10792 ^ x121 ;
  assign n10620 = n9997 ^ n9991 ;
  assign n10621 = ~n10014 & ~n10620 ;
  assign n10622 = n10621 ^ n9991 ;
  assign n10623 = n10006 & n10622 ;
  assign n10624 = n10623 ^ n9923 ;
  assign n10611 = n10013 ^ n10000 ;
  assign n10608 = n10017 ^ n9954 ;
  assign n10609 = n10016 & ~n10608 ;
  assign n10610 = n10609 ^ n10014 ;
  assign n10612 = n10611 ^ n10610 ;
  assign n10607 = n9991 ^ n9923 ;
  assign n10613 = n10612 ^ n10607 ;
  assign n10863 = n10624 ^ n10613 ;
  assign n10614 = n10613 ^ n10610 ;
  assign n10864 = n10863 ^ n10614 ;
  assign n10865 = n10614 ^ n10004 ;
  assign n10866 = n10865 ^ n10614 ;
  assign n10867 = ~n10864 & n10866 ;
  assign n10868 = n10867 ^ n10614 ;
  assign n10869 = n9922 & ~n10868 ;
  assign n10599 = ~n9923 & ~n9954 ;
  assign n10600 = n10001 & n10599 ;
  assign n10861 = n10600 ^ n8235 ;
  assign n10862 = n10861 ^ n10613 ;
  assign n10870 = n10869 ^ n10862 ;
  assign n10853 = n10613 ^ n10600 ;
  assign n10602 = n9998 ^ n9954 ;
  assign n10603 = n10602 ^ n10599 ;
  assign n10604 = n10603 ^ n9923 ;
  assign n10605 = ~n9991 & ~n10604 ;
  assign n10606 = n10605 ^ n10006 ;
  assign n10854 = n10853 ^ n10606 ;
  assign n10855 = n10854 ^ n10600 ;
  assign n10856 = n10600 ^ n9922 ;
  assign n10857 = n10856 ^ n10600 ;
  assign n10858 = n10855 & ~n10857 ;
  assign n10859 = n10858 ^ n10600 ;
  assign n10860 = ~n10004 & n10859 ;
  assign n10871 = n10870 ^ n10860 ;
  assign n10872 = n10871 ^ x115 ;
  assign n10166 = ~n10081 & n10165 ;
  assign n10844 = n10204 ^ n10166 ;
  assign n10829 = n10456 ^ n10187 ;
  assign n10830 = ~n10080 & ~n10181 ;
  assign n10831 = ~n10178 & ~n10830 ;
  assign n10832 = n10829 & n10831 ;
  assign n10833 = n10832 ^ n10830 ;
  assign n10845 = n10844 ^ n10833 ;
  assign n10846 = n10845 ^ n10451 ;
  assign n10835 = n10184 ^ n10115 ;
  assign n10836 = n10835 ^ n10169 ;
  assign n10837 = n10836 ^ n10833 ;
  assign n10834 = n10833 ^ n10172 ;
  assign n10838 = n10837 ^ n10834 ;
  assign n10839 = n10837 ^ n10078 ;
  assign n10840 = n10839 ^ n10837 ;
  assign n10841 = ~n10838 & n10840 ;
  assign n10842 = n10841 ^ n10837 ;
  assign n10843 = n10077 & n10842 ;
  assign n10847 = n10846 ^ n10843 ;
  assign n10822 = n10204 ^ n10078 ;
  assign n10823 = n10822 ^ n10204 ;
  assign n10824 = n10204 ^ n10156 ;
  assign n10825 = n10824 ^ n10204 ;
  assign n10826 = n10823 & n10825 ;
  assign n10827 = n10826 ^ n10204 ;
  assign n10828 = n10202 & ~n10827 ;
  assign n10848 = n10847 ^ n10828 ;
  assign n10849 = ~n10440 & ~n10848 ;
  assign n10850 = ~n10475 & n10849 ;
  assign n10851 = n10850 ^ n8260 ;
  assign n10852 = n10851 ^ x114 ;
  assign n6910 = n6909 ^ x94 ;
  assign n7633 = n7611 ^ n7596 ;
  assign n7629 = ~n7594 & n7625 ;
  assign n7632 = n7613 & ~n7629 ;
  assign n7634 = n7633 ^ n7632 ;
  assign n7635 = n7634 ^ n7604 ;
  assign n7636 = n7635 ^ n7598 ;
  assign n7637 = n7636 ^ n7615 ;
  assign n7638 = n7637 ^ n7634 ;
  assign n7639 = n7374 & ~n7638 ;
  assign n7640 = n7639 ^ n7635 ;
  assign n7641 = n7626 & n7640 ;
  assign n7642 = n7641 ^ n7634 ;
  assign n7628 = n7600 ^ n7578 ;
  assign n7630 = n7629 ^ n7628 ;
  assign n7631 = n7624 & ~n7630 ;
  assign n7643 = n7642 ^ n7631 ;
  assign n7627 = n7605 & ~n7626 ;
  assign n7644 = n7643 ^ n7627 ;
  assign n7645 = n7594 ^ n7582 ;
  assign n7646 = ~n7398 & n7645 ;
  assign n7647 = n7646 ^ n7594 ;
  assign n7648 = n7647 ^ n7374 ;
  assign n7649 = n7648 ^ n7647 ;
  assign n7651 = ~n7398 & n7650 ;
  assign n7652 = n7651 ^ n7647 ;
  assign n7653 = n7649 & n7652 ;
  assign n7654 = n7653 ^ n7647 ;
  assign n7655 = ~n7644 & n7654 ;
  assign n7656 = n7655 ^ n7644 ;
  assign n7657 = ~n7622 & ~n7656 ;
  assign n7658 = n7657 ^ n6935 ;
  assign n7659 = n7658 ^ x101 ;
  assign n8355 = ~n6910 & ~n7659 ;
  assign n8356 = n8355 ^ n7659 ;
  assign n7974 = n7973 ^ x116 ;
  assign n7338 = n7337 ^ n6941 ;
  assign n7339 = n7338 ^ x76 ;
  assign n8349 = n7974 ^ n7339 ;
  assign n8348 = ~n7339 & ~n7974 ;
  assign n8350 = n8349 ^ n8348 ;
  assign n8351 = n8350 ^ n7339 ;
  assign n8352 = n6910 & ~n8351 ;
  assign n8353 = ~n7659 & n8352 ;
  assign n8346 = n6910 & ~n7339 ;
  assign n8347 = ~n7659 & n8346 ;
  assign n8354 = n8353 ^ n8347 ;
  assign n8357 = n8356 ^ n8354 ;
  assign n8215 = n8214 ^ x125 ;
  assign n8343 = n8342 ^ x67 ;
  assign n8358 = n8215 & n8343 ;
  assign n8359 = n8358 ^ n8215 ;
  assign n8360 = ~n8357 & n8359 ;
  assign n7975 = n7659 & n7974 ;
  assign n7976 = ~n7339 & n7975 ;
  assign n7977 = ~n6910 & n7976 ;
  assign n8344 = n8343 ^ n8215 ;
  assign n8345 = n7977 & ~n8344 ;
  assign n8361 = n8360 ^ n8345 ;
  assign n8390 = n7977 ^ n7976 ;
  assign n8396 = n8390 ^ n8346 ;
  assign n8362 = ~n7974 & n8346 ;
  assign n8397 = n8396 ^ n8362 ;
  assign n8388 = n8353 ^ n8352 ;
  assign n8391 = n8390 ^ n8388 ;
  assign n8392 = n8391 ^ n8347 ;
  assign n8393 = n8392 ^ n8346 ;
  assign n8394 = n8393 ^ n8352 ;
  assign n8368 = ~n8350 & n8355 ;
  assign n8389 = n8388 ^ n8368 ;
  assign n8395 = n8394 ^ n8389 ;
  assign n8398 = n8397 ^ n8395 ;
  assign n8399 = n8215 & n8398 ;
  assign n8364 = n8348 & n8355 ;
  assign n8369 = n8368 ^ n8364 ;
  assign n8366 = ~n8351 & n8355 ;
  assign n8367 = n8366 ^ n8355 ;
  assign n8370 = n8369 ^ n8367 ;
  assign n8403 = n8399 ^ n8370 ;
  assign n8363 = n8362 ^ n8348 ;
  assign n8400 = n8363 ^ n8356 ;
  assign n8401 = n8400 ^ n7974 ;
  assign n8402 = ~n8215 & n8401 ;
  assign n8404 = n8403 ^ n8402 ;
  assign n8405 = ~n8344 & n8404 ;
  assign n8406 = n8405 ^ n8399 ;
  assign n8379 = n8352 ^ n8351 ;
  assign n8380 = n8379 ^ n8366 ;
  assign n8373 = n7976 ^ n7975 ;
  assign n8374 = ~n6910 & n8373 ;
  assign n8375 = n8374 ^ n8373 ;
  assign n8376 = n8375 ^ n8362 ;
  assign n8377 = n8376 ^ n8357 ;
  assign n8365 = n8364 ^ n8363 ;
  assign n8371 = n8370 ^ n8365 ;
  assign n8372 = n8371 ^ n8353 ;
  assign n8378 = n8377 ^ n8372 ;
  assign n8381 = n8380 ^ n8378 ;
  assign n8382 = n8381 ^ n8377 ;
  assign n8383 = n8377 ^ n8215 ;
  assign n8384 = n8383 ^ n8377 ;
  assign n8385 = n8382 & ~n8384 ;
  assign n8386 = n8385 ^ n8377 ;
  assign n8387 = n8343 & ~n8386 ;
  assign n8407 = n8406 ^ n8387 ;
  assign n8408 = ~n8361 & ~n8407 ;
  assign n8410 = n8374 ^ n8365 ;
  assign n8409 = n8380 ^ n8368 ;
  assign n8411 = n8410 ^ n8409 ;
  assign n8412 = n8410 ^ n8343 ;
  assign n8413 = n8412 ^ n8410 ;
  assign n8414 = ~n8411 & n8413 ;
  assign n8415 = n8414 ^ n8410 ;
  assign n8416 = n8215 & n8415 ;
  assign n8417 = n8408 & ~n8416 ;
  assign n8418 = n8417 ^ n7033 ;
  assign n10794 = n8418 ^ x97 ;
  assign n8705 = n8704 ^ x120 ;
  assign n8710 = n8709 ^ n6661 ;
  assign n8711 = ~n6872 & n8710 ;
  assign n8730 = n6872 ^ n6690 ;
  assign n8731 = n8730 ^ n6885 ;
  assign n8732 = n8731 ^ n8709 ;
  assign n8733 = n6680 & ~n8732 ;
  assign n8734 = n8733 ^ n6872 ;
  assign n8735 = n6874 ^ n6680 ;
  assign n8736 = ~n8734 & ~n8735 ;
  assign n8712 = n6878 ^ n6696 ;
  assign n8718 = n8717 ^ n8712 ;
  assign n8719 = ~n5380 & ~n8718 ;
  assign n8720 = n8719 ^ n6696 ;
  assign n8721 = n8720 ^ n6856 ;
  assign n8722 = n8721 ^ n8720 ;
  assign n8723 = n8720 ^ n6683 ;
  assign n8724 = n8723 ^ n6668 ;
  assign n8725 = n8724 ^ n8720 ;
  assign n8726 = ~n8722 & ~n8725 ;
  assign n8727 = n8726 ^ n8720 ;
  assign n8728 = ~n6862 & ~n8727 ;
  assign n8729 = n8728 ^ n8720 ;
  assign n8737 = n8736 ^ n8729 ;
  assign n8738 = ~n6907 & ~n8737 ;
  assign n8739 = ~n8711 & n8738 ;
  assign n8740 = n6862 ^ n6684 ;
  assign n8741 = n6681 ^ n6200 ;
  assign n8742 = n8741 ^ n6684 ;
  assign n8743 = ~n5380 & n8742 ;
  assign n8744 = n8743 ^ n6685 ;
  assign n8745 = n8740 & n8744 ;
  assign n8746 = n8745 ^ n6684 ;
  assign n8747 = n8739 & ~n8746 ;
  assign n8748 = ~n8707 & n8747 ;
  assign n8749 = n8748 ^ n6017 ;
  assign n8750 = n8749 ^ x64 ;
  assign n8751 = ~n8705 & ~n8750 ;
  assign n8753 = n8751 ^ n8705 ;
  assign n8759 = n8753 ^ n8750 ;
  assign n8635 = n8634 ^ x89 ;
  assign n8650 = n7902 ^ n7890 ;
  assign n8651 = n8650 ^ n7882 ;
  assign n8652 = n8651 ^ n8648 ;
  assign n8647 = n8646 ^ n7961 ;
  assign n8649 = n8648 ^ n8647 ;
  assign n8653 = n8652 ^ n8649 ;
  assign n8654 = n8649 ^ n8648 ;
  assign n8655 = n8654 ^ n7725 ;
  assign n8656 = ~n7945 & n8655 ;
  assign n8657 = n8656 ^ n7725 ;
  assign n8658 = ~n8653 & ~n8657 ;
  assign n8659 = n8658 ^ n8652 ;
  assign n8660 = ~n7907 & n8659 ;
  assign n8661 = n7893 & n8660 ;
  assign n8643 = n7926 ^ n7910 ;
  assign n8644 = n8643 ^ n7905 ;
  assign n8645 = n7725 & n8644 ;
  assign n8662 = n8661 ^ n8645 ;
  assign n8663 = ~n7945 & ~n8662 ;
  assign n8664 = n8663 ^ n8661 ;
  assign n8636 = n7901 ^ n7889 ;
  assign n8637 = n8636 ^ n7912 ;
  assign n8638 = n7912 ^ n7725 ;
  assign n8639 = n8638 ^ n7912 ;
  assign n8640 = ~n8637 & ~n8639 ;
  assign n8641 = n8640 ^ n7912 ;
  assign n8642 = ~n7688 & n8641 ;
  assign n8665 = n8664 ^ n8642 ;
  assign n8667 = n8666 ^ n8665 ;
  assign n8677 = n8676 ^ n8667 ;
  assign n8678 = n8677 ^ n7951 ;
  assign n8679 = n8678 ^ n6108 ;
  assign n8680 = n8679 ^ x74 ;
  assign n8681 = ~n8635 & n8680 ;
  assign n8682 = n8681 ^ n8680 ;
  assign n8764 = n8682 ^ n8635 ;
  assign n8800 = ~n8759 & n8764 ;
  assign n8588 = n8587 ^ x115 ;
  assign n8460 = n8459 ^ x122 ;
  assign n8589 = n8588 ^ n8460 ;
  assign n8760 = n8682 & ~n8759 ;
  assign n10815 = ~n8589 & n8760 ;
  assign n8770 = n8759 ^ n8705 ;
  assign n8775 = n8764 & ~n8770 ;
  assign n8766 = n8750 ^ n8680 ;
  assign n8767 = n8680 ^ n8635 ;
  assign n8768 = ~n8766 & ~n8767 ;
  assign n8773 = n8768 ^ n8760 ;
  assign n8772 = ~n8705 & n8768 ;
  assign n8774 = n8773 ^ n8772 ;
  assign n8776 = n8775 ^ n8774 ;
  assign n8801 = n8800 ^ n8776 ;
  assign n8791 = ~n8635 & n8766 ;
  assign n8756 = n8750 ^ n8705 ;
  assign n8757 = n8756 ^ n8635 ;
  assign n8758 = n8680 & n8757 ;
  assign n8761 = n8760 ^ n8758 ;
  assign n8754 = n8681 & ~n8753 ;
  assign n8752 = n8682 & n8751 ;
  assign n8755 = n8754 ^ n8752 ;
  assign n8762 = n8761 ^ n8755 ;
  assign n8771 = n8770 ^ n8762 ;
  assign n8777 = n8776 ^ n8771 ;
  assign n8778 = n8777 ^ n8774 ;
  assign n8769 = n8768 ^ n8682 ;
  assign n8779 = n8778 ^ n8769 ;
  assign n8780 = n8779 ^ n8751 ;
  assign n8765 = n8751 & n8764 ;
  assign n8781 = n8780 ^ n8765 ;
  assign n8792 = n8791 ^ n8781 ;
  assign n8784 = n8764 ^ n8680 ;
  assign n8785 = ~n8753 & ~n8784 ;
  assign n8790 = n8785 ^ n8762 ;
  assign n8793 = n8792 ^ n8790 ;
  assign n8794 = n8793 ^ n8775 ;
  assign n8795 = n8794 ^ n8774 ;
  assign n8796 = n8795 ^ n8760 ;
  assign n8799 = n8796 ^ n8759 ;
  assign n8802 = n8801 ^ n8799 ;
  assign n8803 = n8802 ^ n8785 ;
  assign n8804 = n8803 ^ n8777 ;
  assign n8805 = n8804 ^ n8800 ;
  assign n8788 = n8781 ^ n8772 ;
  assign n8789 = n8788 ^ n8765 ;
  assign n8797 = n8796 ^ n8789 ;
  assign n8798 = n8797 ^ n8761 ;
  assign n8806 = n8805 ^ n8798 ;
  assign n10812 = ~n8588 & n8806 ;
  assign n10550 = n8765 ^ n8754 ;
  assign n10551 = n10550 ^ n8790 ;
  assign n10552 = n10551 ^ n8772 ;
  assign n10553 = n10552 ^ n10550 ;
  assign n10554 = n10550 ^ n8460 ;
  assign n10555 = n10554 ^ n10550 ;
  assign n10556 = n10553 & ~n10555 ;
  assign n10557 = n10556 ^ n10550 ;
  assign n10558 = n8589 & n10557 ;
  assign n10807 = n10558 ^ n10550 ;
  assign n10574 = n8785 ^ n8774 ;
  assign n10575 = n8774 ^ n8588 ;
  assign n10576 = n10575 ^ n8774 ;
  assign n10577 = n10574 & ~n10576 ;
  assign n10578 = n10577 ^ n8774 ;
  assign n10579 = ~n8460 & n10578 ;
  assign n10808 = n10807 ^ n10579 ;
  assign n10801 = n8778 ^ n8755 ;
  assign n10802 = n8755 ^ n8588 ;
  assign n10803 = n10802 ^ n8755 ;
  assign n10804 = ~n10801 & ~n10803 ;
  assign n10805 = n10804 ^ n8755 ;
  assign n10806 = ~n8460 & n10805 ;
  assign n10809 = n10808 ^ n10806 ;
  assign n8782 = n8460 & ~n8588 ;
  assign n8783 = ~n8781 & n8782 ;
  assign n10810 = n10809 ^ n8783 ;
  assign n10798 = n8794 ^ n8779 ;
  assign n10799 = n10798 ^ n8802 ;
  assign n10800 = n8782 & n10799 ;
  assign n10811 = n10810 ^ n10800 ;
  assign n10813 = n10812 ^ n10811 ;
  assign n8808 = n8782 ^ n8460 ;
  assign n10795 = n8794 ^ n8781 ;
  assign n10796 = n10795 ^ n8777 ;
  assign n10797 = n8808 & ~n10796 ;
  assign n10814 = n10813 ^ n10797 ;
  assign n10816 = n10815 ^ n10814 ;
  assign n10817 = ~n8800 & ~n10816 ;
  assign n10818 = n10817 ^ n7687 ;
  assign n10819 = n10818 ^ x88 ;
  assign n10820 = ~n10794 & n10819 ;
  assign n10883 = n10820 ^ n10819 ;
  assign n10884 = n10883 ^ n10794 ;
  assign n10892 = ~n10852 & n10884 ;
  assign n10821 = n10820 ^ n10794 ;
  assign n10893 = n10892 ^ n10821 ;
  assign n10894 = ~n10872 & ~n10893 ;
  assign n10920 = n10894 ^ n10821 ;
  assign n10873 = n10852 & n10872 ;
  assign n10877 = n10873 ^ n10852 ;
  assign n10878 = n10877 ^ n10872 ;
  assign n10887 = ~n10878 & n10884 ;
  assign n10874 = n10873 ^ n10872 ;
  assign n10875 = ~n10821 & n10874 ;
  assign n10919 = n10887 ^ n10875 ;
  assign n10921 = n10920 ^ n10919 ;
  assign n10885 = n10873 & n10884 ;
  assign n10917 = n10885 ^ n10819 ;
  assign n10918 = n10917 ^ n10893 ;
  assign n10922 = n10921 ^ n10918 ;
  assign n10937 = n10922 ^ n10873 ;
  assign n10927 = n10922 ^ n10887 ;
  assign n10903 = n10892 ^ n10887 ;
  assign n10900 = n10820 & n10873 ;
  assign n10897 = n10820 & n10877 ;
  assign n10886 = n10885 ^ n10875 ;
  assign n10888 = n10887 ^ n10886 ;
  assign n10880 = n10872 ^ n10852 ;
  assign n10881 = ~n10819 & ~n10880 ;
  assign n10882 = n10881 ^ n10821 ;
  assign n10889 = n10888 ^ n10882 ;
  assign n10879 = n10820 & ~n10878 ;
  assign n10890 = n10889 ^ n10879 ;
  assign n10891 = n10890 ^ n10878 ;
  assign n10895 = n10894 ^ n10891 ;
  assign n10898 = n10897 ^ n10895 ;
  assign n10899 = n10898 ^ n10879 ;
  assign n10901 = n10900 ^ n10899 ;
  assign n10896 = n10895 ^ n10820 ;
  assign n10902 = n10901 ^ n10896 ;
  assign n10904 = n10903 ^ n10902 ;
  assign n10876 = n10875 ^ n10874 ;
  assign n10905 = n10904 ^ n10876 ;
  assign n10928 = n10927 ^ n10905 ;
  assign n10926 = n10887 ^ n10879 ;
  assign n10929 = n10928 ^ n10926 ;
  assign n10930 = n10929 ^ n10819 ;
  assign n10931 = n10930 ^ n10882 ;
  assign n10924 = n10872 ^ n10794 ;
  assign n10925 = n10924 ^ n10852 ;
  assign n10932 = n10931 ^ n10925 ;
  assign n10923 = n10922 ^ n10900 ;
  assign n10933 = n10932 ^ n10923 ;
  assign n10934 = n10933 ^ n10885 ;
  assign n10938 = n10937 ^ n10934 ;
  assign n10939 = n10938 ^ n10932 ;
  assign n10940 = n10939 ^ n10921 ;
  assign n10941 = n10940 ^ n10879 ;
  assign n13151 = n10941 ^ n10898 ;
  assign n13162 = n13151 ^ n10922 ;
  assign n13163 = ~n10793 & n13162 ;
  assign n13164 = n13163 ^ n10922 ;
  assign n10972 = n10889 ^ n10887 ;
  assign n10973 = n10972 ^ n10894 ;
  assign n12668 = n10973 ^ n10918 ;
  assign n13148 = n12668 ^ n10928 ;
  assign n13149 = n10793 & n13148 ;
  assign n13150 = n13149 ^ n10928 ;
  assign n13172 = n13164 ^ n13150 ;
  assign n10974 = n10973 ^ n10903 ;
  assign n10975 = n10974 ^ n10905 ;
  assign n9228 = ~n8850 & n9227 ;
  assign n9214 = n9209 ^ n9143 ;
  assign n9215 = n9143 ^ n8850 ;
  assign n9216 = n9215 ^ n9143 ;
  assign n9217 = ~n9214 & n9216 ;
  assign n9218 = n9217 ^ n9143 ;
  assign n9219 = ~n9014 & ~n9218 ;
  assign n9186 = ~n9135 & ~n9185 ;
  assign n9191 = ~n9186 & ~n9190 ;
  assign n9181 = n9153 & ~n9180 ;
  assign n9167 = n9164 ^ n9148 ;
  assign n9171 = n9170 ^ n9167 ;
  assign n9172 = n9171 ^ n9164 ;
  assign n9173 = n9164 ^ n9014 ;
  assign n9174 = n9173 ^ n9164 ;
  assign n9175 = n9172 & n9174 ;
  assign n9176 = n9175 ^ n9164 ;
  assign n9177 = n8850 & n9176 ;
  assign n9159 = n9158 ^ n9131 ;
  assign n9160 = n9157 & n9159 ;
  assign n9161 = n9160 ^ n9131 ;
  assign n9162 = ~n9015 & n9161 ;
  assign n9165 = n9164 ^ n9162 ;
  assign n9178 = n9177 ^ n9165 ;
  assign n9182 = n9181 ^ n9178 ;
  assign n9154 = n9153 ^ n9135 ;
  assign n9155 = n9152 & n9154 ;
  assign n9183 = n9182 ^ n9155 ;
  assign n9150 = n9149 ^ n9142 ;
  assign n9151 = n9150 ^ n9140 ;
  assign n9184 = n9183 ^ n9151 ;
  assign n9192 = n9191 ^ n9184 ;
  assign n9220 = n9219 ^ n9192 ;
  assign n9221 = n9220 ^ n9213 ;
  assign n9201 = n9188 ^ n9164 ;
  assign n9206 = n9201 & n9205 ;
  assign n9207 = n9206 ^ n9188 ;
  assign n9208 = n9015 & n9207 ;
  assign n9222 = n9221 ^ n9208 ;
  assign n9223 = n9222 ^ n7084 ;
  assign n9193 = n9192 ^ n9183 ;
  assign n9194 = n9193 ^ n9141 ;
  assign n9195 = n9194 ^ n9193 ;
  assign n9196 = n9193 ^ n8850 ;
  assign n9197 = n9196 ^ n9193 ;
  assign n9198 = n9195 & ~n9197 ;
  assign n9199 = n9198 ^ n9193 ;
  assign n9200 = ~n9015 & n9199 ;
  assign n9224 = n9223 ^ n9200 ;
  assign n9229 = n9228 ^ n9224 ;
  assign n10907 = n9229 ^ x82 ;
  assign n10976 = n10907 ^ n10905 ;
  assign n10977 = n10976 ^ n10905 ;
  assign n10978 = ~n10975 & n10977 ;
  assign n10979 = n10978 ^ n10905 ;
  assign n10980 = n10793 & n10979 ;
  assign n13173 = n13172 ^ n10980 ;
  assign n13174 = n13173 ^ n9792 ;
  assign n13165 = n13164 ^ n10901 ;
  assign n13166 = n13165 ^ n10890 ;
  assign n13167 = n13166 ^ n10933 ;
  assign n13168 = n13167 ^ n13164 ;
  assign n13169 = n10793 & n13168 ;
  assign n13170 = n13169 ^ n13165 ;
  assign n13171 = ~n10907 & ~n13170 ;
  assign n13175 = n13174 ^ n13171 ;
  assign n10948 = n10907 ^ n10793 ;
  assign n13160 = n10903 ^ n10885 ;
  assign n13161 = n10948 & n13160 ;
  assign n13176 = n13175 ^ n13161 ;
  assign n10966 = n10902 ^ n10889 ;
  assign n13153 = n13150 ^ n10966 ;
  assign n13152 = n13151 ^ n13150 ;
  assign n13154 = n13153 ^ n13152 ;
  assign n13157 = n10793 & n13154 ;
  assign n13158 = n13157 ^ n13153 ;
  assign n13159 = n10907 & n13158 ;
  assign n13177 = n13176 ^ n13159 ;
  assign n13178 = n13177 ^ x125 ;
  assign n13179 = n13147 & ~n13178 ;
  assign n13180 = n13179 ^ n13178 ;
  assign n13181 = n13180 ^ n13147 ;
  assign n10267 = n10266 ^ n9832 ;
  assign n10268 = n9832 ^ n9728 ;
  assign n10269 = n10268 ^ n9832 ;
  assign n10270 = ~n10267 & ~n10269 ;
  assign n10271 = n10270 ^ n9832 ;
  assign n10272 = ~n9727 & ~n10271 ;
  assign n11093 = ~n9729 & n9842 ;
  assign n9834 = n9727 & n9728 ;
  assign n11089 = n9830 ^ n9812 ;
  assign n11090 = n11089 ^ n9840 ;
  assign n11091 = n9834 & n11090 ;
  assign n11082 = n9805 ^ n9795 ;
  assign n11083 = n11082 ^ n9844 ;
  assign n11084 = ~n9727 & n11083 ;
  assign n11081 = n11080 ^ n9807 ;
  assign n11085 = n11084 ^ n11081 ;
  assign n11092 = n11091 ^ n11085 ;
  assign n11094 = n11093 ^ n11092 ;
  assign n11086 = n11085 ^ n9841 ;
  assign n10263 = n9727 & n9841 ;
  assign n11087 = n11086 ^ n10263 ;
  assign n11088 = n9728 & ~n11087 ;
  assign n11095 = n11094 ^ n11088 ;
  assign n11076 = n9832 ^ n9829 ;
  assign n11077 = n9860 & ~n11076 ;
  assign n11078 = n11077 ^ n9829 ;
  assign n11079 = n9729 & n11078 ;
  assign n11096 = n11095 ^ n11079 ;
  assign n11069 = n9815 ^ n9728 ;
  assign n11070 = n9812 ^ n9727 ;
  assign n11071 = n9812 ^ n9728 ;
  assign n11072 = n11071 ^ n9812 ;
  assign n11073 = n11070 & n11072 ;
  assign n11074 = n11073 ^ n9812 ;
  assign n11075 = ~n11069 & ~n11074 ;
  assign n11097 = n11096 ^ n11075 ;
  assign n11098 = ~n10272 & n11097 ;
  assign n11099 = n11098 ^ n7848 ;
  assign n11100 = n11099 ^ x106 ;
  assign n10515 = n8416 ^ n8360 ;
  assign n10497 = n8390 ^ n8357 ;
  assign n10498 = n10497 ^ n7975 ;
  assign n10499 = n10498 ^ n8410 ;
  assign n10500 = n10499 ^ n7659 ;
  assign n10494 = n8391 ^ n8375 ;
  assign n10495 = n10494 ^ n8372 ;
  assign n10484 = n8370 ^ n8366 ;
  assign n10485 = n10484 ^ n8359 ;
  assign n10486 = n8358 ^ n8343 ;
  assign n10487 = n10486 ^ n8376 ;
  assign n10488 = n8376 ^ n8359 ;
  assign n10489 = n10488 ^ n8376 ;
  assign n10490 = ~n10487 & ~n10489 ;
  assign n10491 = n10490 ^ n8376 ;
  assign n10492 = n10485 & n10491 ;
  assign n10493 = n10492 ^ n10484 ;
  assign n10496 = n10495 ^ n10493 ;
  assign n10501 = n10500 ^ n10496 ;
  assign n10502 = n10501 ^ n10493 ;
  assign n10503 = ~n8215 & ~n10502 ;
  assign n10504 = n10503 ^ n10496 ;
  assign n10516 = n10515 ^ n10504 ;
  assign n10517 = n10516 ^ n7475 ;
  assign n10506 = n8380 ^ n8377 ;
  assign n10507 = n10506 ^ n8372 ;
  assign n10512 = ~n8215 & ~n10507 ;
  assign n10505 = n10504 ^ n10493 ;
  assign n10513 = n10512 ^ n10505 ;
  assign n10514 = ~n8343 & n10513 ;
  assign n10518 = n10517 ^ n10514 ;
  assign n11101 = n10518 ^ x99 ;
  assign n11102 = ~n11100 & ~n11101 ;
  assign n11180 = n11102 ^ n11101 ;
  assign n11213 = n11180 ^ n11100 ;
  assign n11214 = n11213 ^ n11101 ;
  assign n11021 = n9130 ^ n9127 ;
  assign n11022 = n11021 ^ n9139 ;
  assign n11023 = n9014 & ~n11022 ;
  assign n11024 = n11023 ^ n9148 ;
  assign n11025 = ~n9015 & n11024 ;
  assign n11005 = n9141 ^ n9123 ;
  assign n11006 = n11005 ^ n9169 ;
  assign n10993 = n9153 ^ n9143 ;
  assign n10994 = ~n9186 & ~n10993 ;
  assign n10992 = n9179 ^ n9139 ;
  assign n10995 = n10994 ^ n10992 ;
  assign n10996 = n9135 ^ n9130 ;
  assign n10997 = n10996 ^ n9186 ;
  assign n10998 = n10997 ^ n10996 ;
  assign n10999 = n10996 ^ n9139 ;
  assign n11000 = n10999 ^ n10996 ;
  assign n11001 = n10998 & n11000 ;
  assign n11002 = n11001 ^ n10996 ;
  assign n11003 = n10995 & ~n11002 ;
  assign n10990 = n9208 ^ n9179 ;
  assign n10991 = n10990 ^ n9162 ;
  assign n11004 = n11003 ^ n10991 ;
  assign n11007 = n11006 ^ n11004 ;
  assign n11018 = n11007 ^ n9219 ;
  assign n11008 = n11007 ^ n9201 ;
  assign n11009 = n11008 ^ n11004 ;
  assign n11010 = n11009 ^ n9150 ;
  assign n11011 = n11010 ^ n9201 ;
  assign n11012 = n11011 ^ n11009 ;
  assign n11013 = n11009 ^ n9014 ;
  assign n11014 = n11013 ^ n11009 ;
  assign n11015 = n11012 & n11014 ;
  assign n11016 = n11015 ^ n11009 ;
  assign n11017 = ~n9015 & n11016 ;
  assign n11019 = n11018 ^ n11017 ;
  assign n10989 = n9158 & n9179 ;
  assign n11020 = n11019 ^ n10989 ;
  assign n11026 = n11025 ^ n11020 ;
  assign n11027 = ~n10659 & ~n11026 ;
  assign n11028 = n11027 ^ n8928 ;
  assign n11029 = n11028 ^ x123 ;
  assign n10198 = n10197 ^ n10153 ;
  assign n10199 = n10167 & ~n10198 ;
  assign n10200 = n10199 ^ n10166 ;
  assign n11031 = ~n10200 & ~n10440 ;
  assign n10236 = n10192 ^ n10179 ;
  assign n10237 = n10179 ^ n10077 ;
  assign n10238 = n10237 ^ n10179 ;
  assign n10239 = n10236 & n10238 ;
  assign n10240 = n10239 ^ n10179 ;
  assign n10241 = n10078 & n10240 ;
  assign n11039 = n10188 ^ n10162 ;
  assign n11040 = n10080 & n11039 ;
  assign n11041 = n10830 ^ n10190 ;
  assign n11042 = n10178 ^ n10159 ;
  assign n11043 = n11042 ^ n10198 ;
  assign n11044 = n10080 & ~n11043 ;
  assign n11045 = n11044 ^ n10167 ;
  assign n11046 = ~n11041 & n11045 ;
  assign n11047 = ~n11040 & ~n11046 ;
  assign n11032 = n10469 ^ n10191 ;
  assign n11033 = n11032 ^ n10175 ;
  assign n11034 = n10175 ^ n10078 ;
  assign n11035 = n11034 ^ n10175 ;
  assign n11036 = n11033 & ~n11035 ;
  assign n11037 = n11036 ^ n10175 ;
  assign n11038 = ~n10202 & n11037 ;
  assign n11048 = n11047 ^ n11038 ;
  assign n11051 = ~n10078 & n10183 ;
  assign n11052 = n11051 ^ n10186 ;
  assign n11053 = n10202 & n11052 ;
  assign n11054 = n11053 ^ n10186 ;
  assign n11055 = n11048 & n11054 ;
  assign n11056 = n11055 ^ n11048 ;
  assign n11057 = ~n10241 & n11056 ;
  assign n11058 = n11031 & n11057 ;
  assign n11059 = n11058 ^ n7724 ;
  assign n11060 = n11059 ^ x73 ;
  assign n10601 = n10004 ^ n9922 ;
  assign n10615 = ~n10004 & n10614 ;
  assign n10616 = n10615 ^ n10610 ;
  assign n10617 = n10616 ^ n10606 ;
  assign n10618 = n10617 ^ n9922 ;
  assign n10619 = n10618 ^ n10617 ;
  assign n10625 = n10624 ^ n10616 ;
  assign n10626 = n10625 ^ n10617 ;
  assign n10627 = n10619 & ~n10626 ;
  assign n10628 = n10627 ^ n10617 ;
  assign n10629 = n10601 & ~n10628 ;
  assign n10630 = n10629 ^ n10616 ;
  assign n10631 = ~n10600 & ~n10630 ;
  assign n10632 = n10631 ^ n7397 ;
  assign n10988 = n10632 ^ x104 ;
  assign n11062 = n11060 ^ n10988 ;
  assign n11061 = n10988 & n11060 ;
  assign n11063 = n11062 ^ n11061 ;
  assign n11064 = n11029 & ~n11063 ;
  assign n11065 = n11064 ^ n11029 ;
  assign n11030 = n10988 & n11029 ;
  assign n11066 = n11065 ^ n11030 ;
  assign n11125 = n9440 & n9497 ;
  assign n11120 = n9454 ^ n9434 ;
  assign n11121 = n11120 ^ n9454 ;
  assign n11122 = n9473 & ~n10740 ;
  assign n11123 = ~n11121 & n11122 ;
  assign n11124 = n11123 ^ n11120 ;
  assign n11126 = n11125 ^ n11124 ;
  assign n11141 = n11140 ^ n11126 ;
  assign n9500 = n9474 ^ n9436 ;
  assign n9501 = n9436 ^ n9303 ;
  assign n9502 = n9501 ^ n9436 ;
  assign n9503 = ~n9500 & n9502 ;
  assign n9504 = n9503 ^ n9436 ;
  assign n9505 = n9304 & n9504 ;
  assign n11142 = n11141 ^ n9505 ;
  assign n11143 = n11142 ^ n10768 ;
  assign n11127 = n11126 ^ n9465 ;
  assign n11128 = n11127 ^ n9484 ;
  assign n11129 = n11128 ^ n11126 ;
  assign n11130 = n11126 ^ n9303 ;
  assign n11131 = n11130 ^ n11126 ;
  assign n11132 = n11129 & ~n11131 ;
  assign n11133 = n11132 ^ n11126 ;
  assign n11134 = n9270 & n11133 ;
  assign n11144 = n11143 ^ n11134 ;
  assign n11111 = n10742 ^ n9460 ;
  assign n9477 = n9476 ^ n9474 ;
  assign n11113 = n11112 ^ n9477 ;
  assign n11114 = n11113 ^ n10740 ;
  assign n11115 = n10740 ^ n9460 ;
  assign n11116 = n11115 ^ n10740 ;
  assign n11117 = ~n11114 & ~n11116 ;
  assign n11118 = n11117 ^ n10740 ;
  assign n11119 = n11111 & ~n11118 ;
  assign n11145 = n11144 ^ n11119 ;
  assign n11110 = n9475 & ~n10740 ;
  assign n11146 = n11145 ^ n11110 ;
  assign n11104 = n9486 ^ n9447 ;
  assign n11105 = n9486 ^ n9270 ;
  assign n11106 = n11105 ^ n9486 ;
  assign n11107 = n11104 & n11106 ;
  assign n11108 = n11107 ^ n9486 ;
  assign n11109 = n9304 & n11108 ;
  assign n11147 = n11146 ^ n11109 ;
  assign n11148 = ~n10744 & n11147 ;
  assign n11149 = n11148 ^ n8889 ;
  assign n11150 = n11149 ^ x113 ;
  assign n11170 = n11066 & n11150 ;
  assign n11155 = ~n11029 & n11150 ;
  assign n11156 = ~n11063 & n11155 ;
  assign n11151 = ~n11060 & ~n11150 ;
  assign n11152 = n10988 & n11151 ;
  assign n11153 = n11152 ^ n11151 ;
  assign n11154 = n11153 ^ n11063 ;
  assign n11157 = n11156 ^ n11154 ;
  assign n11171 = n11170 ^ n11157 ;
  assign n11168 = n11030 & n11151 ;
  assign n11165 = ~n11029 & n11061 ;
  assign n11166 = n11165 ^ n11061 ;
  assign n11167 = n11166 ^ n11030 ;
  assign n11169 = n11168 ^ n11167 ;
  assign n11172 = n11171 ^ n11169 ;
  assign n11164 = n11155 ^ n11150 ;
  assign n11173 = n11172 ^ n11164 ;
  assign n11187 = n11173 ^ n11166 ;
  assign n12738 = n11187 ^ n11168 ;
  assign n13215 = ~n11214 & ~n12738 ;
  assign n11188 = n11061 & n11155 ;
  assign n11204 = n11188 ^ n11165 ;
  assign n11189 = n11188 ^ n11168 ;
  assign n11190 = n11189 ^ n11187 ;
  assign n11191 = n11190 ^ n11169 ;
  assign n13207 = n11204 ^ n11191 ;
  assign n11067 = n11063 ^ n10988 ;
  assign n11068 = n11067 ^ n11066 ;
  assign n11159 = n11068 & ~n11150 ;
  assign n11199 = n11159 ^ n11068 ;
  assign n11200 = n11199 ^ n11156 ;
  assign n11181 = n11170 ^ n11066 ;
  assign n12463 = n11200 ^ n11181 ;
  assign n12743 = n12463 ^ n11157 ;
  assign n13208 = n13207 ^ n12743 ;
  assign n13209 = n11100 & n13208 ;
  assign n11198 = n11188 ^ n11155 ;
  assign n11201 = n11200 ^ n11198 ;
  assign n13205 = n12743 ^ n11201 ;
  assign n11158 = n11157 ^ n11064 ;
  assign n11163 = n11158 ^ n11153 ;
  assign n13194 = n11171 ^ n11163 ;
  assign n13195 = n13194 ^ n11181 ;
  assign n13192 = n11170 ^ n11158 ;
  assign n11185 = n11168 ^ n11152 ;
  assign n12433 = n11185 ^ n11159 ;
  assign n13193 = n13192 ^ n12433 ;
  assign n13196 = n13195 ^ n13193 ;
  assign n13197 = ~n11100 & ~n13196 ;
  assign n13198 = n13197 ^ n13195 ;
  assign n13206 = n13205 ^ n13198 ;
  assign n13210 = n13209 ^ n13206 ;
  assign n13211 = n11101 & ~n13210 ;
  assign n13203 = n11100 & n11204 ;
  assign n13182 = n11185 ^ n11173 ;
  assign n13199 = n13198 ^ n13182 ;
  assign n11162 = n11101 ^ n11100 ;
  assign n11228 = n11172 ^ n11171 ;
  assign n11229 = n11228 ^ n11171 ;
  assign n11230 = n11171 ^ n11100 ;
  assign n11231 = n11230 ^ n11171 ;
  assign n11232 = ~n11229 & ~n11231 ;
  assign n11233 = n11232 ^ n11171 ;
  assign n11234 = ~n11162 & ~n11233 ;
  assign n13200 = n13199 ^ n11234 ;
  assign n13201 = n13200 ^ n9758 ;
  assign n13202 = n13201 ^ n11201 ;
  assign n13204 = n13203 ^ n13202 ;
  assign n13212 = n13211 ^ n13204 ;
  assign n13190 = n11159 ^ n11156 ;
  assign n13191 = ~n11213 & n13190 ;
  assign n13213 = n13212 ^ n13191 ;
  assign n13183 = n13182 ^ n11189 ;
  assign n13184 = n13183 ^ n13182 ;
  assign n13185 = n13182 ^ n11101 ;
  assign n13186 = n13185 ^ n13182 ;
  assign n13187 = n13184 & ~n13186 ;
  assign n13188 = n13187 ^ n13182 ;
  assign n13189 = ~n11162 & ~n13188 ;
  assign n13214 = n13213 ^ n13189 ;
  assign n13216 = n13215 ^ n13214 ;
  assign n13217 = n13216 ^ x76 ;
  assign n10026 = n10022 ^ n10004 ;
  assign n10027 = n10026 ^ n10025 ;
  assign n10028 = n10027 ^ n10003 ;
  assign n10029 = n10028 ^ n6440 ;
  assign n11664 = n10029 ^ x69 ;
  assign n11688 = n8374 ^ n8364 ;
  assign n11689 = n11688 ^ n8376 ;
  assign n11690 = n11689 ^ n8397 ;
  assign n11691 = ~n8215 & n11690 ;
  assign n11692 = n11691 ^ n11688 ;
  assign n11678 = n8394 ^ n8364 ;
  assign n11679 = n8364 ^ n8215 ;
  assign n11680 = n11679 ^ n8364 ;
  assign n11681 = n11678 & n11680 ;
  assign n11682 = n11681 ^ n8364 ;
  assign n11683 = ~n8344 & n11682 ;
  assign n11701 = n11692 ^ n11683 ;
  assign n11702 = n11701 ^ n8416 ;
  assign n11703 = n11702 ^ n8068 ;
  assign n11694 = n8380 & ~n10486 ;
  assign n11695 = n8359 ^ n7977 ;
  assign n11696 = n11695 ^ n8371 ;
  assign n11697 = ~n11694 & n11696 ;
  assign n11693 = n11692 ^ n8366 ;
  assign n11698 = n11697 ^ n11693 ;
  assign n11685 = n8357 ^ n8352 ;
  assign n11686 = n11685 ^ n8397 ;
  assign n11687 = n8343 & ~n11686 ;
  assign n11699 = n11698 ^ n11687 ;
  assign n11700 = n8344 & n11699 ;
  assign n11704 = n11703 ^ n11700 ;
  assign n11684 = n8358 & ~n10497 ;
  assign n11705 = n11704 ^ n11684 ;
  assign n11671 = n8354 ^ n7977 ;
  assign n11670 = n8409 ^ n7977 ;
  assign n11672 = n11671 ^ n11670 ;
  assign n11673 = n11671 ^ n8215 ;
  assign n11674 = n11673 ^ n11671 ;
  assign n11675 = ~n11672 & ~n11674 ;
  assign n11676 = n11675 ^ n11671 ;
  assign n11677 = ~n8343 & n11676 ;
  assign n11709 = n11705 ^ n11677 ;
  assign n11710 = n11709 ^ x125 ;
  assign n11718 = ~n8588 & n8797 ;
  assign n11719 = n11718 ^ n8796 ;
  assign n10563 = n8785 & n10558 ;
  assign n10564 = n10563 ^ n8460 ;
  assign n10565 = ~n8806 & ~n10564 ;
  assign n10566 = n10565 ^ n8460 ;
  assign n11728 = n11719 ^ n10566 ;
  assign n10545 = n8776 ^ n8588 ;
  assign n10546 = n10545 ^ n8776 ;
  assign n10547 = n8801 & ~n10546 ;
  assign n10548 = n10547 ^ n8776 ;
  assign n10549 = n8460 & n10548 ;
  assign n11729 = n11728 ^ n10549 ;
  assign n10521 = n8765 & n8782 ;
  assign n10522 = n10521 ^ n8783 ;
  assign n11730 = n11729 ^ n10522 ;
  assign n11731 = n11730 ^ n10806 ;
  assign n11732 = n11731 ^ n8040 ;
  assign n10531 = n8791 ^ n8750 ;
  assign n10532 = n8756 ^ n8680 ;
  assign n10533 = n10532 ^ n8635 ;
  assign n10534 = n10531 & n10533 ;
  assign n11720 = n11719 ^ n10534 ;
  assign n8786 = n8785 ^ n8754 ;
  assign n11721 = n11720 ^ n8786 ;
  assign n11722 = n11721 ^ n11719 ;
  assign n11725 = n8588 & n11722 ;
  assign n11726 = n11725 ^ n11719 ;
  assign n11727 = n8460 & ~n11726 ;
  assign n11733 = n11732 ^ n11727 ;
  assign n11711 = n8793 ^ n8460 ;
  assign n11712 = n11711 ^ n8793 ;
  assign n11713 = n8793 ^ n8758 ;
  assign n11714 = n11713 ^ n8793 ;
  assign n11715 = n11712 & n11714 ;
  assign n11716 = n11715 ^ n8793 ;
  assign n11717 = ~n8588 & ~n11716 ;
  assign n11734 = n11733 ^ n11717 ;
  assign n11735 = n11734 ^ x110 ;
  assign n11736 = ~n11710 & ~n11735 ;
  assign n11742 = n11736 ^ n11710 ;
  assign n11666 = n11263 ^ x108 ;
  assign n9870 = n9834 ^ n9727 ;
  assign n10309 = n9861 & n9870 ;
  assign n10300 = n10299 ^ n9842 ;
  assign n10276 = n9844 ^ n9829 ;
  assign n10277 = n10276 ^ n9828 ;
  assign n10278 = n10277 ^ n9844 ;
  assign n10279 = ~n9728 & n10278 ;
  assign n10280 = n10279 ^ n10276 ;
  assign n10282 = n10280 ^ n9814 ;
  assign n10283 = n10282 ^ n9838 ;
  assign n10281 = n10280 ^ n9815 ;
  assign n10284 = n10283 ^ n10281 ;
  assign n10273 = n9815 ^ n9810 ;
  assign n10274 = n10273 ^ n9831 ;
  assign n10275 = ~n9728 & n10274 ;
  assign n10285 = n10284 ^ n10275 ;
  assign n10286 = n10285 ^ n10272 ;
  assign n10301 = n10300 ^ n10286 ;
  assign n10306 = n10301 ^ n5379 ;
  assign n10302 = n10301 ^ n10300 ;
  assign n10303 = n10302 ^ n10272 ;
  assign n10304 = n10303 ^ n10280 ;
  assign n10305 = ~n9729 & n10304 ;
  assign n10307 = n10306 ^ n10305 ;
  assign n10264 = n10263 ^ n9842 ;
  assign n10265 = n9728 & n10264 ;
  assign n10308 = n10307 ^ n10265 ;
  assign n10310 = n10309 ^ n10308 ;
  assign n11667 = n10310 ^ x83 ;
  assign n11668 = n11666 & n11667 ;
  assign n11669 = n11668 ^ n11667 ;
  assign n11750 = n11669 ^ n11666 ;
  assign n11751 = ~n11742 & ~n11750 ;
  assign n11739 = n11668 ^ n11666 ;
  assign n11740 = n11736 & n11739 ;
  assign n12155 = n11751 ^ n11740 ;
  assign n11771 = n11736 & ~n11750 ;
  assign n11737 = n11736 ^ n11735 ;
  assign n11754 = n11668 & ~n11737 ;
  assign n11738 = n11669 & ~n11737 ;
  assign n11768 = n11754 ^ n11738 ;
  assign n11766 = ~n11737 & ~n11750 ;
  assign n11767 = n11766 ^ n11737 ;
  assign n11769 = n11768 ^ n11767 ;
  assign n11772 = n11771 ^ n11769 ;
  assign n11756 = n11668 & n11736 ;
  assign n11743 = n11742 ^ n11735 ;
  assign n11749 = n11739 & ~n11743 ;
  assign n11752 = n11751 ^ n11749 ;
  assign n11757 = n11756 ^ n11752 ;
  assign n11745 = n11668 & ~n11742 ;
  assign n11744 = n11669 & ~n11743 ;
  assign n11746 = n11745 ^ n11744 ;
  assign n11758 = n11757 ^ n11746 ;
  assign n11755 = n11754 ^ n11744 ;
  assign n11759 = n11758 ^ n11755 ;
  assign n11753 = n11752 ^ n11668 ;
  assign n11760 = n11759 ^ n11753 ;
  assign n11764 = n11760 ^ n11744 ;
  assign n11763 = n11749 ^ n11743 ;
  assign n11765 = n11764 ^ n11763 ;
  assign n11773 = n11772 ^ n11765 ;
  assign n11774 = n11773 ^ n11740 ;
  assign n11775 = n11774 ^ n11756 ;
  assign n11776 = n11775 ^ n11736 ;
  assign n11770 = n11769 ^ n11765 ;
  assign n11777 = n11776 ^ n11770 ;
  assign n12156 = n12155 ^ n11777 ;
  assign n11663 = n11320 ^ x86 ;
  assign n12157 = n11777 ^ n11663 ;
  assign n12158 = n12157 ^ n11777 ;
  assign n12159 = n12156 & n12158 ;
  assign n12160 = n12159 ^ n11777 ;
  assign n12161 = n11664 & n12160 ;
  assign n11781 = n11771 ^ n11749 ;
  assign n11782 = n11781 ^ n11740 ;
  assign n11783 = n11782 ^ n11739 ;
  assign n11784 = n11783 ^ n11772 ;
  assign n11785 = n11784 ^ n11771 ;
  assign n11786 = n11785 ^ n11749 ;
  assign n11778 = n11777 ^ n11764 ;
  assign n11761 = n11760 ^ n11738 ;
  assign n11762 = n11761 ^ n11669 ;
  assign n11779 = n11778 ^ n11762 ;
  assign n11787 = n11786 ^ n11779 ;
  assign n11788 = ~n11663 & ~n11787 ;
  assign n11789 = n11788 ^ n11785 ;
  assign n12162 = n12161 ^ n11789 ;
  assign n11793 = n11663 & ~n11664 ;
  assign n12152 = n11779 & n11793 ;
  assign n12147 = n11754 ^ n11664 ;
  assign n12148 = n12147 ^ n11754 ;
  assign n12149 = n11768 & ~n12148 ;
  assign n12150 = n12149 ^ n11754 ;
  assign n12151 = ~n11663 & n12150 ;
  assign n12153 = n12152 ^ n12151 ;
  assign n11794 = n11793 ^ n11664 ;
  assign n11819 = n11794 ^ n11663 ;
  assign n12142 = n11819 ^ n11664 ;
  assign n12143 = n11761 & n12142 ;
  assign n12140 = n11784 ^ n11765 ;
  assign n12141 = n11819 & n12140 ;
  assign n12144 = n12143 ^ n12141 ;
  assign n12154 = n12153 ^ n12144 ;
  assign n12163 = n12162 ^ n12154 ;
  assign n11795 = n11770 & ~n11794 ;
  assign n12164 = n12163 ^ n11795 ;
  assign n12165 = n12164 ^ n8214 ;
  assign n12133 = n11766 ^ n11745 ;
  assign n12134 = n12133 ^ n11772 ;
  assign n12135 = n11772 ^ n11663 ;
  assign n12136 = n12135 ^ n11772 ;
  assign n12137 = ~n12134 & n12136 ;
  assign n12138 = n12137 ^ n11772 ;
  assign n12139 = n11664 & ~n12138 ;
  assign n12166 = n12165 ^ n12139 ;
  assign n11807 = n11777 ^ n11761 ;
  assign n12131 = n11807 ^ n11770 ;
  assign n12132 = n11793 & n12131 ;
  assign n12167 = n12166 ^ n12132 ;
  assign n11665 = n11664 ^ n11663 ;
  assign n12123 = n11789 ^ n11755 ;
  assign n12126 = n12123 ^ n11759 ;
  assign n12127 = n12126 ^ n12123 ;
  assign n12128 = ~n11663 & n12127 ;
  assign n12129 = n12128 ^ n12123 ;
  assign n12130 = ~n11665 & ~n12129 ;
  assign n12168 = n12167 ^ n12130 ;
  assign n13218 = n12168 ^ x126 ;
  assign n13219 = ~n13217 & n13218 ;
  assign n13220 = n13219 ^ n13218 ;
  assign n13221 = n13181 & n13220 ;
  assign n9723 = ~n9684 & n9701 ;
  assign n9717 = n9673 ^ n9631 ;
  assign n9688 = n9687 ^ n9568 ;
  assign n9653 = n9652 ^ n9626 ;
  assign n9654 = n9653 ^ n9650 ;
  assign n9689 = n9688 ^ n9654 ;
  assign n9668 = n9626 ^ n9590 ;
  assign n9669 = n9668 ^ n9636 ;
  assign n9690 = n9689 ^ n9669 ;
  assign n9718 = n9717 ^ n9690 ;
  assign n9675 = n9674 ^ n9669 ;
  assign n9716 = n9715 ^ n9675 ;
  assign n9719 = n9718 ^ n9716 ;
  assign n9720 = n9719 ^ n9671 ;
  assign n9721 = ~n9538 & ~n9720 ;
  assign n9693 = n9689 ^ n9537 ;
  assign n9694 = n9693 ^ n9689 ;
  assign n9695 = ~n9690 & n9694 ;
  assign n9696 = n9695 ^ n9689 ;
  assign n9697 = n9538 & ~n9696 ;
  assign n9685 = n9673 & ~n9684 ;
  assign n9676 = n9675 ^ n9631 ;
  assign n9677 = n9676 ^ n9675 ;
  assign n9678 = n9675 ^ n9536 ;
  assign n9679 = n9678 ^ n9675 ;
  assign n9680 = n9677 & ~n9679 ;
  assign n9681 = n9680 ^ n9675 ;
  assign n9682 = n9538 & n9681 ;
  assign n9686 = n9685 ^ n9682 ;
  assign n9698 = n9697 ^ n9686 ;
  assign n9712 = n9711 ^ n9698 ;
  assign n9713 = n9712 ^ n6855 ;
  assign n9663 = n9640 ^ n9633 ;
  assign n9664 = n9663 ^ n9647 ;
  assign n9666 = n9665 ^ n9664 ;
  assign n9667 = n9662 & ~n9666 ;
  assign n9714 = n9713 ^ n9667 ;
  assign n9722 = n9721 ^ n9714 ;
  assign n9724 = n9723 ^ n9722 ;
  assign n9657 = n9650 ^ n9536 ;
  assign n9658 = n9657 ^ n9650 ;
  assign n9659 = ~n9654 & n9658 ;
  assign n9660 = n9659 ^ n9650 ;
  assign n9661 = n9538 & ~n9660 ;
  assign n9725 = n9724 ^ n9661 ;
  assign n9726 = n9725 ^ x107 ;
  assign n9230 = n9229 ^ x90 ;
  assign n11590 = n9726 ^ n9230 ;
  assign n9468 = n9467 ^ n9457 ;
  assign n9506 = n9487 ^ n9468 ;
  assign n9507 = n9506 ^ n9505 ;
  assign n9499 = n9498 ^ n7250 ;
  assign n9508 = n9507 ^ n9499 ;
  assign n9488 = n9487 ^ n9440 ;
  assign n9490 = n9489 ^ n9488 ;
  assign n9491 = n9490 ^ n9487 ;
  assign n9492 = n9487 ^ n9303 ;
  assign n9493 = n9492 ^ n9487 ;
  assign n9494 = n9491 & n9493 ;
  assign n9495 = n9494 ^ n9487 ;
  assign n9496 = n9270 & n9495 ;
  assign n9509 = n9508 ^ n9496 ;
  assign n9478 = n9477 ^ n9472 ;
  assign n9479 = n9472 ^ n9270 ;
  assign n9480 = n9479 ^ n9472 ;
  assign n9481 = ~n9478 & ~n9480 ;
  assign n9482 = n9481 ^ n9472 ;
  assign n9483 = ~n9303 & n9482 ;
  assign n9510 = n9509 ^ n9483 ;
  assign n9444 = n9443 ^ n9440 ;
  assign n9448 = n9447 ^ n9444 ;
  assign n9437 = n9436 ^ n9434 ;
  assign n9445 = n9444 ^ n9437 ;
  assign n9446 = n9303 & n9445 ;
  assign n9449 = n9448 ^ n9446 ;
  assign n9451 = n9450 ^ n9449 ;
  assign n9469 = n9468 ^ n9451 ;
  assign n9470 = ~n9304 & n9469 ;
  assign n9511 = n9510 ^ n9470 ;
  assign n9512 = n9511 ^ x89 ;
  assign n9871 = n9816 & n9870 ;
  assign n9846 = n9807 ^ n9805 ;
  assign n9848 = n9847 ^ n9846 ;
  assign n9849 = ~n9728 & n9848 ;
  assign n9866 = n9849 ^ n7290 ;
  assign n9867 = n9866 ^ n9865 ;
  assign n9845 = n9844 ^ n9806 ;
  assign n9850 = n9849 ^ n9845 ;
  assign n9801 = n9800 ^ n9795 ;
  assign n9851 = n9850 ^ n9801 ;
  assign n9852 = n9851 ^ n9806 ;
  assign n9853 = n9852 ^ n9850 ;
  assign n9854 = n9850 ^ n9728 ;
  assign n9855 = n9854 ^ n9850 ;
  assign n9856 = n9853 & n9855 ;
  assign n9857 = n9856 ^ n9850 ;
  assign n9858 = n9729 & n9857 ;
  assign n9868 = n9867 ^ n9858 ;
  assign n9833 = n9832 ^ n9828 ;
  assign n9837 = ~n9833 & n9834 ;
  assign n9869 = n9868 ^ n9837 ;
  assign n9872 = n9871 ^ n9869 ;
  assign n9835 = n9834 ^ n9728 ;
  assign n9836 = ~n9833 & n9835 ;
  assign n9873 = n9872 ^ n9836 ;
  assign n9819 = n9818 ^ n9812 ;
  assign n9808 = n9807 ^ n9801 ;
  assign n9820 = n9819 ^ n9808 ;
  assign n9821 = n9808 ^ n9728 ;
  assign n9822 = n9821 ^ n9808 ;
  assign n9823 = ~n9820 & ~n9822 ;
  assign n9824 = n9823 ^ n9808 ;
  assign n9825 = ~n9729 & n9824 ;
  assign n9874 = n9873 ^ n9825 ;
  assign n9875 = n9874 ^ x80 ;
  assign n9877 = ~n9726 & n9875 ;
  assign n9909 = n9877 ^ n9230 ;
  assign n9891 = n9230 & n9875 ;
  assign n9908 = n9891 ^ n9726 ;
  assign n9910 = n9909 ^ n9908 ;
  assign n9911 = n9512 & n9910 ;
  assign n9912 = n9911 ^ n9908 ;
  assign n11591 = n11590 ^ n9912 ;
  assign n9883 = n9230 & ~n9512 ;
  assign n9884 = n9883 ^ n9230 ;
  assign n9885 = n9884 ^ n9512 ;
  assign n9886 = ~n9877 & ~n9885 ;
  assign n9887 = n9886 ^ n9512 ;
  assign n11592 = n11591 ^ n9887 ;
  assign n9876 = n9875 ^ n9726 ;
  assign n9878 = n9877 ^ n9876 ;
  assign n9890 = n9878 ^ n9230 ;
  assign n9892 = n9891 ^ n9890 ;
  assign n11587 = n9892 ^ n9726 ;
  assign n9902 = n9875 ^ n9512 ;
  assign n9903 = n9512 ^ n9230 ;
  assign n9904 = ~n9875 & ~n9903 ;
  assign n9905 = n9904 ^ n9726 ;
  assign n9906 = n9902 & n9905 ;
  assign n11588 = n11587 ^ n9906 ;
  assign n11584 = n9230 & n9878 ;
  assign n11589 = n11588 ^ n11584 ;
  assign n11593 = n11592 ^ n11589 ;
  assign n11594 = n11593 ^ n9512 ;
  assign n11585 = n11584 ^ n9877 ;
  assign n11586 = n11585 ^ n9885 ;
  assign n11595 = n11594 ^ n11586 ;
  assign n8419 = n8418 ^ x112 ;
  assign n11603 = n11594 ^ n11592 ;
  assign n11604 = ~n8419 & ~n11603 ;
  assign n11605 = n11604 ^ n11592 ;
  assign n9879 = n9878 ^ n9875 ;
  assign n9880 = ~n9512 & n9879 ;
  assign n9881 = n9880 ^ n9875 ;
  assign n9882 = ~n9230 & n9881 ;
  assign n9888 = n9887 ^ n9882 ;
  assign n9889 = n9888 ^ n9885 ;
  assign n11599 = n9908 ^ n9889 ;
  assign n11597 = n11588 ^ n9883 ;
  assign n11596 = n9904 ^ n9880 ;
  assign n11598 = n11597 ^ n11596 ;
  assign n11600 = n11599 ^ n11598 ;
  assign n11601 = n8419 & n11600 ;
  assign n11602 = n11601 ^ n11598 ;
  assign n11606 = n11605 ^ n11602 ;
  assign n8811 = n8806 ^ n8772 ;
  assign n8812 = n8811 ^ n8754 ;
  assign n8809 = n8765 & n8808 ;
  assign n8787 = n8786 ^ n8783 ;
  assign n8807 = n8806 ^ n8787 ;
  assign n8810 = n8809 ^ n8807 ;
  assign n8813 = n8812 ^ n8810 ;
  assign n8814 = n8813 ^ n8775 ;
  assign n8815 = n8814 ^ n8810 ;
  assign n8816 = n8810 ^ n8588 ;
  assign n8817 = n8816 ^ n8810 ;
  assign n8818 = n8815 & ~n8817 ;
  assign n8819 = n8818 ^ n8810 ;
  assign n8820 = ~n8460 & n8819 ;
  assign n8821 = n8820 ^ n8810 ;
  assign n8763 = ~n8589 & n8762 ;
  assign n8822 = n8821 ^ n8763 ;
  assign n8823 = n8774 ^ n8460 ;
  assign n8824 = n8823 ^ n8774 ;
  assign n8825 = n8800 ^ n8777 ;
  assign n8826 = n8825 ^ n8774 ;
  assign n8827 = n8824 & ~n8826 ;
  assign n8828 = n8827 ^ n8774 ;
  assign n8829 = n8588 & n8828 ;
  assign n8830 = n8829 ^ n8774 ;
  assign n8831 = ~n8822 & ~n8830 ;
  assign n8832 = n8589 & n8831 ;
  assign n8833 = n8779 ^ n8775 ;
  assign n8834 = n8833 ^ n8805 ;
  assign n8835 = ~n8460 & n8834 ;
  assign n8836 = n8835 ^ n8793 ;
  assign n8837 = n8832 & ~n8836 ;
  assign n8838 = n8837 ^ n8831 ;
  assign n8839 = n8760 ^ n8460 ;
  assign n8840 = n8839 ^ n8760 ;
  assign n8843 = n8775 & n8840 ;
  assign n8844 = n8843 ^ n8760 ;
  assign n8845 = ~n8588 & n8844 ;
  assign n8846 = n8838 & ~n8845 ;
  assign n8847 = n8846 ^ n6198 ;
  assign n8848 = n8847 ^ x65 ;
  assign n11607 = n11605 ^ n8848 ;
  assign n11608 = n11607 ^ n11605 ;
  assign n11609 = ~n11606 & ~n11608 ;
  assign n11610 = n11609 ^ n11605 ;
  assign n11611 = n11595 & ~n11610 ;
  assign n11612 = n11611 ^ n8704 ;
  assign n13222 = n11612 ^ x108 ;
  assign n11829 = n11059 ^ x122 ;
  assign n11830 = n10818 ^ x66 ;
  assign n11898 = n11829 & ~n11830 ;
  assign n11907 = n11898 ^ n11829 ;
  assign n11839 = ~n8371 & n11694 ;
  assign n11842 = n11839 ^ n8392 ;
  assign n11837 = n8365 ^ n8357 ;
  assign n11838 = n11837 ^ n8409 ;
  assign n11840 = ~n8359 & ~n11839 ;
  assign n11841 = ~n11838 & n11840 ;
  assign n11843 = n11842 ^ n11841 ;
  assign n11852 = n11843 ^ n8361 ;
  assign n11846 = n8394 ^ n8375 ;
  assign n11844 = n8368 ^ n8363 ;
  assign n11845 = n8358 & n11844 ;
  assign n11847 = n11846 ^ n11845 ;
  assign n11848 = n11847 ^ n8397 ;
  assign n11849 = n11848 ^ n11843 ;
  assign n11834 = n10484 ^ n8374 ;
  assign n11835 = n11834 ^ n8397 ;
  assign n11836 = ~n8215 & n11835 ;
  assign n11850 = n11849 ^ n11836 ;
  assign n11851 = ~n8344 & ~n11850 ;
  assign n11853 = n11852 ^ n11851 ;
  assign n11854 = ~n11683 & n11853 ;
  assign n11855 = n11854 ^ n7813 ;
  assign n11856 = n11855 ^ x98 ;
  assign n10426 = n9641 & n9662 ;
  assign n10429 = n10428 ^ n10426 ;
  assign n11872 = n9685 ^ n9626 ;
  assign n11865 = n9699 ^ n9637 ;
  assign n11866 = n9537 & n11865 ;
  assign n11867 = n11866 ^ n9647 ;
  assign n11873 = n11872 ^ n11867 ;
  assign n11868 = n11867 ^ n9626 ;
  assign n10433 = n9648 ^ n9626 ;
  assign n11860 = n10433 ^ n9688 ;
  assign n10395 = n9718 ^ n9643 ;
  assign n10394 = n9699 ^ n9641 ;
  assign n10396 = n10395 ^ n10394 ;
  assign n11861 = n11860 ^ n10396 ;
  assign n11859 = n9587 ^ n9568 ;
  assign n11862 = n11861 ^ n11859 ;
  assign n11869 = n11868 ^ n11862 ;
  assign n11857 = n9700 ^ n9643 ;
  assign n11858 = n11857 ^ n9669 ;
  assign n11863 = n11862 ^ n11858 ;
  assign n11864 = ~n9537 & ~n11863 ;
  assign n11870 = n11869 ^ n11864 ;
  assign n11871 = n9536 & n11870 ;
  assign n11874 = n11873 ^ n11871 ;
  assign n11875 = ~n10429 & n11874 ;
  assign n11876 = ~n9697 & n11875 ;
  assign n11878 = n9538 & ~n9719 ;
  assign n11879 = n11876 & n11878 ;
  assign n11877 = n11876 ^ n7874 ;
  assign n11880 = n11879 ^ n11877 ;
  assign n11881 = n11880 ^ x120 ;
  assign n11882 = n11856 & n11881 ;
  assign n11890 = n11882 ^ n11881 ;
  assign n11831 = n11099 ^ x81 ;
  assign n11832 = n10792 ^ x72 ;
  assign n11833 = n11831 & n11832 ;
  assign n11886 = n11833 ^ n11831 ;
  assign n11918 = n11886 ^ n11832 ;
  assign n11935 = n11890 & ~n11918 ;
  assign n12213 = n11907 & n11935 ;
  assign n11887 = n11882 ^ n11856 ;
  assign n11888 = n11887 ^ n11881 ;
  assign n11930 = ~n11888 & ~n11918 ;
  assign n11919 = n11918 ^ n11831 ;
  assign n11920 = n11887 & n11919 ;
  assign n11899 = n11832 ^ n11831 ;
  assign n11900 = n11887 ^ n11832 ;
  assign n11901 = n11899 & ~n11900 ;
  assign n11902 = n11901 ^ n11886 ;
  assign n11921 = n11920 ^ n11902 ;
  assign n11917 = n11882 & n11886 ;
  assign n11922 = n11921 ^ n11917 ;
  assign n11891 = n11833 & n11890 ;
  assign n11926 = n11922 ^ n11891 ;
  assign n11883 = n11833 & n11882 ;
  assign n11927 = n11926 ^ n11883 ;
  assign n11889 = n11886 & ~n11888 ;
  assign n11923 = n11889 ^ n11886 ;
  assign n11924 = n11923 ^ n11922 ;
  assign n11903 = n11833 & n11887 ;
  assign n11925 = n11924 ^ n11903 ;
  assign n11928 = n11927 ^ n11925 ;
  assign n11916 = n11889 ^ n11831 ;
  assign n11929 = n11928 ^ n11916 ;
  assign n11931 = n11930 ^ n11929 ;
  assign n11967 = n11930 ^ n11829 ;
  assign n11968 = n11967 ^ n11930 ;
  assign n11969 = n11931 & ~n11968 ;
  assign n11970 = n11969 ^ n11930 ;
  assign n11971 = ~n11830 & n11970 ;
  assign n12214 = n12213 ^ n11971 ;
  assign n12250 = n11920 ^ n11917 ;
  assign n12251 = n11920 ^ n11830 ;
  assign n12252 = n12251 ^ n11920 ;
  assign n12253 = n12250 & n12252 ;
  assign n12254 = n12253 ^ n11920 ;
  assign n12255 = ~n11829 & n12254 ;
  assign n12256 = n12255 ^ n11925 ;
  assign n11952 = n11830 ^ n11829 ;
  assign n11983 = n11935 ^ n11883 ;
  assign n11984 = n11983 ^ n11929 ;
  assign n12240 = ~n11830 & n11984 ;
  assign n12241 = n12240 ^ n11929 ;
  assign n11990 = n11921 ^ n11883 ;
  assign n11942 = n11890 & n11919 ;
  assign n11943 = n11942 ^ n11921 ;
  assign n11944 = n11943 ^ n11935 ;
  assign n11904 = n11903 ^ n11887 ;
  assign n11905 = n11904 ^ n11902 ;
  assign n11985 = n11944 ^ n11905 ;
  assign n11986 = n11985 ^ n11891 ;
  assign n11932 = n11889 ^ n11888 ;
  assign n11933 = n11932 ^ n11931 ;
  assign n11987 = n11986 ^ n11933 ;
  assign n11988 = n11987 ^ n11900 ;
  assign n11989 = n11988 ^ n11984 ;
  assign n11991 = n11990 ^ n11989 ;
  assign n11982 = n11922 ^ n11882 ;
  assign n11992 = n11991 ^ n11982 ;
  assign n12242 = n12241 ^ n11992 ;
  assign n12243 = n12242 ^ n12241 ;
  assign n12246 = ~n11830 & ~n12243 ;
  assign n12247 = n12246 ^ n12241 ;
  assign n12248 = ~n11952 & n12247 ;
  assign n12249 = n12248 ^ n12241 ;
  assign n12257 = n12256 ^ n12249 ;
  assign n12258 = n12257 ^ n11989 ;
  assign n11934 = n11933 ^ n11905 ;
  assign n12259 = n12258 ^ n11934 ;
  assign n12233 = n11928 ^ n11829 ;
  assign n12234 = n12233 ^ n11928 ;
  assign n12235 = n11943 ^ n11925 ;
  assign n12236 = n12235 ^ n11928 ;
  assign n12237 = ~n12234 & n12236 ;
  assign n12238 = n12237 ^ n11928 ;
  assign n12239 = ~n11952 & n12238 ;
  assign n12260 = n12259 ^ n12239 ;
  assign n12231 = n11930 ^ n11920 ;
  assign n12232 = n11907 & n12231 ;
  assign n12261 = n12260 ^ n12232 ;
  assign n12223 = n11989 ^ n11942 ;
  assign n12224 = n12223 ^ n11992 ;
  assign n12225 = n12224 ^ n11989 ;
  assign n12226 = n11989 ^ n11830 ;
  assign n12227 = n12226 ^ n11989 ;
  assign n12228 = ~n12225 & n12227 ;
  assign n12229 = n12228 ^ n11989 ;
  assign n12230 = ~n11829 & ~n12229 ;
  assign n12262 = n12261 ^ n12230 ;
  assign n12215 = n11934 ^ n11917 ;
  assign n11892 = n11891 ^ n11889 ;
  assign n12216 = n12215 ^ n11892 ;
  assign n12217 = n12216 ^ n11934 ;
  assign n12218 = n11934 ^ n11830 ;
  assign n12219 = n12218 ^ n11934 ;
  assign n12220 = n12217 & ~n12219 ;
  assign n12221 = n12220 ^ n11934 ;
  assign n12222 = ~n11952 & ~n12221 ;
  assign n12263 = n12262 ^ n12222 ;
  assign n12264 = ~n12214 & ~n12263 ;
  assign n12265 = n12264 ^ n7973 ;
  assign n13223 = n12265 ^ x94 ;
  assign n13224 = ~n13222 & n13223 ;
  assign n13225 = n13224 ^ n13223 ;
  assign n13226 = n13225 ^ n13222 ;
  assign n13227 = n13226 ^ n13223 ;
  assign n13228 = n13221 & ~n13227 ;
  assign n13232 = n13181 ^ n13178 ;
  assign n13263 = n13219 & n13232 ;
  assign n13235 = n13219 ^ n13217 ;
  assign n13242 = n13235 ^ n13218 ;
  assign n13246 = n13179 & n13242 ;
  assign n13239 = n13232 & ~n13235 ;
  assign n13240 = n13239 ^ n13235 ;
  assign n13237 = ~n13180 & ~n13235 ;
  assign n13236 = n13179 & ~n13235 ;
  assign n13238 = n13237 ^ n13236 ;
  assign n13241 = n13240 ^ n13238 ;
  assign n13247 = n13246 ^ n13241 ;
  assign n13245 = n13181 & n13242 ;
  assign n13248 = n13247 ^ n13245 ;
  assign n13244 = n13232 & n13242 ;
  assign n13249 = n13248 ^ n13244 ;
  assign n13243 = n13242 ^ n13241 ;
  assign n13250 = n13249 ^ n13243 ;
  assign n13260 = n13250 ^ n13244 ;
  assign n13259 = ~n13180 & n13220 ;
  assign n13261 = n13260 ^ n13259 ;
  assign n13257 = n13244 ^ n13237 ;
  assign n13258 = n13257 ^ n13180 ;
  assign n13262 = n13261 ^ n13258 ;
  assign n13264 = n13263 ^ n13262 ;
  assign n13254 = n13246 ^ n13221 ;
  assign n13255 = n13254 ^ n13181 ;
  assign n13256 = n13255 ^ n13248 ;
  assign n13265 = n13264 ^ n13256 ;
  assign n13251 = n13250 ^ n13246 ;
  assign n13252 = n13251 ^ n13236 ;
  assign n13253 = n13252 ^ n13245 ;
  assign n13266 = n13265 ^ n13253 ;
  assign n13230 = n13218 ^ n13147 ;
  assign n13231 = ~n13217 & ~n13230 ;
  assign n13233 = n13232 ^ n13231 ;
  assign n13234 = n13233 ^ n13220 ;
  assign n13267 = n13266 ^ n13234 ;
  assign n13268 = n13267 ^ n13259 ;
  assign n13229 = n13221 ^ n13220 ;
  assign n13269 = n13268 ^ n13229 ;
  assign n13270 = n13269 ^ n13264 ;
  assign n13271 = n13270 ^ n13248 ;
  assign n13272 = n13222 & ~n13271 ;
  assign n13273 = n13272 ^ n13248 ;
  assign n13274 = n13223 & ~n13273 ;
  assign n13275 = n13226 & n13260 ;
  assign n13304 = n13224 & ~n13268 ;
  assign n13276 = n13265 ^ n13219 ;
  assign n13277 = n13276 ^ n13256 ;
  assign n13300 = n13277 ^ n13239 ;
  assign n13301 = ~n13222 & ~n13300 ;
  assign n13284 = n13267 ^ n13264 ;
  assign n13296 = ~n13227 & n13284 ;
  assign n13290 = n13259 ^ n13239 ;
  assign n13291 = n13239 ^ n13223 ;
  assign n13292 = n13291 ^ n13239 ;
  assign n13293 = n13290 & n13292 ;
  assign n13294 = n13293 ^ n13239 ;
  assign n13295 = n13222 & n13294 ;
  assign n13297 = n13296 ^ n13295 ;
  assign n13281 = n13223 ^ n13222 ;
  assign n13285 = n13284 ^ n13247 ;
  assign n13282 = n13250 ^ n13236 ;
  assign n13286 = n13285 ^ n13282 ;
  assign n13287 = n13223 & ~n13286 ;
  assign n13283 = n13282 ^ n13237 ;
  assign n13288 = n13287 ^ n13283 ;
  assign n13289 = ~n13281 & n13288 ;
  assign n13298 = n13297 ^ n13289 ;
  assign n13279 = n13254 ^ n13236 ;
  assign n13280 = n13226 & n13279 ;
  assign n13299 = n13298 ^ n13280 ;
  assign n13302 = n13301 ^ n13299 ;
  assign n13278 = ~n13223 & ~n13277 ;
  assign n13303 = n13302 ^ n13278 ;
  assign n13305 = n13304 ^ n13303 ;
  assign n13306 = ~n13275 & ~n13305 ;
  assign n13307 = ~n13274 & n13306 ;
  assign n13308 = ~n13228 & n13307 ;
  assign n13309 = n13308 ^ n10310 ;
  assign n13310 = n13309 ^ x69 ;
  assign n10633 = n10632 ^ x116 ;
  assign n10669 = n10668 ^ x102 ;
  assign n10437 = n9662 & n9699 ;
  assign n10434 = n10433 ^ n9673 ;
  assign n10435 = n9683 & ~n10434 ;
  assign n10407 = n9652 ^ n9641 ;
  assign n10408 = n10407 ^ n9702 ;
  assign n10409 = n10408 ^ n9537 ;
  assign n10399 = n10395 ^ n9536 ;
  assign n10400 = n10399 ^ n10395 ;
  assign n10401 = ~n10396 & n10400 ;
  assign n10402 = n10401 ^ n10395 ;
  assign n10403 = ~n9537 & ~n10402 ;
  assign n10410 = n10409 ^ n10403 ;
  assign n10404 = n9651 ^ n9629 ;
  assign n10405 = n10404 ^ n9700 ;
  assign n10406 = n9684 & ~n10405 ;
  assign n10411 = n10410 ^ n10406 ;
  assign n10412 = n10411 ^ n10403 ;
  assign n10413 = n10412 ^ n9537 ;
  assign n10414 = n10413 ^ n10412 ;
  assign n10415 = n10412 ^ n9715 ;
  assign n10416 = n10415 ^ n10412 ;
  assign n10417 = n10414 & n10416 ;
  assign n10418 = n10417 ^ n10412 ;
  assign n10419 = n9536 & n10418 ;
  assign n10420 = n10419 ^ n10411 ;
  assign n10421 = n10420 ^ n10403 ;
  assign n10422 = n9689 ^ n9674 ;
  assign n10423 = n9704 & ~n10422 ;
  assign n10424 = ~n10421 & n10423 ;
  assign n10425 = n10424 ^ n10420 ;
  assign n10430 = n10429 ^ n10425 ;
  assign n10431 = n10430 ^ n9697 ;
  assign n10432 = n10431 ^ n7449 ;
  assign n10436 = n10435 ^ n10432 ;
  assign n10438 = n10437 ^ n10436 ;
  assign n10439 = n10438 ^ x70 ;
  assign n10479 = n10478 ^ x67 ;
  assign n10480 = ~n10439 & n10479 ;
  assign n10481 = n10480 ^ n10479 ;
  assign n10570 = n8808 & n8812 ;
  assign n10530 = n8793 ^ n8777 ;
  assign n10567 = n10566 ^ n10530 ;
  assign n10568 = n10567 ^ n10549 ;
  assign n10535 = n10534 ^ n10530 ;
  assign n10536 = n10535 ^ n8775 ;
  assign n10537 = n10536 ^ n10530 ;
  assign n10538 = n10530 ^ n8460 ;
  assign n10539 = n10538 ^ n10530 ;
  assign n10540 = n10537 & ~n10539 ;
  assign n10541 = n10540 ^ n10530 ;
  assign n10542 = n8589 & n10541 ;
  assign n10569 = n10568 ^ n10542 ;
  assign n10571 = n10570 ^ n10569 ;
  assign n10523 = n8779 ^ n8762 ;
  assign n10524 = n10523 ^ n8804 ;
  assign n10525 = n8804 ^ n8460 ;
  assign n10526 = n10525 ^ n8804 ;
  assign n10527 = n10524 & ~n10526 ;
  assign n10528 = n10527 ^ n8804 ;
  assign n10529 = ~n8588 & ~n10528 ;
  assign n10572 = n10571 ^ n10529 ;
  assign n10573 = ~n10522 & n10572 ;
  assign n10580 = ~n8845 & ~n10579 ;
  assign n10581 = n10573 & n10580 ;
  assign n10582 = n10581 ^ n7518 ;
  assign n10583 = n10582 ^ x84 ;
  assign n10696 = n10481 & n10583 ;
  assign n10519 = n10518 ^ x77 ;
  assign n10584 = ~n10519 & ~n10583 ;
  assign n10585 = n10584 ^ n10583 ;
  assign n10674 = n10481 & ~n10585 ;
  assign n10675 = n10674 ^ n10481 ;
  assign n10697 = n10696 ^ n10675 ;
  assign n10698 = n10697 ^ n10584 ;
  assign n10482 = n10481 ^ n10439 ;
  assign n10483 = n10482 ^ n10479 ;
  assign n10588 = n10584 ^ n10519 ;
  assign n10678 = ~n10483 & ~n10588 ;
  assign n10586 = ~n10483 & ~n10585 ;
  assign n10596 = n10586 ^ n10482 ;
  assign n10593 = n10482 & ~n10585 ;
  assign n10589 = n10482 & ~n10588 ;
  assign n10594 = n10593 ^ n10589 ;
  assign n10591 = n10482 & n10584 ;
  assign n10592 = n10591 ^ n10586 ;
  assign n10595 = n10594 ^ n10592 ;
  assign n10597 = n10596 ^ n10595 ;
  assign n10685 = n10678 ^ n10597 ;
  assign n10520 = ~n10483 & n10519 ;
  assign n10587 = n10586 ^ n10520 ;
  assign n10689 = n10685 ^ n10587 ;
  assign n10688 = n10595 ^ n10479 ;
  assign n10690 = n10689 ^ n10688 ;
  assign n10691 = n10690 ^ n10591 ;
  assign n10699 = n10698 ^ n10691 ;
  assign n10679 = n10678 ^ n10593 ;
  assign n10680 = n10679 ^ n10588 ;
  assign n10676 = n10480 & ~n10588 ;
  assign n10677 = n10676 ^ n10594 ;
  assign n10681 = n10680 ^ n10677 ;
  assign n10682 = n10681 ^ n10675 ;
  assign n11541 = n10699 ^ n10682 ;
  assign n11542 = n10669 & n11541 ;
  assign n11543 = n11542 ^ n10682 ;
  assign n11544 = n10633 & ~n11543 ;
  assign n11506 = n10669 ^ n10633 ;
  assign n11531 = n10674 ^ n10520 ;
  assign n11525 = n10696 ^ n10688 ;
  assign n11520 = n10691 ^ n10688 ;
  assign n11521 = n10691 ^ n10633 ;
  assign n11522 = n11506 & ~n11521 ;
  assign n11523 = n11522 ^ n10633 ;
  assign n11524 = n11520 & ~n11523 ;
  assign n11526 = n11525 ^ n11524 ;
  assign n11537 = n11531 ^ n11526 ;
  assign n10673 = n10480 & ~n10585 ;
  assign n11533 = n10673 ^ n10591 ;
  assign n11534 = n11533 ^ n10587 ;
  assign n11532 = n11531 ^ n10676 ;
  assign n11535 = n11534 ^ n11532 ;
  assign n11536 = ~n10669 & n11535 ;
  assign n11538 = n11537 ^ n11536 ;
  assign n11539 = n11506 & ~n11538 ;
  assign n10713 = n10697 ^ n10673 ;
  assign n11513 = n10713 ^ n10674 ;
  assign n11514 = n10674 ^ n10669 ;
  assign n11515 = n11514 ^ n10674 ;
  assign n11516 = n11513 & ~n11515 ;
  assign n11517 = n11516 ^ n10674 ;
  assign n11518 = ~n11506 & n11517 ;
  assign n10670 = ~n10633 & ~n10669 ;
  assign n10686 = n10670 & n10685 ;
  assign n11519 = n11518 ^ n10686 ;
  assign n11527 = n11526 ^ n11519 ;
  assign n10711 = n10676 ^ n10669 ;
  assign n11509 = n10711 ^ n10676 ;
  assign n11510 = n10677 & ~n11509 ;
  assign n11511 = n11510 ^ n10676 ;
  assign n11512 = n11506 & n11511 ;
  assign n11528 = n11527 ^ n11512 ;
  assign n10709 = n10670 ^ n10633 ;
  assign n10693 = n10585 ^ n10519 ;
  assign n10694 = n10480 & ~n10693 ;
  assign n10701 = n10694 ^ n10681 ;
  assign n11504 = n10701 ^ n10691 ;
  assign n11505 = ~n10709 & n11504 ;
  assign n11529 = n11528 ^ n11505 ;
  assign n11530 = n11529 ^ n8459 ;
  assign n11540 = n11539 ^ n11530 ;
  assign n11545 = n11544 ^ n11540 ;
  assign n11546 = n11545 ^ x98 ;
  assign n11581 = n11580 ^ x120 ;
  assign n11613 = n11612 ^ x96 ;
  assign n11823 = n11752 & n11793 ;
  assign n11820 = n11784 ^ n11766 ;
  assign n11821 = n11819 & ~n11820 ;
  assign n11796 = n11756 ^ n11668 ;
  assign n11797 = ~n11663 & n11796 ;
  assign n11798 = n11797 ^ n11778 ;
  assign n11814 = n11798 ^ n11789 ;
  assign n11808 = n11807 ^ n11756 ;
  assign n11809 = n11756 ^ n11663 ;
  assign n11810 = n11809 ^ n11756 ;
  assign n11811 = n11808 & ~n11810 ;
  assign n11812 = n11811 ^ n11756 ;
  assign n11813 = n11665 & n11812 ;
  assign n11815 = n11814 ^ n11813 ;
  assign n11799 = n11798 ^ n11756 ;
  assign n11800 = n11799 ^ n11775 ;
  assign n11801 = n11800 ^ n11799 ;
  assign n11804 = n11663 & n11801 ;
  assign n11805 = n11804 ^ n11799 ;
  assign n11806 = n11664 & n11805 ;
  assign n11816 = n11815 ^ n11806 ;
  assign n11817 = n11816 ^ n11795 ;
  assign n11818 = n11817 ^ n8634 ;
  assign n11822 = n11821 ^ n11818 ;
  assign n11824 = n11823 ^ n11822 ;
  assign n11780 = n11779 ^ n11740 ;
  assign n11790 = n11789 ^ n11780 ;
  assign n11741 = n11740 ^ n11738 ;
  assign n11747 = n11746 ^ n11741 ;
  assign n11748 = n11663 & n11747 ;
  assign n11791 = n11790 ^ n11748 ;
  assign n11792 = ~n11665 & ~n11791 ;
  assign n11825 = n11824 ^ n11792 ;
  assign n11826 = n11825 ^ x65 ;
  assign n12010 = ~n11613 & n11826 ;
  assign n12051 = n12010 ^ n11826 ;
  assign n9921 = n9725 ^ x75 ;
  assign n10311 = n10310 ^ x93 ;
  assign n10381 = ~n9921 & ~n10311 ;
  assign n10382 = n10381 ^ n9921 ;
  assign n10030 = n10029 ^ x94 ;
  assign n10058 = n10047 ^ n9169 ;
  assign n10061 = n10058 ^ n10055 ;
  assign n10056 = n9135 ^ n9134 ;
  assign n10057 = n10056 ^ n9125 ;
  assign n10059 = n10058 ^ n10057 ;
  assign n10060 = n8850 & n10059 ;
  assign n10062 = n10061 ^ n10060 ;
  assign n10063 = n10062 ^ n10055 ;
  assign n10048 = n10047 ^ n9148 ;
  assign n10049 = ~n8850 & n10048 ;
  assign n10064 = n10063 ^ n10049 ;
  assign n10065 = ~n9014 & n10064 ;
  assign n10066 = n10065 ^ n10062 ;
  assign n10044 = ~n9014 & ~n9147 ;
  assign n10042 = n9143 ^ n9137 ;
  assign n10043 = n10042 ^ n9169 ;
  assign n10045 = n10044 ^ n10043 ;
  assign n10046 = n8850 & ~n10045 ;
  assign n10067 = n10066 ^ n10046 ;
  assign n10041 = n9132 & ~n9180 ;
  assign n10068 = n10067 ^ n10041 ;
  assign n10036 = n10032 ^ n8850 ;
  assign n10037 = n10036 ^ n10032 ;
  assign n10038 = n10033 & n10037 ;
  assign n10039 = n10038 ^ n10032 ;
  assign n10040 = n9015 & n10039 ;
  assign n10069 = n10068 ^ n10040 ;
  assign n10070 = ~n9208 & ~n10069 ;
  assign n10071 = n10070 ^ n6656 ;
  assign n10072 = n10071 ^ x124 ;
  assign n10073 = n10030 & n10072 ;
  assign n10074 = n10073 ^ n10030 ;
  assign n10075 = n10074 ^ n10072 ;
  assign n10224 = n10186 ^ n10159 ;
  assign n10225 = ~n10078 & n10224 ;
  assign n10219 = n10195 & n10218 ;
  assign n10220 = n10219 ^ n10188 ;
  assign n10221 = n10202 & n10220 ;
  assign n10222 = n10221 ^ n10188 ;
  assign n10214 = n10159 ^ n10154 ;
  assign n10215 = n10214 ^ n10162 ;
  assign n10223 = n10222 ^ n10215 ;
  assign n10226 = n10225 ^ n10223 ;
  assign n10227 = n10226 ^ n10222 ;
  assign n10230 = n10227 ^ n10174 ;
  assign n10231 = n10230 ^ n10227 ;
  assign n10232 = ~n10078 & n10231 ;
  assign n10233 = n10232 ^ n10227 ;
  assign n10234 = ~n10077 & n10233 ;
  assign n10235 = n10234 ^ n10226 ;
  assign n10242 = ~n10235 & ~n10241 ;
  assign n10201 = n10200 ^ n5929 ;
  assign n10213 = n10212 ^ n10201 ;
  assign n10243 = n10242 ^ n10213 ;
  assign n10244 = n10243 ^ x76 ;
  assign n10245 = n8847 ^ x117 ;
  assign n10246 = ~n10244 & n10245 ;
  assign n10247 = n10246 ^ n10244 ;
  assign n10248 = n10247 ^ n10245 ;
  assign n10249 = n10248 ^ n10244 ;
  assign n10319 = ~n10075 & n10249 ;
  assign n10256 = n10074 & n10248 ;
  assign n10320 = n10319 ^ n10256 ;
  assign n10261 = n10073 & n10246 ;
  assign n10338 = n10320 ^ n10261 ;
  assign n10332 = n10246 ^ n10072 ;
  assign n10335 = n10244 ^ n10072 ;
  assign n10333 = n10245 ^ n10030 ;
  assign n10334 = n10333 ^ n10246 ;
  assign n10336 = n10335 ^ n10334 ;
  assign n10337 = ~n10332 & ~n10336 ;
  assign n10339 = n10338 ^ n10337 ;
  assign n10255 = n10073 & n10248 ;
  assign n10340 = n10339 ^ n10255 ;
  assign n10329 = n10073 & n10249 ;
  assign n10330 = n10329 ^ n10319 ;
  assign n10076 = n10075 ^ n10030 ;
  assign n10250 = n10076 & n10249 ;
  assign n10328 = n10250 ^ n10249 ;
  assign n10331 = n10330 ^ n10328 ;
  assign n10341 = n10340 ^ n10331 ;
  assign n10342 = n10341 ^ n10072 ;
  assign n10321 = n10074 & n10246 ;
  assign n10251 = n10076 & n10246 ;
  assign n10324 = n10321 ^ n10251 ;
  assign n10323 = n10261 ^ n10246 ;
  assign n10325 = n10324 ^ n10323 ;
  assign n10322 = n10321 ^ n10320 ;
  assign n10326 = n10325 ^ n10322 ;
  assign n10253 = ~n10075 & n10248 ;
  assign n10318 = n10255 ^ n10253 ;
  assign n10327 = n10326 ^ n10318 ;
  assign n10343 = n10342 ^ n10327 ;
  assign n10257 = n10256 ^ n10255 ;
  assign n10254 = n10253 ^ n10248 ;
  assign n10258 = n10257 ^ n10254 ;
  assign n11658 = n10343 ^ n10258 ;
  assign n11659 = ~n10382 & ~n11658 ;
  assign n11660 = n11659 ^ n8749 ;
  assign n10383 = n10382 ^ n10311 ;
  assign n10371 = n10329 ^ n10325 ;
  assign n11614 = n10383 ^ n10371 ;
  assign n11615 = n10381 ^ n10371 ;
  assign n11616 = n11615 ^ n10381 ;
  assign n11617 = n10337 ^ n10335 ;
  assign n11618 = n11617 ^ n10381 ;
  assign n11619 = ~n11616 & ~n11618 ;
  assign n11620 = n11619 ^ n10381 ;
  assign n11621 = ~n11614 & n11620 ;
  assign n11622 = n11621 ^ n10383 ;
  assign n11629 = n10383 ^ n10381 ;
  assign n11643 = n10311 & n10320 ;
  assign n11644 = n11643 ^ n10256 ;
  assign n11645 = n11629 & n11644 ;
  assign n11631 = n10339 ^ n10253 ;
  assign n11632 = n11631 ^ n10258 ;
  assign n10252 = n10251 ^ n10250 ;
  assign n11630 = n10261 ^ n10252 ;
  assign n11633 = n11632 ^ n11630 ;
  assign n11634 = n11632 ^ n10311 ;
  assign n11635 = n11634 ^ n11632 ;
  assign n11636 = n11633 & n11635 ;
  assign n11637 = n11636 ^ n11632 ;
  assign n11638 = n11629 & n11637 ;
  assign n11646 = n11645 ^ n11638 ;
  assign n11626 = n10261 ^ n10253 ;
  assign n11623 = n10325 ^ n10253 ;
  assign n10357 = n10321 ^ n10250 ;
  assign n11624 = n11623 ^ n10357 ;
  assign n11625 = n9921 & n11624 ;
  assign n11627 = n11626 ^ n11625 ;
  assign n11628 = ~n10311 & n11627 ;
  assign n11647 = n11646 ^ n11628 ;
  assign n11648 = ~n9921 & ~n11647 ;
  assign n10259 = n10258 ^ n10076 ;
  assign n10260 = n10259 ^ n10252 ;
  assign n10344 = n10343 ^ n10260 ;
  assign n10345 = n10344 ^ n10340 ;
  assign n10346 = n10345 ^ n10257 ;
  assign n11653 = ~n10311 & ~n10346 ;
  assign n11654 = n11653 ^ n10257 ;
  assign n11655 = n11648 & n11654 ;
  assign n11656 = n11655 ^ n11647 ;
  assign n11657 = n11622 & ~n11656 ;
  assign n11661 = n11660 ^ n11657 ;
  assign n11662 = n11661 ^ x105 ;
  assign n11975 = n11905 ^ n11883 ;
  assign n11936 = n11923 ^ n11903 ;
  assign n11937 = n11936 ^ n11935 ;
  assign n11938 = n11937 ^ n11934 ;
  assign n11939 = n11830 & ~n11938 ;
  assign n11940 = n11939 ^ n11923 ;
  assign n11976 = n11975 ^ n11940 ;
  assign n11908 = n11907 ^ n11830 ;
  assign n11909 = n11908 ^ n11829 ;
  assign n11972 = n11933 ^ n11903 ;
  assign n11973 = ~n11909 & ~n11972 ;
  assign n11974 = n11973 ^ n11971 ;
  assign n11977 = n11976 ^ n11974 ;
  assign n11953 = n11942 ^ n11929 ;
  assign n11954 = ~n11830 & n11953 ;
  assign n11955 = n11954 ^ n11929 ;
  assign n11956 = n11955 ^ n11917 ;
  assign n11957 = n11956 ^ n11883 ;
  assign n11958 = n11957 ^ n11955 ;
  assign n11961 = n11830 & n11958 ;
  assign n11962 = n11961 ^ n11955 ;
  assign n11963 = n11952 & n11962 ;
  assign n11964 = n11963 ^ n11955 ;
  assign n11978 = n11977 ^ n11964 ;
  assign n11941 = n11940 ^ n11903 ;
  assign n11945 = n11944 ^ n11941 ;
  assign n11946 = n11945 ^ n11940 ;
  assign n11949 = n11830 & n11946 ;
  assign n11950 = n11949 ^ n11940 ;
  assign n11951 = n11829 & n11950 ;
  assign n11979 = n11978 ^ n11951 ;
  assign n11906 = n11905 ^ n11898 ;
  assign n11910 = n11909 ^ n11901 ;
  assign n11911 = n11901 ^ n11898 ;
  assign n11912 = n11911 ^ n11901 ;
  assign n11913 = n11910 & ~n11912 ;
  assign n11914 = n11913 ^ n11901 ;
  assign n11915 = n11906 & n11914 ;
  assign n11980 = n11979 ^ n11915 ;
  assign n11884 = n11883 ^ n11830 ;
  assign n11885 = n11884 ^ n11883 ;
  assign n11895 = n11885 & n11892 ;
  assign n11896 = n11895 ^ n11883 ;
  assign n11897 = ~n11829 & n11896 ;
  assign n11981 = n11980 ^ n11897 ;
  assign n11993 = n11992 ^ n11920 ;
  assign n11994 = n11993 ^ n11942 ;
  assign n11995 = n11942 ^ n11830 ;
  assign n11996 = n11995 ^ n11942 ;
  assign n11997 = ~n11994 & n11996 ;
  assign n11998 = n11997 ^ n11942 ;
  assign n11999 = n11829 & n11998 ;
  assign n12000 = ~n11981 & ~n11999 ;
  assign n12001 = n12000 ^ n8679 ;
  assign n12002 = n12001 ^ x115 ;
  assign n12007 = ~n11662 & ~n12002 ;
  assign n12011 = n12010 ^ n11613 ;
  assign n12032 = n12011 ^ n11826 ;
  assign n12033 = n12007 & n12032 ;
  assign n11827 = n11826 ^ n11662 ;
  assign n12024 = n11662 ^ n11613 ;
  assign n12025 = ~n11827 & ~n12024 ;
  assign n12026 = n12025 ^ n11613 ;
  assign n12027 = n12002 & ~n12026 ;
  assign n12008 = n12007 ^ n12002 ;
  assign n12009 = n12008 ^ n11662 ;
  assign n12018 = ~n12009 & n12010 ;
  assign n12028 = n12027 ^ n12018 ;
  assign n12014 = n12007 ^ n11662 ;
  assign n12015 = ~n12011 & ~n12014 ;
  assign n12019 = n12018 ^ n12015 ;
  assign n12017 = n12007 & n12010 ;
  assign n12020 = n12019 ^ n12017 ;
  assign n12021 = n12020 ^ n12010 ;
  assign n12013 = ~n12008 & n12010 ;
  assign n12016 = n12015 ^ n12013 ;
  assign n12022 = n12021 ^ n12016 ;
  assign n12012 = ~n12009 & ~n12011 ;
  assign n12023 = n12022 ^ n12012 ;
  assign n12029 = n12028 ^ n12023 ;
  assign n12037 = n12033 ^ n12029 ;
  assign n12003 = n12002 ^ n11613 ;
  assign n12004 = ~n11827 & n12003 ;
  assign n12034 = n12033 ^ n12004 ;
  assign n12035 = n12034 ^ n12019 ;
  assign n12036 = n12035 ^ n12033 ;
  assign n12038 = n12037 ^ n12036 ;
  assign n12031 = n12025 ^ n12015 ;
  assign n12039 = n12038 ^ n12031 ;
  assign n12043 = n12039 ^ n12017 ;
  assign n12042 = n12033 ^ n12007 ;
  assign n12044 = n12043 ^ n12042 ;
  assign n12052 = n12051 ^ n12044 ;
  assign n12053 = n12052 ^ n12038 ;
  assign n12054 = n12053 ^ n12039 ;
  assign n11828 = n11827 ^ n11613 ;
  assign n12005 = n12004 ^ n11828 ;
  assign n12048 = n12002 ^ n11826 ;
  assign n12049 = ~n12005 & ~n12048 ;
  assign n12050 = n12049 ^ n12033 ;
  assign n12055 = n12054 ^ n12050 ;
  assign n13344 = n12055 ^ n12035 ;
  assign n13345 = n13344 ^ n12017 ;
  assign n13346 = ~n11581 & n13345 ;
  assign n13335 = n12043 ^ n12015 ;
  assign n13347 = n13346 ^ n13335 ;
  assign n13348 = ~n11546 & n13347 ;
  assign n12056 = n12055 ^ n12029 ;
  assign n12057 = n12056 ^ n12053 ;
  assign n12058 = n12053 ^ n11581 ;
  assign n12059 = n12058 ^ n12053 ;
  assign n12060 = n12057 & n12059 ;
  assign n12061 = n12060 ^ n12053 ;
  assign n12062 = n11546 & n12061 ;
  assign n13336 = n13335 ^ n12062 ;
  assign n12089 = ~n12008 & ~n12011 ;
  assign n12090 = n12089 ^ n12022 ;
  assign n13329 = n12090 ^ n12033 ;
  assign n13330 = n12033 ^ n11581 ;
  assign n13331 = n13330 ^ n12033 ;
  assign n13332 = n13329 & ~n13331 ;
  assign n13333 = n13332 ^ n12033 ;
  assign n13334 = ~n11546 & n13333 ;
  assign n13337 = n13336 ^ n13334 ;
  assign n12063 = n11581 ^ n11546 ;
  assign n12076 = n12015 ^ n11546 ;
  assign n12077 = n12076 ^ n12015 ;
  assign n13326 = n12016 & n12077 ;
  assign n13327 = n13326 ^ n12015 ;
  assign n13328 = ~n12063 & n13327 ;
  assign n13338 = n13337 ^ n13328 ;
  assign n12109 = n12027 ^ n12009 ;
  assign n12110 = n12109 ^ n12022 ;
  assign n11582 = n11546 & n11581 ;
  assign n12071 = n11582 ^ n11581 ;
  assign n12111 = n12071 ^ n11546 ;
  assign n12112 = ~n12110 & ~n12111 ;
  assign n12102 = n12039 ^ n11581 ;
  assign n12103 = n12102 ^ n12039 ;
  assign n12106 = n12054 & ~n12103 ;
  assign n12107 = n12106 ^ n12039 ;
  assign n12108 = ~n11546 & n12107 ;
  assign n12113 = n12112 ^ n12108 ;
  assign n13339 = n13338 ^ n12113 ;
  assign n12030 = n12029 ^ n12013 ;
  assign n12040 = n12039 ^ n12030 ;
  assign n12006 = n12005 ^ n11613 ;
  assign n12041 = n12040 ^ n12006 ;
  assign n12045 = n12044 ^ n12041 ;
  assign n12087 = ~n12045 & n12071 ;
  assign n12081 = n12035 ^ n12012 ;
  assign n12082 = n12012 ^ n11546 ;
  assign n12083 = n12082 ^ n12012 ;
  assign n12084 = n12081 & ~n12083 ;
  assign n12085 = n12084 ^ n12012 ;
  assign n12086 = n12063 & n12085 ;
  assign n12088 = n12087 ^ n12086 ;
  assign n13340 = n13339 ^ n12088 ;
  assign n13341 = n13340 ^ n8847 ;
  assign n13317 = n12110 ^ n12044 ;
  assign n13316 = n12055 ^ n12036 ;
  assign n13318 = n13317 ^ n13316 ;
  assign n13319 = n13316 ^ n11581 ;
  assign n13320 = n13319 ^ n13316 ;
  assign n13321 = ~n13318 & n13320 ;
  assign n13322 = n13321 ^ n13316 ;
  assign n13323 = n11546 & n13322 ;
  assign n13342 = n13341 ^ n13323 ;
  assign n13313 = n12089 ^ n12023 ;
  assign n13314 = n13313 ^ n12027 ;
  assign n13315 = n12071 & n13314 ;
  assign n13343 = n13342 ^ n13315 ;
  assign n13349 = n13348 ^ n13343 ;
  assign n13350 = n13349 ^ x93 ;
  assign n12832 = n11545 ^ x73 ;
  assign n12377 = n11659 ^ n10253 ;
  assign n12360 = n10338 ^ n10250 ;
  assign n12367 = n12360 ^ n10340 ;
  assign n10358 = n10357 ^ n10331 ;
  assign n12361 = n10358 ^ n10319 ;
  assign n12362 = n12361 ^ n12360 ;
  assign n10317 = n10311 ^ n9921 ;
  assign n12363 = n12360 ^ n9921 ;
  assign n12364 = n10317 & n12363 ;
  assign n12365 = n12364 ^ n9921 ;
  assign n12366 = n12362 & n12365 ;
  assign n12368 = n12367 ^ n12366 ;
  assign n12378 = n12377 ^ n12368 ;
  assign n10262 = n10261 ^ n10260 ;
  assign n10314 = n10262 & ~n10311 ;
  assign n10315 = n10314 ^ n10261 ;
  assign n10316 = ~n9921 & n10315 ;
  assign n12379 = n12378 ^ n10316 ;
  assign n12380 = n12379 ^ n11645 ;
  assign n12371 = n10252 ^ n10247 ;
  assign n12372 = n12371 ^ n10344 ;
  assign n12373 = n12372 ^ n10371 ;
  assign n12374 = ~n10311 & n12373 ;
  assign n12369 = n12368 ^ n10247 ;
  assign n12370 = n12369 ^ n10344 ;
  assign n12375 = n12374 ^ n12370 ;
  assign n12376 = n11629 & n12375 ;
  assign n12381 = n12380 ^ n12376 ;
  assign n12354 = n10311 ^ n10253 ;
  assign n12355 = n12354 ^ n10253 ;
  assign n12357 = n10325 & n12355 ;
  assign n12358 = n12357 ^ n10253 ;
  assign n12359 = ~n9921 & n12358 ;
  assign n12382 = n12381 ^ n12359 ;
  assign n12383 = n12382 ^ n10251 ;
  assign n12384 = n12383 ^ n12382 ;
  assign n10347 = n10256 ^ n10247 ;
  assign n10348 = n10347 ^ n10346 ;
  assign n12385 = n12384 ^ n10348 ;
  assign n12386 = ~n9921 & n12385 ;
  assign n12387 = n12386 ^ n12383 ;
  assign n12398 = n12387 ^ n9041 ;
  assign n12388 = n12387 ^ n12382 ;
  assign n12389 = n12388 ^ n12387 ;
  assign n12390 = n10344 ^ n10331 ;
  assign n12391 = ~n10311 & ~n12390 ;
  assign n12392 = n12391 ^ n10331 ;
  assign n12395 = ~n12389 & ~n12392 ;
  assign n12396 = n12395 ^ n12387 ;
  assign n12397 = n10317 & ~n12396 ;
  assign n12399 = n12398 ^ n12397 ;
  assign n12833 = n12399 ^ x64 ;
  assign n12834 = ~n12832 & ~n12833 ;
  assign n12905 = n12834 ^ n12832 ;
  assign n11365 = n11362 ^ n11336 ;
  assign n11366 = n11365 ^ n11357 ;
  assign n11363 = n11362 ^ n11360 ;
  assign n11364 = n11363 ^ n11335 ;
  assign n11367 = n11366 ^ n11364 ;
  assign n12498 = n11367 & n11372 ;
  assign n12499 = ~n11577 & n12498 ;
  assign n12500 = n12499 ^ n11577 ;
  assign n12868 = n12500 ^ n9085 ;
  assign n11370 = n11265 & ~n11360 ;
  assign n11368 = n11367 ^ n11327 ;
  assign n11369 = ~n11266 & n11368 ;
  assign n11371 = n11370 ^ n11369 ;
  assign n12869 = n12868 ^ n11371 ;
  assign n12492 = n11266 ^ n11264 ;
  assign n12493 = n11346 ^ n11329 ;
  assign n12494 = n12492 & ~n12493 ;
  assign n12479 = n11264 ^ n11239 ;
  assign n12836 = n11359 ^ n11264 ;
  assign n12837 = n12836 ^ n11359 ;
  assign n11378 = n11377 ^ n11351 ;
  assign n12846 = n11378 ^ n11346 ;
  assign n12847 = n11265 & ~n12846 ;
  assign n12840 = n11345 ^ n11264 ;
  assign n12841 = n12840 ^ n11345 ;
  assign n12842 = n11366 & ~n12841 ;
  assign n12843 = n12842 ^ n11345 ;
  assign n12844 = ~n12479 & ~n12843 ;
  assign n12845 = n12844 ^ n11328 ;
  assign n12848 = n12847 ^ n12845 ;
  assign n12849 = n12848 ^ n11331 ;
  assign n12850 = n12849 ^ n12848 ;
  assign n12851 = n12850 ^ n11359 ;
  assign n12852 = ~n12837 & n12851 ;
  assign n12853 = n12852 ^ n11359 ;
  assign n12854 = ~n12479 & n12853 ;
  assign n12855 = n12854 ^ n12849 ;
  assign n12856 = n12855 ^ n11354 ;
  assign n12857 = n12856 ^ n11354 ;
  assign n12858 = n12857 ^ n12856 ;
  assign n12859 = n12857 ^ n12492 ;
  assign n12860 = n12859 ^ n12857 ;
  assign n12861 = n12857 ^ n12848 ;
  assign n12862 = n12861 ^ n12857 ;
  assign n12863 = n12860 & n12862 ;
  assign n12864 = n12858 & n12863 ;
  assign n12865 = n12864 ^ n12858 ;
  assign n12866 = n12865 ^ n12856 ;
  assign n12867 = ~n12494 & n12866 ;
  assign n12870 = n12869 ^ n12867 ;
  assign n12871 = n12870 ^ x90 ;
  assign n10956 = n10900 ^ n10793 ;
  assign n10957 = n10956 ^ n10900 ;
  assign n10960 = ~n10923 & ~n10957 ;
  assign n10961 = n10960 ^ n10900 ;
  assign n10962 = ~n10948 & n10961 ;
  assign n12654 = n10793 & n10904 ;
  assign n12655 = n12654 ^ n10903 ;
  assign n12657 = n12655 ^ n10885 ;
  assign n12656 = n12655 ^ n10933 ;
  assign n12658 = n12657 ^ n12656 ;
  assign n12661 = n10793 & ~n12658 ;
  assign n12662 = n12661 ^ n12657 ;
  assign n12663 = n10907 & n12662 ;
  assign n12664 = n12663 ^ n12655 ;
  assign n12872 = ~n10962 & ~n12664 ;
  assign n10913 = n10793 & ~n10907 ;
  assign n10963 = n10913 & ~n10940 ;
  assign n12891 = n10963 ^ n10940 ;
  assign n10906 = n10905 ^ n10902 ;
  assign n10910 = n10906 & n10907 ;
  assign n10911 = n10910 ^ n10902 ;
  assign n10912 = ~n10793 & n10911 ;
  assign n12892 = n12891 ^ n10912 ;
  assign n12888 = n10927 ^ n10889 ;
  assign n12889 = n12888 ^ n10941 ;
  assign n12890 = n10948 & ~n12889 ;
  assign n12893 = n12892 ^ n12890 ;
  assign n12887 = ~n10793 & ~n10889 ;
  assign n12894 = n12893 ^ n12887 ;
  assign n12880 = n10940 ^ n10793 ;
  assign n12881 = n12880 ^ n10940 ;
  assign n12882 = n10940 ^ n10897 ;
  assign n12883 = n12882 ^ n10940 ;
  assign n12884 = ~n12881 & n12883 ;
  assign n12885 = n12884 ^ n10940 ;
  assign n12886 = n10907 & ~n12885 ;
  assign n12895 = n12894 ^ n12886 ;
  assign n12873 = n10898 ^ n10886 ;
  assign n12874 = n12873 ^ n10898 ;
  assign n12875 = n10898 ^ n10793 ;
  assign n12876 = n12875 ^ n10898 ;
  assign n12877 = n12874 & n12876 ;
  assign n12878 = n12877 ^ n10898 ;
  assign n12879 = ~n10948 & n12878 ;
  assign n12896 = n12895 ^ n12879 ;
  assign n12897 = ~n10980 & n12896 ;
  assign n12898 = n12872 & n12897 ;
  assign n12899 = n12898 ^ n9120 ;
  assign n12900 = n12899 ^ x112 ;
  assign n12901 = n12871 & n12900 ;
  assign n12902 = n12901 ^ n12900 ;
  assign n12903 = n12902 ^ n12871 ;
  assign n12915 = n12903 ^ n12900 ;
  assign n12931 = ~n12905 & n12915 ;
  assign n12829 = n11825 ^ x114 ;
  assign n12464 = n12463 ^ n11204 ;
  assign n12453 = n11199 ^ n11158 ;
  assign n12444 = n11187 ^ n11185 ;
  assign n12445 = n12444 ^ n11169 ;
  assign n12446 = n12445 ^ n11201 ;
  assign n12454 = n12453 ^ n12446 ;
  assign n12447 = n11169 ^ n11162 ;
  assign n12448 = ~n12446 & n12447 ;
  assign n12452 = n11100 & n12448 ;
  assign n12455 = n12454 ^ n12452 ;
  assign n12465 = n12464 ^ n12455 ;
  assign n12459 = n11168 ^ n11159 ;
  assign n12460 = n12459 ^ n11200 ;
  assign n12461 = n12460 ^ n11165 ;
  assign n12462 = ~n11100 & n12461 ;
  assign n12466 = n12465 ^ n12462 ;
  assign n12467 = ~n11162 & n12466 ;
  assign n12442 = n11170 & ~n11213 ;
  assign n11174 = n11173 ^ n11163 ;
  assign n11175 = n11173 ^ n11100 ;
  assign n11176 = n11175 ^ n11173 ;
  assign n11177 = n11174 & n11176 ;
  assign n11178 = n11177 ^ n11173 ;
  assign n11179 = ~n11162 & ~n11178 ;
  assign n12443 = n12442 ^ n11179 ;
  assign n12449 = n12448 ^ n12443 ;
  assign n11222 = n11187 ^ n11163 ;
  assign n11223 = n11187 ^ n11100 ;
  assign n11224 = n11223 ^ n11187 ;
  assign n11225 = n11222 & ~n11224 ;
  assign n11226 = n11225 ^ n11187 ;
  assign n11227 = ~n11162 & ~n11226 ;
  assign n12450 = n12449 ^ n11227 ;
  assign n12451 = n12450 ^ n9013 ;
  assign n12456 = n12455 ^ n12451 ;
  assign n12436 = n11157 ^ n11100 ;
  assign n12437 = n12436 ^ n11157 ;
  assign n12438 = n11171 ^ n11157 ;
  assign n12439 = n12437 & n12438 ;
  assign n12440 = n12439 ^ n11157 ;
  assign n12441 = ~n11101 & ~n12440 ;
  assign n12457 = n12456 ^ n12441 ;
  assign n11197 = n11173 ^ n11168 ;
  assign n11202 = n11201 ^ n11197 ;
  assign n12434 = n12433 ^ n11202 ;
  assign n12435 = ~n11214 & ~n12434 ;
  assign n12458 = n12457 ^ n12435 ;
  assign n12468 = n12467 ^ n12458 ;
  assign n12830 = n12468 ^ x123 ;
  assign n12950 = n12829 & ~n12830 ;
  assign n12951 = n12950 ^ n12829 ;
  assign n13351 = n12931 & n12951 ;
  assign n12916 = n12834 & n12915 ;
  assign n12970 = n12916 & n12951 ;
  assign n13352 = n13351 ^ n12970 ;
  assign n12835 = n12834 ^ n12833 ;
  assign n12920 = n12835 ^ n12832 ;
  assign n12924 = ~n12903 & ~n12920 ;
  assign n12987 = n12924 & n12950 ;
  assign n12967 = ~n12835 & n12915 ;
  assign n12906 = n12902 & ~n12905 ;
  assign n12981 = n12967 ^ n12906 ;
  assign n12982 = n12906 ^ n12830 ;
  assign n12983 = n12982 ^ n12906 ;
  assign n12984 = n12981 & ~n12983 ;
  assign n12985 = n12984 ^ n12906 ;
  assign n12986 = n12829 & n12985 ;
  assign n12988 = n12987 ^ n12986 ;
  assign n12917 = n12834 & ~n12871 ;
  assign n12918 = n12917 ^ n12834 ;
  assign n12919 = n12918 ^ n12916 ;
  assign n12932 = n12931 ^ n12919 ;
  assign n13353 = n12932 & n12950 ;
  assign n12904 = ~n12835 & ~n12903 ;
  assign n12952 = n12951 ^ n12830 ;
  assign n12953 = n12952 ^ n12829 ;
  assign n12980 = n12904 & ~n12953 ;
  assign n13354 = n13353 ^ n12980 ;
  assign n12831 = n12830 ^ n12829 ;
  assign n12921 = n12901 & ~n12920 ;
  assign n12954 = n12921 ^ n12920 ;
  assign n12927 = n12902 & ~n12920 ;
  assign n12928 = n12927 ^ n12924 ;
  assign n12955 = n12954 ^ n12928 ;
  assign n12958 = n12927 ^ n12829 ;
  assign n12959 = n12958 ^ n12927 ;
  assign n12962 = ~n12955 & ~n12959 ;
  assign n12963 = n12962 ^ n12927 ;
  assign n12964 = n12831 & n12963 ;
  assign n12965 = n12964 ^ n12927 ;
  assign n12922 = n12921 ^ n12919 ;
  assign n12913 = n12901 & ~n12905 ;
  assign n12914 = n12913 ^ n12901 ;
  assign n12923 = n12922 ^ n12914 ;
  assign n13376 = n12923 & n12952 ;
  assign n12969 = n12931 & ~n12953 ;
  assign n13356 = n12969 ^ n12919 ;
  assign n12998 = ~n12903 & ~n12905 ;
  assign n12935 = n12927 ^ n12904 ;
  assign n12936 = n12935 ^ n12923 ;
  assign n12937 = n12936 ^ n12913 ;
  assign n12933 = n12924 ^ n12906 ;
  assign n12934 = n12933 ^ n12932 ;
  assign n12938 = n12937 ^ n12934 ;
  assign n12930 = n12905 ^ n12903 ;
  assign n12939 = n12938 ^ n12930 ;
  assign n12929 = n12928 ^ n12916 ;
  assign n12940 = n12939 ^ n12929 ;
  assign n12925 = n12924 ^ n12923 ;
  assign n12926 = n12925 ^ n12834 ;
  assign n12941 = n12940 ^ n12926 ;
  assign n12999 = n12998 ^ n12941 ;
  assign n13357 = n13356 ^ n12999 ;
  assign n13355 = n12906 & n12952 ;
  assign n13358 = n13357 ^ n13355 ;
  assign n12942 = n12941 ^ n12935 ;
  assign n13372 = n13358 ^ n12942 ;
  assign n12907 = n12906 ^ n12904 ;
  assign n12912 = n12907 ^ n12902 ;
  assign n12943 = n12942 ^ n12912 ;
  assign n13369 = n12943 ^ n12917 ;
  assign n12960 = n12955 ^ n12927 ;
  assign n13370 = n13369 ^ n12960 ;
  assign n13371 = n12830 & ~n13370 ;
  assign n13373 = n13372 ^ n13371 ;
  assign n13374 = n12829 & n13373 ;
  assign n13365 = n12967 ^ n12921 ;
  assign n13366 = n12952 & n13365 ;
  assign n13359 = n12925 ^ n12913 ;
  assign n13360 = n12913 ^ n12829 ;
  assign n13361 = n13360 ^ n12913 ;
  assign n13362 = n13359 & ~n13361 ;
  assign n13363 = n13362 ^ n12913 ;
  assign n13364 = ~n12830 & n13363 ;
  assign n13367 = n13366 ^ n13364 ;
  assign n13368 = n13367 ^ n13358 ;
  assign n13375 = n13374 ^ n13368 ;
  assign n13377 = n13376 ^ n13375 ;
  assign n13378 = ~n12965 & ~n13377 ;
  assign n13379 = ~n13354 & n13378 ;
  assign n13380 = ~n12988 & n13379 ;
  assign n13381 = ~n13352 & n13380 ;
  assign n13382 = n13381 ^ n10071 ;
  assign n13383 = n13382 ^ x100 ;
  assign n13384 = n13350 & n13383 ;
  assign n13385 = n13384 ^ n13350 ;
  assign n13460 = n13385 ^ n13383 ;
  assign n10384 = n10348 & ~n10383 ;
  assign n10365 = n10330 ^ n10324 ;
  assign n10366 = n10365 ^ n10343 ;
  assign n10367 = n10366 ^ n10339 ;
  assign n10359 = n10358 ^ n10251 ;
  assign n10360 = n10359 ^ n10311 ;
  assign n10361 = n10317 ^ n10311 ;
  assign n10362 = n10360 & ~n10361 ;
  assign n10363 = n10362 ^ n10311 ;
  assign n10364 = n10249 & ~n10363 ;
  assign n10368 = n10367 ^ n10364 ;
  assign n10377 = n10368 ^ n10327 ;
  assign n10349 = n10348 ^ n10253 ;
  assign n10373 = n10349 ^ n10256 ;
  assign n10374 = n10373 ^ n10258 ;
  assign n10370 = n10327 ^ n10251 ;
  assign n10372 = n10371 ^ n10370 ;
  assign n10375 = n10374 ^ n10372 ;
  assign n10376 = n10311 & n10375 ;
  assign n10378 = n10377 ^ n10376 ;
  assign n10379 = ~n9921 & ~n10378 ;
  assign n10369 = n10368 ^ n10258 ;
  assign n10380 = n10379 ^ n10369 ;
  assign n10385 = n10384 ^ n10380 ;
  assign n10350 = n10349 ^ n10258 ;
  assign n10351 = n10350 ^ n10258 ;
  assign n10352 = n10258 ^ n9921 ;
  assign n10353 = n10352 ^ n10258 ;
  assign n10354 = n10351 & n10353 ;
  assign n10355 = n10354 ^ n10258 ;
  assign n10356 = n10317 & n10355 ;
  assign n10386 = n10385 ^ n10356 ;
  assign n10387 = ~n10316 & n10386 ;
  assign n10388 = n10387 ^ n6909 ;
  assign n10389 = n10388 ^ x78 ;
  assign n10683 = n10682 ^ n10673 ;
  assign n10671 = n10670 ^ n10669 ;
  assign n10684 = ~n10671 & ~n10681 ;
  assign n10687 = n10686 ^ n10684 ;
  assign n10714 = n10713 ^ n10694 ;
  assign n10717 = n10714 ^ n10676 ;
  assign n10700 = n10699 ^ n10674 ;
  assign n10712 = n10700 ^ n10593 ;
  assign n10715 = n10714 ^ n10712 ;
  assign n10716 = n10633 & ~n10715 ;
  assign n10718 = n10717 ^ n10716 ;
  assign n10719 = n10711 & n10718 ;
  assign n10720 = n10719 ^ n10676 ;
  assign n10710 = n10595 & ~n10709 ;
  assign n10721 = n10720 ^ n10710 ;
  assign n10702 = n10701 ^ n10700 ;
  assign n10692 = n10691 ^ n10597 ;
  assign n10695 = n10694 ^ n10692 ;
  assign n10703 = n10702 ^ n10695 ;
  assign n10704 = n10695 ^ n10633 ;
  assign n10705 = n10704 ^ n10695 ;
  assign n10706 = ~n10703 & ~n10705 ;
  assign n10707 = n10706 ^ n10695 ;
  assign n10708 = ~n10669 & ~n10707 ;
  assign n10722 = n10721 ^ n10708 ;
  assign n10723 = n10670 ^ n10586 ;
  assign n10724 = n10723 ^ n10722 ;
  assign n10672 = n10671 ^ n10633 ;
  assign n10725 = n10690 ^ n10672 ;
  assign n10726 = ~n10670 & ~n10725 ;
  assign n10727 = n10726 ^ n10690 ;
  assign n10728 = n10724 & n10727 ;
  assign n10729 = n10728 ^ n10670 ;
  assign n10730 = ~n10722 & ~n10729 ;
  assign n10731 = ~n10687 & n10730 ;
  assign n10732 = ~n10671 & n10731 ;
  assign n10733 = ~n10683 & n10732 ;
  assign n10734 = n10733 ^ n10731 ;
  assign n10737 = n10734 ^ n9269 ;
  assign n10590 = n10589 ^ n10587 ;
  assign n10598 = n10597 ^ n10590 ;
  assign n10735 = ~n10672 & n10734 ;
  assign n10736 = n10598 & n10735 ;
  assign n10738 = n10737 ^ n10736 ;
  assign n10739 = n10738 ^ x75 ;
  assign n10970 = n10900 & n10948 ;
  assign n10914 = n10913 ^ n10793 ;
  assign n10967 = n10914 & ~n10966 ;
  assign n10964 = n10963 ^ n10962 ;
  assign n10935 = n10934 ^ n10793 ;
  assign n10936 = n10935 ^ n10934 ;
  assign n10942 = n10933 & ~n10941 ;
  assign n10943 = n10942 ^ n10934 ;
  assign n10944 = n10936 & ~n10943 ;
  assign n10945 = n10944 ^ n10934 ;
  assign n10946 = n10907 & ~n10945 ;
  assign n10947 = n10946 ^ n10933 ;
  assign n10951 = ~n10793 & ~n10931 ;
  assign n10952 = n10951 ^ n10882 ;
  assign n10953 = ~n10948 & ~n10952 ;
  assign n10954 = n10953 ^ n10882 ;
  assign n10955 = n10947 & n10954 ;
  assign n10965 = n10964 ^ n10955 ;
  assign n10968 = n10967 ^ n10965 ;
  assign n10915 = n10914 ^ n10907 ;
  assign n10916 = n10898 & n10915 ;
  assign n10969 = n10968 ^ n10916 ;
  assign n10971 = n10970 ^ n10969 ;
  assign n10981 = n10971 & ~n10980 ;
  assign n10982 = ~n10912 & n10981 ;
  assign n10983 = n10982 ^ n8342 ;
  assign n10984 = n10983 ^ x100 ;
  assign n10985 = ~n10739 & ~n10984 ;
  assign n10986 = n10985 ^ n10739 ;
  assign n10987 = n10986 ^ n10984 ;
  assign n11103 = n11068 & n11102 ;
  assign n11219 = ~n11100 & n11159 ;
  assign n11215 = n11200 ^ n11170 ;
  assign n11216 = ~n11214 & n11215 ;
  assign n11205 = n11204 ^ n11201 ;
  assign n11184 = n11166 ^ n11157 ;
  assign n11186 = n11185 ^ n11184 ;
  assign n11192 = n11191 ^ n11186 ;
  assign n11193 = n11100 & n11192 ;
  assign n11194 = n11193 ^ n11191 ;
  assign n11206 = n11205 ^ n11194 ;
  assign n11203 = n11202 ^ n11199 ;
  assign n11207 = n11206 ^ n11203 ;
  assign n11208 = n11207 ^ n11194 ;
  assign n11209 = n11100 & ~n11208 ;
  assign n11210 = n11209 ^ n11206 ;
  assign n11211 = ~n11162 & ~n11210 ;
  assign n11182 = n11181 ^ n11156 ;
  assign n11183 = ~n11180 & n11182 ;
  assign n11195 = n11194 ^ n11183 ;
  assign n11196 = n11195 ^ n11179 ;
  assign n11212 = n11211 ^ n11196 ;
  assign n11217 = n11216 ^ n11212 ;
  assign n11160 = n11159 ^ n11158 ;
  assign n11161 = ~n11101 & ~n11160 ;
  assign n11218 = n11217 ^ n11161 ;
  assign n11220 = n11219 ^ n11218 ;
  assign n11221 = ~n11103 & n11220 ;
  assign n11235 = ~n11227 & ~n11234 ;
  assign n11236 = n11221 & n11235 ;
  assign n11237 = n11236 ^ n10146 ;
  assign n11238 = n11237 ^ x102 ;
  assign n11415 = n11414 ^ n10114 ;
  assign n11405 = n11361 ^ n11343 ;
  assign n11397 = n11342 ^ n11325 ;
  assign n11396 = n11363 ^ n11351 ;
  assign n11398 = n11397 ^ n11396 ;
  assign n11399 = n11239 & ~n11398 ;
  assign n11400 = n11399 ^ n11397 ;
  assign n11408 = n11405 ^ n11400 ;
  assign n11404 = n11349 ^ n11336 ;
  assign n11406 = n11405 ^ n11404 ;
  assign n11407 = ~n11239 & n11406 ;
  assign n11409 = n11408 ^ n11407 ;
  assign n11410 = n11264 & n11409 ;
  assign n11379 = n11378 ^ n11357 ;
  assign n11401 = n11400 ^ n11379 ;
  assign n11402 = n11401 ^ n11395 ;
  assign n11382 = n11332 ^ n11239 ;
  assign n11383 = n11382 ^ n11332 ;
  assign n11386 = ~n11333 & ~n11383 ;
  assign n11387 = n11386 ^ n11332 ;
  assign n11388 = ~n11373 & n11387 ;
  assign n11403 = n11402 ^ n11388 ;
  assign n11411 = n11410 ^ n11403 ;
  assign n11374 = n11367 ^ n11329 ;
  assign n11375 = n11374 ^ n11343 ;
  assign n11380 = n11379 ^ n11375 ;
  assign n11381 = n11373 & n11380 ;
  assign n11412 = n11411 ^ n11381 ;
  assign n11413 = ~n11371 & n11412 ;
  assign n11416 = n11415 ^ n11413 ;
  assign n11417 = n11416 ^ x117 ;
  assign n11418 = n11238 & ~n11417 ;
  assign n11424 = n11418 ^ n11238 ;
  assign n11436 = ~n10987 & n11424 ;
  assign n11421 = n10985 ^ n10984 ;
  assign n11426 = n11418 & ~n11421 ;
  assign n11425 = ~n11421 & n11424 ;
  assign n11427 = n11426 ^ n11425 ;
  assign n11419 = n11418 ^ n11417 ;
  assign n11422 = ~n11419 & ~n11421 ;
  assign n11423 = n11422 ^ n11421 ;
  assign n11428 = n11427 ^ n11423 ;
  assign n11437 = n11436 ^ n11428 ;
  assign n11435 = n10985 & ~n11419 ;
  assign n11438 = n11437 ^ n11435 ;
  assign n11439 = n11438 ^ n11424 ;
  assign n11434 = ~n10985 & n11424 ;
  assign n11440 = n11439 ^ n11434 ;
  assign n11480 = n11440 ^ n11438 ;
  assign n11455 = ~n10986 & n11418 ;
  assign n11450 = n11424 ^ n11417 ;
  assign n11451 = n10985 & n11450 ;
  assign n11471 = n11455 ^ n11451 ;
  assign n11488 = n11480 ^ n11471 ;
  assign n11489 = n11488 ^ n10739 ;
  assign n11457 = ~n10987 & n11450 ;
  assign n11458 = n11457 ^ n11426 ;
  assign n11459 = n11458 ^ n10987 ;
  assign n11446 = n11436 ^ n11426 ;
  assign n11420 = ~n10987 & ~n11419 ;
  assign n11447 = n11446 ^ n11420 ;
  assign n11460 = n11459 ^ n11447 ;
  assign n11461 = n11460 ^ n11426 ;
  assign n11456 = n11455 ^ n11418 ;
  assign n11462 = n11461 ^ n11456 ;
  assign n11453 = n11436 ^ n11425 ;
  assign n11454 = n11453 ^ n11434 ;
  assign n11463 = n11462 ^ n11454 ;
  assign n11449 = ~n10986 & ~n11419 ;
  assign n11470 = n11463 ^ n11449 ;
  assign n11487 = n11470 ^ n11435 ;
  assign n11490 = n11489 ^ n11487 ;
  assign n13420 = n11490 ^ n11436 ;
  assign n8849 = n8848 ^ n8419 ;
  assign n9907 = n9906 ^ n9903 ;
  assign n9913 = n9912 ^ n9907 ;
  assign n9914 = ~n8419 & ~n9913 ;
  assign n9915 = n9914 ^ n9912 ;
  assign n9893 = n9892 ^ n9889 ;
  assign n9894 = n9893 ^ n9726 ;
  assign n9895 = n9894 ^ n9893 ;
  assign n9896 = n9893 ^ n9891 ;
  assign n9897 = n9896 ^ n9893 ;
  assign n9898 = n9895 & n9897 ;
  assign n9899 = n9898 ^ n9893 ;
  assign n9900 = n8419 & n9899 ;
  assign n9901 = n9900 ^ n9888 ;
  assign n9916 = n9915 ^ n9901 ;
  assign n9917 = ~n8849 & n9916 ;
  assign n9918 = n9917 ^ n9915 ;
  assign n9919 = n9918 ^ n9386 ;
  assign n9920 = n9919 ^ x124 ;
  assign n13405 = ~n9920 & n11455 ;
  assign n13421 = n13420 ^ n13405 ;
  assign n13417 = n11480 ^ n11436 ;
  assign n11452 = n11451 ^ n11449 ;
  assign n13418 = n13417 ^ n11452 ;
  assign n13419 = ~n9920 & n13418 ;
  assign n13422 = n13421 ^ n13419 ;
  assign n13423 = n10389 & n13422 ;
  assign n10390 = ~n9920 & n10389 ;
  assign n10391 = n10390 ^ n9920 ;
  assign n10392 = n10391 ^ n10389 ;
  assign n13413 = n11487 ^ n11437 ;
  assign n13414 = n10392 & ~n13413 ;
  assign n13407 = ~n10391 & n11435 ;
  assign n11465 = n11460 ^ n11422 ;
  assign n11497 = n10392 & ~n11465 ;
  assign n13408 = n13407 ^ n11497 ;
  assign n10393 = n10392 ^ n9920 ;
  assign n11429 = n11428 ^ n11420 ;
  assign n11430 = n10393 & ~n11429 ;
  assign n13403 = n11465 ^ n11430 ;
  assign n13404 = n13403 ^ n11463 ;
  assign n13406 = n13405 ^ n13404 ;
  assign n13409 = n13408 ^ n13406 ;
  assign n13410 = n13409 ^ n10243 ;
  assign n13395 = n10389 ^ n9920 ;
  assign n13396 = n11463 ^ n10389 ;
  assign n13397 = n13396 ^ n11463 ;
  assign n13400 = n11458 & n13397 ;
  assign n13401 = n13400 ^ n11463 ;
  assign n13402 = n13395 & ~n13401 ;
  assign n13411 = n13410 ^ n13402 ;
  assign n13388 = n11465 ^ n11429 ;
  assign n13389 = n13388 ^ n11465 ;
  assign n13390 = n11465 ^ n9920 ;
  assign n13391 = n13390 ^ n11465 ;
  assign n13392 = n13389 & ~n13391 ;
  assign n13393 = n13392 ^ n11465 ;
  assign n13394 = ~n10389 & n13393 ;
  assign n13412 = n13411 ^ n13394 ;
  assign n13415 = n13414 ^ n13412 ;
  assign n13386 = n11457 ^ n11425 ;
  assign n13387 = ~n9920 & n13386 ;
  assign n13416 = n13415 ^ n13387 ;
  assign n13424 = n13423 ^ n13416 ;
  assign n13425 = n13424 ^ x83 ;
  assign n12737 = ~n11103 & ~n12443 ;
  assign n12768 = n11162 & n11204 ;
  assign n12739 = n12738 ^ n11201 ;
  assign n12740 = n12739 ^ n11100 ;
  assign n12741 = n12463 ^ n11171 ;
  assign n12742 = n12741 ^ n11100 ;
  assign n12744 = n12743 ^ n11101 ;
  assign n12747 = ~n12741 & n12744 ;
  assign n12748 = n12747 ^ n11101 ;
  assign n12749 = n12742 & ~n12748 ;
  assign n12750 = n12749 ^ n11100 ;
  assign n12751 = n12453 ^ n11183 ;
  assign n12752 = n12751 ^ n11171 ;
  assign n12753 = ~n12750 & n12752 ;
  assign n12756 = ~n12740 & ~n12753 ;
  assign n12757 = n12756 ^ n11100 ;
  assign n12758 = n11189 ^ n11181 ;
  assign n12759 = n12758 ^ n11166 ;
  assign n12760 = n11100 & n12759 ;
  assign n12761 = n12760 ^ n12445 ;
  assign n12762 = n11101 & ~n12761 ;
  assign n12764 = n12762 ^ n11101 ;
  assign n12763 = n12762 ^ n12753 ;
  assign n12765 = n12764 ^ n12763 ;
  assign n12766 = ~n12757 & ~n12765 ;
  assign n12767 = n12766 ^ n12764 ;
  assign n12771 = n12768 ^ n12767 ;
  assign n12772 = n12737 & n12771 ;
  assign n12773 = n12772 ^ n9378 ;
  assign n12774 = n12773 ^ x122 ;
  assign n12495 = n12494 ^ n11369 ;
  assign n12480 = n11405 ^ n11377 ;
  assign n12481 = n12480 ^ n11557 ;
  assign n12482 = n11239 & ~n12481 ;
  assign n12483 = n12482 ^ n11558 ;
  assign n12496 = n12495 ^ n12483 ;
  assign n12497 = n12496 ^ n11388 ;
  assign n12501 = n12500 ^ n12497 ;
  assign n12502 = n12501 ^ n9623 ;
  assign n12484 = n12483 ^ n11355 ;
  assign n12485 = n12484 ^ n11356 ;
  assign n12486 = n12485 ^ n12484 ;
  assign n12487 = n12484 ^ n11264 ;
  assign n12488 = n12487 ^ n12484 ;
  assign n12489 = n12486 & ~n12488 ;
  assign n12490 = n12489 ^ n12484 ;
  assign n12491 = ~n12479 & n12490 ;
  assign n12503 = n12502 ^ n12491 ;
  assign n12736 = n12503 ^ x104 ;
  assign n12423 = n11929 ^ n11922 ;
  assign n12413 = ~n11830 & ~n11991 ;
  assign n12414 = n12413 ^ n11989 ;
  assign n12424 = n12423 ^ n12414 ;
  assign n12419 = n11903 ^ n11892 ;
  assign n12420 = n12419 ^ n11921 ;
  assign n12421 = n12420 ^ n11929 ;
  assign n12422 = n11830 & n12421 ;
  assign n12425 = n12424 ^ n12422 ;
  assign n12426 = n11829 & ~n12425 ;
  assign n12415 = n12414 ^ n12214 ;
  assign n12403 = ~n11829 & ~n11987 ;
  assign n12404 = n12403 ^ n11933 ;
  assign n12416 = n12415 ^ n12404 ;
  assign n12417 = n12416 ^ n12255 ;
  assign n12418 = n12417 ^ n11999 ;
  assign n12427 = n12426 ^ n12418 ;
  assign n12406 = n12404 ^ n11989 ;
  assign n12401 = n11930 ^ n11924 ;
  assign n12402 = n12401 ^ n11933 ;
  assign n12405 = n12404 ^ n12402 ;
  assign n12407 = n12406 ^ n12405 ;
  assign n12410 = ~n11829 & n12407 ;
  assign n12411 = n12410 ^ n12406 ;
  assign n12412 = ~n11830 & n12411 ;
  assign n12428 = n12427 ^ n12412 ;
  assign n12429 = ~n12249 & ~n12428 ;
  assign n12430 = n12429 ^ n9535 ;
  assign n12652 = n12430 ^ x82 ;
  assign n12649 = n10687 ^ n9990 ;
  assign n12641 = n10696 ^ n10679 ;
  assign n12642 = n12641 ^ n11534 ;
  assign n12632 = n10690 ^ n10586 ;
  assign n12635 = n12632 ^ n10694 ;
  assign n12631 = n10699 ^ n10594 ;
  assign n12633 = n12632 ^ n12631 ;
  assign n12634 = ~n10669 & n12633 ;
  assign n12636 = n12635 ^ n12634 ;
  assign n12181 = n10713 ^ n10685 ;
  assign n12639 = n12636 ^ n12181 ;
  assign n12640 = n12639 ^ n12636 ;
  assign n12643 = n12642 ^ n12640 ;
  assign n12644 = n10669 & n12643 ;
  assign n12645 = n12644 ^ n12639 ;
  assign n12646 = n11506 & ~n12645 ;
  assign n12637 = n12636 ^ n11518 ;
  assign n12192 = n11541 ^ n10699 ;
  assign n12193 = n12192 ^ n10590 ;
  assign n12194 = n12193 ^ n10699 ;
  assign n12195 = n10699 ^ n10669 ;
  assign n12196 = n12195 ^ n10699 ;
  assign n12197 = n12194 & n12196 ;
  assign n12198 = n12197 ^ n10699 ;
  assign n12199 = n10633 & ~n12198 ;
  assign n12638 = n12637 ^ n12199 ;
  assign n12647 = n12646 ^ n12638 ;
  assign n12648 = ~n11512 & n12647 ;
  assign n12650 = n12649 ^ n12648 ;
  assign n12651 = n12650 ^ x72 ;
  assign n12677 = ~n10793 & ~n10920 ;
  assign n12669 = n10938 ^ n10903 ;
  assign n12670 = n12669 ^ n10794 ;
  assign n12671 = n12670 ^ n10903 ;
  assign n12672 = n10903 ^ n10793 ;
  assign n12673 = n12672 ^ n10903 ;
  assign n12674 = n12671 & n12673 ;
  assign n12675 = n12674 ^ n10903 ;
  assign n12676 = n12668 & ~n12675 ;
  assign n12678 = n12677 ^ n12676 ;
  assign n12679 = n10948 & ~n12678 ;
  assign n12680 = n12679 ^ n12677 ;
  assign n12665 = n10905 ^ n10890 ;
  assign n12666 = n12665 ^ n10900 ;
  assign n12667 = n10915 & ~n12666 ;
  assign n12681 = n12680 ^ n12667 ;
  assign n12682 = ~n12664 & ~n12681 ;
  assign n12683 = n10948 ^ n10897 ;
  assign n12688 = n10941 ^ n10933 ;
  assign n12685 = n10973 ^ n10940 ;
  assign n12684 = n10920 ^ n10902 ;
  assign n12686 = n12685 ^ n12684 ;
  assign n12689 = n12688 ^ n12686 ;
  assign n12690 = ~n10907 & ~n12689 ;
  assign n12687 = n12686 ^ n10897 ;
  assign n12691 = n12690 ^ n12687 ;
  assign n12692 = ~n12683 & ~n12691 ;
  assign n12693 = n12692 ^ n10897 ;
  assign n12694 = n12682 & ~n12693 ;
  assign n12695 = n12694 ^ n9302 ;
  assign n12696 = n12695 ^ x99 ;
  assign n12777 = ~n12651 & ~n12696 ;
  assign n12711 = n10250 ^ n9921 ;
  assign n12712 = n10311 ^ n10250 ;
  assign n12713 = n10341 ^ n10311 ;
  assign n12714 = ~n12712 & ~n12713 ;
  assign n12715 = n12714 ^ n10311 ;
  assign n12716 = n12711 & n12715 ;
  assign n12709 = n10371 & ~n10382 ;
  assign n12701 = n10261 ^ n10256 ;
  assign n12702 = n12701 ^ n10374 ;
  assign n12699 = n10339 ^ n10254 ;
  assign n12700 = ~n9921 & n12699 ;
  assign n12703 = n12702 ^ n12700 ;
  assign n12705 = n12701 ^ n9921 ;
  assign n12704 = n12701 ^ n10311 ;
  assign n12706 = n12705 ^ n12704 ;
  assign n12707 = ~n12703 & ~n12706 ;
  assign n12708 = n12707 ^ n12704 ;
  assign n12710 = n12709 ^ n12708 ;
  assign n12717 = n12716 ^ n12710 ;
  assign n12718 = n12717 ^ n10324 ;
  assign n12697 = n12392 ^ n10324 ;
  assign n12698 = n11629 & n12697 ;
  assign n12719 = n12718 ^ n12698 ;
  assign n12720 = n10344 ^ n10325 ;
  assign n12721 = ~n9921 & ~n12720 ;
  assign n12722 = n12721 ^ n10325 ;
  assign n12723 = n12722 ^ n10311 ;
  assign n12724 = n12723 ^ n12722 ;
  assign n12725 = ~n9921 & n10330 ;
  assign n12726 = n12725 ^ n12722 ;
  assign n12727 = ~n12724 & n12726 ;
  assign n12728 = n12727 ^ n12722 ;
  assign n12729 = n12719 & ~n12728 ;
  assign n12730 = n12729 ^ n9953 ;
  assign n12731 = n12730 ^ x81 ;
  assign n12778 = n12777 ^ n12731 ;
  assign n12732 = n12696 & ~n12731 ;
  assign n12775 = n12732 ^ n12696 ;
  assign n12776 = n12775 ^ n12651 ;
  assign n12779 = n12778 ^ n12776 ;
  assign n12780 = ~n12652 & n12779 ;
  assign n13443 = n12780 ^ n12732 ;
  assign n12786 = n12731 ^ n12652 ;
  assign n12787 = n12786 ^ n12696 ;
  assign n12793 = n12732 & ~n12787 ;
  assign n13444 = n13443 ^ n12793 ;
  assign n12782 = n12696 ^ n12651 ;
  assign n13445 = n13444 ^ n12782 ;
  assign n12783 = n12731 ^ n12651 ;
  assign n12792 = n12786 ^ n12651 ;
  assign n12794 = n12787 ^ n12731 ;
  assign n12795 = n12794 ^ n12793 ;
  assign n12796 = ~n12792 & ~n12795 ;
  assign n12791 = n12775 ^ n12731 ;
  assign n12797 = n12796 ^ n12791 ;
  assign n12798 = n12797 ^ n12794 ;
  assign n12799 = n12798 ^ n12786 ;
  assign n12788 = ~n12731 & ~n12787 ;
  assign n12789 = n12788 ^ n12787 ;
  assign n12653 = n12651 & n12652 ;
  assign n12733 = n12653 & ~n12732 ;
  assign n12790 = n12789 ^ n12733 ;
  assign n12800 = n12799 ^ n12790 ;
  assign n12801 = n12800 ^ n12651 ;
  assign n12804 = n12783 & n12801 ;
  assign n12805 = n12804 ^ n12652 ;
  assign n12806 = n12782 & n12805 ;
  assign n12807 = n12806 ^ n12801 ;
  assign n13440 = n12807 ^ n12733 ;
  assign n13441 = n13440 ^ n12652 ;
  assign n13427 = ~n12652 & ~n12783 ;
  assign n13442 = n13441 ^ n13427 ;
  assign n13446 = n13445 ^ n13442 ;
  assign n13447 = n12736 & n13446 ;
  assign n13448 = n13447 ^ n13445 ;
  assign n13428 = n13427 ^ n12786 ;
  assign n12781 = n12780 ^ n12778 ;
  assign n13429 = n13428 ^ n12781 ;
  assign n13426 = n12782 ^ n12731 ;
  assign n13430 = n13429 ^ n13426 ;
  assign n13431 = n13430 ^ n12787 ;
  assign n13432 = n13431 ^ n12652 ;
  assign n13433 = n13432 ^ n12788 ;
  assign n13434 = n13433 ^ n13430 ;
  assign n13435 = ~n12651 & ~n13434 ;
  assign n13436 = n13435 ^ n13431 ;
  assign n13437 = ~n12736 & n13436 ;
  assign n13438 = n13437 ^ n13430 ;
  assign n13449 = n13448 ^ n13438 ;
  assign n13450 = ~n12774 & n13449 ;
  assign n13439 = n13438 ^ n12774 ;
  assign n13451 = n13450 ^ n13439 ;
  assign n13452 = n13451 ^ n10029 ;
  assign n13453 = n13452 ^ x70 ;
  assign n13454 = ~n13425 & n13453 ;
  assign n13455 = n13454 ^ n13453 ;
  assign n13457 = n13455 ^ n13425 ;
  assign n13468 = n13457 ^ n13453 ;
  assign n13469 = ~n13460 & ~n13468 ;
  assign n13467 = n13454 & ~n13460 ;
  assign n13470 = n13469 ^ n13467 ;
  assign n13463 = ~n13350 & n13455 ;
  assign n13464 = n13383 & n13463 ;
  assign n13465 = n13464 ^ n13463 ;
  assign n15477 = n13470 ^ n13465 ;
  assign n15478 = n15477 ^ n13460 ;
  assign n15479 = n15478 ^ n13465 ;
  assign n12400 = n12399 ^ x113 ;
  assign n12431 = n12430 ^ x74 ;
  assign n12578 = ~n12400 & ~n12431 ;
  assign n12579 = n12578 ^ n12431 ;
  assign n12469 = n12468 ^ x80 ;
  assign n12473 = n11602 ^ n9585 ;
  assign n12470 = n11605 ^ n11595 ;
  assign n12471 = n12470 ^ n11602 ;
  assign n12472 = ~n8848 & ~n12471 ;
  assign n12474 = n12473 ^ n12472 ;
  assign n12475 = n12474 ^ x107 ;
  assign n12476 = n12469 & n12475 ;
  assign n12477 = n12476 ^ n12469 ;
  assign n12504 = n12503 ^ x89 ;
  assign n12520 = n11793 ^ n11764 ;
  assign n12523 = n11782 ^ n11664 ;
  assign n12524 = ~n11665 & ~n12523 ;
  assign n12525 = n12524 ^ n11664 ;
  assign n12526 = n11739 & ~n12525 ;
  assign n12521 = n11782 ^ n11766 ;
  assign n12527 = n12526 ^ n12521 ;
  assign n12530 = ~n12520 & ~n12527 ;
  assign n12531 = n12530 ^ n11793 ;
  assign n12507 = n11779 ^ n11756 ;
  assign n12534 = n12507 ^ n11663 ;
  assign n12532 = n12507 ^ n11794 ;
  assign n12533 = n12532 ^ n12527 ;
  assign n12535 = n12534 ^ n12533 ;
  assign n12536 = n12531 & n12535 ;
  assign n12537 = n12536 ^ n12534 ;
  assign n12538 = n12537 ^ n12161 ;
  assign n12508 = n11754 ^ n11746 ;
  assign n12509 = n12508 ^ n11785 ;
  assign n12510 = ~n11663 & n12509 ;
  assign n12511 = n12510 ^ n11746 ;
  assign n12539 = n12538 ^ n12511 ;
  assign n12513 = n12511 ^ n12140 ;
  assign n12512 = n12511 ^ n12507 ;
  assign n12514 = n12513 ^ n12512 ;
  assign n12517 = ~n11663 & n12514 ;
  assign n12518 = n12517 ^ n12513 ;
  assign n12519 = n11664 & n12518 ;
  assign n12540 = n12539 ^ n12519 ;
  assign n12541 = ~n12151 & n12540 ;
  assign n12505 = n11795 ^ n9567 ;
  assign n12506 = n12505 ^ n12143 ;
  assign n12542 = n12541 ^ n12506 ;
  assign n12543 = n12542 ^ x106 ;
  assign n12544 = ~n12504 & n12543 ;
  assign n12549 = n12544 ^ n12543 ;
  assign n12550 = n12549 ^ n12504 ;
  assign n12581 = n12477 & n12550 ;
  assign n12562 = n12476 & n12544 ;
  assign n12595 = n12581 ^ n12562 ;
  assign n12478 = n12477 ^ n12475 ;
  assign n12551 = ~n12478 & n12550 ;
  assign n12548 = ~n12478 & n12544 ;
  assign n12552 = n12551 ^ n12548 ;
  assign n12593 = n12581 ^ n12552 ;
  assign n12590 = n12543 ^ n12504 ;
  assign n12591 = ~n12475 & ~n12590 ;
  assign n12592 = n12591 ^ n12475 ;
  assign n12594 = n12593 ^ n12592 ;
  assign n12596 = n12595 ^ n12594 ;
  assign n12589 = n12477 & n12549 ;
  assign n12597 = n12596 ^ n12589 ;
  assign n13136 = n12597 ^ n12469 ;
  assign n13137 = ~n12579 & ~n13136 ;
  assign n12587 = n12579 ^ n12400 ;
  assign n12611 = n12591 ^ n12504 ;
  assign n12612 = ~n12469 & n12611 ;
  assign n13134 = ~n12587 & n12612 ;
  assign n12554 = n12476 & n12550 ;
  assign n12563 = n12562 ^ n12554 ;
  assign n12560 = n12476 & n12549 ;
  assign n12561 = n12560 ^ n12476 ;
  assign n12564 = n12563 ^ n12561 ;
  assign n12545 = n12544 ^ n12504 ;
  assign n12546 = ~n12478 & ~n12545 ;
  assign n12547 = n12546 ^ n12478 ;
  assign n12553 = n12552 ^ n12547 ;
  assign n12580 = n12564 ^ n12553 ;
  assign n12582 = n12581 ^ n12580 ;
  assign n12583 = ~n12578 & n12582 ;
  assign n13126 = n12583 ^ n12560 ;
  assign n13131 = n12578 & n12597 ;
  assign n13132 = n13131 ^ n12400 ;
  assign n13133 = ~n13126 & ~n13132 ;
  assign n13135 = n13134 ^ n13133 ;
  assign n13138 = n13137 ^ n13135 ;
  assign n13124 = n12589 ^ n12563 ;
  assign n13125 = ~n12587 & n13124 ;
  assign n13139 = n13138 ^ n13125 ;
  assign n13140 = n13139 ^ n12546 ;
  assign n12588 = n12562 ^ n12477 ;
  assign n12598 = n12597 ^ n12588 ;
  assign n12599 = n12598 ^ n12545 ;
  assign n12556 = n12476 ^ n12475 ;
  assign n12557 = n12549 & n12556 ;
  assign n12558 = n12557 ^ n12548 ;
  assign n12559 = n12558 ^ n12546 ;
  assign n12565 = n12564 ^ n12559 ;
  assign n12566 = n12565 ^ n12558 ;
  assign n12600 = n12599 ^ n12566 ;
  assign n13119 = n12546 ^ n12400 ;
  assign n13120 = n13119 ^ n12546 ;
  assign n13121 = n12600 & ~n13120 ;
  assign n13122 = n13121 ^ n12546 ;
  assign n13123 = n12431 & n13122 ;
  assign n13141 = n13140 ^ n13123 ;
  assign n13142 = n13141 ^ n12552 ;
  assign n12432 = n12431 ^ n12400 ;
  assign n12610 = n12600 ^ n12557 ;
  assign n13111 = n12610 ^ n12594 ;
  assign n13112 = ~n12431 & ~n13111 ;
  assign n13113 = n13112 ^ n12594 ;
  assign n12613 = n12612 ^ n12559 ;
  assign n12614 = n12613 ^ n12552 ;
  assign n12615 = n12614 ^ n12556 ;
  assign n12616 = n12615 ^ n12610 ;
  assign n13114 = n13113 ^ n12616 ;
  assign n13115 = ~n12432 & ~n13114 ;
  assign n13116 = n13115 ^ n12616 ;
  assign n13143 = n13142 ^ n13116 ;
  assign n13144 = n13143 ^ n9725 ;
  assign n13106 = n12552 ^ n12400 ;
  assign n13107 = n13106 ^ n12552 ;
  assign n13108 = n12614 & ~n13107 ;
  assign n13109 = n13108 ^ n12552 ;
  assign n13110 = ~n12432 & n13109 ;
  assign n13145 = n13144 ^ n13110 ;
  assign n13146 = n13145 ^ x118 ;
  assign n15480 = n13465 ^ n13146 ;
  assign n15481 = n15480 ^ n13465 ;
  assign n15482 = ~n15479 & ~n15481 ;
  assign n15483 = n15482 ^ n13465 ;
  assign n15484 = ~n13310 & n15483 ;
  assign n13461 = n13460 ^ n13350 ;
  assign n13462 = n13457 & n13461 ;
  assign n15270 = n13310 ^ n13146 ;
  assign n15271 = n13462 & n15270 ;
  assign n15981 = n13470 ^ n13462 ;
  assign n13484 = n13385 & n13454 ;
  assign n13481 = n13469 ^ n13464 ;
  assign n13479 = n13384 & ~n13468 ;
  assign n13482 = n13481 ^ n13479 ;
  assign n13485 = n13484 ^ n13482 ;
  assign n13458 = n13384 & n13457 ;
  assign n13473 = n13458 ^ n13457 ;
  assign n13466 = n13465 ^ n13460 ;
  assign n13471 = n13470 ^ n13466 ;
  assign n13472 = n13471 ^ n13462 ;
  assign n13474 = n13473 ^ n13472 ;
  assign n13486 = n13485 ^ n13474 ;
  assign n13456 = n13385 & n13455 ;
  assign n13487 = n13486 ^ n13456 ;
  assign n13483 = n13482 ^ n13385 ;
  assign n13488 = n13487 ^ n13483 ;
  assign n13489 = n13488 ^ n13484 ;
  assign n13477 = n13350 & n13425 ;
  assign n13459 = n13458 ^ n13456 ;
  assign n13475 = n13474 ^ n13459 ;
  assign n13478 = n13477 ^ n13475 ;
  assign n13480 = n13479 ^ n13478 ;
  assign n13490 = n13489 ^ n13480 ;
  assign n13476 = n13475 ^ n13350 ;
  assign n13491 = n13490 ^ n13476 ;
  assign n15469 = n13491 ^ n13475 ;
  assign n15982 = n15981 ^ n15469 ;
  assign n13492 = n13491 ^ n13488 ;
  assign n13493 = n13492 ^ n13484 ;
  assign n13498 = n13493 ^ n13467 ;
  assign n13499 = n13498 ^ n13454 ;
  assign n13500 = n13499 ^ n13488 ;
  assign n13509 = n13500 ^ n13456 ;
  assign n15985 = n15982 ^ n13509 ;
  assign n15455 = n13467 ^ n13464 ;
  assign n13532 = n13500 ^ n13470 ;
  assign n13533 = n13532 ^ n13488 ;
  assign n13531 = n13492 ^ n13479 ;
  assign n13534 = n13533 ^ n13531 ;
  assign n13530 = n13489 ^ n13425 ;
  assign n13535 = n13534 ^ n13530 ;
  assign n15980 = n15455 ^ n13535 ;
  assign n15983 = n15982 ^ n15980 ;
  assign n15984 = ~n13310 & n15983 ;
  assign n15986 = n15985 ^ n15984 ;
  assign n15987 = ~n15270 & ~n15986 ;
  assign n15988 = n15987 ^ n13509 ;
  assign n13311 = n13146 & n13310 ;
  assign n13312 = n13311 ^ n13310 ;
  assign n13507 = n13312 ^ n13146 ;
  assign n13539 = n13507 ^ n13310 ;
  assign n15979 = n13490 & n13539 ;
  assign n15989 = n15988 ^ n15979 ;
  assign n15972 = n13492 ^ n13478 ;
  assign n15971 = n13485 ^ n13465 ;
  assign n15973 = n15972 ^ n15971 ;
  assign n15974 = n15972 ^ n13310 ;
  assign n15975 = n15974 ^ n15972 ;
  assign n15976 = ~n15973 & n15975 ;
  assign n15977 = n15976 ^ n15972 ;
  assign n15978 = ~n13146 & ~n15977 ;
  assign n15990 = n15989 ^ n15978 ;
  assign n15991 = ~n15271 & n15990 ;
  assign n15992 = ~n15484 & n15991 ;
  assign n15286 = n13535 ^ n13474 ;
  assign n15287 = n13310 & ~n15286 ;
  assign n15288 = n15287 ^ n13474 ;
  assign n15297 = n15270 & ~n15288 ;
  assign n15969 = n15297 ^ n15288 ;
  assign n15970 = n15969 ^ n12730 ;
  assign n15993 = n15992 ^ n15970 ;
  assign n15994 = n15993 ^ x114 ;
  assign n13935 = n12927 & n12950 ;
  assign n13936 = n13935 ^ n12969 ;
  assign n12956 = ~n12953 & ~n12955 ;
  assign n12908 = n12830 & n12907 ;
  assign n12909 = n12908 ^ n12906 ;
  assign n12910 = n12909 ^ n12829 ;
  assign n12911 = n12910 ^ n12909 ;
  assign n12946 = ~n12911 & n12943 ;
  assign n12947 = n12946 ^ n12909 ;
  assign n12948 = ~n12831 & n12947 ;
  assign n12949 = n12948 ^ n12909 ;
  assign n12957 = n12956 ^ n12949 ;
  assign n13954 = n12951 & n12998 ;
  assign n12975 = n12941 ^ n12917 ;
  assign n13944 = n12975 ^ n12943 ;
  assign n13945 = n13944 ^ n12921 ;
  assign n13948 = n13945 ^ n12919 ;
  assign n13000 = n12999 ^ n12916 ;
  assign n13943 = n13000 ^ n12927 ;
  assign n13946 = n13945 ^ n13943 ;
  assign n13947 = n12830 & n13946 ;
  assign n13949 = n13948 ^ n13947 ;
  assign n13950 = n12831 & n13949 ;
  assign n13941 = n13366 ^ n12919 ;
  assign n13942 = n13941 ^ n12986 ;
  assign n13951 = n13950 ^ n13942 ;
  assign n13938 = n12955 ^ n12904 ;
  assign n13939 = n13938 ^ n12925 ;
  assign n13940 = n12951 & ~n13939 ;
  assign n13952 = n13951 ^ n13940 ;
  assign n13937 = n12933 & ~n12953 ;
  assign n13953 = n13952 ^ n13937 ;
  assign n13955 = n13954 ^ n13953 ;
  assign n13956 = n12916 ^ n12913 ;
  assign n13957 = n12916 ^ n12830 ;
  assign n13958 = n13957 ^ n12916 ;
  assign n13959 = n13956 & n13958 ;
  assign n13960 = n13959 ^ n12916 ;
  assign n13961 = ~n12829 & n13960 ;
  assign n13962 = ~n13955 & ~n13961 ;
  assign n13963 = ~n12957 & n13962 ;
  assign n13964 = ~n13354 & n13963 ;
  assign n13965 = ~n13936 & n13964 ;
  assign n13966 = ~n12970 & n13965 ;
  assign n13967 = n13966 ^ n9229 ;
  assign n13968 = n13967 ^ x123 ;
  assign n13655 = n10738 ^ x85 ;
  assign n13656 = n12695 ^ x67 ;
  assign n13657 = ~n13655 & ~n13656 ;
  assign n13648 = n9919 ^ x86 ;
  assign n13587 = n12140 ^ n11766 ;
  assign n13613 = n13587 ^ n11749 ;
  assign n13585 = n11779 ^ n11764 ;
  assign n13586 = n13585 ^ n11769 ;
  assign n13588 = n13587 ^ n13586 ;
  assign n13589 = n11663 & ~n13588 ;
  assign n13590 = n13589 ^ n13585 ;
  assign n13599 = n13590 ^ n12153 ;
  assign n13600 = n13599 ^ n11813 ;
  assign n13591 = n13590 ^ n11777 ;
  assign n13592 = n13591 ^ n11754 ;
  assign n13593 = n13592 ^ n13590 ;
  assign n13596 = n11663 & n13593 ;
  assign n13597 = n13596 ^ n13590 ;
  assign n13598 = n11665 & n13597 ;
  assign n13601 = n13600 ^ n13598 ;
  assign n13614 = n11793 & ~n13601 ;
  assign n13615 = n13613 & n13614 ;
  assign n13611 = n12144 ^ n9343 ;
  assign n13612 = n13611 ^ n13601 ;
  assign n13616 = n13615 ^ n13612 ;
  assign n13606 = n11745 ^ n11663 ;
  assign n13607 = n13606 ^ n11745 ;
  assign n13608 = n11777 & n13607 ;
  assign n13609 = n13608 ^ n11745 ;
  assign n13610 = n11664 & n13609 ;
  assign n13617 = n13616 ^ n13610 ;
  assign n13579 = n12155 ^ n11772 ;
  assign n13580 = n13579 ^ n11740 ;
  assign n13581 = n11740 ^ n11664 ;
  assign n13582 = n13581 ^ n11740 ;
  assign n13583 = ~n13580 & ~n13582 ;
  assign n13584 = n13583 ^ n11740 ;
  assign n13602 = ~n11663 & ~n13601 ;
  assign n13603 = n13584 & n13602 ;
  assign n13618 = n13617 ^ n13603 ;
  assign n13619 = n13618 ^ x68 ;
  assign n13644 = ~n11829 & ~n12414 ;
  assign n13636 = n11973 ^ n11909 ;
  assign n13633 = n11989 ^ n11905 ;
  assign n13634 = n11907 & ~n13633 ;
  assign n13631 = n11921 ^ n11892 ;
  assign n13632 = n11829 & n13631 ;
  assign n13635 = n13634 ^ n13632 ;
  assign n13637 = n13636 ^ n13635 ;
  assign n13638 = n13637 ^ n11964 ;
  assign n13639 = n13638 ^ n11999 ;
  assign n13640 = n13639 ^ n12249 ;
  assign n13641 = n13640 ^ n9430 ;
  assign n13624 = n11935 ^ n11909 ;
  assign n13625 = n11908 ^ n11889 ;
  assign n13628 = ~n11935 & ~n13625 ;
  assign n13629 = n13628 ^ n11908 ;
  assign n13630 = ~n13624 & n13629 ;
  assign n13642 = n13641 ^ n13630 ;
  assign n13620 = n12402 ^ n11934 ;
  assign n13621 = n12219 & n13620 ;
  assign n13622 = n13621 ^ n11934 ;
  assign n13623 = n11952 & ~n13622 ;
  assign n13643 = n13642 ^ n13623 ;
  assign n13645 = n13644 ^ n13643 ;
  assign n13646 = n13645 ^ x116 ;
  assign n13673 = n13619 & n13646 ;
  assign n13676 = n13673 ^ n13619 ;
  assign n13677 = n13648 & n13676 ;
  assign n13662 = ~n13619 & n13648 ;
  assign n13675 = n13662 ^ n13648 ;
  assign n13678 = n13677 ^ n13675 ;
  assign n13682 = n13678 ^ n13673 ;
  assign n13647 = n12773 ^ x109 ;
  assign n13649 = ~n13647 & n13648 ;
  assign n13650 = n13649 ^ n13647 ;
  assign n13651 = n13650 ^ n13648 ;
  assign n13652 = n13646 & n13651 ;
  assign n13653 = ~n13619 & n13652 ;
  assign n13654 = n13653 ^ n13652 ;
  assign n13683 = n13682 ^ n13654 ;
  assign n13667 = ~n13619 & ~n13650 ;
  assign n13681 = n13667 ^ n13650 ;
  assign n13684 = n13683 ^ n13681 ;
  assign n13898 = n13657 & ~n13684 ;
  assign n13658 = n13657 ^ n13656 ;
  assign n13668 = n13646 & n13667 ;
  assign n13669 = n13668 ^ n13667 ;
  assign n13670 = ~n13658 & n13669 ;
  assign n13899 = n13898 ^ n13670 ;
  assign n13659 = n13658 ^ n13655 ;
  assign n13722 = n13683 ^ n13668 ;
  assign n13674 = n13649 & n13673 ;
  assign n13928 = n13722 ^ n13674 ;
  assign n13698 = n13652 ^ n13651 ;
  assign n13680 = n13677 ^ n13676 ;
  assign n13685 = n13684 ^ n13680 ;
  assign n13699 = n13698 ^ n13685 ;
  assign n13663 = n13647 & n13662 ;
  assign n13693 = ~n13646 & n13663 ;
  assign n13700 = n13699 ^ n13693 ;
  assign n13679 = n13678 ^ n13674 ;
  assign n13686 = n13685 ^ n13679 ;
  assign n13701 = n13700 ^ n13686 ;
  assign n13694 = n13693 ^ n13663 ;
  assign n13695 = n13694 ^ n13652 ;
  assign n13697 = n13695 ^ n13647 ;
  assign n13702 = n13701 ^ n13697 ;
  assign n13717 = n13702 ^ n13677 ;
  assign n13925 = n13717 ^ n13683 ;
  assign n13926 = n13925 ^ n13646 ;
  assign n13664 = n13663 ^ n13662 ;
  assign n13665 = n13646 & n13664 ;
  assign n13706 = n13665 ^ n13664 ;
  assign n13707 = n13706 ^ n13684 ;
  assign n13708 = n13707 ^ n13683 ;
  assign n13709 = n13708 ^ n13669 ;
  assign n13703 = n13702 ^ n13694 ;
  assign n13704 = n13703 ^ n13699 ;
  assign n13705 = n13704 ^ n13653 ;
  assign n13710 = n13709 ^ n13705 ;
  assign n13927 = n13926 ^ n13710 ;
  assign n13929 = n13928 ^ n13927 ;
  assign n13930 = ~n13659 & ~n13929 ;
  assign n13915 = n13658 ^ n13652 ;
  assign n13916 = n13915 ^ n13702 ;
  assign n13917 = n13683 ^ n13658 ;
  assign n13739 = n13684 ^ n13674 ;
  assign n13740 = n13739 ^ n13665 ;
  assign n13918 = n13917 ^ n13740 ;
  assign n13919 = ~n13916 & n13918 ;
  assign n13660 = n13659 ^ n13656 ;
  assign n13911 = n13702 ^ n13693 ;
  assign n13912 = n13911 ^ n13653 ;
  assign n13913 = ~n13660 & n13912 ;
  assign n13732 = n13706 ^ n13699 ;
  assign n13733 = n13699 ^ n13655 ;
  assign n13734 = n13733 ^ n13699 ;
  assign n13735 = ~n13732 & n13734 ;
  assign n13736 = n13735 ^ n13699 ;
  assign n13737 = n13656 & ~n13736 ;
  assign n13910 = n13737 ^ n13658 ;
  assign n13914 = n13913 ^ n13910 ;
  assign n13920 = n13919 ^ n13914 ;
  assign n13901 = n13699 ^ n13679 ;
  assign n13902 = n13901 ^ n13694 ;
  assign n13718 = n13717 ^ n13668 ;
  assign n13719 = n13718 ^ n13654 ;
  assign n13720 = n13719 ^ n13669 ;
  assign n13903 = n13902 ^ n13720 ;
  assign n13900 = n13708 ^ n13679 ;
  assign n13904 = n13903 ^ n13900 ;
  assign n13905 = n13900 ^ n13656 ;
  assign n13906 = n13905 ^ n13900 ;
  assign n13907 = n13904 & ~n13906 ;
  assign n13908 = n13907 ^ n13900 ;
  assign n13909 = ~n13655 & ~n13908 ;
  assign n13924 = n13920 ^ n13909 ;
  assign n13931 = n13930 ^ n13924 ;
  assign n13932 = ~n13899 & n13931 ;
  assign n13933 = n13932 ^ n10792 ;
  assign n13934 = n13933 ^ x97 ;
  assign n14094 = n13968 ^ n13934 ;
  assign n14028 = n11471 ^ n11435 ;
  assign n14029 = n14028 ^ n11490 ;
  assign n14030 = n10393 & n14029 ;
  assign n14016 = n11452 ^ n11434 ;
  assign n14019 = n14016 ^ n11461 ;
  assign n14020 = n14019 ^ n11463 ;
  assign n14021 = n14020 ^ n11490 ;
  assign n14022 = n14021 ^ n14016 ;
  assign n14023 = ~n10389 & n14022 ;
  assign n14024 = n14023 ^ n14019 ;
  assign n14025 = n9920 & ~n14024 ;
  assign n14026 = n14025 ^ n11420 ;
  assign n14017 = n14016 ^ n11420 ;
  assign n14018 = ~n10390 & n14017 ;
  assign n14027 = n14026 ^ n14018 ;
  assign n14031 = n14030 ^ n14027 ;
  assign n11464 = n11463 ^ n11452 ;
  assign n14009 = n13386 ^ n11464 ;
  assign n14010 = n14009 ^ n13386 ;
  assign n14011 = n13386 ^ n10389 ;
  assign n14012 = n14011 ^ n13386 ;
  assign n14013 = ~n14010 & n14012 ;
  assign n14014 = n14013 ^ n13386 ;
  assign n14015 = n13395 & n14014 ;
  assign n14032 = n14031 ^ n14015 ;
  assign n14008 = ~n10391 & n11458 ;
  assign n14033 = n14032 ^ n14008 ;
  assign n11431 = n10393 ^ n10391 ;
  assign n11481 = n11480 ^ n11422 ;
  assign n11482 = n11422 ^ n10389 ;
  assign n11483 = n11482 ^ n11422 ;
  assign n11484 = n11481 & ~n11483 ;
  assign n11485 = n11484 ^ n11422 ;
  assign n11486 = n11431 & n11485 ;
  assign n14034 = n14033 ^ n11486 ;
  assign n14035 = n14034 ^ n13408 ;
  assign n14036 = n14035 ^ n11430 ;
  assign n14037 = n14036 ^ n10851 ;
  assign n14038 = n14037 ^ x90 ;
  assign n12169 = n12168 ^ x101 ;
  assign n12170 = n10983 ^ x110 ;
  assign n12171 = ~n12169 & n12170 ;
  assign n12172 = n12171 ^ n12170 ;
  assign n12173 = n12172 ^ n12169 ;
  assign n12206 = n10690 ^ n10674 ;
  assign n12207 = n12206 ^ n10598 ;
  assign n12208 = ~n10669 & ~n12207 ;
  assign n12200 = n10679 ^ n10673 ;
  assign n12209 = n12208 ^ n12200 ;
  assign n12210 = n11506 & n12209 ;
  assign n12201 = n12200 ^ n11543 ;
  assign n12202 = n12201 ^ n12199 ;
  assign n12203 = n12202 ^ n11505 ;
  assign n12204 = n12203 ^ n7658 ;
  assign n12183 = n10676 ^ n10592 ;
  assign n12184 = n12183 ^ n10701 ;
  assign n12185 = n12184 ^ n11543 ;
  assign n12182 = n12181 ^ n10699 ;
  assign n12186 = n12185 ^ n12182 ;
  assign n12187 = n12185 ^ n10669 ;
  assign n12188 = n12187 ^ n12185 ;
  assign n12189 = ~n12186 & n12188 ;
  assign n12190 = n12189 ^ n12185 ;
  assign n12191 = ~n10633 & n12190 ;
  assign n12205 = n12204 ^ n12191 ;
  assign n12211 = n12210 ^ n12205 ;
  assign n12212 = n12211 ^ x77 ;
  assign n12266 = n12265 ^ x92 ;
  assign n12267 = ~n12212 & n12266 ;
  assign n12174 = n10388 ^ x70 ;
  assign n12175 = n9901 ^ n8848 ;
  assign n12176 = n12175 ^ n9917 ;
  assign n12177 = n12176 ^ n7338 ;
  assign n12178 = n12177 ^ x83 ;
  assign n12179 = n12174 & n12178 ;
  assign n12180 = n12179 ^ n12174 ;
  assign n12283 = n12180 ^ n12178 ;
  assign n12303 = n12267 & ~n12283 ;
  assign n12270 = n12267 ^ n12212 ;
  assign n12279 = n12179 ^ n12178 ;
  assign n12285 = ~n12270 & n12279 ;
  assign n12319 = n12303 ^ n12285 ;
  assign n12347 = n12319 ^ n12174 ;
  assign n12292 = n12266 ^ n12212 ;
  assign n12298 = n12292 ^ n12174 ;
  assign n12287 = n12212 ^ n12178 ;
  assign n12294 = n12266 ^ n12174 ;
  assign n12295 = n12178 & n12294 ;
  assign n12296 = n12295 ^ n12174 ;
  assign n12297 = n12287 & n12296 ;
  assign n12299 = n12298 ^ n12297 ;
  assign n12288 = ~n12174 & n12287 ;
  assign n12293 = n12292 ^ n12288 ;
  assign n12300 = n12299 ^ n12293 ;
  assign n12290 = n12287 ^ n12174 ;
  assign n12275 = n12179 & ~n12270 ;
  assign n12291 = n12290 ^ n12275 ;
  assign n12301 = n12300 ^ n12291 ;
  assign n12268 = n12267 ^ n12266 ;
  assign n12280 = n12268 ^ n12212 ;
  assign n12281 = n12279 & n12280 ;
  assign n12302 = n12301 ^ n12281 ;
  assign n12304 = n12303 ^ n12302 ;
  assign n12305 = n12304 ^ n12283 ;
  assign n12348 = n12347 ^ n12305 ;
  assign n12286 = n12285 ^ n12281 ;
  assign n12289 = n12288 ^ n12286 ;
  assign n12306 = n12305 ^ n12289 ;
  assign n12307 = n12306 ^ n12302 ;
  assign n12284 = n12268 & ~n12283 ;
  assign n12308 = n12307 ^ n12284 ;
  assign n12309 = n12308 ^ n12305 ;
  assign n12349 = n12348 ^ n12309 ;
  assign n12350 = n12173 & n12349 ;
  assign n12336 = n12299 ^ n12174 ;
  assign n12310 = n12309 ^ n12303 ;
  assign n12274 = n12179 & n12268 ;
  assign n12276 = n12275 ^ n12274 ;
  assign n12272 = n12179 & n12267 ;
  assign n12273 = n12272 ^ n12179 ;
  assign n12277 = n12276 ^ n12273 ;
  assign n12269 = n12180 & n12268 ;
  assign n12278 = n12277 ^ n12269 ;
  assign n12282 = n12281 ^ n12278 ;
  assign n12311 = n12310 ^ n12282 ;
  assign n12337 = n12336 ^ n12311 ;
  assign n14039 = n12173 & n12337 ;
  assign n14040 = ~n12350 & ~n14039 ;
  assign n12312 = n12296 ^ n12284 ;
  assign n12313 = n12312 ^ n12311 ;
  assign n12271 = n12270 ^ n12269 ;
  assign n12314 = n12313 ^ n12271 ;
  assign n12338 = n12337 ^ n12314 ;
  assign n12335 = n12269 ^ n12180 ;
  assign n12339 = n12338 ^ n12335 ;
  assign n12340 = n12339 ^ n12304 ;
  assign n12341 = n12304 ^ n12170 ;
  assign n12342 = n12341 ^ n12304 ;
  assign n12343 = n12340 & ~n12342 ;
  assign n12344 = n12343 ^ n12304 ;
  assign n12345 = n12169 & n12344 ;
  assign n14053 = n12284 ^ n12272 ;
  assign n14054 = n12170 & n14053 ;
  assign n14055 = n14054 ^ n12272 ;
  assign n14052 = n12314 ^ n12274 ;
  assign n14058 = n14055 ^ n14052 ;
  assign n14049 = ~n12170 & ~n12300 ;
  assign n14050 = n14049 ^ n12299 ;
  assign n14045 = n12275 ^ n12272 ;
  assign n14046 = n14045 ^ n12339 ;
  assign n14047 = n12170 & n14046 ;
  assign n14048 = n14047 ^ n12275 ;
  assign n14051 = n14050 ^ n14048 ;
  assign n14059 = n14058 ^ n14051 ;
  assign n14041 = n12301 ^ n12274 ;
  assign n14042 = n14041 ^ n12277 ;
  assign n14043 = n14042 ^ n12314 ;
  assign n14044 = ~n12170 & n14043 ;
  assign n14060 = n14059 ^ n14044 ;
  assign n14061 = n12169 & ~n14060 ;
  assign n14062 = n14061 ^ n14050 ;
  assign n14063 = ~n12345 & n14062 ;
  assign n14064 = n14040 & n14063 ;
  assign n14065 = n14064 ^ n8418 ;
  assign n14066 = n14065 ^ x73 ;
  assign n14067 = ~n14038 & ~n14066 ;
  assign n14068 = n14067 ^ n14066 ;
  assign n14069 = n14068 ^ n14038 ;
  assign n13989 = n11546 & n12012 ;
  assign n13974 = n12090 ^ n12019 ;
  assign n13975 = n13974 ^ n12110 ;
  assign n13976 = ~n11546 & ~n13975 ;
  assign n13986 = n13976 ^ n12108 ;
  assign n13979 = n12027 ^ n11828 ;
  assign n13977 = n12056 ^ n12043 ;
  assign n13978 = n13977 ^ n13976 ;
  assign n13980 = n13979 ^ n13978 ;
  assign n13981 = n13978 ^ n11546 ;
  assign n13982 = n13981 ^ n13978 ;
  assign n13983 = n13980 & n13982 ;
  assign n13984 = n13983 ^ n13978 ;
  assign n13985 = ~n11581 & n13984 ;
  assign n13987 = n13986 ^ n13985 ;
  assign n13971 = n12053 ^ n12036 ;
  assign n13972 = n13971 ^ n12029 ;
  assign n13973 = n11582 & n13972 ;
  assign n13988 = n13987 ^ n13973 ;
  assign n13990 = n13989 ^ n13988 ;
  assign n13991 = ~n13328 & ~n13990 ;
  assign n13969 = n12013 & ~n12111 ;
  assign n12075 = n12055 ^ n12015 ;
  assign n12078 = n12075 & ~n12077 ;
  assign n12079 = n12078 ^ n12015 ;
  assign n12080 = n11581 & n12079 ;
  assign n13970 = n13969 ^ n12080 ;
  assign n13992 = n13991 ^ n13970 ;
  assign n13993 = ~n12044 & n13992 ;
  assign n13994 = n13993 ^ n10818 ;
  assign n13995 = n13994 ^ x64 ;
  assign n12812 = n12788 ^ n12652 ;
  assign n12813 = n12651 & n12812 ;
  assign n12814 = n12813 ^ n12787 ;
  assign n13998 = n12814 ^ n12781 ;
  assign n13999 = n12736 & ~n13998 ;
  assign n14000 = n13999 ^ n12781 ;
  assign n14004 = n14000 ^ n10871 ;
  assign n14001 = n14000 ^ n13440 ;
  assign n12816 = n12799 ^ n12651 ;
  assign n12734 = n12653 & ~n12696 ;
  assign n12808 = n12807 ^ n12734 ;
  assign n13996 = n12816 ^ n12808 ;
  assign n13997 = n12736 & n13996 ;
  assign n14002 = n14001 ^ n13997 ;
  assign n14003 = n12774 & n14002 ;
  assign n14005 = n14004 ^ n14003 ;
  assign n14006 = n14005 ^ x120 ;
  assign n14007 = ~n13995 & n14006 ;
  assign n14071 = n14007 ^ n14006 ;
  assign n14072 = n14071 ^ n13995 ;
  assign n14109 = ~n14069 & n14072 ;
  assign n14097 = ~n14068 & n14071 ;
  assign n14079 = n14007 & n14067 ;
  assign n14070 = n14007 & ~n14069 ;
  assign n14084 = n14079 ^ n14070 ;
  assign n14077 = n14067 ^ n14038 ;
  assign n14082 = n14007 & ~n14077 ;
  assign n14083 = n14082 ^ n14007 ;
  assign n14085 = n14084 ^ n14083 ;
  assign n14106 = n14097 ^ n14085 ;
  assign n14107 = n14106 ^ n14068 ;
  assign n14073 = n14072 ^ n14006 ;
  assign n14074 = ~n14068 & ~n14073 ;
  assign n14108 = n14107 ^ n14074 ;
  assign n14110 = n14109 ^ n14108 ;
  assign n14095 = n14072 & ~n14077 ;
  assign n14105 = n14095 ^ n14072 ;
  assign n14111 = n14110 ^ n14105 ;
  assign n14112 = n14111 ^ n14079 ;
  assign n14664 = n14112 ^ n14082 ;
  assign n14081 = n14067 & ~n14073 ;
  assign n14104 = n14081 ^ n14067 ;
  assign n14113 = n14112 ^ n14104 ;
  assign n14649 = n14113 ^ n14108 ;
  assign n14121 = n14070 ^ n14069 ;
  assign n14086 = n14085 ^ n14081 ;
  assign n14087 = n14086 ^ n14082 ;
  assign n14078 = ~n14073 & ~n14077 ;
  assign n14080 = n14079 ^ n14078 ;
  assign n14088 = n14087 ^ n14080 ;
  assign n14075 = n14074 ^ n14070 ;
  assign n14076 = n14075 ^ n13995 ;
  assign n14089 = n14088 ^ n14076 ;
  assign n14120 = n14109 ^ n14089 ;
  assign n14122 = n14121 ^ n14120 ;
  assign n14661 = n14649 ^ n14122 ;
  assign n14662 = n14661 ^ n14110 ;
  assign n14665 = n14664 ^ n14662 ;
  assign n14666 = ~n13934 & n14665 ;
  assign n14658 = n14084 ^ n14081 ;
  assign n14659 = n14658 ^ n14097 ;
  assign n14660 = n14659 ^ n14074 ;
  assign n14663 = n14662 ^ n14660 ;
  assign n14667 = n14666 ^ n14663 ;
  assign n14668 = n14094 & ~n14667 ;
  assign n14656 = ~n13968 & n14082 ;
  assign n14650 = n14649 ^ n14085 ;
  assign n14123 = n14122 ^ n14113 ;
  assign n14119 = n14097 ^ n14071 ;
  assign n14124 = n14123 ^ n14119 ;
  assign n14137 = n14124 ^ n14108 ;
  assign n14647 = n14137 ^ n14111 ;
  assign n14651 = n14650 ^ n14647 ;
  assign n14652 = n13934 & ~n14651 ;
  assign n14648 = n14647 ^ n14095 ;
  assign n14653 = n14652 ^ n14648 ;
  assign n14654 = ~n14094 & ~n14653 ;
  assign n14642 = n13934 & n13968 ;
  assign n14643 = n14089 ^ n14078 ;
  assign n14644 = n14642 & ~n14643 ;
  assign n14645 = n14644 ^ n14084 ;
  assign n14140 = n14122 ^ n14078 ;
  assign n14141 = n14078 ^ n13934 ;
  assign n14142 = n14141 ^ n14078 ;
  assign n14143 = n14140 & ~n14142 ;
  assign n14144 = n14143 ^ n14078 ;
  assign n14145 = n14094 & n14144 ;
  assign n14646 = n14645 ^ n14145 ;
  assign n14655 = n14654 ^ n14646 ;
  assign n14657 = n14656 ^ n14655 ;
  assign n14669 = n14668 ^ n14657 ;
  assign n14672 = n14109 ^ n13968 ;
  assign n14673 = n14672 ^ n14109 ;
  assign n14674 = ~n14120 & ~n14673 ;
  assign n14675 = n14674 ^ n14109 ;
  assign n14676 = ~n13934 & n14675 ;
  assign n14677 = ~n14669 & ~n14676 ;
  assign n14678 = n14677 ^ n12695 ;
  assign n16031 = n14678 ^ x96 ;
  assign n12735 = n12734 ^ n12733 ;
  assign n12809 = n12808 ^ n12781 ;
  assign n12810 = n12774 & ~n12809 ;
  assign n12811 = n12810 ^ n12808 ;
  assign n12817 = n12816 ^ n12811 ;
  assign n12815 = n12814 ^ n12811 ;
  assign n12818 = n12817 ^ n12815 ;
  assign n12819 = n12817 ^ n12774 ;
  assign n12820 = n12819 ^ n12817 ;
  assign n12821 = n12818 & n12820 ;
  assign n12822 = n12821 ^ n12817 ;
  assign n12823 = n12736 & n12822 ;
  assign n12824 = n12823 ^ n12811 ;
  assign n12825 = ~n12735 & n12824 ;
  assign n12826 = n12825 ^ n10632 ;
  assign n12827 = n12826 ^ x92 ;
  assign n12966 = ~n12957 & ~n12965 ;
  assign n12968 = n12967 ^ n12925 ;
  assign n12989 = n12988 ^ n12980 ;
  assign n12976 = n12975 ^ n12913 ;
  assign n12990 = n12989 ^ n12976 ;
  assign n12977 = n12976 ^ n12922 ;
  assign n12971 = n12900 ^ n12832 ;
  assign n12972 = n12971 ^ n12922 ;
  assign n12973 = n12972 ^ n12939 ;
  assign n12974 = ~n12829 & ~n12973 ;
  assign n12978 = n12977 ^ n12974 ;
  assign n12979 = n12831 & n12978 ;
  assign n12991 = n12990 ^ n12979 ;
  assign n12992 = n12991 ^ n12970 ;
  assign n12993 = n12992 ^ n12969 ;
  assign n12994 = n12951 & ~n12993 ;
  assign n12995 = n12968 & n12994 ;
  assign n12996 = n12995 ^ n12993 ;
  assign n12997 = ~n12830 & ~n12996 ;
  assign n13001 = n13000 ^ n12923 ;
  assign n13002 = n12923 ^ n12829 ;
  assign n13003 = n13002 ^ n12923 ;
  assign n13004 = n13001 & n13003 ;
  assign n13005 = n13004 ^ n12923 ;
  assign n13006 = n12997 & n13005 ;
  assign n13007 = n13006 ^ n12996 ;
  assign n13008 = n12966 & ~n13007 ;
  assign n13009 = n13008 ^ n10668 ;
  assign n13010 = n13009 ^ x78 ;
  assign n13056 = n12827 & n13010 ;
  assign n13057 = n13056 ^ n12827 ;
  assign n13058 = n13057 ^ n13010 ;
  assign n13059 = n13058 ^ n12827 ;
  assign n11491 = n11490 ^ n11446 ;
  assign n11492 = n11446 ^ n10389 ;
  assign n11493 = n11492 ^ n11446 ;
  assign n11494 = n11491 & ~n11493 ;
  assign n11495 = n11494 ^ n11446 ;
  assign n11496 = n11431 & n11495 ;
  assign n11498 = n11497 ^ n11496 ;
  assign n11499 = n11498 ^ n11486 ;
  assign n11432 = n11417 ^ n10739 ;
  assign n11433 = n11432 ^ n11425 ;
  assign n11441 = n11440 ^ n11433 ;
  assign n11442 = n10389 & n11441 ;
  assign n11443 = n11442 ^ n11425 ;
  assign n11444 = n11431 & n11443 ;
  assign n11445 = n11444 ^ n11425 ;
  assign n11472 = n11471 ^ n11470 ;
  assign n11466 = n11465 ^ n11428 ;
  assign n11467 = n11466 ^ n11464 ;
  assign n11468 = ~n10389 & ~n11467 ;
  assign n11473 = n11472 ^ n11468 ;
  assign n11448 = n11447 ^ n11435 ;
  assign n11469 = n11468 ^ n11448 ;
  assign n11474 = n11473 ^ n11469 ;
  assign n11475 = ~n10389 & ~n11474 ;
  assign n11476 = n11475 ^ n11473 ;
  assign n11477 = n9920 & ~n11476 ;
  assign n11478 = n11477 ^ n11468 ;
  assign n11479 = ~n11445 & ~n11478 ;
  assign n11500 = n11499 ^ n11479 ;
  assign n11501 = n11500 ^ n11430 ;
  assign n11502 = n11501 ^ n10478 ;
  assign n11503 = n11502 ^ x110 ;
  assign n12094 = n12022 ^ n12018 ;
  assign n12095 = n12094 ^ n12039 ;
  assign n12096 = ~n11546 & n12095 ;
  assign n12091 = n12090 ^ n12017 ;
  assign n12092 = n12091 ^ n12088 ;
  assign n12093 = n12092 ^ n12080 ;
  assign n12097 = n12096 ^ n12093 ;
  assign n12114 = n12113 ^ n12097 ;
  assign n12098 = n12097 ^ n12088 ;
  assign n12099 = n12098 ^ n12080 ;
  assign n12074 = n11546 & n12040 ;
  assign n12100 = n12099 ^ n12074 ;
  assign n12101 = n12063 & n12100 ;
  assign n12115 = n12114 ^ n12101 ;
  assign n12072 = n12023 ^ n12017 ;
  assign n12073 = n12071 & n12072 ;
  assign n12116 = n12115 ^ n12073 ;
  assign n12066 = n12036 ^ n11581 ;
  assign n12067 = n12066 ^ n12036 ;
  assign n12068 = n12038 & ~n12067 ;
  assign n12069 = n12068 ^ n12036 ;
  assign n12070 = ~n12063 & n12069 ;
  assign n12117 = n12116 ^ n12070 ;
  assign n12118 = n12117 ^ n12062 ;
  assign n12119 = n12118 ^ n10582 ;
  assign n11583 = n11582 ^ n11546 ;
  assign n12046 = n12045 ^ n12035 ;
  assign n12047 = n11583 & ~n12046 ;
  assign n12120 = n12119 ^ n12047 ;
  assign n12121 = n12120 ^ x91 ;
  assign n12122 = ~n11503 & ~n12121 ;
  assign n13023 = n12122 ^ n12121 ;
  assign n12351 = n12350 ^ n10518 ;
  assign n12315 = n12173 & n12314 ;
  assign n12317 = n12170 ^ n12169 ;
  assign n12320 = n12319 ^ n12274 ;
  assign n12321 = n12320 ^ n12272 ;
  assign n12318 = n12313 ^ n12290 ;
  assign n12322 = n12321 ^ n12318 ;
  assign n12323 = n12170 & n12322 ;
  assign n12324 = n12323 ^ n12321 ;
  assign n12325 = n12324 ^ n12299 ;
  assign n12326 = n12325 ^ n12309 ;
  assign n12327 = n12326 ^ n12276 ;
  assign n12328 = n12327 ^ n12324 ;
  assign n12329 = n12170 & ~n12328 ;
  assign n12330 = n12329 ^ n12325 ;
  assign n12331 = ~n12317 & ~n12330 ;
  assign n12332 = n12331 ^ n12324 ;
  assign n12316 = n12170 & n12278 ;
  assign n12333 = n12332 ^ n12316 ;
  assign n12334 = ~n12315 & ~n12333 ;
  assign n12346 = n12334 & ~n12345 ;
  assign n12352 = n12351 ^ n12346 ;
  assign n12353 = n12352 ^ x116 ;
  assign n12617 = n12616 ^ n12600 ;
  assign n12618 = n12432 & n12617 ;
  assign n12584 = n12560 ^ n12477 ;
  assign n12585 = n12584 ^ n12583 ;
  assign n12586 = n12579 & ~n12585 ;
  assign n12603 = n12594 ^ n12583 ;
  assign n12608 = n12586 & n12603 ;
  assign n12567 = ~n12431 & n12566 ;
  assign n12568 = n12567 ^ n12558 ;
  assign n12570 = n12568 ^ n12552 ;
  assign n12555 = n12554 ^ n12553 ;
  assign n12569 = n12568 ^ n12555 ;
  assign n12571 = n12570 ^ n12569 ;
  assign n12572 = n12570 ^ n12400 ;
  assign n12573 = n12572 ^ n12570 ;
  assign n12574 = ~n12571 & ~n12573 ;
  assign n12575 = n12574 ^ n12570 ;
  assign n12576 = n12432 & n12575 ;
  assign n12577 = n12576 ^ n12568 ;
  assign n12604 = n12603 ^ n12577 ;
  assign n12601 = n12600 ^ n12551 ;
  assign n12602 = ~n12587 & n12601 ;
  assign n12605 = n12604 ^ n12602 ;
  assign n12609 = n12608 ^ n12605 ;
  assign n12619 = n12618 ^ n12609 ;
  assign n12620 = n12619 ^ n12602 ;
  assign n12621 = n12620 ^ n12577 ;
  assign n12622 = n12598 ^ n12589 ;
  assign n12623 = n12622 ^ n12595 ;
  assign n12624 = n12431 & ~n12623 ;
  assign n12625 = ~n12621 & n12624 ;
  assign n12626 = n12625 ^ n12619 ;
  assign n12627 = n12626 ^ n10438 ;
  assign n12628 = n12627 ^ x109 ;
  assign n12629 = ~n12353 & ~n12628 ;
  assign n13050 = n12629 ^ n12628 ;
  assign n13051 = ~n13023 & ~n13050 ;
  assign n13011 = n12629 ^ n12353 ;
  assign n13024 = ~n13011 & ~n13023 ;
  assign n13073 = n13051 ^ n13024 ;
  assign n13045 = n12629 & ~n13023 ;
  assign n13013 = n12122 ^ n11503 ;
  assign n13020 = n12629 & ~n13013 ;
  assign n13014 = n13011 ^ n12628 ;
  assign n13015 = ~n13013 & ~n13014 ;
  assign n13021 = n13020 ^ n13015 ;
  assign n13046 = n13045 ^ n13021 ;
  assign n12630 = n12122 & n12629 ;
  assign n13043 = n13015 ^ n12630 ;
  assign n13044 = n13043 ^ n12629 ;
  assign n13047 = n13046 ^ n13044 ;
  assign n13041 = n13013 ^ n12121 ;
  assign n13042 = ~n13014 & ~n13041 ;
  assign n13048 = n13047 ^ n13042 ;
  assign n13029 = n13015 ^ n13013 ;
  assign n13026 = ~n12628 & ~n13013 ;
  assign n13030 = n13029 ^ n13026 ;
  assign n13027 = n13026 ^ n13020 ;
  assign n13012 = n12122 & ~n13011 ;
  assign n13028 = n13027 ^ n13012 ;
  assign n13031 = n13030 ^ n13028 ;
  assign n13032 = n13031 ^ n13027 ;
  assign n13025 = n13024 ^ n13011 ;
  assign n13033 = n13032 ^ n13025 ;
  assign n13049 = n13048 ^ n13033 ;
  assign n13072 = n13049 ^ n13041 ;
  assign n13074 = n13073 ^ n13072 ;
  assign n13075 = n13074 ^ n13045 ;
  assign n13071 = n13049 ^ n11503 ;
  assign n13076 = n13075 ^ n13071 ;
  assign n15125 = n13059 & ~n13076 ;
  assign n13019 = n13010 ^ n12827 ;
  assign n16053 = ~n13019 & n13042 ;
  assign n13034 = n12628 ^ n12353 ;
  assign n13035 = n11503 & n13034 ;
  assign n13036 = n13035 ^ n12353 ;
  assign n13037 = n13036 ^ n12628 ;
  assign n13038 = n13037 ^ n13031 ;
  assign n15797 = n13038 ^ n13030 ;
  assign n16043 = n15797 ^ n12827 ;
  assign n16045 = n15797 ^ n13026 ;
  assign n16044 = n15797 ^ n13043 ;
  assign n16046 = n16045 ^ n16044 ;
  assign n16047 = n16045 ^ n13010 ;
  assign n16048 = n16047 ^ n16045 ;
  assign n16049 = n16046 & n16048 ;
  assign n16050 = n16049 ^ n16045 ;
  assign n16051 = ~n16043 & ~n16050 ;
  assign n16052 = n16051 ^ n12827 ;
  assign n16054 = n16053 ^ n16052 ;
  assign n16035 = n13076 ^ n13045 ;
  assign n16036 = n16035 ^ n13024 ;
  assign n16037 = n16036 ^ n13047 ;
  assign n16034 = n12628 ^ n11503 ;
  assign n16038 = n16037 ^ n16034 ;
  assign n16033 = n12121 & ~n13036 ;
  assign n16039 = n16038 ^ n16033 ;
  assign n16040 = n13010 & ~n16039 ;
  assign n16041 = n16040 ^ n16037 ;
  assign n16042 = n12827 & ~n16041 ;
  assign n16055 = n16054 ^ n16042 ;
  assign n16056 = ~n15125 & n16055 ;
  assign n16057 = n13047 ^ n13033 ;
  assign n16058 = ~n12827 & n16057 ;
  assign n16059 = n16058 ^ n13072 ;
  assign n16061 = n16059 ^ n16045 ;
  assign n16060 = n16059 ^ n16036 ;
  assign n16062 = n16061 ^ n16060 ;
  assign n16065 = ~n12827 & ~n16062 ;
  assign n16066 = n16065 ^ n16061 ;
  assign n16067 = ~n13010 & ~n16066 ;
  assign n16068 = n16067 ^ n16059 ;
  assign n16069 = n16056 & n16068 ;
  assign n16070 = n16069 ^ n12650 ;
  assign n16071 = n16070 ^ x105 ;
  assign n16072 = ~n16031 & ~n16071 ;
  assign n14207 = n11446 ^ n11422 ;
  assign n14208 = n10392 & n14207 ;
  assign n14203 = n11457 ^ n11422 ;
  assign n14204 = n10393 & n14203 ;
  assign n14198 = n11488 ^ n11454 ;
  assign n14194 = n11451 ^ n11425 ;
  assign n14195 = n14194 ^ n11437 ;
  assign n14196 = n14195 ^ n11440 ;
  assign n14197 = n10389 & n14196 ;
  assign n14199 = n14198 ^ n14197 ;
  assign n14200 = n14199 ^ n11460 ;
  assign n14201 = n14200 ^ n11428 ;
  assign n14205 = n14204 ^ n14201 ;
  assign n14191 = n11490 ^ n11425 ;
  assign n14192 = n14191 ^ n11462 ;
  assign n14193 = n14192 ^ n11449 ;
  assign n14202 = n14201 ^ n14193 ;
  assign n14206 = n14205 ^ n14202 ;
  assign n14209 = n14208 ^ n14206 ;
  assign n14210 = n11452 ^ n11429 ;
  assign n14211 = n11452 ^ n10389 ;
  assign n14212 = n14211 ^ n11452 ;
  assign n14213 = ~n14210 & n14212 ;
  assign n14214 = n14213 ^ n11452 ;
  assign n14215 = n14209 & ~n14214 ;
  assign n14216 = n14215 ^ n14205 ;
  assign n14217 = n11431 & ~n14216 ;
  assign n14218 = n14217 ^ n14205 ;
  assign n14219 = ~n14008 & ~n14218 ;
  assign n14220 = ~n11496 & n14219 ;
  assign n14221 = n14220 ^ n11059 ;
  assign n14807 = n14221 ^ x98 ;
  assign n14808 = n13994 ^ x107 ;
  assign n14809 = ~n14807 & n14808 ;
  assign n14810 = n14809 ^ n14808 ;
  assign n14852 = n12614 ^ n12560 ;
  assign n14850 = n12563 ^ n12548 ;
  assign n14853 = n14852 ^ n14850 ;
  assign n14854 = n12431 & n14853 ;
  assign n14849 = n12622 ^ n12559 ;
  assign n14851 = n14850 ^ n14849 ;
  assign n14855 = n14854 ^ n14851 ;
  assign n14856 = ~n12432 & ~n14855 ;
  assign n14857 = n14856 ^ n12559 ;
  assign n14848 = ~n12431 & ~n12553 ;
  assign n14858 = n14857 ^ n14848 ;
  assign n13127 = n12578 ^ n12400 ;
  assign n14846 = n12589 ^ n12564 ;
  assign n14847 = ~n13127 & n14846 ;
  assign n14859 = n14858 ^ n14847 ;
  assign n14845 = n12432 & n12595 ;
  assign n14860 = n14859 ^ n14845 ;
  assign n14861 = n12616 ^ n12431 ;
  assign n14862 = n14861 ^ n12616 ;
  assign n13562 = n12564 ^ n12554 ;
  assign n14863 = n12400 & n13562 ;
  assign n14864 = n14863 ^ n12616 ;
  assign n14865 = ~n14862 & n14864 ;
  assign n14866 = n14865 ^ n12616 ;
  assign n14867 = ~n14860 & n14866 ;
  assign n14868 = n14867 ^ n14860 ;
  assign n14869 = ~n12602 & ~n14868 ;
  assign n14870 = n14869 ^ n11880 ;
  assign n14844 = ~n12432 & ~n13113 ;
  assign n14873 = n14870 ^ n14844 ;
  assign n14874 = n14873 ^ x96 ;
  assign n14287 = n13273 ^ n13221 ;
  assign n14284 = n13249 ^ n13233 ;
  assign n14285 = ~n13222 & ~n14284 ;
  assign n14286 = n14285 ^ n13249 ;
  assign n14288 = n14287 ^ n14286 ;
  assign n14289 = n14288 ^ n13237 ;
  assign n14290 = n14289 ^ n13221 ;
  assign n14291 = n14290 ^ n14288 ;
  assign n14292 = n14288 ^ n13222 ;
  assign n14293 = n14292 ^ n14288 ;
  assign n14294 = n14291 & ~n14293 ;
  assign n14295 = n14294 ^ n14288 ;
  assign n14296 = n13223 & n14295 ;
  assign n14297 = n14296 ^ n14286 ;
  assign n13787 = n13260 ^ n13223 ;
  assign n13788 = n13787 ^ n13260 ;
  assign n13789 = n13261 & ~n13788 ;
  assign n13790 = n13789 ^ n13260 ;
  assign n13791 = ~n13281 & n13790 ;
  assign n14310 = n14297 ^ n13791 ;
  assign n14305 = n13259 ^ n13222 ;
  assign n14306 = n14305 ^ n13259 ;
  assign n14307 = n13270 & ~n14306 ;
  assign n14308 = n14307 ^ n13259 ;
  assign n14309 = n13281 & n14308 ;
  assign n14311 = n14310 ^ n14309 ;
  assign n13763 = n13277 ^ n13269 ;
  assign n14282 = n13763 ^ n13223 ;
  assign n14283 = n14282 ^ n13763 ;
  assign n14298 = n13238 & n14297 ;
  assign n14299 = n14298 ^ n13763 ;
  assign n14300 = n14283 & n14299 ;
  assign n14301 = n14300 ^ n13763 ;
  assign n14302 = n13222 & n14301 ;
  assign n14312 = n14311 ^ n14302 ;
  assign n14313 = n14312 ^ n13228 ;
  assign n14314 = n14313 ^ n11099 ;
  assign n14875 = n14314 ^ x122 ;
  assign n14876 = n14874 & ~n14875 ;
  assign n14877 = n14876 ^ n14874 ;
  assign n14878 = n14877 ^ n14875 ;
  assign n14879 = n14878 ^ n14874 ;
  assign n14812 = n13933 ^ x113 ;
  assign n14831 = n12171 ^ n12169 ;
  assign n14407 = n12348 ^ n12306 ;
  assign n14832 = n14407 ^ n12319 ;
  assign n14399 = n12339 ^ n12274 ;
  assign n14827 = n14399 ^ n12275 ;
  assign n14833 = n14832 ^ n14827 ;
  assign n14834 = ~n14831 & ~n14833 ;
  assign n14828 = n14827 ^ n12337 ;
  assign n14829 = n12172 & n14828 ;
  assign n14822 = n12302 ^ n12278 ;
  assign n14823 = n14822 ^ n12338 ;
  assign n14824 = n12171 & n14823 ;
  assign n14821 = n12170 & n12309 ;
  assign n14825 = n14824 ^ n14821 ;
  assign n14814 = n12306 ^ n12301 ;
  assign n14815 = n14814 ^ n12311 ;
  assign n14816 = n12311 ^ n12170 ;
  assign n14817 = n14816 ^ n12311 ;
  assign n14818 = ~n14815 & n14817 ;
  assign n14819 = n14818 ^ n12311 ;
  assign n14820 = n12169 & n14819 ;
  assign n14826 = n14825 ^ n14820 ;
  assign n14830 = n14829 ^ n14826 ;
  assign n14835 = n14834 ^ n14830 ;
  assign n14391 = n14054 ^ n12284 ;
  assign n14836 = n14835 ^ n14391 ;
  assign n14837 = n14836 ^ n14039 ;
  assign n14813 = n12169 & n14053 ;
  assign n14838 = n14837 ^ n14813 ;
  assign n14839 = ~n12315 & ~n14838 ;
  assign n14840 = n14839 ^ n11855 ;
  assign n14841 = n14840 ^ x74 ;
  assign n14842 = ~n14812 & ~n14841 ;
  assign n14886 = n14842 ^ n14812 ;
  assign n14895 = ~n14879 & ~n14886 ;
  assign n14892 = n14842 & n14877 ;
  assign n14888 = n14886 ^ n14841 ;
  assign n14889 = n14878 & ~n14888 ;
  assign n14887 = n14878 & ~n14886 ;
  assign n14890 = n14889 ^ n14887 ;
  assign n14843 = n14842 ^ n14841 ;
  assign n14884 = ~n14843 & n14878 ;
  assign n14885 = n14884 ^ n14878 ;
  assign n14891 = n14890 ^ n14885 ;
  assign n14893 = n14892 ^ n14891 ;
  assign n14882 = n14842 & n14876 ;
  assign n14883 = n14882 ^ n14842 ;
  assign n14894 = n14893 ^ n14883 ;
  assign n14896 = n14895 ^ n14894 ;
  assign n14880 = ~n14843 & ~n14879 ;
  assign n14881 = n14880 ^ n14879 ;
  assign n14897 = n14896 ^ n14881 ;
  assign n15250 = n14810 & ~n14897 ;
  assign n14914 = n14876 & ~n14888 ;
  assign n14915 = n14914 ^ n14892 ;
  assign n16010 = n14915 ^ n14884 ;
  assign n14902 = ~n14843 & n14876 ;
  assign n14916 = n14915 ^ n14902 ;
  assign n14912 = n14875 ^ n14812 ;
  assign n14913 = n14874 & n14912 ;
  assign n14917 = n14916 ^ n14913 ;
  assign n14903 = n14902 ^ n14895 ;
  assign n14904 = n14903 ^ n14880 ;
  assign n14900 = n14895 ^ n14884 ;
  assign n14901 = n14900 ^ n14843 ;
  assign n14905 = n14904 ^ n14901 ;
  assign n14918 = n14917 ^ n14905 ;
  assign n16011 = n16010 ^ n14918 ;
  assign n16012 = n16011 ^ n16010 ;
  assign n16013 = n16010 ^ n14808 ;
  assign n16014 = n16013 ^ n16010 ;
  assign n16015 = ~n16012 & ~n16014 ;
  assign n16016 = n16015 ^ n16010 ;
  assign n16017 = n14807 & n16016 ;
  assign n16018 = n16017 ^ n14914 ;
  assign n14910 = n14808 ^ n14807 ;
  assign n14960 = n14905 ^ n14887 ;
  assign n16002 = n14960 ^ n14892 ;
  assign n16003 = n16002 ^ n14915 ;
  assign n16004 = n16003 ^ n14892 ;
  assign n16005 = n14892 ^ n14807 ;
  assign n16006 = n16005 ^ n14892 ;
  assign n16007 = ~n16004 & ~n16006 ;
  assign n16008 = n16007 ^ n14892 ;
  assign n16009 = n14910 & n16008 ;
  assign n16019 = n16018 ^ n16009 ;
  assign n14948 = n14810 & n14887 ;
  assign n16020 = n16019 ^ n14948 ;
  assign n14811 = n14810 ^ n14807 ;
  assign n14899 = n14811 ^ n14808 ;
  assign n15856 = n14882 & ~n14899 ;
  assign n14937 = n14891 ^ n14880 ;
  assign n14938 = n14807 & n14937 ;
  assign n14939 = n14938 ^ n14880 ;
  assign n14936 = n14917 ^ n14884 ;
  assign n14940 = n14939 ^ n14936 ;
  assign n14941 = n14940 ^ n14939 ;
  assign n14942 = n14939 ^ n14807 ;
  assign n14943 = n14942 ^ n14939 ;
  assign n14944 = n14941 & ~n14943 ;
  assign n14945 = n14944 ^ n14939 ;
  assign n14946 = n14808 & n14945 ;
  assign n14947 = n14946 ^ n14939 ;
  assign n15857 = n15856 ^ n14947 ;
  assign n16021 = n16020 ^ n15857 ;
  assign n14928 = n14918 ^ n14892 ;
  assign n14929 = n14928 ^ n14877 ;
  assign n14926 = n14882 ^ n14876 ;
  assign n14925 = n14914 ^ n14902 ;
  assign n14927 = n14926 ^ n14925 ;
  assign n14930 = n14929 ^ n14927 ;
  assign n14931 = n14929 ^ n14807 ;
  assign n14932 = n14931 ^ n14929 ;
  assign n14933 = ~n14930 & ~n14932 ;
  assign n14934 = n14933 ^ n14929 ;
  assign n14935 = ~n14910 & ~n14934 ;
  assign n16022 = n16021 ^ n14935 ;
  assign n16023 = n16022 ^ n14896 ;
  assign n14898 = n14811 & ~n14897 ;
  assign n16024 = n16023 ^ n14898 ;
  assign n15230 = n14902 ^ n14807 ;
  assign n15231 = n15230 ^ n14902 ;
  assign n15242 = n14925 & n15231 ;
  assign n15243 = n15242 ^ n14902 ;
  assign n15244 = n14910 & n15243 ;
  assign n16025 = n16024 ^ n15244 ;
  assign n15245 = n14918 ^ n14889 ;
  assign n15246 = ~n14899 & ~n15245 ;
  assign n14971 = n14897 ^ n14880 ;
  assign n14972 = n14880 ^ n14807 ;
  assign n14973 = n14972 ^ n14880 ;
  assign n14974 = ~n14971 & ~n14973 ;
  assign n14975 = n14974 ^ n14880 ;
  assign n14976 = n14808 & n14975 ;
  assign n15247 = n15246 ^ n14976 ;
  assign n16026 = n16025 ^ n15247 ;
  assign n15995 = n14896 ^ n14891 ;
  assign n15996 = n15995 ^ n14876 ;
  assign n15997 = n15996 ^ n14896 ;
  assign n15998 = n15997 ^ n14925 ;
  assign n15999 = n14807 & n15998 ;
  assign n16000 = n15999 ^ n15995 ;
  assign n16001 = ~n14910 & n16000 ;
  assign n16027 = n16026 ^ n16001 ;
  assign n16028 = ~n15250 & ~n16027 ;
  assign n16029 = n16028 ^ n12430 ;
  assign n16030 = n16029 ^ x115 ;
  assign n16032 = ~n16030 & ~n16031 ;
  assign n16073 = n16072 ^ n16032 ;
  assign n16074 = n15994 & n16073 ;
  assign n13577 = n11502 ^ x85 ;
  assign n13574 = n12562 & n12578 ;
  assign n13571 = n12594 ^ n12562 ;
  assign n13572 = ~n12431 & ~n13571 ;
  assign n13569 = ~n12622 & ~n13127 ;
  assign n13566 = n12563 ^ n12476 ;
  assign n13567 = n12432 & n13566 ;
  assign n13563 = n13562 ^ n12593 ;
  assign n13564 = n12578 & n13563 ;
  assign n13556 = n12559 ^ n12478 ;
  assign n13557 = n13556 ^ n12612 ;
  assign n13550 = n12595 ^ n12560 ;
  assign n13551 = n13550 ^ n12555 ;
  assign n13552 = n12431 & ~n13551 ;
  assign n13553 = n13552 ^ n13116 ;
  assign n13558 = n13557 ^ n13553 ;
  assign n13559 = n13558 ^ n13116 ;
  assign n13560 = n12432 & ~n13559 ;
  assign n13554 = n12602 ^ n11263 ;
  assign n13555 = n13554 ^ n13553 ;
  assign n13561 = n13560 ^ n13555 ;
  assign n13565 = n13564 ^ n13561 ;
  assign n13568 = n13567 ^ n13565 ;
  assign n13570 = n13569 ^ n13568 ;
  assign n13573 = n13572 ^ n13570 ;
  assign n13575 = n13574 ^ n13573 ;
  assign n13576 = n13575 ^ x94 ;
  assign n13578 = n13577 ^ n13576 ;
  assign n13750 = n13009 ^ x76 ;
  assign n13796 = n13450 ^ n13448 ;
  assign n13797 = n13796 ^ n11293 ;
  assign n13798 = n13797 ^ x67 ;
  assign n13804 = ~n13750 & ~n13798 ;
  assign n13661 = n13654 & ~n13660 ;
  assign n13666 = ~n13660 & n13665 ;
  assign n13671 = n13670 ^ n13666 ;
  assign n13672 = n13656 ^ n13655 ;
  assign n13729 = ~n13672 & n13693 ;
  assign n13711 = n13710 ^ n13646 ;
  assign n13696 = n13695 ^ n13669 ;
  assign n13712 = n13711 ^ n13696 ;
  assign n13713 = n13655 & ~n13712 ;
  assign n13714 = n13713 ^ n13696 ;
  assign n13725 = n13720 ^ n13714 ;
  assign n13716 = n13702 ^ n13686 ;
  assign n13721 = n13720 ^ n13716 ;
  assign n13723 = n13722 ^ n13721 ;
  assign n13724 = ~n13655 & ~n13723 ;
  assign n13726 = n13725 ^ n13724 ;
  assign n13727 = n13656 & n13726 ;
  assign n13687 = n13686 ^ n13665 ;
  assign n13688 = n13665 ^ n13655 ;
  assign n13689 = n13688 ^ n13665 ;
  assign n13690 = ~n13687 & n13689 ;
  assign n13691 = n13690 ^ n13665 ;
  assign n13692 = ~n13672 & n13691 ;
  assign n13715 = n13714 ^ n13692 ;
  assign n13728 = n13727 ^ n13715 ;
  assign n13730 = n13729 ^ n13728 ;
  assign n13731 = ~n13671 & ~n13730 ;
  assign n13738 = n13731 & ~n13737 ;
  assign n13743 = ~n13689 & ~n13740 ;
  assign n13744 = n13743 ^ n13665 ;
  assign n13745 = ~n13656 & n13744 ;
  assign n13746 = n13738 & ~n13745 ;
  assign n13747 = ~n13661 & n13746 ;
  assign n13748 = n13747 ^ n11320 ;
  assign n13749 = n13748 ^ x117 ;
  assign n13783 = ~n13247 & ~n13281 ;
  assign n13776 = ~n13222 & n13245 ;
  assign n13777 = n13776 ^ n13275 ;
  assign n13767 = n13296 ^ n13281 ;
  assign n13768 = n13767 ^ n13296 ;
  assign n13769 = ~n13226 & ~n13263 ;
  assign n13770 = n13769 ^ n13268 ;
  assign n13771 = ~n13221 & ~n13770 ;
  assign n13772 = n13768 & n13771 ;
  assign n13773 = n13772 ^ n13767 ;
  assign n13778 = n13777 ^ n13773 ;
  assign n13752 = n13281 ^ n13236 ;
  assign n13753 = n13239 ^ n13236 ;
  assign n13754 = n13753 ^ n13223 ;
  assign n13755 = n13754 ^ n13753 ;
  assign n13756 = n13281 ^ n13245 ;
  assign n13757 = n13756 ^ n13753 ;
  assign n13758 = ~n13755 & ~n13757 ;
  assign n13759 = n13758 ^ n13753 ;
  assign n13760 = n13752 & n13759 ;
  assign n13761 = n13760 ^ n13236 ;
  assign n13779 = n13778 ^ n13761 ;
  assign n13766 = n13270 ^ n13256 ;
  assign n13774 = n13222 & n13773 ;
  assign n13775 = n13766 & n13774 ;
  assign n13780 = n13779 ^ n13775 ;
  assign n13764 = n13763 ^ n13262 ;
  assign n13765 = n13225 & ~n13764 ;
  assign n13781 = n13780 ^ n13765 ;
  assign n13751 = ~n13222 & n13237 ;
  assign n13782 = n13781 ^ n13751 ;
  assign n13784 = n13783 ^ n13782 ;
  assign n13792 = ~n13784 & ~n13791 ;
  assign n13793 = n13792 ^ n11287 ;
  assign n13794 = n13793 ^ x124 ;
  assign n13802 = n13749 & ~n13794 ;
  assign n13810 = n13802 ^ n13794 ;
  assign n13815 = n13804 & ~n13810 ;
  assign n13805 = n13804 ^ n13798 ;
  assign n13811 = n13810 ^ n13749 ;
  assign n13814 = ~n13805 & n13811 ;
  assign n13816 = n13815 ^ n13814 ;
  assign n13812 = n13811 ^ n13794 ;
  assign n13813 = ~n13805 & n13812 ;
  assign n13817 = n13816 ^ n13813 ;
  assign n13808 = ~n13794 & ~n13798 ;
  assign n13809 = n13808 ^ n13805 ;
  assign n13818 = n13817 ^ n13809 ;
  assign n13819 = n13818 ^ n13813 ;
  assign n13795 = ~n13750 & ~n13794 ;
  assign n13853 = n13819 ^ n13795 ;
  assign n13844 = n13794 ^ n13750 ;
  assign n13845 = n13808 ^ n13749 ;
  assign n13846 = ~n13844 & n13845 ;
  assign n13836 = n13804 & n13811 ;
  assign n13806 = n13805 ^ n13750 ;
  assign n13823 = ~n13806 & ~n13810 ;
  assign n13839 = n13836 ^ n13823 ;
  assign n13840 = n13839 ^ n13815 ;
  assign n13835 = ~n13805 & ~n13810 ;
  assign n13837 = n13836 ^ n13835 ;
  assign n13838 = n13837 ^ n13810 ;
  assign n13841 = n13840 ^ n13838 ;
  assign n13847 = n13846 ^ n13841 ;
  assign n13854 = n13853 ^ n13847 ;
  assign n13887 = n13854 ^ n13812 ;
  assign n13807 = n13802 & ~n13806 ;
  assign n13820 = n13819 ^ n13807 ;
  assign n13799 = n13798 ^ n13795 ;
  assign n13800 = n13749 & n13799 ;
  assign n13801 = n13800 ^ n13749 ;
  assign n13803 = n13802 ^ n13801 ;
  assign n13821 = n13820 ^ n13803 ;
  assign n13875 = n13821 ^ n13813 ;
  assign n13888 = n13887 ^ n13875 ;
  assign n13868 = n13836 ^ n13811 ;
  assign n13824 = n13806 ^ n13798 ;
  assign n13825 = n13811 & ~n13824 ;
  assign n13826 = n13825 ^ n13814 ;
  assign n13869 = n13868 ^ n13826 ;
  assign n13889 = n13888 ^ n13869 ;
  assign n13890 = n13869 ^ n13577 ;
  assign n13891 = n13890 ^ n13869 ;
  assign n13892 = ~n13889 & ~n13891 ;
  assign n13893 = n13892 ^ n13869 ;
  assign n13894 = n13578 & n13893 ;
  assign n16109 = n13894 ^ n12503 ;
  assign n13870 = n13576 & n13577 ;
  assign n13871 = n13870 ^ n13576 ;
  assign n13872 = n13869 & n13871 ;
  assign n13873 = n13576 & ~n13872 ;
  assign n13874 = n13802 & ~n13805 ;
  assign n13876 = n13875 ^ n13874 ;
  assign n13877 = n13876 ^ n13801 ;
  assign n13878 = n13877 ^ n13874 ;
  assign n13879 = n13878 ^ n13841 ;
  assign n13880 = n13878 ^ n13577 ;
  assign n13881 = n13880 ^ n13878 ;
  assign n13882 = n13879 & n13881 ;
  assign n13883 = n13882 ^ n13878 ;
  assign n13884 = n13873 & ~n13883 ;
  assign n13885 = n13884 ^ n13872 ;
  assign n16102 = n13869 ^ n13819 ;
  assign n16103 = n16102 ^ n13835 ;
  assign n16104 = n13577 & ~n16103 ;
  assign n15343 = n13869 ^ n13846 ;
  assign n15342 = n13839 ^ n13835 ;
  assign n15344 = n15343 ^ n15342 ;
  assign n16095 = n15344 ^ n13840 ;
  assign n16096 = n16095 ^ n13888 ;
  assign n16097 = n13577 & n16096 ;
  assign n16098 = n16097 ^ n15344 ;
  assign n16101 = n16098 ^ n13817 ;
  assign n16105 = n16104 ^ n16101 ;
  assign n16106 = n13576 & ~n16105 ;
  assign n15357 = n13854 ^ n13821 ;
  assign n15358 = n15357 ^ n13877 ;
  assign n15359 = n13877 ^ n13576 ;
  assign n15360 = n15359 ^ n13877 ;
  assign n15361 = n15358 & n15360 ;
  assign n15362 = n15361 ^ n13877 ;
  assign n15363 = n13577 & ~n15362 ;
  assign n16099 = n16098 ^ n15363 ;
  assign n15620 = n13841 ^ n13819 ;
  assign n15621 = n13819 ^ n13577 ;
  assign n15622 = n15621 ^ n13819 ;
  assign n15623 = n15620 & ~n15622 ;
  assign n15624 = n15623 ^ n13819 ;
  assign n15625 = n13578 & ~n15624 ;
  assign n16100 = n16099 ^ n15625 ;
  assign n16107 = n16106 ^ n16100 ;
  assign n16108 = ~n13885 & n16107 ;
  assign n16110 = n16109 ^ n16108 ;
  assign n16111 = n16110 ^ x72 ;
  assign n16080 = n16071 ^ n16030 ;
  assign n16076 = n16030 ^ n15994 ;
  assign n16077 = n16076 ^ n16031 ;
  assign n16078 = n16072 ^ n16030 ;
  assign n16079 = n16077 & n16078 ;
  assign n16081 = n16080 ^ n16079 ;
  assign n16083 = n16031 ^ n16030 ;
  assign n16084 = n16071 ^ n16031 ;
  assign n16087 = ~n16083 & n16084 ;
  assign n16088 = n16087 ^ n16031 ;
  assign n16089 = ~n16077 & n16088 ;
  assign n16118 = n16081 & ~n16089 ;
  assign n14167 = n12352 ^ x104 ;
  assign n14315 = n14314 ^ x82 ;
  assign n14168 = ~n12949 & ~n13936 ;
  assign n14180 = n12921 ^ n12917 ;
  assign n14181 = n14180 ^ n12938 ;
  assign n14182 = ~n12829 & n14181 ;
  assign n14179 = n12938 ^ n12934 ;
  assign n14183 = n14182 ^ n14179 ;
  assign n14184 = ~n12830 & n14183 ;
  assign n14177 = n12829 & n12938 ;
  assign n14175 = n13367 ^ n12934 ;
  assign n14176 = n14175 ^ n13961 ;
  assign n14178 = n14177 ^ n14176 ;
  assign n14185 = n14184 ^ n14178 ;
  assign n14169 = n12999 ^ n12940 ;
  assign n14170 = n12940 ^ n12830 ;
  assign n14171 = n14170 ^ n12940 ;
  assign n14172 = n14169 & n14171 ;
  assign n14173 = n14172 ^ n12940 ;
  assign n14174 = n12829 & n14173 ;
  assign n14186 = n14185 ^ n14174 ;
  assign n14187 = ~n13352 & ~n14186 ;
  assign n14188 = n14168 & n14187 ;
  assign n14189 = n14188 ^ n11028 ;
  assign n14190 = n14189 ^ x99 ;
  assign n14222 = n14221 ^ x114 ;
  assign n14223 = n14190 & n14222 ;
  assign n14329 = n14223 ^ n14190 ;
  assign n14224 = n13718 ^ n13656 ;
  assign n14225 = n14224 ^ n13655 ;
  assign n14234 = n13656 ^ n13652 ;
  assign n14235 = n13686 ^ n13652 ;
  assign n14236 = n14235 ^ n13701 ;
  assign n14237 = n14236 ^ n14235 ;
  assign n14238 = n14235 ^ n13655 ;
  assign n14239 = n14238 ^ n14235 ;
  assign n14240 = n14237 & n14239 ;
  assign n14241 = n14240 ^ n14235 ;
  assign n14242 = ~n14234 & n14241 ;
  assign n14243 = n14242 ^ n13656 ;
  assign n14229 = n13705 ^ n13655 ;
  assign n14230 = n14229 ^ n13705 ;
  assign n14231 = n13710 & n14230 ;
  assign n14232 = n14231 ^ n13705 ;
  assign n14233 = n13656 & ~n14232 ;
  assign n14244 = n14243 ^ n14233 ;
  assign n14226 = ~n13659 & n13703 ;
  assign n14245 = n14244 ^ n14226 ;
  assign n14246 = ~n14225 & n14245 ;
  assign n14247 = n14246 ^ n14245 ;
  assign n14250 = n14246 ^ n13674 ;
  assign n14251 = n14250 ^ n14246 ;
  assign n14252 = n14246 ^ n13656 ;
  assign n14253 = n14252 ^ n14246 ;
  assign n14254 = n14251 & ~n14253 ;
  assign n14255 = n14247 & n14254 ;
  assign n14256 = n14255 ^ n14247 ;
  assign n14257 = n14256 ^ n14245 ;
  assign n14258 = n13672 & n14257 ;
  assign n14259 = n14258 ^ n14245 ;
  assign n14260 = ~n13655 & n14259 ;
  assign n14261 = n13706 ^ n13656 ;
  assign n14262 = n14261 ^ n13706 ;
  assign n14263 = n13706 ^ n13668 ;
  assign n14264 = n14263 ^ n13706 ;
  assign n14265 = ~n14262 & n14264 ;
  assign n14266 = n14265 ^ n13706 ;
  assign n14267 = n14260 & n14266 ;
  assign n14268 = n14267 ^ n14259 ;
  assign n14269 = ~n13692 & n14268 ;
  assign n14270 = ~n13661 & ~n13899 ;
  assign n14271 = n14269 & n14270 ;
  assign n14272 = n14271 ^ n11149 ;
  assign n14273 = n14272 ^ x89 ;
  assign n14274 = n12826 ^ x80 ;
  assign n14275 = n14273 & n14274 ;
  assign n14334 = n14275 ^ n14274 ;
  assign n14335 = n14329 & n14334 ;
  assign n14277 = n14223 ^ n14222 ;
  assign n14321 = n14277 ^ n14190 ;
  assign n14327 = n14275 & ~n14321 ;
  assign n15025 = n14335 ^ n14327 ;
  assign n14339 = ~n14321 & n14334 ;
  assign n14338 = n14223 & n14334 ;
  assign n14340 = n14339 ^ n14338 ;
  assign n14330 = n14275 & n14329 ;
  assign n14341 = n14340 ^ n14330 ;
  assign n14331 = n14330 ^ n14275 ;
  assign n14336 = n14335 ^ n14331 ;
  assign n14337 = n14336 ^ n14274 ;
  assign n14342 = n14341 ^ n14337 ;
  assign n14375 = n14342 ^ n14330 ;
  assign n14376 = n14375 ^ n14338 ;
  assign n15026 = n15025 ^ n14376 ;
  assign n15027 = n14315 & n15026 ;
  assign n14278 = n14275 ^ n14273 ;
  assign n14279 = n14278 ^ n14274 ;
  assign n14280 = n14277 & ~n14279 ;
  assign n15028 = n15027 ^ n14280 ;
  assign n15029 = n14167 & n15028 ;
  assign n14325 = n14223 & ~n14279 ;
  assign n14991 = n14167 & n14315 ;
  assign n14995 = n14991 ^ n14315 ;
  assign n15022 = n14995 ^ n14167 ;
  assign n15023 = n14325 & ~n15022 ;
  assign n14372 = n14315 ^ n14167 ;
  assign n15003 = n14336 ^ n14167 ;
  assign n14276 = n14223 & n14275 ;
  assign n15000 = n14330 ^ n14276 ;
  assign n15001 = n15000 ^ n14336 ;
  assign n15002 = n14315 & ~n15001 ;
  assign n15004 = n15003 ^ n15002 ;
  assign n15005 = n15004 ^ n14315 ;
  assign n15006 = n15005 ^ n15004 ;
  assign n15007 = n15005 ^ n14341 ;
  assign n15008 = n15007 ^ n15005 ;
  assign n15009 = n15005 ^ n14276 ;
  assign n15010 = n15009 ^ n15005 ;
  assign n15011 = ~n15008 & ~n15010 ;
  assign n15012 = ~n15006 & n15011 ;
  assign n15013 = n15012 ^ n15006 ;
  assign n15014 = n15013 ^ n15004 ;
  assign n15015 = ~n14372 & n15014 ;
  assign n15016 = n15015 ^ n15004 ;
  assign n14346 = ~n14279 & ~n14321 ;
  assign n14347 = n14346 ^ n14279 ;
  assign n14345 = n14325 ^ n14280 ;
  assign n14348 = n14347 ^ n14345 ;
  assign n14323 = n14223 & n14278 ;
  assign n14996 = n14348 ^ n14323 ;
  assign n14997 = n14996 ^ n14346 ;
  assign n14328 = n14327 ^ n14276 ;
  assign n14332 = n14331 ^ n14328 ;
  assign n14998 = n14997 ^ n14332 ;
  assign n14999 = n14995 & ~n14998 ;
  assign n15017 = n15016 ^ n14999 ;
  assign n14992 = n14991 ^ n14167 ;
  assign n14322 = n14278 & ~n14321 ;
  assign n14324 = n14323 ^ n14322 ;
  assign n14361 = n14324 ^ n14278 ;
  assign n14343 = n14342 ^ n14277 ;
  assign n14333 = n14332 ^ n14280 ;
  assign n14344 = n14343 ^ n14333 ;
  assign n14362 = n14361 ^ n14344 ;
  assign n14993 = n14362 ^ n14347 ;
  assign n14994 = n14992 & ~n14993 ;
  assign n15018 = n15017 ^ n14994 ;
  assign n15019 = n15018 ^ n14280 ;
  assign n14349 = n14348 ^ n14344 ;
  assign n14350 = n14349 ^ n14339 ;
  assign n14351 = ~n14315 & ~n14350 ;
  assign n14352 = n14351 ^ n14339 ;
  assign n14326 = n14325 ^ n14324 ;
  assign n14353 = n14352 ^ n14326 ;
  assign n14354 = n14353 ^ n14352 ;
  assign n14357 = n14315 & n14354 ;
  assign n14358 = n14357 ^ n14352 ;
  assign n14359 = n14167 & n14358 ;
  assign n14360 = n14359 ^ n14352 ;
  assign n15020 = n15019 ^ n14360 ;
  assign n15021 = n15020 ^ n12773 ;
  assign n15024 = n15023 ^ n15021 ;
  assign n15030 = n15029 ^ n15024 ;
  assign n15968 = n15030 ^ x90 ;
  assign n16223 = n16118 ^ n15968 ;
  assign n16112 = n16071 ^ n15994 ;
  assign n16113 = n16084 ^ n15994 ;
  assign n16114 = ~n16076 & n16113 ;
  assign n16115 = n16114 ^ n16030 ;
  assign n16116 = n16112 & ~n16115 ;
  assign n16117 = n16116 ^ n16084 ;
  assign n16119 = n16118 ^ n16117 ;
  assign n16120 = n15968 & n16119 ;
  assign n16121 = n16120 ^ n16118 ;
  assign n16224 = n16223 ^ n16121 ;
  assign n16225 = n16224 ^ n16117 ;
  assign n16090 = n16089 ^ n16031 ;
  assign n16227 = n16225 ^ n16090 ;
  assign n16226 = n16225 ^ n16081 ;
  assign n16228 = n16227 ^ n16226 ;
  assign n16229 = n16227 ^ n15968 ;
  assign n16230 = n16229 ^ n16227 ;
  assign n16231 = ~n16228 & n16230 ;
  assign n16232 = n16231 ^ n16227 ;
  assign n16233 = ~n16111 & ~n16232 ;
  assign n16234 = n16233 ^ n16225 ;
  assign n16235 = ~n16074 & n16234 ;
  assign n16236 = n16235 ^ n12826 ;
  assign n17495 = n16236 ^ x113 ;
  assign n14784 = n13349 ^ x106 ;
  assign n14680 = n14065 ^ x88 ;
  assign n14749 = n13967 ^ x66 ;
  assign n14738 = n13684 ^ n13668 ;
  assign n14739 = ~n13658 & ~n14738 ;
  assign n14724 = n13674 ^ n13650 ;
  assign n14725 = n13655 & ~n14724 ;
  assign n14723 = n13925 ^ n13669 ;
  assign n14726 = n14725 ^ n14723 ;
  assign n14729 = n14726 ^ n13705 ;
  assign n14732 = n14729 ^ n13647 ;
  assign n14733 = n14732 ^ n14729 ;
  assign n14734 = n13655 & n14733 ;
  assign n14735 = n14734 ^ n14729 ;
  assign n14736 = ~n13656 & ~n14735 ;
  assign n14727 = n14726 ^ n13661 ;
  assign n14728 = n14727 ^ n13913 ;
  assign n14737 = n14736 ^ n14728 ;
  assign n14740 = n14739 ^ n14737 ;
  assign n14741 = n14740 ^ n13706 ;
  assign n14722 = n13657 & n13679 ;
  assign n14742 = n14741 ^ n14722 ;
  assign n14715 = n13706 ^ n13659 ;
  assign n14716 = n13902 ^ n13657 ;
  assign n14719 = ~n13659 & n14716 ;
  assign n14720 = n14719 ^ n13657 ;
  assign n14721 = ~n14715 & ~n14720 ;
  assign n14743 = n14742 ^ n14721 ;
  assign n14744 = ~n13671 & ~n14743 ;
  assign n14745 = ~n13745 & n14744 ;
  assign n14746 = n14745 ^ n9511 ;
  assign n14747 = n14746 ^ x65 ;
  assign n14681 = ~n13228 & ~n13777 ;
  assign n14696 = n13262 ^ n13227 ;
  assign n14697 = n14696 ^ n13267 ;
  assign n14698 = n14697 ^ n13276 ;
  assign n14699 = ~n13769 & ~n14698 ;
  assign n14700 = n14699 ^ n13269 ;
  assign n14708 = n14700 ^ n13295 ;
  assign n14701 = n14700 ^ n13266 ;
  assign n14702 = n14701 ^ n13256 ;
  assign n14703 = n14702 ^ n14700 ;
  assign n14704 = n14703 ^ n13284 ;
  assign n14705 = ~n13222 & ~n14704 ;
  assign n14706 = n14705 ^ n14701 ;
  assign n14707 = n13223 & ~n14706 ;
  assign n14709 = n14708 ^ n14707 ;
  assign n14688 = n13257 ^ n13236 ;
  assign n14689 = n14688 ^ n13259 ;
  assign n14690 = n14689 ^ n13236 ;
  assign n14691 = n13236 ^ n13223 ;
  assign n14692 = n14691 ^ n13236 ;
  assign n14693 = n14690 & ~n14692 ;
  assign n14694 = n14693 ^ n13236 ;
  assign n14695 = ~n13222 & n14694 ;
  assign n14710 = n14709 ^ n14695 ;
  assign n14682 = n13251 ^ n13241 ;
  assign n14683 = n13241 ^ n13223 ;
  assign n14684 = n14683 ^ n13241 ;
  assign n14685 = ~n14682 & n14684 ;
  assign n14686 = n14685 ^ n13241 ;
  assign n14687 = n13281 & ~n14686 ;
  assign n14711 = n14710 ^ n14687 ;
  assign n14712 = n14681 & n14711 ;
  assign n14713 = n14712 ^ n9874 ;
  assign n14714 = n14713 ^ x121 ;
  assign n14778 = n14747 ^ n14714 ;
  assign n14779 = ~n14749 & ~n14778 ;
  assign n14780 = n14779 ^ n14747 ;
  assign n14748 = n13145 ^ x112 ;
  assign n14753 = n14748 ^ n14747 ;
  assign n14754 = n14753 ^ n14749 ;
  assign n14750 = n14749 ^ n14748 ;
  assign n14751 = ~n14747 & ~n14750 ;
  assign n14752 = n14751 ^ n14749 ;
  assign n14755 = n14754 ^ n14752 ;
  assign n14756 = ~n14714 & ~n14755 ;
  assign n14757 = n14749 ^ n14714 ;
  assign n14758 = n14749 ^ n14747 ;
  assign n14759 = n14758 ^ n14748 ;
  assign n14760 = n14759 ^ n14758 ;
  assign n14761 = n14758 ^ n14714 ;
  assign n14762 = n14761 ^ n14749 ;
  assign n14763 = n14760 & ~n14762 ;
  assign n14764 = n14763 ^ n14749 ;
  assign n14765 = n14749 & n14764 ;
  assign n14766 = n14757 & n14765 ;
  assign n14767 = n14766 ^ n14763 ;
  assign n14768 = n14767 ^ n14748 ;
  assign n14769 = n14768 ^ n14757 ;
  assign n14770 = ~n14756 & ~n14769 ;
  assign n14781 = n14780 ^ n14770 ;
  assign n14782 = n14781 ^ n14758 ;
  assign n14774 = n14748 ^ n14714 ;
  assign n14791 = n14782 ^ n14774 ;
  assign n14788 = n14753 ^ n14714 ;
  assign n14786 = n14779 ^ n14714 ;
  assign n14787 = n14750 & ~n14786 ;
  assign n14789 = n14788 ^ n14787 ;
  assign n14790 = n14789 ^ n14770 ;
  assign n14792 = n14791 ^ n14790 ;
  assign n14793 = n14792 ^ n14754 ;
  assign n14794 = n14793 ^ n14752 ;
  assign n14795 = n14794 ^ n14793 ;
  assign n14796 = n14793 ^ n14714 ;
  assign n14797 = n14796 ^ n14793 ;
  assign n14798 = n14795 & n14797 ;
  assign n14799 = n14798 ^ n14793 ;
  assign n14800 = n14680 & n14799 ;
  assign n14801 = n14800 ^ n14792 ;
  assign n14772 = ~n14714 & ~n14749 ;
  assign n14775 = ~n14772 & ~n14774 ;
  assign n14771 = n14770 ^ n14749 ;
  assign n14773 = n14772 ^ n14771 ;
  assign n14776 = n14775 ^ n14773 ;
  assign n14777 = n14680 & ~n14776 ;
  assign n14783 = n14782 ^ n14777 ;
  assign n14802 = n14801 ^ n14783 ;
  assign n14803 = n14784 & n14802 ;
  assign n14785 = n14784 ^ n14783 ;
  assign n14804 = n14803 ^ n14785 ;
  assign n14805 = n14804 ^ n9919 ;
  assign n15453 = n14805 ^ x92 ;
  assign n15456 = n13462 ^ n13457 ;
  assign n13494 = n13493 ^ n13458 ;
  assign n15457 = n15456 ^ n13494 ;
  assign n15458 = n15457 ^ n15455 ;
  assign n15459 = n13310 & n15458 ;
  assign n15454 = n13472 ^ n13457 ;
  assign n15460 = n15459 ^ n15454 ;
  assign n15485 = n15460 ^ n15297 ;
  assign n15486 = n15485 ^ n15484 ;
  assign n13536 = n13146 & n13535 ;
  assign n15487 = n15486 ^ n13536 ;
  assign n13540 = n13462 & n13539 ;
  assign n15488 = n15487 ^ n13540 ;
  assign n13501 = n13500 ^ n13480 ;
  assign n13502 = n13480 ^ n13310 ;
  assign n13503 = n13502 ^ n13480 ;
  assign n13504 = n13501 & n13503 ;
  assign n13505 = n13504 ^ n13480 ;
  assign n13506 = ~n13146 & ~n13505 ;
  assign n15489 = n15488 ^ n13506 ;
  assign n15490 = n15489 ^ n10388 ;
  assign n15470 = n15469 ^ n13481 ;
  assign n15468 = n13470 ^ n13456 ;
  assign n15471 = n15470 ^ n15468 ;
  assign n15472 = n15468 ^ n13310 ;
  assign n15473 = n15472 ^ n15468 ;
  assign n15474 = n15471 & n15473 ;
  assign n15475 = n15474 ^ n15468 ;
  assign n15476 = ~n13146 & n15475 ;
  assign n15491 = n15490 ^ n15476 ;
  assign n15461 = n15460 ^ n13498 ;
  assign n15462 = n15461 ^ n15460 ;
  assign n15465 = ~n13310 & n15462 ;
  assign n15466 = n15465 ^ n15460 ;
  assign n15467 = n15270 & ~n15466 ;
  assign n15492 = n15491 ^ n15467 ;
  assign n15493 = n15492 ^ x109 ;
  assign n15494 = ~n15453 & ~n15493 ;
  assign n15495 = n15494 ^ n15453 ;
  assign n14103 = n13934 & n14080 ;
  assign n15577 = n14103 ^ n14087 ;
  assign n15578 = ~n14094 & n15577 ;
  assign n15572 = n14110 ^ n14080 ;
  assign n14090 = n14089 ^ n14075 ;
  assign n14091 = n13968 & ~n14090 ;
  assign n14092 = n14091 ^ n14075 ;
  assign n15573 = n15572 ^ n14092 ;
  assign n15571 = n13968 & ~n14662 ;
  assign n15574 = n15573 ^ n15571 ;
  assign n15575 = ~n13934 & ~n15574 ;
  assign n14098 = n14097 ^ n14080 ;
  assign n14099 = ~n13934 & n14098 ;
  assign n14100 = n14099 ^ n14097 ;
  assign n14101 = n13968 & n14100 ;
  assign n14096 = ~n14094 & n14095 ;
  assign n14102 = n14101 ^ n14096 ;
  assign n15569 = n14102 ^ n10983 ;
  assign n15566 = n14092 ^ n14080 ;
  assign n15567 = n15566 ^ n14676 ;
  assign n15558 = n14122 ^ n13934 ;
  assign n15568 = n15567 ^ n15558 ;
  assign n15570 = n15569 ^ n15568 ;
  assign n15576 = n15575 ^ n15570 ;
  assign n15579 = n15578 ^ n15576 ;
  assign n15563 = n14642 ^ n13934 ;
  assign n15564 = n14113 ^ n14095 ;
  assign n15565 = n15563 & ~n15564 ;
  assign n15580 = n15579 ^ n15565 ;
  assign n15559 = n15558 ^ n14122 ;
  assign n15560 = n14137 & n15559 ;
  assign n15561 = n15560 ^ n14122 ;
  assign n15562 = n13968 & ~n15561 ;
  assign n15581 = n15580 ^ n15562 ;
  assign n14154 = n14085 ^ n13968 ;
  assign n15548 = n14642 ^ n14094 ;
  assign n15549 = n15548 ^ n14085 ;
  assign n15550 = n15549 ^ n14094 ;
  assign n15553 = ~n14154 & n15550 ;
  assign n15554 = n15553 ^ n14094 ;
  assign n15555 = n14111 & n15554 ;
  assign n15582 = n15581 ^ n15555 ;
  assign n15583 = n15582 ^ x68 ;
  assign n13822 = n13821 ^ n13807 ;
  assign n15584 = n13870 ^ n13577 ;
  assign n15585 = ~n13822 & n15584 ;
  assign n15586 = n15584 ^ n13576 ;
  assign n15587 = n13888 ^ n13878 ;
  assign n15588 = ~n15586 & n15587 ;
  assign n15605 = n13870 & ~n13876 ;
  assign n15595 = n13835 ^ n13577 ;
  assign n15598 = n13825 ^ n13810 ;
  assign n15599 = n15598 ^ n13835 ;
  assign n15600 = n15599 ^ n13888 ;
  assign n15601 = n13576 & n15600 ;
  assign n15596 = n13835 ^ n13815 ;
  assign n15597 = n15596 ^ n13825 ;
  assign n15602 = n15601 ^ n15597 ;
  assign n15603 = n15595 & ~n15602 ;
  assign n15604 = n15603 ^ n13577 ;
  assign n15606 = n15605 ^ n15604 ;
  assign n15589 = n13820 ^ n13814 ;
  assign n15590 = n15589 ^ n13810 ;
  assign n15591 = n15590 ^ n13823 ;
  assign n15592 = ~n13576 & n15591 ;
  assign n15593 = n15592 ^ n13820 ;
  assign n15594 = ~n13577 & ~n15593 ;
  assign n15607 = n15606 ^ n15594 ;
  assign n15608 = ~n13894 & ~n15607 ;
  assign n15609 = ~n15588 & n15608 ;
  assign n15610 = ~n15585 & n15609 ;
  assign n15611 = n13854 ^ n13576 ;
  assign n15612 = n15611 ^ n13854 ;
  assign n15613 = n13854 ^ n13839 ;
  assign n15614 = n15613 ^ n13854 ;
  assign n15615 = n15612 & n15614 ;
  assign n15616 = n15615 ^ n13854 ;
  assign n15617 = n13578 & n15616 ;
  assign n15618 = n15617 ^ n13854 ;
  assign n15619 = n15610 & ~n15618 ;
  assign n15626 = n15619 & ~n15625 ;
  assign n15627 = ~n13872 & n15626 ;
  assign n15628 = n15627 ^ n11416 ;
  assign n15629 = n15628 ^ x85 ;
  assign n15630 = ~n15583 & n15629 ;
  assign n15541 = n14341 & n14991 ;
  assign n15539 = n14323 & n14995 ;
  assign n15529 = n14362 ^ n14223 ;
  assign n15530 = n15529 ^ n14323 ;
  assign n15527 = n14274 ^ n14273 ;
  assign n15528 = n15527 ^ n14222 ;
  assign n15531 = n15530 ^ n15528 ;
  assign n15532 = n15531 ^ n14372 ;
  assign n15533 = ~n14344 & ~n15532 ;
  assign n15534 = n15533 ^ n14372 ;
  assign n15535 = n15022 ^ n14344 ;
  assign n15536 = n15534 & ~n15535 ;
  assign n15523 = n15022 ^ n14362 ;
  assign n15506 = n14375 ^ n14335 ;
  assign n15507 = n15506 ^ n14276 ;
  assign n15513 = n15507 ^ n14346 ;
  assign n15504 = n14348 ^ n14328 ;
  assign n15505 = n15504 ^ n14338 ;
  assign n15508 = n15507 ^ n15505 ;
  assign n15509 = n15505 ^ n14315 ;
  assign n15510 = ~n14372 & n15509 ;
  assign n15511 = n15510 ^ n14315 ;
  assign n15512 = ~n15508 & n15511 ;
  assign n15514 = n15513 ^ n15512 ;
  assign n15524 = n15523 ^ n15514 ;
  assign n15525 = n15524 ^ n11237 ;
  assign n14281 = n14280 ^ n14276 ;
  assign n14318 = n14281 & n14315 ;
  assign n14319 = n14318 ^ n14280 ;
  assign n14320 = n14167 & n14319 ;
  assign n15526 = n15525 ^ n14320 ;
  assign n15537 = n15536 ^ n15526 ;
  assign n15515 = n15514 ^ n14322 ;
  assign n15516 = n15515 ^ n14347 ;
  assign n15517 = n15516 ^ n15514 ;
  assign n15518 = n15514 ^ n14315 ;
  assign n15519 = n15518 ^ n15514 ;
  assign n15520 = ~n15517 & n15519 ;
  assign n15521 = n15520 ^ n15514 ;
  assign n15522 = ~n14372 & n15521 ;
  assign n15538 = n15537 ^ n15522 ;
  assign n15540 = n15539 ^ n15538 ;
  assign n15542 = n15541 ^ n15540 ;
  assign n15497 = n14362 ^ n14315 ;
  assign n15498 = n15497 ^ n14362 ;
  assign n15499 = n14362 ^ n14325 ;
  assign n15500 = n15499 ^ n14362 ;
  assign n15501 = ~n15498 & n15500 ;
  assign n15502 = n15501 ^ n14362 ;
  assign n15503 = n14167 & n15502 ;
  assign n15543 = n15542 ^ n15503 ;
  assign n15544 = n15543 ^ x70 ;
  assign n13054 = n13038 ^ n12630 ;
  assign n13053 = n13012 ^ n12122 ;
  assign n13055 = n13054 ^ n13053 ;
  assign n15136 = n13073 ^ n13055 ;
  assign n15134 = n13048 ^ n12630 ;
  assign n13039 = n13038 ^ n13033 ;
  assign n15135 = n15134 ^ n13039 ;
  assign n15137 = n15136 ^ n15135 ;
  assign n15138 = n13057 & n15137 ;
  assign n15127 = n13073 ^ n13039 ;
  assign n15124 = n13028 & n13057 ;
  assign n15126 = n15125 ^ n15124 ;
  assign n15128 = n15127 ^ n15126 ;
  assign n15121 = n13045 ^ n13033 ;
  assign n15122 = n15121 ^ n13073 ;
  assign n15123 = n13059 & n15122 ;
  assign n15129 = n15128 ^ n15123 ;
  assign n15113 = n13042 ^ n13039 ;
  assign n15114 = n15113 ^ n13010 ;
  assign n15115 = n15114 ^ n15113 ;
  assign n15116 = n15113 ^ n13047 ;
  assign n15117 = n15116 ^ n15113 ;
  assign n15118 = ~n15115 & n15117 ;
  assign n15119 = n15118 ^ n15113 ;
  assign n15120 = ~n12827 & ~n15119 ;
  assign n15130 = n15129 ^ n15120 ;
  assign n15131 = n15130 ^ n13055 ;
  assign n13091 = ~n13010 & ~n13032 ;
  assign n13092 = n13091 ^ n13027 ;
  assign n13077 = n13076 ^ n13072 ;
  assign n13078 = n13077 ^ n13045 ;
  assign n13093 = n13092 ^ n13078 ;
  assign n13094 = n13093 ^ n13092 ;
  assign n13095 = n13092 ^ n12827 ;
  assign n13096 = n13095 ^ n13092 ;
  assign n13097 = n13094 & n13096 ;
  assign n13098 = n13097 ^ n13092 ;
  assign n13099 = n13019 & n13098 ;
  assign n13100 = n13099 ^ n13092 ;
  assign n15132 = n15131 ^ n13100 ;
  assign n15133 = n15132 ^ n10738 ;
  assign n15139 = n15138 ^ n15133 ;
  assign n15106 = n13021 ^ n12827 ;
  assign n15107 = n15106 ^ n13021 ;
  assign n15108 = n13054 ^ n13020 ;
  assign n15109 = n15108 ^ n13021 ;
  assign n15110 = ~n15107 & ~n15109 ;
  assign n15111 = n15110 ^ n13021 ;
  assign n15112 = n13010 & n15111 ;
  assign n15140 = n15139 ^ n15112 ;
  assign n15545 = n15140 ^ x110 ;
  assign n15546 = ~n15544 & n15545 ;
  assign n15547 = n15546 ^ n15544 ;
  assign n15644 = n15547 ^ n15545 ;
  assign n15645 = n15630 & n15644 ;
  assign n15639 = n15630 ^ n15583 ;
  assign n15640 = ~n15547 & ~n15639 ;
  assign n15641 = n15640 ^ n15547 ;
  assign n15632 = n15630 ^ n15629 ;
  assign n15633 = n15632 ^ n15583 ;
  assign n15634 = ~n15547 & n15633 ;
  assign n15631 = ~n15547 & n15630 ;
  assign n15635 = n15634 ^ n15631 ;
  assign n15642 = n15641 ^ n15635 ;
  assign n15646 = n15645 ^ n15642 ;
  assign n15647 = n15646 ^ n15634 ;
  assign n15648 = n15647 ^ n15640 ;
  assign n15637 = n15629 ^ n15544 ;
  assign n15638 = ~n15545 & ~n15637 ;
  assign n15643 = n15642 ^ n15638 ;
  assign n15649 = n15648 ^ n15643 ;
  assign n15660 = n15649 ^ n15642 ;
  assign n15652 = n15546 ^ n15545 ;
  assign n15654 = n15632 & n15652 ;
  assign n15659 = n15654 ^ n15632 ;
  assign n15661 = n15660 ^ n15659 ;
  assign n15656 = n15546 & n15630 ;
  assign n15685 = n15661 ^ n15656 ;
  assign n15668 = n15546 & n15633 ;
  assign n15684 = n15668 ^ n15546 ;
  assign n15686 = n15685 ^ n15684 ;
  assign n17122 = ~n15495 & ~n15686 ;
  assign n15496 = n15495 ^ n15493 ;
  assign n15653 = ~n15639 & n15652 ;
  assign n17119 = n15661 ^ n15653 ;
  assign n17120 = ~n15496 & ~n17119 ;
  assign n15683 = n15493 ^ n15453 ;
  assign n15662 = n15649 ^ n15646 ;
  assign n15663 = n15662 ^ n15631 ;
  assign n15664 = n15663 ^ n15661 ;
  assign n15657 = n15656 ^ n15654 ;
  assign n15658 = n15657 ^ n15629 ;
  assign n15665 = n15664 ^ n15658 ;
  assign n15666 = n15665 ^ n15652 ;
  assign n15655 = n15654 ^ n15653 ;
  assign n15667 = n15666 ^ n15655 ;
  assign n15669 = n15668 ^ n15667 ;
  assign n15670 = n15669 ^ n15633 ;
  assign n15671 = n15670 ^ n15648 ;
  assign n15672 = n15671 ^ n15645 ;
  assign n15651 = n15642 ^ n15640 ;
  assign n15673 = n15672 ^ n15651 ;
  assign n17104 = n15673 ^ n15665 ;
  assign n17106 = n17104 ^ n15660 ;
  assign n17105 = n17104 ^ n15673 ;
  assign n17107 = n17106 ^ n17105 ;
  assign n17108 = n17106 ^ n15493 ;
  assign n17109 = n17108 ^ n17106 ;
  assign n17110 = ~n17107 & n17109 ;
  assign n17111 = n17110 ^ n17106 ;
  assign n17112 = n15683 & ~n17111 ;
  assign n17113 = n17112 ^ n17104 ;
  assign n17095 = n15644 ^ n15631 ;
  assign n17096 = n17095 ^ n15672 ;
  assign n17097 = ~n15453 & ~n17096 ;
  assign n17098 = n17097 ^ n15648 ;
  assign n17114 = n17113 ^ n17098 ;
  assign n15674 = n15673 ^ n15660 ;
  assign n15675 = n15674 ^ n15644 ;
  assign n15676 = n15675 ^ n15646 ;
  assign n15694 = n15496 ^ n15453 ;
  assign n16304 = n15676 & ~n15694 ;
  assign n17115 = n17114 ^ n16304 ;
  assign n15713 = n15668 ^ n15653 ;
  assign n15733 = n15713 ^ n15657 ;
  assign n15734 = n15657 ^ n15493 ;
  assign n15735 = n15734 ^ n15657 ;
  assign n15736 = n15733 & ~n15735 ;
  assign n15737 = n15736 ^ n15657 ;
  assign n15738 = ~n15453 & n15737 ;
  assign n17116 = n17115 ^ n15738 ;
  assign n17117 = n17116 ^ n14221 ;
  assign n17100 = n15673 ^ n15667 ;
  assign n17099 = n17098 ^ n15638 ;
  assign n17101 = n17100 ^ n17099 ;
  assign n17091 = n15632 ^ n15546 ;
  assign n17092 = n17091 ^ n15648 ;
  assign n17093 = n17092 ^ n15667 ;
  assign n17094 = n15453 & ~n17093 ;
  assign n17102 = n17101 ^ n17094 ;
  assign n17103 = ~n15493 & ~n17102 ;
  assign n17118 = n17117 ^ n17103 ;
  assign n17121 = n17120 ^ n17118 ;
  assign n17123 = n17122 ^ n17121 ;
  assign n17496 = n17123 ^ x82 ;
  assign n17497 = n17495 & n17496 ;
  assign n13101 = n13100 ^ n11545 ;
  assign n13016 = n13015 ^ n13012 ;
  assign n13017 = n13010 & n13016 ;
  assign n12828 = n12630 & ~n12827 ;
  assign n13018 = n13017 ^ n12828 ;
  assign n13087 = n13074 ^ n13030 ;
  assign n13088 = n13056 & n13087 ;
  assign n13060 = ~n13055 & n13059 ;
  assign n13065 = n13060 ^ n13047 ;
  assign n13052 = n13051 ^ n13049 ;
  assign n13061 = n13060 ^ n13052 ;
  assign n13022 = n13021 ^ n12630 ;
  assign n13040 = n13039 ^ n13022 ;
  assign n13062 = n13061 ^ n13040 ;
  assign n13063 = ~n13010 & ~n13062 ;
  assign n13064 = n13063 ^ n13061 ;
  assign n13066 = n13065 ^ n13064 ;
  assign n13067 = n13066 ^ n13010 ;
  assign n13068 = n13067 ^ n13066 ;
  assign n13069 = n13066 ^ n13047 ;
  assign n13070 = n13069 ^ n13066 ;
  assign n13079 = n13078 ^ n13066 ;
  assign n13080 = n13079 ^ n13066 ;
  assign n13081 = ~n13070 & n13080 ;
  assign n13082 = ~n13068 & n13081 ;
  assign n13083 = n13082 ^ n13068 ;
  assign n13084 = n13083 ^ n13067 ;
  assign n13085 = ~n13019 & n13084 ;
  assign n13086 = n13085 ^ n13064 ;
  assign n13089 = n13088 ^ n13086 ;
  assign n13090 = ~n13018 & ~n13089 ;
  assign n13102 = n13101 ^ n13090 ;
  assign n13103 = n13102 ^ x106 ;
  assign n13544 = ~n13487 & n13539 ;
  assign n13523 = n13477 ^ n13383 ;
  assign n13524 = n13477 ^ n13350 ;
  assign n13525 = n13524 ^ n13453 ;
  assign n13526 = n13311 & n13525 ;
  assign n13527 = ~n13523 & n13526 ;
  assign n13528 = n13527 ^ n13472 ;
  assign n13517 = n13474 ^ n13471 ;
  assign n13518 = n13471 ^ n13146 ;
  assign n13519 = n13518 ^ n13471 ;
  assign n13520 = n13517 & n13519 ;
  assign n13521 = n13520 ^ n13471 ;
  assign n13522 = n13310 & ~n13521 ;
  assign n13529 = n13528 ^ n13522 ;
  assign n13537 = n13536 ^ n13529 ;
  assign n13508 = n13507 ^ n13472 ;
  assign n13510 = n13509 ^ n13492 ;
  assign n13511 = n13510 ^ n13311 ;
  assign n13514 = ~n13507 & n13511 ;
  assign n13515 = n13514 ^ n13311 ;
  assign n13516 = n13508 & ~n13515 ;
  assign n13538 = n13537 ^ n13516 ;
  assign n13541 = n13540 ^ n13538 ;
  assign n13542 = n13541 ^ n13506 ;
  assign n13543 = n13542 ^ n12399 ;
  assign n13545 = n13544 ^ n13543 ;
  assign n13495 = n13494 ^ n13465 ;
  assign n13496 = n13495 ^ n13469 ;
  assign n13497 = n13312 & n13496 ;
  assign n13546 = n13545 ^ n13497 ;
  assign n13547 = n13546 ^ x97 ;
  assign n13548 = n13103 & n13547 ;
  assign n13549 = n13548 ^ n13103 ;
  assign n13895 = n13894 ^ n12870 ;
  assign n13855 = n13854 ^ n13819 ;
  assign n13856 = n13855 ^ n13815 ;
  assign n13857 = n13856 ^ n13800 ;
  assign n13858 = n13800 ^ n13577 ;
  assign n13859 = n13858 ^ n13800 ;
  assign n13860 = ~n13857 & ~n13859 ;
  assign n13861 = n13860 ^ n13800 ;
  assign n13862 = ~n13576 & n13861 ;
  assign n13863 = n13862 ^ n13841 ;
  assign n13852 = n13578 & n13837 ;
  assign n13864 = n13863 ^ n13852 ;
  assign n13842 = n13841 ^ n13577 ;
  assign n13843 = n13842 ^ n13841 ;
  assign n13849 = n13843 & n13846 ;
  assign n13850 = n13849 ^ n13841 ;
  assign n13851 = n13576 & ~n13850 ;
  assign n13865 = n13864 ^ n13851 ;
  assign n13827 = n13826 ^ n13823 ;
  assign n13866 = n13865 ^ n13827 ;
  assign n13828 = n13827 ^ n13822 ;
  assign n13829 = n13828 ^ n13827 ;
  assign n13830 = n13827 ^ n13576 ;
  assign n13831 = n13830 ^ n13827 ;
  assign n13832 = ~n13829 & n13831 ;
  assign n13833 = n13832 ^ n13827 ;
  assign n13834 = n13578 & n13833 ;
  assign n13867 = n13866 ^ n13834 ;
  assign n13886 = n13867 & ~n13885 ;
  assign n13896 = n13895 ^ n13886 ;
  assign n13897 = n13896 ^ x123 ;
  assign n14093 = n13934 & n14092 ;
  assign n14114 = n14113 ^ n14080 ;
  assign n14115 = n14114 ^ n14100 ;
  assign n14116 = n14115 ^ n14103 ;
  assign n14117 = n14094 & ~n14116 ;
  assign n14118 = n14117 ^ n14113 ;
  assign n14125 = n14124 ^ n14109 ;
  assign n14126 = n14125 ^ n14085 ;
  assign n14129 = n14111 ^ n13934 ;
  assign n14130 = n14129 ^ n14111 ;
  assign n14131 = ~n14126 & n14130 ;
  assign n14132 = n14131 ^ n14111 ;
  assign n14133 = ~n13968 & ~n14132 ;
  assign n14146 = n14145 ^ n14133 ;
  assign n14136 = n14089 ^ n14081 ;
  assign n14138 = n14137 ^ n14136 ;
  assign n14139 = ~n13934 & ~n14138 ;
  assign n14147 = n14146 ^ n14139 ;
  assign n14134 = n14082 ^ n14075 ;
  assign n14135 = n14134 ^ n14109 ;
  assign n14148 = n14147 ^ n14135 ;
  assign n14149 = n14148 ^ n14133 ;
  assign n14150 = ~n14094 & n14149 ;
  assign n14151 = n14150 ^ n14147 ;
  assign n14155 = n14154 ^ n14085 ;
  assign n14156 = n14106 & n14155 ;
  assign n14157 = n14156 ^ n14085 ;
  assign n14158 = ~n13934 & n14157 ;
  assign n14159 = ~n14151 & ~n14158 ;
  assign n14160 = n14118 & n14159 ;
  assign n14161 = ~n14102 & n14160 ;
  assign n14162 = ~n14093 & n14161 ;
  assign n14163 = n14162 ^ n12899 ;
  assign n14164 = n14163 ^ x80 ;
  assign n14165 = n13897 & n14164 ;
  assign n14166 = n14165 ^ n13897 ;
  assign n14387 = n13452 ^ x108 ;
  assign n14390 = n13575 ^ x84 ;
  assign n14417 = n12337 ^ n12277 ;
  assign n14418 = ~n12169 & n14417 ;
  assign n14394 = ~n12169 & ~n12308 ;
  assign n14395 = n14394 ^ n12284 ;
  assign n14416 = n14395 ^ n12275 ;
  assign n14419 = n14418 ^ n14416 ;
  assign n14420 = n12170 & n14419 ;
  assign n14414 = n12172 & n12269 ;
  assign n14400 = n14399 ^ n12338 ;
  assign n14397 = n12303 ^ n12288 ;
  assign n14398 = n14397 ^ n12301 ;
  assign n14401 = n14400 ^ n14398 ;
  assign n14402 = n12170 & n14401 ;
  assign n14403 = n14402 ^ n14400 ;
  assign n14405 = n14403 ^ n12286 ;
  assign n14406 = n14405 ^ n12302 ;
  assign n14408 = n14407 ^ n14406 ;
  assign n14409 = n14408 ^ n14403 ;
  assign n14410 = n12170 & ~n14409 ;
  assign n14411 = n14410 ^ n14405 ;
  assign n14412 = n12169 & n14411 ;
  assign n14396 = n14395 ^ n12350 ;
  assign n14404 = n14403 ^ n14396 ;
  assign n14413 = n14412 ^ n14404 ;
  assign n14415 = n14414 ^ n14413 ;
  assign n14421 = n14420 ^ n14415 ;
  assign n14422 = n14421 ^ n14391 ;
  assign n14392 = n14391 ^ n14048 ;
  assign n14393 = n12169 & n14392 ;
  assign n14423 = n14422 ^ n14393 ;
  assign n14424 = ~n12315 & ~n14039 ;
  assign n14425 = ~n14423 & n14424 ;
  assign n14426 = n14425 ^ n11709 ;
  assign n14427 = n14426 ^ x101 ;
  assign n14428 = ~n14390 & n14427 ;
  assign n14429 = n14428 ^ n14427 ;
  assign n14448 = n12012 & ~n12111 ;
  assign n14443 = n13334 ^ n12086 ;
  assign n14438 = n12056 ^ n12033 ;
  assign n14439 = n14438 ^ n12019 ;
  assign n14440 = ~n12111 & ~n14439 ;
  assign n14441 = n14440 ^ n12020 ;
  assign n14442 = ~n11546 & ~n14441 ;
  assign n14444 = n14443 ^ n14442 ;
  assign n14437 = ~n12054 & n12071 ;
  assign n14445 = n14444 ^ n14437 ;
  assign n14433 = n12055 ^ n12039 ;
  assign n14434 = n14433 ^ n12023 ;
  assign n14435 = n14434 ^ n12046 ;
  assign n14436 = n11582 & ~n14435 ;
  assign n14446 = n14445 ^ n14436 ;
  assign n14430 = n12049 ^ n11828 ;
  assign n14431 = n14430 ^ n12053 ;
  assign n14432 = n11583 & ~n14431 ;
  assign n14447 = n14446 ^ n14432 ;
  assign n14449 = n14448 ^ n14447 ;
  assign n14450 = ~n13970 & ~n14449 ;
  assign n14451 = n14450 ^ n11734 ;
  assign n14452 = n14451 ^ x86 ;
  assign n14453 = n13309 ^ x126 ;
  assign n14454 = ~n14452 & ~n14453 ;
  assign n14456 = n14454 ^ n14453 ;
  assign n14476 = n14456 ^ n14452 ;
  assign n14487 = n14429 & ~n14476 ;
  assign n14492 = n14487 ^ n14476 ;
  assign n14461 = n14429 ^ n14390 ;
  assign n14478 = n14461 & ~n14476 ;
  assign n14477 = n14428 & ~n14476 ;
  assign n14479 = n14478 ^ n14477 ;
  assign n14493 = n14492 ^ n14479 ;
  assign n14457 = n14428 ^ n14390 ;
  assign n14525 = n14493 ^ n14457 ;
  assign n14482 = n14454 & ~n14457 ;
  assign n14458 = ~n14456 & ~n14457 ;
  assign n14524 = n14482 ^ n14458 ;
  assign n14526 = n14525 ^ n14524 ;
  assign n14527 = n14526 ^ n14479 ;
  assign n14534 = n14527 ^ n14453 ;
  assign n14490 = n14487 ^ n14429 ;
  assign n14462 = ~n14456 & n14461 ;
  assign n14460 = n14428 & ~n14456 ;
  assign n14463 = n14462 ^ n14460 ;
  assign n14459 = n14458 ^ n14456 ;
  assign n14464 = n14463 ^ n14459 ;
  assign n14455 = n14429 & n14454 ;
  assign n14465 = n14464 ^ n14455 ;
  assign n14491 = n14490 ^ n14465 ;
  assign n14494 = n14493 ^ n14491 ;
  assign n14485 = n14476 ^ n14453 ;
  assign n14486 = n14428 & ~n14485 ;
  assign n14488 = n14487 ^ n14486 ;
  assign n14533 = n14494 ^ n14488 ;
  assign n14535 = n14534 ^ n14533 ;
  assign n14536 = n14387 & n14535 ;
  assign n14388 = n13748 ^ x125 ;
  assign n14389 = ~n14387 & n14388 ;
  assign n14518 = n14494 ^ n14478 ;
  assign n14519 = n14518 ^ n14486 ;
  assign n14520 = n14389 & n14519 ;
  assign n14511 = n14389 ^ n14387 ;
  assign n14521 = n14520 ^ n14511 ;
  assign n14528 = n14527 ^ n14491 ;
  assign n14522 = n14493 ^ n14486 ;
  assign n14523 = n14389 & ~n14522 ;
  assign n14529 = n14528 ^ n14523 ;
  assign n14530 = ~n14521 & ~n14529 ;
  assign n14512 = n14482 ^ n14462 ;
  assign n14513 = ~n14511 & n14512 ;
  assign n14467 = n14388 ^ n14387 ;
  assign n14500 = n14487 ^ n14460 ;
  assign n14501 = n14500 ^ n14388 ;
  assign n14502 = n14501 ^ n14500 ;
  assign n14470 = n14428 & n14454 ;
  assign n14481 = n14470 ^ n14455 ;
  assign n14483 = n14482 ^ n14481 ;
  assign n14503 = n14483 ^ n14454 ;
  assign n14504 = n14503 ^ n14487 ;
  assign n14505 = n14504 ^ n14500 ;
  assign n14506 = ~n14502 & n14505 ;
  assign n14507 = n14506 ^ n14500 ;
  assign n14508 = n14467 & n14507 ;
  assign n14509 = n14508 ^ n14487 ;
  assign n14510 = n14509 ^ n14458 ;
  assign n14514 = n14513 ^ n14510 ;
  assign n14515 = n14514 ^ n11825 ;
  assign n14489 = n14488 ^ n14460 ;
  assign n14495 = n14494 ^ n14489 ;
  assign n14480 = n14479 ^ n14462 ;
  assign n14484 = n14483 ^ n14480 ;
  assign n14496 = n14495 ^ n14484 ;
  assign n14497 = n14388 & n14496 ;
  assign n14498 = n14497 ^ n14495 ;
  assign n14499 = n14387 & n14498 ;
  assign n14516 = n14515 ^ n14499 ;
  assign n14468 = n14458 ^ n14388 ;
  assign n14469 = n14468 ^ n14458 ;
  assign n14473 = ~n14469 & n14470 ;
  assign n14474 = n14473 ^ n14458 ;
  assign n14475 = ~n14467 & n14474 ;
  assign n14517 = n14516 ^ n14475 ;
  assign n14531 = n14530 ^ n14517 ;
  assign n14466 = n14389 & ~n14465 ;
  assign n14532 = n14531 ^ n14466 ;
  assign n14537 = n14536 ^ n14532 ;
  assign n14538 = n14537 ^ x82 ;
  assign n14366 = n14347 ^ n14328 ;
  assign n14364 = n14344 ^ n14327 ;
  assign n14365 = n14364 ^ n14341 ;
  assign n14367 = n14366 ^ n14365 ;
  assign n14368 = n14315 & ~n14367 ;
  assign n14369 = n14368 ^ n14365 ;
  assign n14379 = n14369 ^ n14362 ;
  assign n14377 = n14376 ^ n14324 ;
  assign n14378 = ~n14315 & n14377 ;
  assign n14380 = n14379 ^ n14378 ;
  assign n14373 = n14346 ^ n14333 ;
  assign n14374 = n14167 & n14373 ;
  assign n14381 = n14380 ^ n14374 ;
  assign n14382 = ~n14372 & n14381 ;
  assign n14363 = n14362 ^ n14360 ;
  assign n14370 = n14369 ^ n14363 ;
  assign n14371 = n14370 ^ n14320 ;
  assign n14383 = n14382 ^ n14371 ;
  assign n14384 = n14383 ^ n14335 ;
  assign n14385 = n14384 ^ n12468 ;
  assign n14386 = n14385 ^ x120 ;
  assign n14540 = n14538 ^ n14386 ;
  assign n14539 = n14386 & n14538 ;
  assign n14541 = n14540 ^ n14539 ;
  assign n14542 = n14541 ^ n14538 ;
  assign n14543 = n14166 & n14542 ;
  assign n14544 = n13549 & n14543 ;
  assign n17548 = n14544 ^ n14189 ;
  assign n14545 = n13548 ^ n13547 ;
  assign n14546 = n14545 ^ n13103 ;
  assign n14548 = n14166 ^ n14164 ;
  assign n14549 = n14548 ^ n13897 ;
  assign n14566 = ~n14546 & n14549 ;
  assign n14552 = n14166 & n14545 ;
  assign n14550 = n14545 & n14549 ;
  assign n14562 = n14552 ^ n14550 ;
  assign n14553 = n14165 & n14545 ;
  assign n14561 = n14553 ^ n14545 ;
  assign n14563 = n14562 ^ n14561 ;
  assign n14547 = n14166 & ~n14546 ;
  assign n14564 = n14563 ^ n14547 ;
  assign n17501 = n14566 ^ n14564 ;
  assign n17502 = n14538 & n17501 ;
  assign n17503 = n17502 ^ n14566 ;
  assign n14556 = n13549 & n14165 ;
  assign n14555 = n13548 & n14165 ;
  assign n14557 = n14556 ^ n14555 ;
  assign n14554 = n14553 ^ n14165 ;
  assign n14558 = n14557 ^ n14554 ;
  assign n14567 = n14563 ^ n14558 ;
  assign n14568 = n14567 ^ n14566 ;
  assign n14565 = n14564 ^ n14546 ;
  assign n14569 = n14568 ^ n14565 ;
  assign n17506 = n17503 ^ n14569 ;
  assign n17507 = n17506 ^ n17503 ;
  assign n17508 = ~n14538 & ~n17507 ;
  assign n17509 = n17508 ^ n17503 ;
  assign n17510 = n14386 & n17509 ;
  assign n17511 = n17510 ^ n17503 ;
  assign n14551 = n14550 ^ n14547 ;
  assign n17537 = n14553 ^ n14551 ;
  assign n17538 = n17537 ^ n14563 ;
  assign n14575 = n13548 & ~n14548 ;
  assign n14578 = n14575 ^ n14556 ;
  assign n17535 = n14578 ^ n14553 ;
  assign n14581 = n13549 & ~n14548 ;
  assign n14570 = n13548 & n14166 ;
  assign n17534 = n14581 ^ n14570 ;
  assign n17536 = n17535 ^ n17534 ;
  assign n17539 = n17538 ^ n17536 ;
  assign n17540 = n17536 ^ n14538 ;
  assign n17541 = n17540 ^ n17536 ;
  assign n17542 = n17539 & ~n17541 ;
  assign n17543 = n17542 ^ n17536 ;
  assign n17544 = n14386 & n17543 ;
  assign n14571 = n13549 & n14549 ;
  assign n14572 = n14571 ^ n14570 ;
  assign n14573 = n14572 ^ n14555 ;
  assign n14582 = n14581 ^ n14573 ;
  assign n14576 = n14575 ^ n14571 ;
  assign n14574 = n14573 ^ n13548 ;
  assign n14577 = n14576 ^ n14574 ;
  assign n14579 = n14578 ^ n14577 ;
  assign n14580 = n14579 ^ n13103 ;
  assign n14583 = n14582 ^ n14580 ;
  assign n14584 = n14583 ^ n14555 ;
  assign n14585 = n14584 ^ n14569 ;
  assign n17521 = n14585 ^ n14575 ;
  assign n17519 = n14569 ^ n14557 ;
  assign n14614 = n14581 ^ n14577 ;
  assign n17520 = n17519 ^ n14614 ;
  assign n17522 = n17521 ^ n17520 ;
  assign n17523 = n14538 & n17522 ;
  assign n17524 = n17523 ^ n17521 ;
  assign n17525 = ~n14386 & ~n17524 ;
  assign n17526 = n17525 ^ n14566 ;
  assign n17512 = n14566 ^ n14386 ;
  assign n17513 = n17512 ^ n14566 ;
  assign n17516 = n14578 & n17513 ;
  assign n17517 = n17516 ^ n14566 ;
  assign n17518 = ~n14538 & n17517 ;
  assign n17527 = n17526 ^ n17518 ;
  assign n17529 = ~n14540 & n14562 ;
  assign n17530 = ~n17527 & n17529 ;
  assign n17531 = n17530 ^ n17527 ;
  assign n17545 = n17544 ^ n17531 ;
  assign n17528 = n17527 ^ n14541 ;
  assign n17533 = n14558 & ~n17528 ;
  assign n17546 = n17545 ^ n17533 ;
  assign n17547 = ~n17511 & ~n17546 ;
  assign n17549 = n17548 ^ n17547 ;
  assign n17550 = n17549 ^ x96 ;
  assign n15031 = n15030 ^ x77 ;
  assign n15081 = n14482 ^ n14477 ;
  assign n15082 = n15081 ^ n14491 ;
  assign n15036 = n14535 ^ n14493 ;
  assign n15072 = n15036 ^ n14487 ;
  assign n15071 = n14483 ^ n14478 ;
  assign n15073 = n15072 ^ n15071 ;
  assign n15069 = n14526 ^ n14458 ;
  assign n15070 = n15069 ^ n14491 ;
  assign n15074 = n15073 ^ n15070 ;
  assign n15075 = n14388 & n15074 ;
  assign n15076 = n15075 ^ n15073 ;
  assign n15083 = n15082 ^ n15076 ;
  assign n15084 = n14387 & n15083 ;
  assign n15062 = n14503 ^ n14470 ;
  assign n15063 = n14470 ^ n14388 ;
  assign n15064 = n15063 ^ n14470 ;
  assign n15065 = n15062 & n15064 ;
  assign n15066 = n15065 ^ n14470 ;
  assign n15067 = n14467 & n15066 ;
  assign n15053 = n14464 ^ n14463 ;
  assign n15054 = n15053 ^ n14388 ;
  assign n15055 = n15054 ^ n15053 ;
  assign n15056 = n14503 ^ n14463 ;
  assign n15057 = n15056 ^ n15053 ;
  assign n15058 = n15055 & ~n15057 ;
  assign n15059 = n15058 ^ n15053 ;
  assign n15060 = ~n14467 & ~n15059 ;
  assign n15061 = n15060 ^ n14463 ;
  assign n15068 = n15067 ^ n15061 ;
  assign n15077 = n15076 ^ n15068 ;
  assign n15043 = n14388 & n14533 ;
  assign n15044 = n15043 ^ n14494 ;
  assign n15045 = n15044 ^ n14463 ;
  assign n15046 = n15045 ^ n15044 ;
  assign n15049 = n14388 & n15046 ;
  assign n15050 = n15049 ^ n15044 ;
  assign n15051 = ~n14467 & n15050 ;
  assign n15052 = n15051 ^ n15044 ;
  assign n15078 = n15077 ^ n15052 ;
  assign n15037 = n15036 ^ n14526 ;
  assign n15038 = n14526 ^ n14388 ;
  assign n15039 = n15038 ^ n14526 ;
  assign n15040 = ~n15037 & n15039 ;
  assign n15041 = n15040 ^ n14526 ;
  assign n15042 = n14387 & n15041 ;
  assign n15079 = n15078 ^ n15042 ;
  assign n15080 = n15079 ^ n13618 ;
  assign n15085 = n15084 ^ n15080 ;
  assign n15032 = n14511 ^ n14388 ;
  assign n15033 = n14491 ^ n14482 ;
  assign n15034 = n15033 ^ n14535 ;
  assign n15035 = n15032 & ~n15034 ;
  assign n15086 = n15085 ^ n15035 ;
  assign n15087 = n15086 ^ x67 ;
  assign n15088 = n15031 & n15087 ;
  assign n14806 = n14805 ^ x117 ;
  assign n14906 = ~n14899 & ~n14905 ;
  assign n14907 = n14906 ^ n14898 ;
  assign n14908 = n14893 ^ n14842 ;
  assign n14909 = n14810 & n14908 ;
  assign n14969 = n14810 & n14902 ;
  assign n14961 = n14903 ^ n14809 ;
  assign n14962 = n14961 ^ n14929 ;
  assign n14963 = n14962 ^ n14960 ;
  assign n14964 = n14811 & ~n14963 ;
  assign n14965 = n14964 ^ n14809 ;
  assign n14966 = n14927 ^ n14811 ;
  assign n14967 = ~n14965 & n14966 ;
  assign n14955 = n14914 ^ n14894 ;
  assign n14956 = n14955 ^ n14889 ;
  assign n14957 = n14809 & n14956 ;
  assign n14949 = n14929 ^ n14895 ;
  assign n14950 = ~n14899 & ~n14949 ;
  assign n14951 = n14950 ^ n14948 ;
  assign n14952 = n14951 ^ n14947 ;
  assign n14953 = n14952 ^ n14935 ;
  assign n14911 = n14897 ^ n14891 ;
  assign n14919 = n14918 ^ n14911 ;
  assign n14920 = n14918 ^ n14807 ;
  assign n14921 = n14920 ^ n14918 ;
  assign n14922 = n14919 & ~n14921 ;
  assign n14923 = n14922 ^ n14918 ;
  assign n14924 = ~n14910 & ~n14923 ;
  assign n14954 = n14953 ^ n14924 ;
  assign n14958 = n14957 ^ n14954 ;
  assign n14959 = n14958 ^ n14927 ;
  assign n14968 = n14967 ^ n14959 ;
  assign n14970 = n14969 ^ n14968 ;
  assign n14977 = ~n14970 & ~n14976 ;
  assign n14978 = n14893 ^ n14892 ;
  assign n14979 = n14978 ^ n14892 ;
  assign n14980 = n14892 ^ n14808 ;
  assign n14981 = n14980 ^ n14892 ;
  assign n14982 = n14979 & n14981 ;
  assign n14983 = n14982 ^ n14892 ;
  assign n14984 = ~n14807 & n14983 ;
  assign n14985 = n14977 & ~n14984 ;
  assign n14986 = ~n14909 & n14985 ;
  assign n14987 = ~n14907 & n14986 ;
  assign n14988 = n14987 ^ n13645 ;
  assign n14989 = n14988 ^ x84 ;
  assign n14990 = n14806 & ~n14989 ;
  assign n15093 = n14990 ^ n14806 ;
  assign n15094 = n15093 ^ n14989 ;
  assign n15151 = n15088 & n15094 ;
  assign n14679 = n14678 ^ x102 ;
  assign n15141 = n15140 ^ x116 ;
  assign n15178 = n14679 & ~n15141 ;
  assign n15207 = n15178 ^ n14679 ;
  assign n15208 = n15207 ^ n15141 ;
  assign n15209 = n15151 & n15208 ;
  assign n15095 = n15094 ^ n14806 ;
  assign n15096 = n15088 & ~n15095 ;
  assign n15089 = n15088 ^ n15087 ;
  assign n15090 = n15089 ^ n15031 ;
  assign n15091 = n15090 ^ n15087 ;
  assign n15092 = n14990 & n15091 ;
  assign n15217 = n15096 ^ n15092 ;
  assign n15218 = n15208 & n15217 ;
  assign n15156 = n14990 & n15089 ;
  assign n15099 = n15089 & ~n15095 ;
  assign n15164 = n15156 ^ n15099 ;
  assign n15212 = n15156 ^ n14679 ;
  assign n15213 = n15212 ^ n15156 ;
  assign n15214 = n15164 & n15213 ;
  assign n15215 = n15214 ^ n15156 ;
  assign n15216 = ~n15141 & n15215 ;
  assign n15219 = n15218 ^ n15216 ;
  assign n17551 = ~n15209 & ~n15219 ;
  assign n15102 = n15091 & n15093 ;
  assign n15098 = ~n15090 & ~n15095 ;
  assign n15100 = n15099 ^ n15098 ;
  assign n15097 = n15096 ^ n15095 ;
  assign n15101 = n15100 ^ n15097 ;
  assign n15103 = n15102 ^ n15101 ;
  assign n15104 = n15103 ^ n15092 ;
  assign n15105 = n15104 ^ n15091 ;
  assign n15142 = n15141 ^ n15105 ;
  assign n15143 = n15142 ^ n15105 ;
  assign n15144 = ~n15090 & n15094 ;
  assign n15147 = ~n15143 & n15144 ;
  assign n15148 = n15147 ^ n15105 ;
  assign n15149 = ~n14679 & ~n15148 ;
  assign n15150 = n15149 ^ n15105 ;
  assign n17562 = n15156 ^ n15151 ;
  assign n15145 = n15144 ^ n15105 ;
  assign n15153 = n15145 ^ n15094 ;
  assign n15154 = n15153 ^ n15151 ;
  assign n15163 = n15154 ^ n15089 ;
  assign n15165 = n15164 ^ n15163 ;
  assign n15166 = n15165 ^ n15144 ;
  assign n15162 = ~n15090 & n15093 ;
  assign n15167 = n15166 ^ n15162 ;
  assign n15168 = n15167 ^ n15098 ;
  assign n15159 = n15156 ^ n15098 ;
  assign n15160 = n15159 ^ n15102 ;
  assign n15161 = n15160 ^ n15144 ;
  assign n15169 = n15168 ^ n15161 ;
  assign n15157 = n15156 ^ n14990 ;
  assign n15158 = n15157 ^ n14806 ;
  assign n15170 = n15169 ^ n15158 ;
  assign n17563 = n17562 ^ n15170 ;
  assign n17564 = n17563 ^ n15104 ;
  assign n17565 = n17564 ^ n15156 ;
  assign n17566 = n17565 ^ n17563 ;
  assign n17567 = n17563 ^ n15141 ;
  assign n17568 = n17567 ^ n17563 ;
  assign n17569 = ~n17566 & ~n17568 ;
  assign n17570 = n17569 ^ n17563 ;
  assign n17571 = ~n14679 & ~n17570 ;
  assign n17572 = n17571 ^ n15151 ;
  assign n17559 = n15159 ^ n15103 ;
  assign n16706 = n15165 ^ n15154 ;
  assign n17560 = n17559 ^ n16706 ;
  assign n17561 = n15207 & ~n17560 ;
  assign n17573 = n17572 ^ n17561 ;
  assign n15181 = n15141 ^ n14679 ;
  assign n15174 = n15170 ^ n15096 ;
  assign n15173 = n15151 ^ n15088 ;
  assign n15175 = n15174 ^ n15173 ;
  assign n15183 = n15175 ^ n15092 ;
  assign n15184 = n15183 ^ n15157 ;
  assign n15185 = n15184 ^ n15154 ;
  assign n17558 = n15181 & n15185 ;
  assign n17574 = n17573 ^ n17558 ;
  assign n17552 = n15100 ^ n15096 ;
  assign n17553 = n17552 ^ n15162 ;
  assign n17554 = n17553 ^ n15175 ;
  assign n17555 = n14679 & ~n17554 ;
  assign n17556 = n17555 ^ n15100 ;
  assign n17557 = ~n15141 & n17556 ;
  assign n17575 = n17574 ^ n17557 ;
  assign n16713 = ~n15105 & n15208 ;
  assign n17576 = n17575 ^ n16713 ;
  assign n17577 = n15150 & ~n17576 ;
  assign n17578 = n17551 & n17577 ;
  assign n17579 = n17578 ^ n14272 ;
  assign n17580 = n17579 ^ x122 ;
  assign n17581 = n17550 & ~n17580 ;
  assign n17604 = n17581 ^ n17550 ;
  assign n17616 = n17497 & n17604 ;
  assign n17643 = n17616 ^ n17604 ;
  assign n17498 = n17497 ^ n17495 ;
  assign n17499 = n17498 ^ n17496 ;
  assign n17500 = n17499 ^ n17495 ;
  assign n17608 = n17500 & n17604 ;
  assign n17605 = ~n17499 & n17604 ;
  assign n17609 = n17608 ^ n17605 ;
  assign n17644 = n17643 ^ n17609 ;
  assign n15783 = n15032 ^ n14387 ;
  assign n15784 = n14470 ^ n14464 ;
  assign n15785 = n15783 & ~n15784 ;
  assign n15786 = n15785 ^ n14513 ;
  assign n15753 = n14482 ^ n14388 ;
  assign n15754 = n15753 ^ n14482 ;
  assign n15777 = n14524 & ~n15754 ;
  assign n15778 = n15777 ^ n14482 ;
  assign n15779 = n14467 & n15778 ;
  assign n15780 = n15779 ^ n14455 ;
  assign n15770 = n14455 ^ n14388 ;
  assign n15771 = n15770 ^ n14455 ;
  assign n15774 = n14535 & ~n15771 ;
  assign n15775 = n15774 ^ n14455 ;
  assign n15776 = ~n14467 & n15775 ;
  assign n15781 = n15780 ^ n15776 ;
  assign n15758 = n14465 ^ n14429 ;
  assign n15759 = n15758 ^ n14486 ;
  assign n15760 = n15759 ^ n14458 ;
  assign n15761 = n15760 ^ n15758 ;
  assign n15762 = n15758 ^ n14388 ;
  assign n15763 = n15762 ^ n15758 ;
  assign n15764 = n15761 & ~n15763 ;
  assign n15765 = n15764 ^ n15758 ;
  assign n15766 = ~n14467 & ~n15765 ;
  assign n15767 = n15766 ^ n15758 ;
  assign n15752 = n14526 ^ n14482 ;
  assign n15755 = n15752 & n15754 ;
  assign n15756 = n15755 ^ n14482 ;
  assign n15757 = n14387 & n15756 ;
  assign n15768 = n15767 ^ n15757 ;
  assign n15769 = n15768 ^ n14479 ;
  assign n15782 = n15781 ^ n15769 ;
  assign n15787 = n15786 ^ n15782 ;
  assign n15788 = n15787 ^ n15061 ;
  assign n15745 = n14479 ^ n14388 ;
  assign n15746 = n15745 ^ n14479 ;
  assign n15749 = ~n15036 & n15746 ;
  assign n15750 = n15749 ^ n14479 ;
  assign n15751 = n14467 & n15750 ;
  assign n15789 = n15788 ^ n15751 ;
  assign n15790 = ~n15042 & n15789 ;
  assign n15791 = n15790 ^ n12168 ;
  assign n15792 = n15791 ^ x69 ;
  assign n15793 = n15582 ^ x78 ;
  assign n15794 = n15792 & ~n15793 ;
  assign n15795 = n15794 ^ n15792 ;
  assign n15836 = n15492 ^ x101 ;
  assign n15858 = n14925 ^ n14843 ;
  assign n15859 = n15858 ^ n14937 ;
  assign n15860 = n14810 & ~n15859 ;
  assign n15861 = n15860 ^ n14909 ;
  assign n15846 = n14809 & n14904 ;
  assign n15843 = n14902 ^ n14889 ;
  assign n15232 = n14927 ^ n14892 ;
  assign n15844 = n15843 ^ n15232 ;
  assign n15837 = n14955 ^ n14902 ;
  assign n15838 = n14902 ^ n14808 ;
  assign n15839 = n15838 ^ n14902 ;
  assign n15840 = n15837 & ~n15839 ;
  assign n15841 = n15840 ^ n14902 ;
  assign n15842 = n14910 & n15841 ;
  assign n15845 = n15844 ^ n15842 ;
  assign n15847 = n15846 ^ n15845 ;
  assign n15862 = n15861 ^ n15847 ;
  assign n15863 = n15862 ^ n14907 ;
  assign n15864 = n15863 ^ n15857 ;
  assign n15865 = n15864 ^ n14951 ;
  assign n15866 = n15865 ^ n15250 ;
  assign n15867 = n15866 ^ n12265 ;
  assign n15848 = n15847 ^ n14936 ;
  assign n15849 = n15848 ^ n14887 ;
  assign n15850 = n15849 ^ n15847 ;
  assign n15853 = ~n14807 & n15850 ;
  assign n15854 = n15853 ^ n15847 ;
  assign n15855 = ~n14910 & n15854 ;
  assign n15868 = n15867 ^ n15855 ;
  assign n15869 = n15868 ^ x91 ;
  assign n15812 = n13078 ^ n13024 ;
  assign n15813 = n13056 & n15812 ;
  assign n15802 = n13059 ^ n13055 ;
  assign n15803 = n15802 ^ n13060 ;
  assign n15804 = n13058 ^ n13031 ;
  assign n15805 = n15804 ^ n13021 ;
  assign n15806 = ~n15803 & n15805 ;
  assign n15807 = n15806 ^ n13021 ;
  assign n15808 = n15807 ^ n12630 ;
  assign n15800 = n15797 ^ n12630 ;
  assign n15801 = n12827 & n15800 ;
  assign n15809 = n15808 ^ n15801 ;
  assign n15798 = n15797 ^ n13021 ;
  assign n15799 = ~n13010 & n15798 ;
  assign n15810 = n15809 ^ n15799 ;
  assign n15796 = n13057 & ~n13075 ;
  assign n15811 = n15810 ^ n15796 ;
  assign n15814 = n15813 ^ n15811 ;
  assign n15815 = ~n12827 & ~n15814 ;
  assign n15816 = n13048 ^ n11503 ;
  assign n15817 = n15816 ^ n13075 ;
  assign n15818 = ~n13010 & ~n15817 ;
  assign n15819 = n15818 ^ n13048 ;
  assign n15820 = n15815 & n15819 ;
  assign n15821 = n15820 ^ n15814 ;
  assign n15822 = n13019 & ~n15821 ;
  assign n15823 = n13045 ^ n13010 ;
  assign n15824 = n15823 ^ n13045 ;
  assign n15825 = n13046 & ~n15824 ;
  assign n15826 = n15825 ^ n13045 ;
  assign n15827 = n15822 & n15826 ;
  assign n15828 = n15827 ^ n15821 ;
  assign n15829 = ~n15126 & ~n15828 ;
  assign n15830 = n15829 ^ n12211 ;
  assign n15831 = n15830 ^ x108 ;
  assign n15875 = n15869 ^ n15831 ;
  assign n15876 = ~n15869 & ~n15875 ;
  assign n15832 = n14803 ^ n14801 ;
  assign n15833 = n15832 ^ n12177 ;
  assign n15834 = n15833 ^ x118 ;
  assign n15904 = n15876 ^ n15834 ;
  assign n15905 = n15836 & ~n15904 ;
  assign n15835 = ~n15831 & ~n15834 ;
  assign n15879 = n15835 ^ n15834 ;
  assign n15902 = n15836 & ~n15879 ;
  assign n15870 = n15836 & ~n15869 ;
  assign n15882 = n15879 ^ n15831 ;
  assign n15883 = n15870 & ~n15882 ;
  assign n15871 = n15835 & n15870 ;
  assign n15884 = n15883 ^ n15871 ;
  assign n15880 = n15870 & ~n15879 ;
  assign n15881 = n15880 ^ n15870 ;
  assign n15885 = n15884 ^ n15881 ;
  assign n15903 = n15902 ^ n15885 ;
  assign n15906 = n15905 ^ n15903 ;
  assign n16269 = n15795 & n15906 ;
  assign n15877 = n15870 ^ n15869 ;
  assign n15891 = n15877 ^ n15836 ;
  assign n15896 = n15882 ^ n15834 ;
  assign n15897 = n15891 & ~n15896 ;
  assign n15892 = ~n15882 & n15891 ;
  assign n15889 = n15870 ^ n15836 ;
  assign n15890 = ~n15882 & n15889 ;
  assign n15893 = n15892 ^ n15890 ;
  assign n15888 = n15883 ^ n15882 ;
  assign n15894 = n15893 ^ n15888 ;
  assign n15917 = n15897 ^ n15894 ;
  assign n15912 = n15902 ^ n15879 ;
  assign n15886 = n15885 ^ n15871 ;
  assign n15878 = n15877 ^ n15876 ;
  assign n15887 = n15886 ^ n15878 ;
  assign n15895 = n15894 ^ n15887 ;
  assign n15913 = n15912 ^ n15895 ;
  assign n15918 = n15917 ^ n15913 ;
  assign n16299 = n15795 & n15918 ;
  assign n15923 = n15912 ^ n15897 ;
  assign n15899 = n15875 ^ n15834 ;
  assign n15900 = n15899 ^ n15869 ;
  assign n15920 = n15903 ^ n15900 ;
  assign n15908 = n15835 & n15891 ;
  assign n15909 = n15908 ^ n15894 ;
  assign n15907 = n15906 ^ n15884 ;
  assign n15910 = n15909 ^ n15907 ;
  assign n15901 = n15900 ^ n15893 ;
  assign n15911 = n15910 ^ n15901 ;
  assign n15914 = n15913 ^ n15911 ;
  assign n15898 = n15897 ^ n15895 ;
  assign n15915 = n15914 ^ n15898 ;
  assign n15916 = n15915 ^ n15877 ;
  assign n15919 = n15918 ^ n15916 ;
  assign n15921 = n15920 ^ n15919 ;
  assign n15924 = n15923 ^ n15921 ;
  assign n16270 = n15924 ^ n15883 ;
  assign n16271 = n15794 & ~n16270 ;
  assign n15946 = n15919 ^ n15892 ;
  assign n16296 = n15794 & n15946 ;
  assign n16280 = n15903 ^ n15893 ;
  assign n16281 = n16280 ^ n15917 ;
  assign n16277 = n15890 ^ n15880 ;
  assign n16278 = n16277 ^ n15914 ;
  assign n15944 = n15793 ^ n15792 ;
  assign n15953 = n15911 ^ n15793 ;
  assign n15954 = n15953 ^ n15911 ;
  assign n16272 = n15911 ^ n15883 ;
  assign n16273 = n16272 ^ n15911 ;
  assign n16274 = n15954 & n16273 ;
  assign n16275 = n16274 ^ n15911 ;
  assign n16276 = ~n15944 & n16275 ;
  assign n16279 = n16278 ^ n16276 ;
  assign n16282 = n16281 ^ n16279 ;
  assign n16283 = n16282 ^ n16276 ;
  assign n16284 = ~n15792 & n16283 ;
  assign n16285 = n16284 ^ n16279 ;
  assign n15945 = n15902 ^ n15880 ;
  assign n15959 = n15945 ^ n15885 ;
  assign n15960 = n15795 & n15959 ;
  assign n16294 = n16285 ^ n15960 ;
  assign n16286 = n16285 ^ n16276 ;
  assign n15873 = n15836 ^ n15834 ;
  assign n15874 = n15873 ^ n15869 ;
  assign n15922 = n15921 ^ n15874 ;
  assign n16289 = n16286 ^ n15922 ;
  assign n16290 = n16289 ^ n16286 ;
  assign n16291 = ~n15792 & n16290 ;
  assign n16292 = n16291 ^ n16286 ;
  assign n16293 = n15793 & ~n16292 ;
  assign n16295 = n16294 ^ n16293 ;
  assign n16297 = n16296 ^ n16295 ;
  assign n16298 = ~n16271 & n16297 ;
  assign n16300 = n16299 ^ n16298 ;
  assign n16301 = ~n16269 & n16300 ;
  assign n16302 = n16301 ^ n12352 ;
  assign n17493 = n16302 ^ x72 ;
  assign n16814 = n15868 ^ x125 ;
  assign n15305 = n14784 ^ n14680 ;
  assign n15307 = ~n14749 & n14788 ;
  assign n15308 = n15307 ^ n14775 ;
  assign n15309 = n15308 ^ n14789 ;
  assign n15310 = ~n14784 & n15309 ;
  assign n15311 = n15310 ^ n14789 ;
  assign n15306 = n14756 ^ n14754 ;
  assign n15312 = n15311 ^ n15306 ;
  assign n15313 = n15312 ^ n14680 ;
  assign n15314 = n15313 ^ n15312 ;
  assign n15315 = n15311 ^ n14769 ;
  assign n15316 = n15315 ^ n15312 ;
  assign n15317 = n15314 & ~n15316 ;
  assign n15318 = n15317 ^ n15312 ;
  assign n15319 = n15305 & ~n15318 ;
  assign n15320 = n15319 ^ n15311 ;
  assign n15321 = n14770 ^ n14769 ;
  assign n15322 = ~n15320 & n15321 ;
  assign n15323 = n15322 ^ n11612 ;
  assign n16815 = n15323 ^ x76 ;
  assign n16816 = n16814 & n16815 ;
  assign n16742 = n14327 ^ n14278 ;
  assign n16741 = n14348 ^ n14326 ;
  assign n16743 = n16742 ^ n16741 ;
  assign n16744 = n16743 ^ n14326 ;
  assign n16745 = ~n14315 & ~n16744 ;
  assign n16746 = n16745 ^ n16741 ;
  assign n16755 = n16746 ^ n14320 ;
  assign n16748 = n16746 ^ n14997 ;
  assign n16747 = n16746 ^ n15506 ;
  assign n16749 = n16748 ^ n16747 ;
  assign n16752 = n14315 & ~n16749 ;
  assign n16753 = n16752 ^ n16748 ;
  assign n16754 = n14167 & n16753 ;
  assign n16756 = n16755 ^ n16754 ;
  assign n16739 = n14338 ^ n14327 ;
  assign n16740 = n14372 & n16739 ;
  assign n16757 = n16756 ^ n16740 ;
  assign n16738 = ~n15022 & n15506 ;
  assign n16758 = n16757 ^ n16738 ;
  assign n16766 = n14346 ^ n14325 ;
  assign n16767 = n16766 ^ n14332 ;
  assign n16768 = n16767 ^ n14349 ;
  assign n16769 = n14167 & ~n16768 ;
  assign n16770 = n16769 ^ n14332 ;
  assign n16771 = n14315 & n16770 ;
  assign n16772 = n16771 ^ n14339 ;
  assign n16761 = n14339 ^ n14315 ;
  assign n16762 = n16761 ^ n14339 ;
  assign n16763 = n15000 & ~n16762 ;
  assign n16764 = n16763 ^ n14339 ;
  assign n16765 = n14167 & n16764 ;
  assign n16773 = n16772 ^ n16765 ;
  assign n16774 = n16758 & ~n16773 ;
  assign n16775 = n16774 ^ n13216 ;
  assign n16776 = n16775 ^ x75 ;
  assign n16800 = n14644 ^ n14118 ;
  assign n16792 = n14122 ^ n14095 ;
  assign n16791 = n14080 ^ n14070 ;
  assign n16793 = n16792 ^ n16791 ;
  assign n16794 = n16793 ^ n14649 ;
  assign n16795 = ~n13934 & n16794 ;
  assign n16796 = n16795 ^ n14649 ;
  assign n16797 = ~n13968 & n16796 ;
  assign n16789 = n14094 & ~n14124 ;
  assign n16784 = n14113 ^ n14075 ;
  assign n16785 = n13968 & ~n16784 ;
  assign n16778 = n14134 ^ n14095 ;
  assign n14127 = n14126 ^ n14111 ;
  assign n16777 = n14158 ^ n14127 ;
  assign n16779 = n16778 ^ n16777 ;
  assign n16780 = n16779 ^ n14158 ;
  assign n16781 = ~n13968 & n16780 ;
  assign n16782 = n16781 ^ n16777 ;
  assign n16783 = n16782 ^ n14158 ;
  assign n16786 = n16785 ^ n16783 ;
  assign n16787 = ~n13934 & n16786 ;
  assign n16788 = n16787 ^ n16782 ;
  assign n16790 = n16789 ^ n16788 ;
  assign n16798 = n16797 ^ n16790 ;
  assign n16799 = ~n14101 & ~n16798 ;
  assign n16801 = n16800 ^ n16799 ;
  assign n16802 = ~n14676 & ~n16801 ;
  assign n16803 = n16802 ^ n13177 ;
  assign n16804 = n16803 ^ x93 ;
  assign n16805 = n16776 & ~n16804 ;
  assign n16806 = n16805 ^ n16804 ;
  assign n15330 = n13878 ^ n13815 ;
  assign n15331 = n15330 ^ n13869 ;
  assign n15332 = n15331 ^ n13837 ;
  assign n15333 = n15332 ^ n13855 ;
  assign n15334 = n15333 ^ n15331 ;
  assign n15335 = n15331 ^ n13576 ;
  assign n15336 = n15335 ^ n15331 ;
  assign n15337 = ~n15334 & ~n15336 ;
  assign n15338 = n15337 ^ n15331 ;
  assign n15339 = n13578 & ~n15338 ;
  assign n15340 = n15339 ^ n15331 ;
  assign n15341 = n13576 & n15340 ;
  assign n15345 = n15344 ^ n13839 ;
  assign n15346 = n13839 ^ n13577 ;
  assign n15347 = n15346 ^ n13839 ;
  assign n15348 = ~n15345 & ~n15347 ;
  assign n15349 = n15348 ^ n13839 ;
  assign n15350 = n15341 & n15349 ;
  assign n15351 = n15350 ^ n15340 ;
  assign n15356 = n15351 ^ n11580 ;
  assign n15364 = n15363 ^ n15356 ;
  assign n15352 = ~n13577 & ~n13875 ;
  assign n15353 = n15352 ^ n13826 ;
  assign n15354 = ~n13576 & n15353 ;
  assign n15355 = n15351 & n15354 ;
  assign n15365 = n15364 ^ n15355 ;
  assign n16735 = n15365 ^ x100 ;
  assign n16736 = n15791 ^ x94 ;
  assign n16737 = ~n16735 & n16736 ;
  assign n16809 = n16737 ^ n16736 ;
  assign n16830 = n16809 ^ n16735 ;
  assign n16834 = ~n16806 & n16830 ;
  assign n17051 = n16816 & n16834 ;
  assign n16807 = n16737 & ~n16806 ;
  assign n16817 = n16816 ^ n16815 ;
  assign n16819 = n16817 ^ n16814 ;
  assign n17043 = n16807 & ~n16819 ;
  assign n16844 = n16830 ^ n16736 ;
  assign n16869 = n16805 & ~n16844 ;
  assign n17042 = n16817 & n16869 ;
  assign n17044 = n17043 ^ n17042 ;
  assign n16810 = n16805 ^ n16776 ;
  assign n16856 = n16810 & ~n16844 ;
  assign n16833 = n16810 & n16830 ;
  assign n16835 = n16834 ^ n16833 ;
  assign n16831 = n16805 & n16830 ;
  assign n16832 = n16831 ^ n16830 ;
  assign n16836 = n16835 ^ n16832 ;
  assign n17030 = n16856 ^ n16836 ;
  assign n16823 = n16810 ^ n16804 ;
  assign n16845 = n16823 & ~n16844 ;
  assign n17040 = n17030 ^ n16845 ;
  assign n16808 = n16737 & n16805 ;
  assign n17014 = n16809 ^ n16808 ;
  assign n16838 = n16737 & n16823 ;
  assign n17013 = n16838 ^ n16807 ;
  assign n17015 = n17014 ^ n17013 ;
  assign n17016 = n16814 & n17015 ;
  assign n16824 = n16809 & n16823 ;
  assign n16822 = n16805 & n16809 ;
  assign n16825 = n16824 ^ n16822 ;
  assign n16811 = n16809 & n16810 ;
  assign n16821 = n16811 ^ n16809 ;
  assign n16826 = n16825 ^ n16821 ;
  assign n16812 = n16811 ^ n16808 ;
  assign n16827 = n16826 ^ n16812 ;
  assign n17017 = n17016 ^ n16827 ;
  assign n17041 = n17040 ^ n17017 ;
  assign n17045 = n17044 ^ n17041 ;
  assign n17046 = n17045 ^ n14314 ;
  assign n17032 = n16856 ^ n16834 ;
  assign n17031 = n17030 ^ n16869 ;
  assign n17033 = n17032 ^ n17031 ;
  assign n17034 = n17033 ^ n17030 ;
  assign n17035 = n17030 ^ n16815 ;
  assign n17036 = n17035 ^ n17030 ;
  assign n17037 = n17034 & ~n17036 ;
  assign n17038 = n17037 ^ n17030 ;
  assign n17039 = ~n16814 & n17038 ;
  assign n17047 = n17046 ^ n17039 ;
  assign n16848 = n16815 ^ n16814 ;
  assign n17022 = n16845 ^ n16815 ;
  assign n17023 = n17022 ^ n16845 ;
  assign n17024 = n16869 ^ n16833 ;
  assign n17027 = ~n17023 & n17024 ;
  assign n17028 = n17027 ^ n16845 ;
  assign n17029 = n16848 & n17028 ;
  assign n17048 = n17047 ^ n17029 ;
  assign n16862 = ~n16806 & ~n16844 ;
  assign n16878 = n16862 ^ n16836 ;
  assign n17018 = n16878 ^ n16831 ;
  assign n17019 = n17018 ^ n17017 ;
  assign n16852 = n16737 & n16810 ;
  assign n17009 = n16852 ^ n16822 ;
  assign n16813 = n16812 ^ n16807 ;
  assign n16828 = n16827 ^ n16813 ;
  assign n17008 = n16831 ^ n16828 ;
  assign n17010 = n17009 ^ n17008 ;
  assign n17011 = n17010 ^ n16878 ;
  assign n17012 = n16814 & n17011 ;
  assign n17020 = n17019 ^ n17012 ;
  assign n17021 = n16815 & n17020 ;
  assign n17049 = n17048 ^ n17021 ;
  assign n17005 = n16826 ^ n16808 ;
  assign n16839 = n16838 ^ n16811 ;
  assign n17006 = n17005 ^ n16839 ;
  assign n17007 = n16817 & n17006 ;
  assign n17050 = n17049 ^ n17007 ;
  assign n17052 = n17051 ^ n17050 ;
  assign n17494 = n17052 ^ x115 ;
  assign n17674 = n17493 & n17494 ;
  assign n17675 = n17674 ^ n17494 ;
  assign n17582 = n17581 ^ n17580 ;
  assign n17583 = n17582 ^ n17550 ;
  assign n17634 = n17497 & n17583 ;
  assign n19064 = n17634 ^ n17605 ;
  assign n17636 = ~n17499 & ~n17582 ;
  assign n17589 = ~n17499 & n17581 ;
  assign n17590 = n17589 ^ n17581 ;
  assign n17587 = n17497 & n17581 ;
  assign n17586 = n17498 & n17581 ;
  assign n17588 = n17587 ^ n17586 ;
  assign n17591 = n17590 ^ n17588 ;
  assign n17637 = n17636 ^ n17591 ;
  assign n19065 = n19064 ^ n17637 ;
  assign n19066 = n17675 & n19065 ;
  assign n17639 = n17498 & ~n17582 ;
  assign n17665 = n17639 ^ n17493 ;
  assign n17666 = n17665 ^ n17639 ;
  assign n17662 = n17639 ^ n17636 ;
  assign n18110 = n17662 ^ n17639 ;
  assign n18111 = n18110 ^ n17639 ;
  assign n18112 = n17666 & n18111 ;
  assign n18113 = n18112 ^ n17639 ;
  assign n18114 = ~n17494 & n18113 ;
  assign n19057 = n18114 ^ n17586 ;
  assign n17648 = n17498 & n17583 ;
  assign n19055 = n17648 ^ n17616 ;
  assign n19056 = n17674 & n19055 ;
  assign n19058 = n19057 ^ n19056 ;
  assign n19059 = n19058 ^ n18114 ;
  assign n19053 = n17648 ^ n17587 ;
  assign n19054 = ~n17493 & n19053 ;
  assign n19060 = n19059 ^ n19054 ;
  assign n19061 = ~n17494 & n19060 ;
  assign n19062 = n19061 ^ n19058 ;
  assign n17585 = ~n17499 & n17583 ;
  assign n17592 = n17591 ^ n17585 ;
  assign n17584 = n17500 & n17583 ;
  assign n17593 = n17592 ^ n17584 ;
  assign n19051 = n17674 ^ n17493 ;
  assign n19052 = n17593 & n19051 ;
  assign n19063 = n19062 ^ n19052 ;
  assign n19067 = n19066 ^ n19063 ;
  assign n17615 = n17494 ^ n17493 ;
  assign n17618 = n17497 & ~n17582 ;
  assign n17661 = n17618 ^ n17582 ;
  assign n17663 = n17662 ^ n17661 ;
  assign n19045 = n17663 ^ n17608 ;
  assign n19046 = n17608 ^ n17493 ;
  assign n19047 = n19046 ^ n17608 ;
  assign n19048 = ~n19045 & n19047 ;
  assign n19049 = n19048 ^ n17608 ;
  assign n19050 = ~n17615 & n19049 ;
  assign n19068 = n19067 ^ n19050 ;
  assign n19069 = n19068 ^ n17589 ;
  assign n17670 = n17584 & ~n17615 ;
  assign n17664 = n17663 ^ n17639 ;
  assign n17667 = ~n17664 & ~n17666 ;
  assign n17668 = n17667 ^ n17639 ;
  assign n17669 = n17494 & n17668 ;
  assign n17671 = n17670 ^ n17669 ;
  assign n19070 = n19069 ^ n17671 ;
  assign n18127 = n17616 & n17675 ;
  assign n17606 = n17605 ^ n17493 ;
  assign n17607 = n17606 ^ n17605 ;
  assign n17612 = n17607 & n17609 ;
  assign n17613 = n17612 ^ n17605 ;
  assign n17614 = ~n17494 & n17613 ;
  assign n18128 = n18127 ^ n17614 ;
  assign n19071 = n19070 ^ n18128 ;
  assign n17619 = n17618 ^ n17587 ;
  assign n19040 = n17589 ^ n17493 ;
  assign n19041 = n19040 ^ n17589 ;
  assign n19042 = n17619 & n19041 ;
  assign n19043 = n19042 ^ n17589 ;
  assign n19044 = n17615 & n19043 ;
  assign n19072 = n19071 ^ n19044 ;
  assign n19073 = ~n17644 & ~n19072 ;
  assign n19074 = n19073 ^ n14385 ;
  assign n19075 = n19074 ^ x88 ;
  assign n14637 = n13548 & n14543 ;
  assign n14626 = n14614 ^ n14551 ;
  assign n14627 = n14551 ^ n14386 ;
  assign n14628 = n14627 ^ n14551 ;
  assign n14629 = n14626 & n14628 ;
  assign n14630 = n14629 ^ n14551 ;
  assign n14631 = ~n14538 & n14630 ;
  assign n14587 = n14576 ^ n14557 ;
  assign n14588 = n14587 ^ n14567 ;
  assign n14559 = n14558 ^ n14552 ;
  assign n14560 = n14559 ^ n14550 ;
  assign n14586 = n14585 ^ n14560 ;
  assign n14589 = n14588 ^ n14586 ;
  assign n14590 = ~n14538 & ~n14589 ;
  assign n14591 = n14590 ^ n14586 ;
  assign n14632 = n14631 ^ n14591 ;
  assign n14615 = n14614 ^ n14566 ;
  assign n14616 = ~n14386 & n14615 ;
  assign n14617 = n14616 ^ n14566 ;
  assign n14618 = n14617 ^ n14556 ;
  assign n14619 = n14618 ^ n14617 ;
  assign n14620 = n14617 ^ n14538 ;
  assign n14621 = n14620 ^ n14617 ;
  assign n14622 = n14619 & n14621 ;
  assign n14623 = n14622 ^ n14617 ;
  assign n14624 = ~n14540 & n14623 ;
  assign n14625 = n14624 ^ n14617 ;
  assign n14633 = n14632 ^ n14625 ;
  assign n14612 = n14539 & n14572 ;
  assign n14611 = n14543 & ~n14546 ;
  assign n14613 = n14612 ^ n14611 ;
  assign n14634 = n14633 ^ n14613 ;
  assign n14600 = n14563 ^ n14555 ;
  assign n14601 = n14600 ^ n14566 ;
  assign n14602 = n14538 & n14601 ;
  assign n14603 = n14602 ^ n14563 ;
  assign n14606 = n14563 ^ n14538 ;
  assign n14607 = n14606 ^ n14563 ;
  assign n14608 = n14603 & n14607 ;
  assign n14609 = n14608 ^ n14563 ;
  assign n14610 = n14386 & n14609 ;
  assign n14635 = n14634 ^ n14610 ;
  assign n14593 = n14591 ^ n14553 ;
  assign n14592 = n14591 ^ n14551 ;
  assign n14594 = n14593 ^ n14592 ;
  assign n14595 = n14593 ^ n14538 ;
  assign n14596 = n14595 ^ n14593 ;
  assign n14597 = n14594 & n14596 ;
  assign n14598 = n14597 ^ n14593 ;
  assign n14599 = n14386 & ~n14598 ;
  assign n14636 = n14635 ^ n14599 ;
  assign n14638 = n14637 ^ n14636 ;
  assign n14639 = ~n14544 & n14638 ;
  assign n14640 = n14639 ^ n13967 ;
  assign n14641 = n14640 ^ x120 ;
  assign n15228 = ~n14807 & n14890 ;
  assign n15229 = n15228 ^ n14889 ;
  assign n15259 = n15229 ^ n14928 ;
  assign n15260 = n15259 ^ n14903 ;
  assign n15261 = n15260 ^ n14927 ;
  assign n15262 = n15261 ^ n15229 ;
  assign n15263 = ~n14807 & ~n15262 ;
  assign n15264 = n15263 ^ n15259 ;
  assign n15265 = ~n14910 & ~n15264 ;
  assign n15248 = n15247 ^ n14903 ;
  assign n15249 = n15248 ^ n15244 ;
  assign n15251 = n15250 ^ n15249 ;
  assign n15238 = n15232 ^ n14903 ;
  assign n15239 = ~n14807 & n15238 ;
  assign n15252 = n15251 ^ n15239 ;
  assign n15233 = n15232 ^ n14884 ;
  assign n15234 = n15233 ^ n14902 ;
  assign n15235 = ~n15231 & n15234 ;
  assign n15236 = n15235 ^ n14902 ;
  assign n15237 = ~n14910 & n15236 ;
  assign n15253 = n15252 ^ n15237 ;
  assign n15254 = n15253 ^ n15229 ;
  assign n15255 = n15254 ^ n14984 ;
  assign n15256 = n15255 ^ n12001 ;
  assign n15226 = n14929 ^ n14884 ;
  assign n15227 = n14910 & ~n15226 ;
  assign n15257 = n15256 ^ n15227 ;
  assign n15224 = n14891 ^ n14882 ;
  assign n15225 = n14807 & n15224 ;
  assign n15258 = n15257 ^ n15225 ;
  assign n15266 = n15265 ^ n15258 ;
  assign n15267 = n15266 ^ x112 ;
  assign n15268 = n14537 ^ x98 ;
  assign n15269 = n15267 & ~n15268 ;
  assign n15275 = n13531 ^ n13310 ;
  assign n15276 = n15275 ^ n13531 ;
  assign n15277 = n13534 & ~n15276 ;
  assign n15278 = n15277 ^ n13531 ;
  assign n15279 = n13146 & n15278 ;
  assign n15292 = n15279 ^ n13459 ;
  assign n15284 = n13465 ^ n13459 ;
  assign n15285 = n15284 ^ n13481 ;
  assign n15289 = n15288 ^ n15285 ;
  assign n15282 = n13500 ^ n13465 ;
  assign n15283 = ~n13310 & ~n15282 ;
  assign n15290 = n15289 ^ n15283 ;
  assign n15291 = ~n15270 & ~n15290 ;
  assign n15293 = n15292 ^ n15291 ;
  assign n15280 = n13484 ^ n13478 ;
  assign n15281 = n13312 & ~n15280 ;
  assign n15294 = n15293 ^ n15281 ;
  assign n15298 = n15297 ^ n15294 ;
  assign n15272 = ~n13489 & ~n13507 ;
  assign n15299 = n15298 ^ n15272 ;
  assign n15300 = n15299 ^ n15271 ;
  assign n15301 = n15300 ^ n13522 ;
  assign n15302 = n15301 ^ n13506 ;
  assign n15303 = n15302 ^ n11661 ;
  assign n15304 = n15303 ^ x73 ;
  assign n15324 = n15323 ^ x64 ;
  assign n15325 = n15304 & n15324 ;
  assign n15326 = n15325 ^ n15324 ;
  assign n15327 = n15269 & n15326 ;
  assign n15329 = n13102 ^ x66 ;
  assign n15366 = n15365 ^ x88 ;
  assign n15369 = n15326 ^ n15304 ;
  assign n15370 = n15269 ^ n15268 ;
  assign n15371 = n15370 ^ n15267 ;
  assign n15372 = n15371 ^ n15268 ;
  assign n15373 = ~n15369 & n15372 ;
  assign n15409 = n15373 ^ n15269 ;
  assign n15375 = n15372 ^ n15304 ;
  assign n15381 = n15324 ^ n15304 ;
  assign n15382 = n15381 ^ n15267 ;
  assign n15383 = n15382 ^ n15268 ;
  assign n15384 = n15375 & ~n15383 ;
  assign n15401 = n15384 ^ n15324 ;
  assign n15385 = ~n15267 & n15326 ;
  assign n15386 = n15385 ^ n15327 ;
  assign n15391 = n15386 ^ n15375 ;
  assign n15376 = ~n15324 & ~n15375 ;
  assign n15392 = n15391 ^ n15376 ;
  assign n15378 = n15268 ^ n15267 ;
  assign n15389 = n15326 & n15378 ;
  assign n15390 = n15389 ^ n15386 ;
  assign n15393 = n15392 ^ n15390 ;
  assign n15387 = n15386 ^ n15384 ;
  assign n15388 = n15387 ^ n15383 ;
  assign n15394 = n15393 ^ n15388 ;
  assign n15379 = n15378 ^ n15304 ;
  assign n15380 = ~n15324 & n15379 ;
  assign n15395 = n15394 ^ n15380 ;
  assign n15402 = n15401 ^ n15395 ;
  assign n15410 = n15409 ^ n15402 ;
  assign n15406 = n15369 ^ n15324 ;
  assign n15407 = n15269 & n15406 ;
  assign n15403 = n15386 ^ n15326 ;
  assign n15404 = n15403 ^ n15402 ;
  assign n15328 = n15269 & n15325 ;
  assign n15399 = n15389 ^ n15328 ;
  assign n15396 = n15395 ^ n15376 ;
  assign n15374 = n15373 ^ n15369 ;
  assign n15377 = n15376 ^ n15374 ;
  assign n15397 = n15396 ^ n15377 ;
  assign n15398 = n15397 ^ n15373 ;
  assign n15400 = n15399 ^ n15398 ;
  assign n15405 = n15404 ^ n15400 ;
  assign n15408 = n15407 ^ n15405 ;
  assign n15411 = n15410 ^ n15408 ;
  assign n15412 = ~n15366 & ~n15411 ;
  assign n15413 = n15412 ^ n15373 ;
  assign n15414 = n15329 & n15413 ;
  assign n15415 = n15414 ^ n15373 ;
  assign n15419 = n15403 ^ n15390 ;
  assign n15420 = n15419 ^ n15328 ;
  assign n15367 = n15329 & ~n15366 ;
  assign n15428 = n15367 ^ n15329 ;
  assign n15439 = n15420 & n15428 ;
  assign n15422 = n15269 & ~n15369 ;
  assign n15421 = n15420 ^ n15387 ;
  assign n15423 = n15422 ^ n15421 ;
  assign n15424 = n15366 & ~n15423 ;
  assign n15416 = n15407 ^ n15406 ;
  assign n15417 = n15416 ^ n15397 ;
  assign n15418 = n15417 ^ n15393 ;
  assign n15425 = n15424 ^ n15418 ;
  assign n15426 = ~n15329 & n15425 ;
  assign n15427 = n15426 ^ n15417 ;
  assign n15429 = n15367 ^ n15366 ;
  assign n15430 = n15429 ^ n15428 ;
  assign n15431 = n15430 ^ n15402 ;
  assign n15432 = n15422 ^ n15394 ;
  assign n15433 = n15432 ^ n15374 ;
  assign n15434 = n15433 ^ n15407 ;
  assign n15435 = n15434 ^ n15430 ;
  assign n15436 = n15431 & n15435 ;
  assign n15437 = n15436 ^ n15430 ;
  assign n15438 = n15427 & n15437 ;
  assign n15440 = n15439 ^ n15438 ;
  assign n15441 = ~n15415 & n15440 ;
  assign n15368 = n15328 & n15367 ;
  assign n15442 = n15441 ^ n15368 ;
  assign n15443 = ~n15327 & n15442 ;
  assign n15444 = n15422 ^ n15392 ;
  assign n15445 = n15392 ^ n15366 ;
  assign n15446 = n15445 ^ n15392 ;
  assign n15447 = ~n15444 & ~n15446 ;
  assign n15448 = n15447 ^ n15392 ;
  assign n15449 = ~n15329 & ~n15448 ;
  assign n15450 = n15443 & ~n15449 ;
  assign n15451 = n15450 ^ n13994 ;
  assign n15452 = n15451 ^ x97 ;
  assign n15636 = ~n15496 & n15635 ;
  assign n15725 = n15645 ^ n15493 ;
  assign n15726 = n15725 ^ n15645 ;
  assign n15727 = n15672 & ~n15726 ;
  assign n15728 = n15727 ^ n15645 ;
  assign n15729 = n15453 & n15728 ;
  assign n15705 = n15665 ^ n15661 ;
  assign n15706 = n15705 ^ n15546 ;
  assign n15707 = n15493 & n15706 ;
  assign n15708 = n15707 ^ n15685 ;
  assign n15712 = n15708 ^ n15631 ;
  assign n15714 = n15713 ^ n15712 ;
  assign n15715 = n15714 ^ n15708 ;
  assign n15718 = n15493 & ~n15715 ;
  assign n15696 = n15673 ^ n15494 ;
  assign n15697 = n15640 ^ n15453 ;
  assign n15700 = ~n15673 & n15697 ;
  assign n15701 = n15700 ^ n15453 ;
  assign n15702 = n15696 & ~n15701 ;
  assign n15703 = n15702 ^ n15494 ;
  assign n15695 = n15655 & ~n15694 ;
  assign n15704 = n15703 ^ n15695 ;
  assign n15709 = n15708 ^ n15704 ;
  assign n15687 = n15686 ^ n15667 ;
  assign n15688 = n15687 ^ n15651 ;
  assign n15689 = n15651 ^ n15493 ;
  assign n15690 = n15689 ^ n15651 ;
  assign n15691 = n15688 & ~n15690 ;
  assign n15692 = n15691 ^ n15651 ;
  assign n15693 = n15683 & ~n15692 ;
  assign n15710 = n15709 ^ n15693 ;
  assign n15711 = n15710 ^ n15704 ;
  assign n15719 = n15718 ^ n15711 ;
  assign n15720 = n15719 ^ n15693 ;
  assign n15721 = n15683 & ~n15720 ;
  assign n15722 = n15721 ^ n15710 ;
  assign n15730 = n15729 ^ n15722 ;
  assign n15650 = n15649 ^ n15494 ;
  assign n15677 = n15676 ^ n15496 ;
  assign n15680 = ~n15649 & n15677 ;
  assign n15681 = n15680 ^ n15496 ;
  assign n15682 = n15650 & ~n15681 ;
  assign n15731 = n15730 ^ n15682 ;
  assign n15732 = ~n15636 & ~n15731 ;
  assign n15739 = n15732 & ~n15738 ;
  assign n15740 = n15739 ^ n14037 ;
  assign n15741 = n15740 ^ x123 ;
  assign n15742 = ~n15452 & n15741 ;
  assign n15872 = n15795 & n15871 ;
  assign n15929 = n15909 ^ n15906 ;
  assign n15930 = n15929 ^ n15919 ;
  assign n15931 = n15930 ^ n15873 ;
  assign n15932 = ~n15793 & n15931 ;
  assign n15927 = n15919 ^ n15913 ;
  assign n15925 = n15924 ^ n15890 ;
  assign n15926 = n15925 ^ n15894 ;
  assign n15928 = n15927 ^ n15926 ;
  assign n15933 = n15932 ^ n15928 ;
  assign n15961 = n15960 ^ n15933 ;
  assign n15955 = n15945 ^ n15911 ;
  assign n15956 = ~n15954 & n15955 ;
  assign n15957 = n15956 ^ n15911 ;
  assign n15958 = n15944 & n15957 ;
  assign n15962 = n15961 ^ n15958 ;
  assign n15947 = n15946 ^ n15945 ;
  assign n15948 = n15946 ^ n15793 ;
  assign n15949 = n15948 ^ n15946 ;
  assign n15950 = n15947 & n15949 ;
  assign n15951 = n15950 ^ n15946 ;
  assign n15952 = n15944 & n15951 ;
  assign n15963 = n15962 ^ n15952 ;
  assign n15935 = n15893 ^ n15886 ;
  assign n15936 = n15935 ^ n15898 ;
  assign n15937 = n15936 ^ n15933 ;
  assign n15934 = n15933 ^ n15922 ;
  assign n15938 = n15937 ^ n15934 ;
  assign n15939 = n15937 ^ n15793 ;
  assign n15940 = n15939 ^ n15937 ;
  assign n15941 = n15938 & ~n15940 ;
  assign n15942 = n15941 ^ n15937 ;
  assign n15943 = ~n15792 & ~n15942 ;
  assign n15964 = n15963 ^ n15943 ;
  assign n15965 = ~n15872 & n15964 ;
  assign n15966 = n15965 ^ n14065 ;
  assign n15967 = n15966 ^ x106 ;
  assign n16122 = n16121 ^ n14005 ;
  assign n16093 = n16090 ^ n14005 ;
  assign n16082 = n16081 ^ n16074 ;
  assign n16091 = n16090 ^ n16082 ;
  assign n16092 = ~n15968 & n16091 ;
  assign n16094 = n16093 ^ n16092 ;
  assign n16123 = n16122 ^ n16094 ;
  assign n16124 = n16111 & ~n16123 ;
  assign n16125 = n16124 ^ n16094 ;
  assign n16075 = n15968 & n16074 ;
  assign n16126 = n16125 ^ n16075 ;
  assign n16127 = n16126 ^ x88 ;
  assign n16128 = ~n15967 & ~n16127 ;
  assign n16132 = n16128 ^ n15967 ;
  assign n16135 = n16132 ^ n16127 ;
  assign n16143 = n15742 & ~n16135 ;
  assign n16141 = ~n15452 & ~n15967 ;
  assign n15743 = n15742 ^ n15452 ;
  assign n16133 = ~n15743 & ~n16132 ;
  assign n16142 = n16141 ^ n16133 ;
  assign n16144 = n16143 ^ n16142 ;
  assign n16137 = ~n15743 & n16128 ;
  assign n16140 = n16137 ^ n15742 ;
  assign n16145 = n16144 ^ n16140 ;
  assign n16136 = ~n15743 & ~n16135 ;
  assign n16138 = n16137 ^ n16136 ;
  assign n16134 = n16133 ^ n15743 ;
  assign n16139 = n16138 ^ n16134 ;
  assign n16146 = n16145 ^ n16139 ;
  assign n15744 = n15743 ^ n15741 ;
  assign n16129 = n16128 ^ n16127 ;
  assign n16130 = n15744 & ~n16129 ;
  assign n16131 = n16130 ^ n16129 ;
  assign n16147 = n16146 ^ n16131 ;
  assign n15220 = n15219 ^ n15209 ;
  assign n15221 = n15220 ^ n13933 ;
  assign n15182 = n15102 ^ n15100 ;
  assign n15186 = n15185 ^ n15182 ;
  assign n15187 = n15141 & n15186 ;
  assign n15188 = n15187 ^ n15161 ;
  assign n15189 = n15188 ^ n14679 ;
  assign n15190 = n15189 ^ n15188 ;
  assign n15191 = n15188 ^ n15169 ;
  assign n15192 = n15191 ^ n15188 ;
  assign n15193 = n15190 & ~n15192 ;
  assign n15194 = n15193 ^ n15188 ;
  assign n15195 = n15181 & n15194 ;
  assign n15196 = n15195 ^ n15187 ;
  assign n15179 = n15151 ^ n15092 ;
  assign n15180 = n15178 & n15179 ;
  assign n15197 = n15196 ^ n15180 ;
  assign n15152 = n15151 ^ n15101 ;
  assign n15155 = n15154 ^ n15152 ;
  assign n15171 = n15170 ^ n15155 ;
  assign n15172 = ~n15141 & ~n15171 ;
  assign n15176 = n15175 ^ n15172 ;
  assign n15177 = ~n14679 & ~n15176 ;
  assign n15198 = n15197 ^ n15177 ;
  assign n15199 = n15150 & ~n15198 ;
  assign n15200 = n15174 ^ n15162 ;
  assign n15201 = n15162 ^ n15141 ;
  assign n15202 = n15201 ^ n15162 ;
  assign n15203 = ~n15200 & n15202 ;
  assign n15204 = n15203 ^ n15162 ;
  assign n15205 = ~n15181 & n15204 ;
  assign n15206 = n15199 & ~n15205 ;
  assign n15222 = n15221 ^ n15206 ;
  assign n15223 = n15222 ^ x65 ;
  assign n16148 = n16147 ^ n15223 ;
  assign n16149 = n16148 ^ n16147 ;
  assign n16154 = n15744 ^ n15452 ;
  assign n16165 = ~n16135 & n16154 ;
  assign n16157 = n15744 & n16128 ;
  assign n16166 = n16165 ^ n16157 ;
  assign n16167 = n16166 ^ n16147 ;
  assign n16150 = n15742 & n16128 ;
  assign n16151 = n16150 ^ n16137 ;
  assign n16156 = n16151 ^ n16128 ;
  assign n16158 = n16157 ^ n16156 ;
  assign n16168 = n16167 ^ n16158 ;
  assign n16155 = ~n15967 & n16154 ;
  assign n16159 = n16158 ^ n16155 ;
  assign n16162 = n16159 ^ n16130 ;
  assign n16160 = n16159 ^ n16133 ;
  assign n16152 = n16151 ^ n16142 ;
  assign n16153 = n16152 ^ n16132 ;
  assign n16161 = n16160 ^ n16153 ;
  assign n16163 = n16162 ^ n16161 ;
  assign n16164 = n16163 ^ n15452 ;
  assign n16169 = n16168 ^ n16164 ;
  assign n16170 = n16169 ^ n16147 ;
  assign n16171 = n16170 ^ n16147 ;
  assign n16172 = n16171 ^ n16147 ;
  assign n16173 = n16149 & ~n16172 ;
  assign n16174 = n16173 ^ n16147 ;
  assign n16175 = n14641 & n16174 ;
  assign n19138 = n16175 ^ n14163 ;
  assign n16187 = ~n14641 & n15223 ;
  assign n16188 = n16187 ^ n14641 ;
  assign n16218 = ~n16161 & ~n16188 ;
  assign n19130 = n16150 ^ n16139 ;
  assign n19131 = n19130 ^ n16166 ;
  assign n19132 = n15223 & ~n19131 ;
  assign n16177 = n16158 ^ n16133 ;
  assign n19133 = n19132 ^ n16177 ;
  assign n19134 = n14641 & n19133 ;
  assign n16192 = n16188 ^ n15223 ;
  assign n16193 = n16192 ^ n16187 ;
  assign n16202 = n16161 ^ n16145 ;
  assign n16203 = n16161 ^ n15223 ;
  assign n16204 = n16203 ^ n16161 ;
  assign n16205 = ~n16202 & ~n16204 ;
  assign n16206 = n16205 ^ n16161 ;
  assign n16207 = ~n16193 & ~n16206 ;
  assign n19125 = n16207 ^ n16177 ;
  assign n18170 = n16152 ^ n16145 ;
  assign n18171 = n18170 ^ n16139 ;
  assign n18172 = n16139 ^ n15223 ;
  assign n18173 = n18172 ^ n16139 ;
  assign n18174 = ~n18171 & n18173 ;
  assign n18175 = n18174 ^ n16139 ;
  assign n18176 = n14641 & ~n18175 ;
  assign n19126 = n19125 ^ n18176 ;
  assign n18145 = n15223 ^ n14641 ;
  assign n18177 = n16143 ^ n16138 ;
  assign n18178 = n18177 ^ n16143 ;
  assign n18179 = n16143 ^ n15223 ;
  assign n18180 = n18179 ^ n16143 ;
  assign n18181 = n18178 & ~n18180 ;
  assign n18182 = n18181 ^ n16143 ;
  assign n18183 = ~n18145 & n18182 ;
  assign n18184 = n18183 ^ n16143 ;
  assign n19127 = n19126 ^ n18184 ;
  assign n19120 = n16165 ^ n16130 ;
  assign n19118 = n16147 ^ n16130 ;
  assign n19119 = n19118 ^ n16159 ;
  assign n19121 = n19120 ^ n19119 ;
  assign n19122 = n15223 & n19121 ;
  assign n19123 = n19122 ^ n19120 ;
  assign n19124 = ~n14641 & n19123 ;
  assign n19128 = n19127 ^ n19124 ;
  assign n19117 = n16138 & n16193 ;
  assign n19129 = n19128 ^ n19117 ;
  assign n19135 = n19134 ^ n19129 ;
  assign n19116 = ~n16163 & n16192 ;
  assign n19136 = n19135 ^ n19116 ;
  assign n19137 = ~n16218 & ~n19136 ;
  assign n19139 = n19138 ^ n19137 ;
  assign n19140 = n19139 ^ x113 ;
  assign n16820 = n16819 ^ n16815 ;
  assign n16868 = n16820 ^ n16817 ;
  assign n16877 = n16845 ^ n16824 ;
  assign n16879 = n16878 ^ n16877 ;
  assign n16880 = n16878 ^ n16814 ;
  assign n16881 = n16880 ^ n16878 ;
  assign n16882 = n16879 & ~n16881 ;
  assign n16883 = n16882 ^ n16878 ;
  assign n16884 = ~n16868 & n16883 ;
  assign n17261 = n16884 ^ n13309 ;
  assign n17229 = n16831 ^ n16824 ;
  assign n17230 = ~n16815 & n17229 ;
  assign n17231 = n17230 ^ n16831 ;
  assign n17234 = n17231 ^ n17032 ;
  assign n17235 = n17234 ^ n17231 ;
  assign n17236 = n16815 & n17235 ;
  assign n17237 = n17236 ^ n17231 ;
  assign n17238 = ~n16814 & n17237 ;
  assign n17239 = n17238 ^ n17231 ;
  assign n16863 = n16862 ^ n16831 ;
  assign n16864 = n16863 ^ n16834 ;
  assign n17250 = n16869 ^ n16864 ;
  assign n17251 = ~n16815 & n17250 ;
  assign n17252 = n17251 ^ n16835 ;
  assign n17249 = n16828 ^ n16824 ;
  assign n17253 = n17252 ^ n17249 ;
  assign n17245 = n17032 ^ n16824 ;
  assign n17246 = n17245 ^ n16833 ;
  assign n17247 = n17246 ^ n16828 ;
  assign n17248 = ~n16815 & n17247 ;
  assign n17254 = n17253 ^ n17248 ;
  assign n17255 = ~n16814 & n17254 ;
  assign n17256 = n17255 ^ n17252 ;
  assign n17244 = ~n16868 & n17009 ;
  assign n17257 = n17256 ^ n17244 ;
  assign n17242 = n16812 & n16815 ;
  assign n17240 = n16838 ^ n16812 ;
  assign n17241 = n16814 & n17240 ;
  assign n17243 = n17242 ^ n17241 ;
  assign n17258 = n17257 ^ n17243 ;
  assign n17259 = ~n17239 & ~n17258 ;
  assign n17260 = ~n17044 & n17259 ;
  assign n17262 = n17261 ^ n17260 ;
  assign n17871 = n17262 ^ x100 ;
  assign n16365 = n16110 ^ x122 ;
  assign n16368 = n15308 ^ n15306 ;
  assign n16369 = ~n14784 & n16368 ;
  assign n16370 = n16369 ^ n15308 ;
  assign n16379 = n16370 ^ n12474 ;
  assign n16372 = n16370 ^ n14770 ;
  assign n16371 = n16370 ^ n14789 ;
  assign n16373 = n16372 ^ n16371 ;
  assign n16376 = ~n14784 & n16373 ;
  assign n16377 = n16376 ^ n16372 ;
  assign n16378 = n14680 & ~n16377 ;
  assign n16380 = n16379 ^ n16378 ;
  assign n16381 = n16380 ^ x104 ;
  assign n16338 = n14385 ^ x113 ;
  assign n16346 = n14526 ^ n14460 ;
  assign n16347 = n16346 ^ n14455 ;
  assign n16348 = n16347 ^ n15783 ;
  assign n16349 = ~n14511 & ~n16348 ;
  assign n16350 = n16349 ^ n15783 ;
  assign n16353 = n15781 ^ n14387 ;
  assign n16351 = n14486 ^ n14389 ;
  assign n16352 = n16351 ^ n15781 ;
  assign n16354 = n16353 ^ n16352 ;
  assign n16355 = n16350 & ~n16354 ;
  assign n16356 = n16355 ^ n16353 ;
  assign n16357 = n16356 ^ n14509 ;
  assign n16358 = n16357 ^ n15067 ;
  assign n16359 = n16358 ^ n15786 ;
  assign n16360 = n16359 ^ n15052 ;
  assign n16361 = n16360 ^ n15042 ;
  assign n16362 = n16361 ^ n12542 ;
  assign n16339 = n14478 ^ n14389 ;
  assign n16340 = n15032 ^ n14477 ;
  assign n16341 = n15032 ^ n14478 ;
  assign n16342 = n16341 ^ n15032 ;
  assign n16343 = ~n16340 & ~n16342 ;
  assign n16344 = n16343 ^ n15032 ;
  assign n16345 = n16339 & n16344 ;
  assign n16363 = n16362 ^ n16345 ;
  assign n16364 = n16363 ^ x74 ;
  assign n16386 = n16338 & n16364 ;
  assign n16387 = n16386 ^ n16364 ;
  assign n16388 = n16387 ^ n16338 ;
  assign n16389 = ~n16381 & ~n16388 ;
  assign n16390 = n16365 & n16389 ;
  assign n16391 = n16390 ^ n16389 ;
  assign n16334 = n16029 ^ x107 ;
  assign n16335 = n13546 ^ x81 ;
  assign n16336 = ~n16334 & n16335 ;
  assign n16337 = n16336 ^ n16334 ;
  assign n16660 = n16337 ^ n16335 ;
  assign n16666 = n16391 & n16660 ;
  assign n16667 = n16666 ^ n13145 ;
  assign n16366 = n16365 ^ n16364 ;
  assign n16422 = n16366 & ~n16381 ;
  assign n16423 = n16422 ^ n16365 ;
  assign n16424 = n16338 & n16423 ;
  assign n16425 = n16424 ^ n16386 ;
  assign n16393 = ~n16365 & ~n16381 ;
  assign n16404 = n16387 & n16393 ;
  assign n16394 = n16393 ^ n16365 ;
  assign n16395 = n16394 ^ n16381 ;
  assign n16396 = ~n16388 & ~n16395 ;
  assign n16412 = n16404 ^ n16396 ;
  assign n16411 = n16386 & ~n16395 ;
  assign n16413 = n16412 ^ n16411 ;
  assign n16367 = ~n16338 & ~n16366 ;
  assign n16401 = n16391 ^ n16367 ;
  assign n16397 = n16396 ^ n16388 ;
  assign n16398 = n16397 ^ n16389 ;
  assign n16382 = n16381 ^ n16364 ;
  assign n16383 = n16382 ^ n16365 ;
  assign n16384 = n16383 ^ n16338 ;
  assign n16385 = n16367 & ~n16384 ;
  assign n16392 = n16391 ^ n16385 ;
  assign n16399 = n16398 ^ n16392 ;
  assign n16402 = n16401 ^ n16399 ;
  assign n16403 = n16402 ^ n16398 ;
  assign n16405 = n16404 ^ n16403 ;
  assign n16414 = n16413 ^ n16405 ;
  assign n16410 = n16398 ^ n16395 ;
  assign n16415 = n16414 ^ n16410 ;
  assign n16426 = n16425 ^ n16415 ;
  assign n16400 = n16399 ^ n16387 ;
  assign n16406 = n16405 ^ n16400 ;
  assign n16417 = n16406 ^ n16402 ;
  assign n16427 = n16426 ^ n16417 ;
  assign n16428 = n16427 ^ n16394 ;
  assign n16429 = n16428 ^ n16403 ;
  assign n16444 = n16335 ^ n16334 ;
  assign n16460 = ~n16429 & ~n16444 ;
  assign n16408 = n16388 ^ n16364 ;
  assign n16409 = n16393 & n16408 ;
  assign n16454 = n16409 ^ n16390 ;
  assign n16455 = n16390 ^ n16334 ;
  assign n16456 = n16455 ^ n16390 ;
  assign n16457 = n16454 & ~n16456 ;
  assign n16458 = n16457 ^ n16390 ;
  assign n16459 = ~n16335 & n16458 ;
  assign n16461 = n16460 ^ n16459 ;
  assign n16661 = n16403 & n16660 ;
  assign n16648 = ~n16335 & n16427 ;
  assign n16649 = n16648 ^ n16426 ;
  assign n16652 = n16649 ^ n16409 ;
  assign n16653 = n16652 ^ n16649 ;
  assign n16654 = n16335 & n16653 ;
  assign n16655 = n16654 ^ n16649 ;
  assign n16656 = n16334 & n16655 ;
  assign n16657 = n16656 ^ n16649 ;
  assign n16430 = n16429 ^ n16408 ;
  assign n16416 = n16415 ^ n16409 ;
  assign n16431 = n16430 ^ n16416 ;
  assign n16407 = n16406 ^ n16392 ;
  assign n16432 = n16431 ^ n16407 ;
  assign n16636 = n16432 ^ n16396 ;
  assign n16634 = n16411 ^ n16389 ;
  assign n16446 = n16415 ^ n16399 ;
  assign n16635 = n16634 ^ n16446 ;
  assign n16637 = n16636 ^ n16635 ;
  assign n16638 = ~n16334 & ~n16637 ;
  assign n16639 = n16638 ^ n16636 ;
  assign n16658 = n16657 ^ n16639 ;
  assign n16641 = n16639 ^ n16412 ;
  assign n16640 = n16639 ^ n16424 ;
  assign n16642 = n16641 ^ n16640 ;
  assign n16645 = n16334 & n16642 ;
  assign n16646 = n16645 ^ n16641 ;
  assign n16647 = ~n16335 & n16646 ;
  assign n16659 = n16658 ^ n16647 ;
  assign n16662 = n16661 ^ n16659 ;
  assign n16482 = n16411 ^ n16386 ;
  assign n16437 = n16395 ^ n16365 ;
  assign n16438 = n16386 & ~n16437 ;
  assign n16464 = n16438 ^ n16426 ;
  assign n16483 = n16482 ^ n16464 ;
  assign n16633 = ~n16334 & n16483 ;
  assign n16663 = n16662 ^ n16633 ;
  assign n16627 = n16464 ^ n16438 ;
  assign n16628 = n16438 ^ n16335 ;
  assign n16629 = n16628 ^ n16438 ;
  assign n16630 = n16627 & n16629 ;
  assign n16631 = n16630 ^ n16438 ;
  assign n16632 = ~n16444 & n16631 ;
  assign n16664 = n16663 ^ n16632 ;
  assign n16665 = ~n16461 & ~n16664 ;
  assign n16668 = n16667 ^ n16665 ;
  assign n17872 = n16668 ^ x86 ;
  assign n17398 = n16111 ^ n15968 ;
  assign n17403 = n16072 ^ n15994 ;
  assign n17404 = ~n16030 & ~n17403 ;
  assign n17399 = n16090 ^ n16081 ;
  assign n17400 = n17399 ^ n16084 ;
  assign n17391 = n16116 ^ n16082 ;
  assign n17389 = n16115 ^ n16073 ;
  assign n17390 = n17389 ^ n16118 ;
  assign n17392 = n17391 ^ n17390 ;
  assign n17393 = n17392 ^ n16080 ;
  assign n17401 = n17400 ^ n17393 ;
  assign n17402 = n17401 ^ n16084 ;
  assign n17405 = n17404 ^ n17402 ;
  assign n17406 = ~n16111 & ~n17405 ;
  assign n17407 = n17406 ^ n17401 ;
  assign n17394 = n17393 ^ n17390 ;
  assign n17395 = n16111 & n17394 ;
  assign n17396 = n17395 ^ n17390 ;
  assign n17408 = n17407 ^ n17396 ;
  assign n17409 = ~n17398 & n17408 ;
  assign n17397 = n17396 ^ n15968 ;
  assign n17410 = n17409 ^ n17397 ;
  assign n17411 = n17410 ^ n13452 ;
  assign n17867 = n17411 ^ x101 ;
  assign n16927 = ~n15366 & ~n15433 ;
  assign n16499 = n15422 ^ n15373 ;
  assign n16926 = n15329 & n16499 ;
  assign n16928 = n16927 ^ n16926 ;
  assign n16506 = n15366 ^ n15329 ;
  assign n16929 = n15432 ^ n15376 ;
  assign n16930 = n15329 & n16929 ;
  assign n16931 = n16930 ^ n15377 ;
  assign n16932 = n16931 ^ n15366 ;
  assign n16933 = n16932 ^ n16931 ;
  assign n16934 = n16931 ^ n15417 ;
  assign n16935 = n16934 ^ n16931 ;
  assign n16936 = ~n16933 & ~n16935 ;
  assign n16937 = n16936 ^ n16931 ;
  assign n16938 = n16506 & ~n16937 ;
  assign n16939 = n16938 ^ n16931 ;
  assign n16960 = n15432 ^ n15328 ;
  assign n16961 = ~n15429 & n16960 ;
  assign n16521 = n15383 ^ n15380 ;
  assign n16522 = n16521 ^ n15420 ;
  assign n16947 = n16522 ^ n15327 ;
  assign n16948 = n15429 & ~n16947 ;
  assign n16949 = n15402 & n16948 ;
  assign n16950 = n16949 ^ n15445 ;
  assign n16951 = n16950 ^ n15366 ;
  assign n16952 = n16951 ^ n16950 ;
  assign n16953 = n16950 ^ n15419 ;
  assign n16954 = n16953 ^ n15392 ;
  assign n16955 = n16954 ^ n16950 ;
  assign n16956 = ~n16952 & ~n16955 ;
  assign n16957 = n16956 ^ n16950 ;
  assign n16958 = n16506 & ~n16957 ;
  assign n16959 = n16958 ^ n16950 ;
  assign n16962 = n16961 ^ n16959 ;
  assign n16942 = n15407 ^ n15329 ;
  assign n16943 = n16942 ^ n15407 ;
  assign n16944 = n15408 & ~n16943 ;
  assign n16945 = n16944 ^ n15407 ;
  assign n16946 = n15366 & n16945 ;
  assign n16963 = n16962 ^ n16946 ;
  assign n16964 = n16939 & n16963 ;
  assign n16965 = ~n16928 & n16964 ;
  assign n16523 = n16522 ^ n15390 ;
  assign n16524 = ~n15429 & n16523 ;
  assign n16966 = n16965 ^ n16524 ;
  assign n16967 = n16966 ^ n15368 ;
  assign n16968 = n16967 ^ n13349 ;
  assign n17868 = n16968 ^ x124 ;
  assign n17869 = ~n17867 & n17868 ;
  assign n17870 = n17869 ^ n17867 ;
  assign n17840 = n16304 ^ n13424 ;
  assign n17837 = n15494 & ~n15705 ;
  assign n17833 = n15685 ^ n15646 ;
  assign n17834 = ~n15493 & n17833 ;
  assign n17828 = n15686 ^ n15496 ;
  assign n17827 = n15704 ^ n15646 ;
  assign n17829 = n17828 ^ n17827 ;
  assign n17820 = n15655 ^ n15496 ;
  assign n17821 = n15676 ^ n15494 ;
  assign n17824 = ~n15655 & ~n17821 ;
  assign n17825 = n17824 ^ n15494 ;
  assign n17826 = ~n17820 & n17825 ;
  assign n17830 = n17829 ^ n17826 ;
  assign n17813 = n15686 ^ n15453 ;
  assign n17814 = n17813 ^ n15686 ;
  assign n17817 = ~n15647 & n17814 ;
  assign n17818 = n17817 ^ n15686 ;
  assign n17819 = ~n15493 & ~n17818 ;
  assign n17831 = n17830 ^ n17819 ;
  assign n17806 = n15685 ^ n15635 ;
  assign n17807 = n17806 ^ n15649 ;
  assign n17808 = n15649 ^ n15493 ;
  assign n17809 = n17808 ^ n15649 ;
  assign n17810 = ~n17807 & ~n17809 ;
  assign n17811 = n17810 ^ n15649 ;
  assign n17812 = ~n15453 & n17811 ;
  assign n17832 = n17831 ^ n17812 ;
  assign n17835 = n17834 ^ n17832 ;
  assign n17804 = n15669 ^ n15656 ;
  assign n17805 = ~n15495 & n17804 ;
  assign n17836 = n17835 ^ n17805 ;
  assign n17838 = n17837 ^ n17836 ;
  assign n17839 = ~n15636 & n17838 ;
  assign n17841 = n17840 ^ n17839 ;
  assign n17842 = n17841 ^ x118 ;
  assign n17853 = n14577 ^ n14557 ;
  assign n17857 = n17853 ^ n14559 ;
  assign n17854 = n17853 ^ n14573 ;
  assign n17855 = n17854 ^ n17537 ;
  assign n17856 = ~n14386 & n17855 ;
  assign n17858 = n17857 ^ n17856 ;
  assign n17859 = ~n14538 & n17858 ;
  assign n17849 = n17511 ^ n14559 ;
  assign n17850 = n17849 ^ n14625 ;
  assign n17851 = n17850 ^ n14610 ;
  assign n16238 = n14583 ^ n14538 ;
  assign n16239 = n16238 ^ n14583 ;
  assign n16240 = n14583 ^ n14575 ;
  assign n16241 = n16240 ^ n14583 ;
  assign n16242 = n16239 & n16241 ;
  assign n16243 = n16242 ^ n14583 ;
  assign n16244 = ~n14540 & n16243 ;
  assign n17852 = n17851 ^ n16244 ;
  assign n17860 = n17859 ^ n17852 ;
  assign n17843 = n14576 ^ n14552 ;
  assign n17844 = n14576 ^ n14538 ;
  assign n17845 = n17844 ^ n14576 ;
  assign n17846 = n17843 & ~n17845 ;
  assign n17847 = n17846 ^ n14576 ;
  assign n17848 = n14540 & n17847 ;
  assign n17861 = n17860 ^ n17848 ;
  assign n17862 = ~n14544 & ~n17861 ;
  assign n17863 = n17862 ^ n13382 ;
  assign n17864 = n17863 ^ x68 ;
  assign n17865 = n17842 & ~n17864 ;
  assign n17866 = n17865 ^ n17864 ;
  assign n17884 = n17866 ^ n17842 ;
  assign n17920 = ~n17870 & n17884 ;
  assign n17877 = n17864 ^ n17842 ;
  assign n17878 = ~n17870 & n17877 ;
  assign n17876 = n17865 & ~n17868 ;
  assign n17879 = n17878 ^ n17876 ;
  assign n17921 = n17920 ^ n17879 ;
  assign n17894 = n17870 ^ n17868 ;
  assign n17922 = n17921 ^ n17894 ;
  assign n17918 = n17884 & n17894 ;
  assign n17899 = ~n17866 & n17894 ;
  assign n17919 = n17918 ^ n17899 ;
  assign n17923 = n17922 ^ n17919 ;
  assign n17965 = n17923 ^ n17918 ;
  assign n17885 = n17884 ^ n17864 ;
  assign n17917 = ~n17870 & n17885 ;
  assign n17924 = n17923 ^ n17917 ;
  assign n17886 = n17869 & n17885 ;
  assign n17916 = n17886 ^ n17885 ;
  assign n17925 = n17924 ^ n17916 ;
  assign n17966 = n17965 ^ n17925 ;
  assign n17901 = n17865 & n17869 ;
  assign n17926 = n17925 ^ n17901 ;
  assign n17902 = n17901 ^ n17865 ;
  assign n17903 = n17902 ^ n17876 ;
  assign n17927 = n17926 ^ n17903 ;
  assign n17911 = n17869 & n17884 ;
  assign n17895 = n17894 ^ n17867 ;
  assign n17896 = n17884 & n17895 ;
  assign n17905 = n17901 ^ n17896 ;
  assign n17915 = n17911 ^ n17905 ;
  assign n17928 = n17927 ^ n17915 ;
  assign n17914 = n17911 ^ n17895 ;
  assign n17929 = n17928 ^ n17914 ;
  assign n17967 = n17966 ^ n17929 ;
  assign n17968 = ~n17872 & n17967 ;
  assign n17969 = n17968 ^ n17925 ;
  assign n17970 = ~n17871 & n17969 ;
  assign n18521 = n17872 ^ n17871 ;
  assign n18522 = n17872 ^ n17842 ;
  assign n18523 = n18521 & ~n18522 ;
  assign n18524 = ~n17877 & n18523 ;
  assign n18525 = ~n17870 & n18524 ;
  assign n17873 = ~n17871 & ~n17872 ;
  assign n17880 = n17873 ^ n17872 ;
  assign n17881 = n17880 ^ n17871 ;
  assign n18520 = ~n17881 & n17899 ;
  assign n18526 = n18525 ^ n18520 ;
  assign n19141 = ~n17970 & ~n18526 ;
  assign n18896 = n17873 & n17926 ;
  assign n17958 = n17923 ^ n17872 ;
  assign n17959 = n17958 ^ n17923 ;
  assign n17960 = n17924 & n17959 ;
  assign n17961 = n17960 ^ n17923 ;
  assign n17962 = n17871 & n17961 ;
  assign n18897 = n18896 ^ n17962 ;
  assign n19148 = n18521 ^ n17919 ;
  assign n17897 = n17873 ^ n17871 ;
  assign n19153 = n17886 & ~n17897 ;
  assign n19151 = ~n17880 & n17929 ;
  assign n19149 = n17919 ^ n17903 ;
  assign n19150 = n19149 ^ n17911 ;
  assign n19152 = n19151 ^ n19150 ;
  assign n19154 = n19153 ^ n19152 ;
  assign n19155 = n19148 & n19154 ;
  assign n19156 = n19155 ^ n17919 ;
  assign n17904 = n17903 ^ n17886 ;
  assign n17906 = n17905 ^ n17904 ;
  assign n19159 = n17921 ^ n17906 ;
  assign n19160 = ~n17881 & n19159 ;
  assign n19161 = ~n19156 & n19160 ;
  assign n17909 = n17901 ^ n17886 ;
  assign n17910 = n17909 ^ n17869 ;
  assign n17912 = n17911 ^ n17910 ;
  assign n18889 = n17912 ^ n17864 ;
  assign n18890 = n18889 ^ n17906 ;
  assign n17913 = n17912 ^ n17896 ;
  assign n17930 = n17929 ^ n17913 ;
  assign n17933 = n17930 ^ n17876 ;
  assign n17934 = n17933 ^ n17886 ;
  assign n17935 = n17934 ^ n17899 ;
  assign n18891 = n18890 ^ n17935 ;
  assign n18892 = n17871 & ~n18891 ;
  assign n18893 = n18892 ^ n17912 ;
  assign n18894 = ~n18521 & n18893 ;
  assign n19157 = n19156 ^ n18894 ;
  assign n19162 = n19161 ^ n19157 ;
  assign n19163 = n19162 ^ n18894 ;
  assign n19164 = n17921 ^ n17876 ;
  assign n19165 = ~n17880 & n19164 ;
  assign n19166 = ~n19163 & n19165 ;
  assign n19167 = n19166 ^ n19162 ;
  assign n19142 = n17912 ^ n17879 ;
  assign n19143 = n17879 ^ n17872 ;
  assign n19144 = n19143 ^ n17879 ;
  assign n19145 = n19142 & n19144 ;
  assign n19146 = n19145 ^ n17879 ;
  assign n19147 = ~n17871 & n19146 ;
  assign n19168 = n19167 ^ n19147 ;
  assign n19169 = ~n18897 & ~n19168 ;
  assign n19170 = n19141 & n19169 ;
  assign n19171 = n19170 ^ n13546 ;
  assign n19172 = n19171 ^ x65 ;
  assign n16303 = n16302 ^ x84 ;
  assign n16322 = n15673 ^ n15656 ;
  assign n16323 = ~n15683 & n16322 ;
  assign n16315 = n15654 ^ n15647 ;
  assign n16316 = n16315 ^ n15664 ;
  assign n16317 = n15664 ^ n15453 ;
  assign n16318 = n16317 ^ n15664 ;
  assign n16319 = ~n16316 & ~n16318 ;
  assign n16320 = n16319 ^ n15664 ;
  assign n16321 = ~n15493 & ~n16320 ;
  assign n16324 = n16323 ^ n16321 ;
  assign n16307 = n15665 ^ n15493 ;
  assign n16308 = n15655 ^ n15652 ;
  assign n16309 = n16308 ^ n15668 ;
  assign n16310 = n16309 ^ n15665 ;
  assign n16311 = n16310 ^ n15655 ;
  assign n16312 = n15453 & n16311 ;
  assign n16313 = n16312 ^ n16308 ;
  assign n16314 = n16307 & ~n16313 ;
  assign n16325 = n16324 ^ n16314 ;
  assign n16305 = n15676 ^ n15649 ;
  assign n16306 = ~n15495 & n16305 ;
  assign n16326 = n16325 ^ n16306 ;
  assign n16327 = ~n15693 & n16326 ;
  assign n16328 = ~n15636 & n16327 ;
  assign n16329 = ~n16304 & n16328 ;
  assign n16330 = ~n15738 & n16329 ;
  assign n16331 = n16330 ^ n11502 ;
  assign n16332 = n16331 ^ x78 ;
  assign n16333 = ~n16303 & ~n16332 ;
  assign n16545 = n16333 ^ n16303 ;
  assign n16484 = n16483 ^ n16412 ;
  assign n16485 = n16484 ^ n16407 ;
  assign n16480 = n16431 ^ n16402 ;
  assign n16481 = n16480 ^ n16399 ;
  assign n16486 = n16485 ^ n16481 ;
  assign n16487 = ~n16334 & n16486 ;
  assign n16488 = n16487 ^ n16481 ;
  assign n16489 = n16335 & ~n16488 ;
  assign n16474 = n16336 & n16416 ;
  assign n16471 = n16336 & n16390 ;
  assign n16465 = n16464 ^ n16390 ;
  assign n16466 = n16390 ^ n16335 ;
  assign n16467 = n16466 ^ n16390 ;
  assign n16468 = n16465 & ~n16467 ;
  assign n16469 = n16468 ^ n16390 ;
  assign n16470 = n16334 & n16469 ;
  assign n16472 = n16471 ^ n16470 ;
  assign n16462 = n16426 ^ n16404 ;
  assign n16463 = n16462 ^ n16461 ;
  assign n16473 = n16472 ^ n16463 ;
  assign n16475 = n16474 ^ n16473 ;
  assign n16476 = n16475 ^ n12627 ;
  assign n16445 = n16426 ^ n16409 ;
  assign n16447 = n16446 ^ n16445 ;
  assign n16448 = n16447 ^ n16426 ;
  assign n16449 = n16426 ^ n16334 ;
  assign n16450 = n16449 ^ n16426 ;
  assign n16451 = ~n16448 & n16450 ;
  assign n16452 = n16451 ^ n16426 ;
  assign n16453 = n16444 & n16452 ;
  assign n16477 = n16476 ^ n16453 ;
  assign n16435 = n16404 ^ n16335 ;
  assign n16436 = n16435 ^ n16404 ;
  assign n16441 = ~n16436 & n16438 ;
  assign n16442 = n16441 ^ n16404 ;
  assign n16443 = ~n16334 & n16442 ;
  assign n16478 = n16477 ^ n16443 ;
  assign n16433 = n16432 ^ n16391 ;
  assign n16434 = ~n16337 & n16433 ;
  assign n16479 = n16478 ^ n16434 ;
  assign n16490 = n16489 ^ n16479 ;
  assign n16491 = n16490 ^ x77 ;
  assign n16528 = n15417 ^ n15394 ;
  assign n16529 = n15429 ^ n15329 ;
  assign n16530 = ~n16528 & n16529 ;
  assign n16525 = n16524 ^ n15428 ;
  assign n16507 = n15376 ^ n15369 ;
  assign n16508 = n16507 ^ n15395 ;
  assign n16509 = ~n15329 & ~n16508 ;
  assign n16510 = n16509 ^ n15376 ;
  assign n16519 = n16510 ^ n15449 ;
  assign n16512 = n16510 ^ n15387 ;
  assign n16511 = n16510 ^ n15399 ;
  assign n16513 = n16512 ^ n16511 ;
  assign n16516 = ~n15329 & n16513 ;
  assign n16517 = n16516 ^ n16512 ;
  assign n16518 = n16506 & n16517 ;
  assign n16520 = n16519 ^ n16518 ;
  assign n16526 = n16525 ^ n16520 ;
  assign n16500 = n16499 ^ n15392 ;
  assign n16501 = n15392 ^ n15329 ;
  assign n16502 = n16501 ^ n15392 ;
  assign n16503 = ~n16500 & ~n16502 ;
  assign n16504 = n16503 ^ n15392 ;
  assign n16505 = n15366 & ~n16504 ;
  assign n16527 = n16526 ^ n16505 ;
  assign n16531 = n16530 ^ n16527 ;
  assign n16492 = n15428 ^ n15404 ;
  assign n16493 = n15429 ^ n15328 ;
  assign n16494 = n15429 ^ n15404 ;
  assign n16495 = n16494 ^ n15429 ;
  assign n16496 = n16493 & n16495 ;
  assign n16497 = n16496 ^ n15429 ;
  assign n16498 = ~n16492 & ~n16497 ;
  assign n16532 = n16531 ^ n16498 ;
  assign n16533 = n16532 ^ n15368 ;
  assign n16534 = n16533 ^ n12120 ;
  assign n16535 = n16534 ^ x126 ;
  assign n16536 = ~n16491 & n16535 ;
  assign n16546 = n16536 ^ n16535 ;
  assign n16551 = ~n16545 & n16546 ;
  assign n16237 = n16236 ^ x91 ;
  assign n16259 = n14603 ^ n14579 ;
  assign n16260 = n16259 ^ n14550 ;
  assign n16261 = n16260 ^ n14568 ;
  assign n16262 = n16261 ^ n14603 ;
  assign n16263 = n14538 & n16262 ;
  assign n16264 = n16263 ^ n16259 ;
  assign n16265 = ~n14386 & n16264 ;
  assign n16245 = n14569 ^ n14553 ;
  assign n16251 = n16245 ^ n14582 ;
  assign n16252 = n16251 ^ n14556 ;
  assign n16253 = n16252 ^ n14560 ;
  assign n16254 = n16253 ^ n16245 ;
  assign n16255 = ~n14538 & n16254 ;
  assign n16256 = n16255 ^ n16251 ;
  assign n16257 = n14540 & ~n16256 ;
  assign n16246 = n16245 ^ n14603 ;
  assign n16247 = n16246 ^ n14631 ;
  assign n16248 = n16247 ^ n14613 ;
  assign n16249 = n16248 ^ n16244 ;
  assign n16250 = n16249 ^ n13009 ;
  assign n16258 = n16257 ^ n16250 ;
  assign n16266 = n16265 ^ n16258 ;
  assign n16267 = n16266 ^ x109 ;
  assign n16604 = ~n16237 & n16267 ;
  assign n16605 = n16604 ^ n16237 ;
  assign n16616 = n16551 & ~n16605 ;
  assign n16550 = n16536 & ~n16545 ;
  assign n16552 = n16551 ^ n16550 ;
  assign n16547 = n16546 ^ n16491 ;
  assign n16548 = ~n16545 & n16547 ;
  assign n16549 = n16548 ^ n16545 ;
  assign n16553 = n16552 ^ n16549 ;
  assign n16539 = n16333 ^ n16332 ;
  assign n16541 = ~n16491 & ~n16539 ;
  assign n16540 = n16536 & ~n16539 ;
  assign n16542 = n16541 ^ n16540 ;
  assign n16537 = n16536 ^ n16491 ;
  assign n16538 = n16333 & ~n16537 ;
  assign n16543 = n16542 ^ n16538 ;
  assign n16544 = n16543 ^ n16537 ;
  assign n16554 = n16553 ^ n16544 ;
  assign n16569 = n16554 ^ n16548 ;
  assign n16558 = n16539 ^ n16303 ;
  assign n16559 = n16546 & ~n16558 ;
  assign n16570 = n16569 ^ n16559 ;
  assign n16566 = n16536 & ~n16558 ;
  assign n16567 = n16566 ^ n16548 ;
  assign n16568 = n16567 ^ n16558 ;
  assign n16571 = n16570 ^ n16568 ;
  assign n16606 = n16605 ^ n16267 ;
  assign n16617 = n16606 ^ n16237 ;
  assign n16618 = ~n16571 & n16617 ;
  assign n16619 = ~n16616 & ~n16618 ;
  assign n18312 = n16333 & n16536 ;
  assign n16560 = n16559 ^ n16551 ;
  assign n16556 = n16333 & n16546 ;
  assign n16557 = n16556 ^ n16546 ;
  assign n16561 = n16560 ^ n16557 ;
  assign n18321 = n18312 ^ n16561 ;
  assign n18678 = n16540 ^ n16237 ;
  assign n18679 = n18678 ^ n16540 ;
  assign n18680 = n18321 & ~n18679 ;
  assign n18681 = n18680 ^ n16540 ;
  assign n18682 = ~n16267 & n18681 ;
  assign n18683 = n18682 ^ n16540 ;
  assign n18675 = n16552 & n16604 ;
  assign n18684 = n18683 ^ n18675 ;
  assign n16583 = n16571 ^ n16548 ;
  assign n16580 = n16561 ^ n16333 ;
  assign n16579 = n16541 ^ n16332 ;
  assign n16581 = n16580 ^ n16579 ;
  assign n16582 = n16581 ^ n16547 ;
  assign n16584 = n16583 ^ n16582 ;
  assign n18674 = n16584 ^ n16538 ;
  assign n18685 = n18684 ^ n18674 ;
  assign n16268 = n16267 ^ n16237 ;
  assign n18317 = n16556 ^ n16540 ;
  assign n18342 = n18317 ^ n16559 ;
  assign n18343 = n18342 ^ n16538 ;
  assign n18344 = n16538 ^ n16267 ;
  assign n18345 = n18344 ^ n16538 ;
  assign n18346 = n18343 & ~n18345 ;
  assign n18347 = n18346 ^ n16538 ;
  assign n18348 = n16268 & n18347 ;
  assign n18686 = n18685 ^ n18348 ;
  assign n18309 = ~n16553 & n16617 ;
  assign n18308 = n16559 & n16617 ;
  assign n18310 = n18309 ^ n18308 ;
  assign n18687 = n18686 ^ n18310 ;
  assign n18666 = n16581 ^ n16538 ;
  assign n18667 = n18666 ^ n16550 ;
  assign n18668 = n18667 ^ n16538 ;
  assign n18669 = n16538 ^ n16237 ;
  assign n18670 = n18669 ^ n16538 ;
  assign n18671 = ~n18668 & n18670 ;
  assign n18672 = n18671 ^ n16538 ;
  assign n18673 = n16268 & n18672 ;
  assign n18688 = n18687 ^ n18673 ;
  assign n16595 = n16584 ^ n16542 ;
  assign n18326 = n16595 ^ n16566 ;
  assign n18659 = n18326 ^ n16571 ;
  assign n18660 = n18659 ^ n16570 ;
  assign n18661 = n16570 ^ n16267 ;
  assign n18662 = n18661 ^ n16570 ;
  assign n18663 = ~n18660 & n18662 ;
  assign n18664 = n18663 ^ n16570 ;
  assign n18665 = ~n16237 & n18664 ;
  assign n18689 = n18688 ^ n18665 ;
  assign n18322 = n18321 ^ n16551 ;
  assign n18652 = n16584 ^ n16237 ;
  assign n18653 = n18652 ^ n16584 ;
  assign n18656 = n18322 & n18653 ;
  assign n18657 = n18656 ^ n16584 ;
  assign n18658 = n16267 & n18657 ;
  assign n18690 = n18689 ^ n18658 ;
  assign n16607 = n16569 & n16606 ;
  assign n18691 = n18690 ^ n16607 ;
  assign n18692 = n16619 & ~n18691 ;
  assign n18693 = n18692 ^ n13102 ;
  assign n19114 = n18693 ^ x74 ;
  assign n17324 = n16666 ^ n16474 ;
  assign n17321 = n16385 ^ n16384 ;
  assign n17325 = n17324 ^ n17321 ;
  assign n17318 = n16390 ^ n16388 ;
  assign n17319 = n17318 ^ n16385 ;
  assign n17320 = ~n16335 & ~n17319 ;
  assign n17322 = n17321 ^ n17320 ;
  assign n17323 = n16444 & ~n17322 ;
  assign n17326 = n17325 ^ n17323 ;
  assign n17315 = n16464 ^ n16404 ;
  assign n17316 = n17315 ^ n16387 ;
  assign n17317 = n16336 & n17316 ;
  assign n17327 = n17326 ^ n17317 ;
  assign n17328 = n17327 ^ n16391 ;
  assign n17329 = n17328 ^ n16470 ;
  assign n17330 = n17329 ^ n13575 ;
  assign n17310 = n16391 ^ n16335 ;
  assign n17311 = n17310 ^ n16391 ;
  assign n17312 = n16480 & ~n17311 ;
  assign n17313 = n17312 ^ n16391 ;
  assign n17314 = n16334 & n17313 ;
  assign n17331 = n17330 ^ n17314 ;
  assign n17304 = n16404 ^ n16398 ;
  assign n17305 = ~n16436 & ~n17304 ;
  assign n17306 = n17305 ^ n16404 ;
  assign n17307 = ~n16444 & n17306 ;
  assign n17332 = n17331 ^ n17307 ;
  assign n17976 = n17332 ^ x125 ;
  assign n17977 = n16331 ^ x116 ;
  assign n17978 = ~n17976 & n17977 ;
  assign n17979 = n17978 ^ n17976 ;
  assign n17982 = n17409 ^ n17407 ;
  assign n17983 = n17982 ^ n13797 ;
  assign n17984 = n17983 ^ x102 ;
  assign n17375 = n15103 ^ n15099 ;
  assign n17376 = n17375 ^ n15175 ;
  assign n17371 = n15154 ^ n15102 ;
  assign n17372 = n17371 ^ n15166 ;
  assign n17377 = n17376 ^ n17372 ;
  assign n17378 = ~n15141 & n17377 ;
  assign n17367 = n15099 ^ n15090 ;
  assign n17368 = n15141 & ~n17367 ;
  assign n16721 = n15184 ^ n15166 ;
  assign n17369 = n17368 ^ n16721 ;
  assign n17373 = n17372 ^ n17369 ;
  assign n17379 = n17378 ^ n17373 ;
  assign n17380 = ~n14679 & n17379 ;
  assign n17363 = n15096 ^ n15088 ;
  assign n17364 = n17363 ^ n15105 ;
  assign n17365 = n14679 & ~n17364 ;
  assign n17362 = ~n15105 & ~n15141 ;
  assign n17366 = n17365 ^ n17362 ;
  assign n17370 = n17369 ^ n17366 ;
  assign n17381 = n17380 ^ n17370 ;
  assign n16673 = n15208 ^ n14679 ;
  assign n16714 = n15185 & ~n16673 ;
  assign n16715 = n16714 ^ n16713 ;
  assign n17384 = n17381 ^ n16715 ;
  assign n17385 = n17384 ^ n15219 ;
  assign n17386 = n17385 ^ n13748 ;
  assign n17361 = ~n15101 & n15181 ;
  assign n17387 = n17386 ^ n17361 ;
  assign n17985 = n17387 ^ x85 ;
  assign n17986 = ~n17984 & n17985 ;
  assign n18034 = n17986 ^ n17985 ;
  assign n18062 = n18034 ^ n17984 ;
  assign n18018 = n16266 ^ x75 ;
  assign n18043 = n17985 & n18018 ;
  assign n18044 = n18043 ^ n18034 ;
  assign n17987 = n17986 ^ n17984 ;
  assign n17996 = n16878 ^ n16822 ;
  assign n17997 = n17996 ^ n17005 ;
  assign n17998 = n16815 & n17997 ;
  assign n17999 = n17998 ^ n16827 ;
  assign n18000 = n17999 ^ n16807 ;
  assign n18001 = n18000 ^ n16826 ;
  assign n18002 = n18001 ^ n17999 ;
  assign n18005 = ~n16815 & n18002 ;
  assign n18006 = n18005 ^ n17999 ;
  assign n18007 = n16814 & n18006 ;
  assign n18008 = n18007 ^ n17998 ;
  assign n16840 = n16839 ^ n16831 ;
  assign n17994 = n17024 ^ n16840 ;
  assign n17995 = ~n16819 & n17994 ;
  assign n18009 = n18008 ^ n17995 ;
  assign n17993 = n16816 & n16852 ;
  assign n18010 = n18009 ^ n17993 ;
  assign n17990 = ~n17023 & n17032 ;
  assign n17991 = n17990 ^ n16845 ;
  assign n17992 = n16814 & n17991 ;
  assign n18011 = n18010 ^ n17992 ;
  assign n18012 = n18011 ^ n17043 ;
  assign n18013 = ~n17239 & ~n18012 ;
  assign n16870 = n16869 ^ n16852 ;
  assign n16871 = n16869 ^ n16814 ;
  assign n16872 = n16871 ^ n16869 ;
  assign n16873 = n16870 & ~n16872 ;
  assign n16874 = n16873 ^ n16869 ;
  assign n16875 = n16868 & n16874 ;
  assign n18014 = ~n16875 & ~n16884 ;
  assign n18015 = n18013 & n18014 ;
  assign n18016 = n18015 ^ n13793 ;
  assign n18017 = n18016 ^ x92 ;
  assign n18019 = ~n18017 & ~n18018 ;
  assign n18023 = ~n17987 & n18019 ;
  assign n18058 = n18044 ^ n18023 ;
  assign n18059 = n18058 ^ n18019 ;
  assign n18030 = n18019 ^ n18018 ;
  assign n18039 = ~n18030 & n18034 ;
  assign n18028 = n17986 & ~n18017 ;
  assign n18032 = n18028 ^ n17986 ;
  assign n18031 = n17986 & ~n18030 ;
  assign n18033 = n18032 ^ n18031 ;
  assign n18040 = n18039 ^ n18033 ;
  assign n18046 = n18040 ^ n18028 ;
  assign n18060 = n18059 ^ n18046 ;
  assign n18066 = n18062 ^ n18060 ;
  assign n18064 = ~n18030 & n18062 ;
  assign n18020 = n18019 ^ n18017 ;
  assign n18063 = ~n18020 & n18062 ;
  assign n18065 = n18064 ^ n18063 ;
  assign n18067 = n18066 ^ n18065 ;
  assign n19108 = ~n17979 & n18067 ;
  assign n18038 = ~n18020 & n18034 ;
  assign n18041 = n18040 ^ n18038 ;
  assign n17980 = n17978 ^ n17977 ;
  assign n18056 = n17980 ^ n17976 ;
  assign n19106 = n18041 & n18056 ;
  assign n19102 = ~n17976 & n18060 ;
  assign n17981 = n17980 ^ n17979 ;
  assign n19094 = n18065 ^ n18023 ;
  assign n18035 = n18019 & n18034 ;
  assign n18036 = n18035 ^ n18033 ;
  assign n18037 = n18036 ^ n18034 ;
  assign n18042 = n18041 ^ n18037 ;
  assign n18713 = n18042 ^ n18031 ;
  assign n19092 = n18713 ^ n18028 ;
  assign n19098 = n19094 ^ n19092 ;
  assign n19095 = n19094 ^ n18041 ;
  assign n18045 = n18044 ^ n18035 ;
  assign n18047 = n18046 ^ n18045 ;
  assign n19096 = n19095 ^ n18047 ;
  assign n19097 = n17977 & n19096 ;
  assign n19099 = n19098 ^ n19097 ;
  assign n19100 = n17981 & n19099 ;
  assign n18021 = n18020 ^ n18018 ;
  assign n18022 = ~n17987 & ~n18021 ;
  assign n19093 = n19092 ^ n18022 ;
  assign n19101 = n19100 ^ n19093 ;
  assign n19103 = n19102 ^ n19101 ;
  assign n18072 = n17977 ^ n17976 ;
  assign n18025 = ~n17987 & ~n18020 ;
  assign n19085 = n18025 ^ n18022 ;
  assign n19086 = n19085 ^ n18025 ;
  assign n19087 = n18025 ^ n17977 ;
  assign n19088 = n19087 ^ n18025 ;
  assign n19089 = n19086 & ~n19088 ;
  assign n19090 = n19089 ^ n18025 ;
  assign n19091 = n18072 & n19090 ;
  assign n19104 = n19103 ^ n19091 ;
  assign n19105 = n19104 ^ n18035 ;
  assign n19107 = n19106 ^ n19105 ;
  assign n19109 = n19108 ^ n19107 ;
  assign n19078 = n18035 ^ n17980 ;
  assign n18697 = n18067 ^ n18023 ;
  assign n19079 = n18697 ^ n17979 ;
  assign n19080 = n18697 ^ n17980 ;
  assign n19081 = n19080 ^ n18697 ;
  assign n19082 = n19079 & ~n19081 ;
  assign n19083 = n19082 ^ n18697 ;
  assign n19084 = n19078 & n19083 ;
  assign n19110 = n19109 ^ n19084 ;
  assign n18026 = n18025 ^ n17987 ;
  assign n18024 = n18023 ^ n18022 ;
  assign n18027 = n18026 ^ n18024 ;
  assign n18841 = n17981 & ~n18027 ;
  assign n19111 = n19110 ^ n18841 ;
  assign n19112 = n19111 ^ n13896 ;
  assign n19113 = n19112 ^ x120 ;
  assign n19198 = n19114 ^ n19113 ;
  assign n19199 = ~n19172 & n19198 ;
  assign n19115 = ~n19113 & n19114 ;
  assign n19203 = n19199 ^ n19115 ;
  assign n19204 = n19203 ^ n19113 ;
  assign n19175 = n19115 & ~n19172 ;
  assign n19202 = n19175 ^ n19114 ;
  assign n19205 = n19204 ^ n19202 ;
  assign n19206 = n19140 & n19205 ;
  assign n19207 = n19206 ^ n19205 ;
  assign n19180 = ~n19114 & ~n19140 ;
  assign n19208 = n19207 ^ n19180 ;
  assign n19173 = n19140 & ~n19172 ;
  assign n19186 = n19113 & n19173 ;
  assign n19189 = n19114 & n19186 ;
  assign n19190 = n19189 ^ n19186 ;
  assign n19197 = n19190 ^ n19175 ;
  assign n19200 = n19199 ^ n19197 ;
  assign n19179 = ~n19113 & n19172 ;
  assign n19181 = n19179 & n19180 ;
  assign n19201 = n19200 ^ n19181 ;
  assign n19209 = n19208 ^ n19201 ;
  assign n19210 = n19209 ^ n19206 ;
  assign n19176 = n19175 ^ n19115 ;
  assign n19174 = n19115 & n19173 ;
  assign n19177 = n19176 ^ n19174 ;
  assign n19178 = n19177 ^ n19115 ;
  assign n19266 = n19210 ^ n19178 ;
  assign n19267 = n19075 & n19266 ;
  assign n19268 = n19267 ^ n19210 ;
  assign n17412 = n17411 ^ x76 ;
  assign n17388 = n17387 ^ x93 ;
  assign n17417 = n17412 ^ n17388 ;
  assign n17333 = n17332 ^ x83 ;
  assign n17354 = n15329 & ~n16528 ;
  assign n17351 = n15420 & n16529 ;
  assign n17347 = n15433 ^ n15396 ;
  assign n17348 = n15430 & ~n17347 ;
  assign n17342 = n15404 ^ n15392 ;
  assign n17343 = ~n15367 & ~n17342 ;
  assign n17341 = ~n15419 & n16948 ;
  assign n17344 = n17343 ^ n17341 ;
  assign n17345 = ~n15366 & ~n17344 ;
  assign n17338 = n16939 ^ n16505 ;
  assign n17339 = n17338 ^ n15449 ;
  assign n17340 = n17339 ^ n14451 ;
  assign n17346 = n17345 ^ n17340 ;
  assign n17349 = n17348 ^ n17346 ;
  assign n17336 = n15399 ^ n15373 ;
  assign n17337 = n15428 & n17336 ;
  assign n17350 = n17349 ^ n17337 ;
  assign n17352 = n17351 ^ n17350 ;
  assign n17334 = n16528 ^ n15407 ;
  assign n17335 = ~n15366 & ~n17334 ;
  assign n17353 = n17352 ^ n17335 ;
  assign n17355 = n17354 ^ n17353 ;
  assign n17356 = n17355 ^ x117 ;
  assign n17357 = n17333 & n17356 ;
  assign n17263 = n17262 ^ x94 ;
  assign n17264 = n15795 & n15892 ;
  assign n17265 = n15794 ^ n15793 ;
  assign n17266 = ~n15915 & ~n17265 ;
  assign n17275 = n15924 ^ n15792 ;
  assign n17277 = n15924 ^ n15895 ;
  assign n17276 = n15924 ^ n15903 ;
  assign n17278 = n17277 ^ n17276 ;
  assign n17279 = n17277 ^ n15793 ;
  assign n17280 = n17279 ^ n17277 ;
  assign n17281 = n17278 & ~n17280 ;
  assign n17282 = n17281 ^ n17277 ;
  assign n17283 = ~n17275 & n17282 ;
  assign n17284 = n17283 ^ n15792 ;
  assign n17268 = n15925 ^ n15886 ;
  assign n17070 = n15908 ^ n15895 ;
  assign n17267 = n17070 ^ n15946 ;
  assign n17269 = n17268 ^ n17267 ;
  assign n17270 = n17267 ^ n15793 ;
  assign n17271 = n17270 ^ n17267 ;
  assign n17272 = ~n17269 & ~n17271 ;
  assign n17273 = n17272 ^ n17267 ;
  assign n17274 = ~n15792 & n17273 ;
  assign n17285 = n17284 ^ n17274 ;
  assign n17286 = n17285 ^ n16269 ;
  assign n17287 = ~n15872 & ~n17286 ;
  assign n17288 = ~n17266 & n17287 ;
  assign n17289 = ~n17264 & n17288 ;
  assign n17290 = n15909 ^ n15793 ;
  assign n17291 = n17290 ^ n15909 ;
  assign n17294 = ~n15910 & n17291 ;
  assign n17295 = n17294 ^ n15909 ;
  assign n17296 = n15944 & ~n17295 ;
  assign n17297 = n17289 & ~n17296 ;
  assign n17298 = ~n15952 & n17297 ;
  assign n17299 = ~n16299 & n17298 ;
  assign n17300 = n17299 ^ n14426 ;
  assign n17301 = n17300 ^ x69 ;
  assign n17302 = n17263 & ~n17301 ;
  assign n17303 = n17302 ^ n17263 ;
  assign n17420 = n17303 ^ n17301 ;
  assign n17421 = n17420 ^ n17263 ;
  assign n17426 = n17357 & ~n17421 ;
  assign n17453 = n17426 ^ n17357 ;
  assign n17359 = n17302 & n17357 ;
  assign n17358 = n17303 & n17357 ;
  assign n17360 = n17359 ^ n17358 ;
  assign n17454 = n17453 ^ n17360 ;
  assign n17423 = n17357 ^ n17333 ;
  assign n17431 = n17423 ^ n17356 ;
  assign n17449 = n17420 & ~n17431 ;
  assign n17455 = n17454 ^ n17449 ;
  assign n17418 = n17357 ^ n17356 ;
  assign n17419 = n17302 & n17418 ;
  assign n18461 = n17455 ^ n17419 ;
  assign n18462 = n17455 ^ n17388 ;
  assign n18463 = n18462 ^ n17455 ;
  assign n18464 = n18461 & ~n18463 ;
  assign n18465 = n18464 ^ n17455 ;
  assign n18466 = ~n17417 & n18465 ;
  assign n17424 = ~n17421 & n17423 ;
  assign n17422 = n17418 & ~n17421 ;
  assign n17425 = n17424 ^ n17422 ;
  assign n17427 = n17426 ^ n17425 ;
  assign n18615 = n17427 ^ n17359 ;
  assign n17434 = n17356 ^ n17301 ;
  assign n17435 = n17301 ^ n17263 ;
  assign n17436 = ~n17434 & ~n17435 ;
  assign n17437 = n17436 ^ n17358 ;
  assign n17428 = n17427 ^ n17421 ;
  assign n17429 = n17428 ^ n17424 ;
  assign n17438 = n17437 ^ n17429 ;
  assign n17439 = n17438 ^ n17303 ;
  assign n17432 = n17303 & ~n17431 ;
  assign n17433 = n17432 ^ n17358 ;
  assign n17440 = n17439 ^ n17433 ;
  assign n18614 = n17440 ^ n17358 ;
  assign n18616 = n18615 ^ n18614 ;
  assign n18617 = n18615 ^ n17412 ;
  assign n18618 = n18617 ^ n18615 ;
  assign n18619 = ~n18616 & ~n18618 ;
  assign n18620 = n18619 ^ n18615 ;
  assign n18621 = ~n17388 & n18620 ;
  assign n18622 = n18621 ^ n17359 ;
  assign n17465 = n17418 & n17420 ;
  assign n18613 = n17417 & n17465 ;
  assign n18623 = n18622 ^ n18613 ;
  assign n18634 = n17455 ^ n17429 ;
  assign n17443 = n17302 & ~n17431 ;
  assign n17444 = n17443 ^ n17359 ;
  assign n17442 = n17419 ^ n17302 ;
  assign n17445 = n17444 ^ n17442 ;
  assign n17441 = n17440 ^ n17438 ;
  assign n17446 = n17445 ^ n17441 ;
  assign n18629 = n17446 ^ n17443 ;
  assign n18628 = n17263 & ~n17434 ;
  assign n18630 = n18629 ^ n18628 ;
  assign n18631 = n17388 & n18630 ;
  assign n18632 = n18631 ^ n18628 ;
  assign n18635 = n18634 ^ n18632 ;
  assign n17475 = n17445 ^ n17432 ;
  assign n18626 = n17475 ^ n17358 ;
  assign n17413 = ~n17388 & ~n17412 ;
  assign n17414 = n17413 ^ n17388 ;
  assign n17451 = n17414 & ~n17419 ;
  assign n18627 = n18626 ^ n17451 ;
  assign n18633 = n18632 ^ n18627 ;
  assign n18636 = n18635 ^ n18633 ;
  assign n18637 = ~n17388 & n18636 ;
  assign n18638 = n18637 ^ n18633 ;
  assign n18639 = ~n17417 & ~n18638 ;
  assign n18640 = n18639 ^ n18632 ;
  assign n17457 = n17413 ^ n17412 ;
  assign n17466 = n17465 ^ n17420 ;
  assign n17467 = n17466 ^ n17455 ;
  assign n18624 = n17467 ^ n17422 ;
  assign n18625 = ~n17457 & n18624 ;
  assign n18641 = n18640 ^ n18625 ;
  assign n18642 = ~n18623 & ~n18641 ;
  assign n18643 = ~n18466 & n18642 ;
  assign n18646 = n18643 ^ n14537 ;
  assign n17415 = n17414 ^ n17412 ;
  assign n18644 = ~n17428 & n18643 ;
  assign n18645 = ~n17415 & n18644 ;
  assign n18647 = n18646 ^ n18645 ;
  assign n19076 = n18647 ^ x115 ;
  assign n19220 = n19179 ^ n19172 ;
  assign n19244 = n19220 ^ n19113 ;
  assign n19245 = n19244 ^ n19186 ;
  assign n19246 = n19245 ^ n19200 ;
  assign n19187 = n19186 ^ n19173 ;
  assign n19195 = n19187 ^ n19174 ;
  assign n19269 = n19246 ^ n19195 ;
  assign n19270 = n19246 ^ n19076 ;
  assign n19271 = n19270 ^ n19246 ;
  assign n19272 = n19269 & ~n19271 ;
  assign n19273 = n19272 ^ n19246 ;
  assign n19274 = n19075 & n19273 ;
  assign n19275 = ~n19076 & ~n19274 ;
  assign n19276 = n19268 & n19275 ;
  assign n19277 = n19276 ^ n19274 ;
  assign n19224 = ~n19140 & n19176 ;
  assign n20680 = n19224 ^ n19189 ;
  assign n20681 = n20680 ^ n19181 ;
  assign n20682 = n20681 ^ n20680 ;
  assign n20683 = n20680 ^ n19075 ;
  assign n20684 = n20683 ^ n20680 ;
  assign n20685 = n20682 & n20684 ;
  assign n20686 = n20685 ^ n20680 ;
  assign n20687 = n19076 & n20686 ;
  assign n19221 = n19220 ^ n19205 ;
  assign n19222 = n19140 & n19221 ;
  assign n19223 = n19222 ^ n19221 ;
  assign n20671 = n19223 ^ n19175 ;
  assign n20672 = n20671 ^ n19207 ;
  assign n20673 = n19207 ^ n19076 ;
  assign n20674 = n20673 ^ n19207 ;
  assign n20675 = n20672 & ~n20674 ;
  assign n20676 = n20675 ^ n19207 ;
  assign n20677 = ~n19075 & n20676 ;
  assign n19191 = n19181 ^ n19179 ;
  assign n19192 = n19191 ^ n19176 ;
  assign n19228 = n19222 ^ n19192 ;
  assign n20437 = n19228 ^ n19200 ;
  assign n19237 = ~n19075 & n19076 ;
  assign n19247 = n19224 ^ n19176 ;
  assign n19248 = n19247 ^ n19246 ;
  assign n19249 = n19248 ^ n19209 ;
  assign n19250 = n19237 & n19249 ;
  assign n20669 = n20437 ^ n19250 ;
  assign n20446 = n19210 ^ n19174 ;
  assign n20447 = n19076 & n20446 ;
  assign n20448 = n20447 ^ n19210 ;
  assign n19196 = n19195 ^ n19181 ;
  assign n20451 = n20448 ^ n19196 ;
  assign n20452 = n20451 ^ n20448 ;
  assign n20453 = n19076 & n20452 ;
  assign n20454 = n20453 ^ n20448 ;
  assign n20455 = ~n19075 & n20454 ;
  assign n20456 = n20455 ^ n20448 ;
  assign n20670 = n20669 ^ n20456 ;
  assign n20678 = n20677 ^ n20670 ;
  assign n19077 = n19076 ^ n19075 ;
  assign n20433 = n19247 ^ n19223 ;
  assign n19226 = n19207 ^ n19190 ;
  assign n20436 = n20433 ^ n19226 ;
  assign n20438 = n20437 ^ n20436 ;
  assign n20663 = n20438 ^ n20437 ;
  assign n20664 = n20437 ^ n19075 ;
  assign n20665 = n20664 ^ n20437 ;
  assign n20666 = n20663 & n20665 ;
  assign n20667 = n20666 ^ n20437 ;
  assign n20668 = n19077 & n20667 ;
  assign n20679 = n20678 ^ n20668 ;
  assign n20688 = n20687 ^ n20679 ;
  assign n20689 = ~n19277 & ~n20688 ;
  assign n20690 = n20689 ^ n16266 ;
  assign n20691 = n20690 ^ x77 ;
  assign n18410 = n17425 ^ n17421 ;
  assign n18411 = n17413 & ~n18410 ;
  assign n18422 = n17455 ^ n17425 ;
  assign n18423 = n18422 ^ n17359 ;
  assign n18421 = n17454 ^ n17446 ;
  assign n18424 = n18423 ^ n18421 ;
  assign n18425 = n17388 & n18424 ;
  assign n18426 = n18425 ^ n18421 ;
  assign n18456 = n18426 ^ n17465 ;
  assign n18453 = n17449 ^ n17425 ;
  assign n18454 = ~n17414 & n18453 ;
  assign n18434 = n17475 ^ n17359 ;
  assign n18435 = n17388 & ~n18434 ;
  assign n18436 = n18435 ^ n17359 ;
  assign n18437 = n18436 ^ n17388 ;
  assign n18438 = n18437 ^ n17412 ;
  assign n18439 = n18438 ^ n18436 ;
  assign n18440 = n17440 ^ n17412 ;
  assign n18441 = n18440 ^ n18436 ;
  assign n18445 = n18441 ^ n17412 ;
  assign n18446 = n18445 ^ n18441 ;
  assign n18447 = ~n17438 & ~n18446 ;
  assign n18448 = n18440 & n18447 ;
  assign n18449 = n18448 ^ n18440 ;
  assign n18450 = n18449 ^ n18436 ;
  assign n18451 = ~n18439 & ~n18450 ;
  assign n18452 = n18451 ^ n18437 ;
  assign n18455 = n18454 ^ n18452 ;
  assign n18457 = n18456 ^ n18455 ;
  assign n18419 = n17443 ^ n17358 ;
  assign n18420 = n18419 ^ n17419 ;
  assign n18427 = n18426 ^ n18420 ;
  assign n18428 = n18427 ^ n18426 ;
  assign n18431 = n17388 & n18428 ;
  assign n18432 = n18431 ^ n18426 ;
  assign n18433 = ~n17417 & n18432 ;
  assign n18458 = n18457 ^ n18433 ;
  assign n18412 = n17465 ^ n17433 ;
  assign n18413 = n18412 ^ n17465 ;
  assign n18414 = n17465 ^ n17412 ;
  assign n18415 = n18414 ^ n17465 ;
  assign n18416 = n18413 & ~n18415 ;
  assign n18417 = n18416 ^ n17465 ;
  assign n18418 = ~n17388 & n18417 ;
  assign n18459 = n18458 ^ n18418 ;
  assign n18460 = ~n18411 & ~n18459 ;
  assign n17468 = n17467 ^ n17426 ;
  assign n17469 = n17426 ^ n17388 ;
  assign n17470 = n17469 ^ n17426 ;
  assign n17471 = n17468 & ~n17470 ;
  assign n17472 = n17471 ^ n17426 ;
  assign n17473 = ~n17417 & n17472 ;
  assign n18467 = ~n17473 & ~n18466 ;
  assign n18468 = n18460 & n18467 ;
  assign n18469 = n18468 ^ n15791 ;
  assign n18470 = n18469 ^ x100 ;
  assign n18185 = n18184 ^ n18176 ;
  assign n18146 = n16170 ^ n16157 ;
  assign n18147 = n18146 ^ n16130 ;
  assign n18148 = n18147 ^ n14641 ;
  assign n18149 = ~n18145 & ~n18148 ;
  assign n18150 = n18149 ^ n14641 ;
  assign n18153 = n16166 ^ n16133 ;
  assign n18154 = n18153 ^ n16150 ;
  assign n18151 = n16150 ^ n16133 ;
  assign n18152 = n18151 ^ n18147 ;
  assign n18155 = n18154 ^ n18152 ;
  assign n18156 = ~n18150 & ~n18155 ;
  assign n18157 = n18156 ^ n18154 ;
  assign n18186 = n18185 ^ n18157 ;
  assign n18159 = n16127 ^ n15967 ;
  assign n18160 = n18159 ^ n16138 ;
  assign n18161 = n18160 ^ n16156 ;
  assign n18162 = n18161 ^ n15741 ;
  assign n18163 = n18162 ^ n18157 ;
  assign n16178 = n16177 ^ n16157 ;
  assign n16179 = n16178 ^ n16162 ;
  assign n18158 = n18157 ^ n16179 ;
  assign n18164 = n18163 ^ n18158 ;
  assign n18165 = n18163 ^ n15223 ;
  assign n18166 = n18165 ^ n18163 ;
  assign n18167 = ~n18164 & n18166 ;
  assign n18168 = n18167 ^ n18163 ;
  assign n18169 = ~n18145 & ~n18168 ;
  assign n18187 = n18186 ^ n18169 ;
  assign n16216 = ~n16139 & n16187 ;
  assign n18188 = n18187 ^ n16216 ;
  assign n18189 = n18188 ^ n16175 ;
  assign n18190 = n18189 ^ n15582 ;
  assign n18144 = ~n16161 & n16192 ;
  assign n18191 = n18190 ^ n18144 ;
  assign n18471 = n18191 ^ x109 ;
  assign n18472 = n18470 & n18471 ;
  assign n17963 = ~n17881 & n17923 ;
  assign n17964 = n17963 ^ n17962 ;
  assign n17971 = n17970 ^ n17964 ;
  assign n17949 = n17928 ^ n17895 ;
  assign n17950 = n17949 ^ n17903 ;
  assign n17951 = n17903 ^ n17872 ;
  assign n17952 = n17951 ^ n17903 ;
  assign n17953 = n17950 & n17952 ;
  assign n17954 = n17953 ^ n17903 ;
  assign n17955 = ~n17871 & n17954 ;
  assign n17972 = n17971 ^ n17955 ;
  assign n17973 = n17972 ^ n15492 ;
  assign n17882 = n17879 & ~n17881 ;
  assign n17874 = ~n17870 & n17873 ;
  assign n17875 = ~n17866 & n17874 ;
  assign n17883 = n17882 ^ n17875 ;
  assign n17931 = n17930 ^ n17886 ;
  assign n17932 = n17897 & ~n17931 ;
  assign n17936 = n17912 ^ n17881 ;
  assign n17937 = n17936 ^ n17868 ;
  assign n17938 = n17937 ^ n17881 ;
  assign n17941 = ~n17897 & ~n17938 ;
  assign n17942 = n17941 ^ n17881 ;
  assign n17943 = n17935 & ~n17942 ;
  assign n17944 = ~n17932 & n17943 ;
  assign n17900 = n17899 ^ n17878 ;
  assign n17907 = n17906 ^ n17900 ;
  assign n17908 = ~n17880 & n17907 ;
  assign n17945 = n17944 ^ n17908 ;
  assign n17898 = n17896 & ~n17897 ;
  assign n17946 = n17945 ^ n17898 ;
  assign n17889 = n17886 ^ n17865 ;
  assign n17890 = n17889 ^ n17886 ;
  assign n17891 = ~n17867 & n17890 ;
  assign n17892 = n17891 ^ n17886 ;
  assign n17893 = n17873 & n17892 ;
  assign n17947 = n17946 ^ n17893 ;
  assign n17948 = ~n17883 & ~n17947 ;
  assign n17974 = n17973 ^ n17948 ;
  assign n18272 = n17974 ^ x69 ;
  assign n16986 = n16483 ^ n16446 ;
  assign n16996 = n16986 ^ n16431 ;
  assign n16995 = n16657 ^ n16459 ;
  assign n16997 = n16996 ^ n16995 ;
  assign n16998 = n16997 ^ n16472 ;
  assign n16987 = n16986 ^ n16405 ;
  assign n16988 = n16987 ^ n16414 ;
  assign n16989 = n16988 ^ n16987 ;
  assign n16990 = n16987 ^ n16335 ;
  assign n16991 = n16990 ^ n16987 ;
  assign n16992 = n16989 & ~n16991 ;
  assign n16993 = n16992 ^ n16987 ;
  assign n16994 = n16444 & ~n16993 ;
  assign n16999 = n16998 ^ n16994 ;
  assign n16978 = n16416 ^ n16408 ;
  assign n16979 = n16978 ^ n16335 ;
  assign n16980 = n16979 ^ n16978 ;
  assign n16981 = n16978 ^ n16406 ;
  assign n16982 = n16981 ^ n16978 ;
  assign n16983 = n16980 & ~n16982 ;
  assign n16984 = n16983 ^ n16978 ;
  assign n16985 = n16334 & n16984 ;
  assign n17000 = n16999 ^ n16985 ;
  assign n17001 = n17000 ^ n16666 ;
  assign n17002 = n17001 ^ n16474 ;
  assign n17003 = n17002 ^ n14873 ;
  assign n17004 = n17003 ^ x64 ;
  assign n17053 = n17052 ^ x90 ;
  assign n17054 = ~n17004 & ~n17053 ;
  assign n17055 = n17054 ^ n17004 ;
  assign n17073 = n16277 ^ n15892 ;
  assign n17071 = n17070 ^ n15927 ;
  assign n17072 = ~n15793 & ~n17071 ;
  assign n17074 = n17073 ^ n17072 ;
  assign n17075 = n15944 & n17074 ;
  assign n17068 = n15795 & ~n15914 ;
  assign n17059 = n15906 ^ n15886 ;
  assign n17060 = n17059 ^ n15927 ;
  assign n17061 = ~n15792 & ~n17060 ;
  assign n17065 = n17061 ^ n15892 ;
  assign n17062 = n17061 ^ n15885 ;
  assign n17057 = n15905 ^ n15875 ;
  assign n17058 = ~n15792 & n17057 ;
  assign n17063 = n17062 ^ n17058 ;
  assign n17064 = n15793 & n17063 ;
  assign n17066 = n17065 ^ n17064 ;
  assign n17067 = n17066 ^ n16277 ;
  assign n17069 = n17068 ^ n17067 ;
  assign n17076 = n17075 ^ n17069 ;
  assign n17056 = n15794 & n15871 ;
  assign n17077 = n17076 ^ n17056 ;
  assign n17078 = ~n15958 & ~n17077 ;
  assign n17079 = ~n16271 & n17078 ;
  assign n17080 = ~n16269 & n17079 ;
  assign n17081 = ~n15872 & n17080 ;
  assign n17082 = n17081 ^ n14840 ;
  assign n17083 = n17082 ^ x107 ;
  assign n17084 = n15222 ^ x81 ;
  assign n17085 = ~n17083 & n17084 ;
  assign n17086 = n17085 ^ n17084 ;
  assign n17087 = n17086 ^ n17083 ;
  assign n17088 = n17087 ^ n17084 ;
  assign n17089 = ~n17055 & ~n17088 ;
  assign n17090 = n15451 ^ x104 ;
  assign n17124 = n17123 ^ x66 ;
  assign n17125 = n17090 & n17124 ;
  assign n17126 = n17125 ^ n17090 ;
  assign n17127 = n17126 ^ n17124 ;
  assign n17128 = n17127 ^ n17090 ;
  assign n17129 = n17089 & n17128 ;
  assign n17132 = n17055 ^ n17053 ;
  assign n17175 = n17132 ^ n17004 ;
  assign n17176 = n17085 & ~n17175 ;
  assign n17155 = n17054 & n17087 ;
  assign n17200 = n17176 ^ n17155 ;
  assign n17201 = n17126 & n17200 ;
  assign n17135 = n17085 & ~n17132 ;
  assign n17133 = n17087 & ~n17132 ;
  assign n17160 = n17135 ^ n17133 ;
  assign n17137 = ~n17088 & ~n17132 ;
  assign n17153 = n17137 ^ n17132 ;
  assign n17161 = n17160 ^ n17153 ;
  assign n17162 = n17161 ^ n17137 ;
  assign n17163 = n17162 ^ n17089 ;
  assign n17164 = n17163 ^ n17160 ;
  assign n17157 = n17084 ^ n17083 ;
  assign n17151 = n17088 ^ n17053 ;
  assign n17152 = n17004 & ~n17151 ;
  assign n17158 = n17157 ^ n17152 ;
  assign n17159 = n17158 ^ n17086 ;
  assign n17165 = n17164 ^ n17159 ;
  assign n17149 = n17054 & n17086 ;
  assign n17156 = n17155 ^ n17149 ;
  assign n17166 = n17165 ^ n17156 ;
  assign n17167 = n17166 ^ n17054 ;
  assign n18273 = n17167 ^ n17156 ;
  assign n17177 = n17176 ^ n17175 ;
  assign n17154 = n17153 ^ n17152 ;
  assign n17168 = n17167 ^ n17154 ;
  assign n17169 = n17168 ^ n17156 ;
  assign n17146 = n17083 ^ n17004 ;
  assign n17147 = n17146 ^ n17084 ;
  assign n17148 = ~n17053 & n17147 ;
  assign n17150 = n17149 ^ n17148 ;
  assign n17170 = n17169 ^ n17150 ;
  assign n17171 = n17170 ^ n17154 ;
  assign n17178 = n17177 ^ n17171 ;
  assign n18274 = n18273 ^ n17178 ;
  assign n18275 = n17125 & ~n18274 ;
  assign n17144 = ~n17055 & n17085 ;
  assign n18276 = n17144 ^ n17133 ;
  assign n18277 = n17126 & n18276 ;
  assign n18278 = n17128 & n17137 ;
  assign n17130 = ~n17055 & n17086 ;
  assign n17196 = n17130 ^ n17055 ;
  assign n17145 = n17144 ^ n17089 ;
  assign n17197 = n17196 ^ n17145 ;
  assign n17198 = n17197 ^ n17135 ;
  assign n18292 = n17126 & ~n17198 ;
  assign n17205 = n17128 ^ n17126 ;
  assign n18289 = n17170 ^ n17165 ;
  assign n18290 = n17205 & ~n18289 ;
  assign n18279 = n17130 ^ n17124 ;
  assign n18280 = n17160 ^ n17130 ;
  assign n18281 = n18280 ^ n17164 ;
  assign n18282 = n18281 ^ n18280 ;
  assign n18283 = n18280 ^ n17090 ;
  assign n18284 = n18283 ^ n18280 ;
  assign n18285 = ~n18282 & n18284 ;
  assign n18286 = n18285 ^ n18280 ;
  assign n18287 = n18279 & ~n18286 ;
  assign n18288 = n18287 ^ n17124 ;
  assign n18291 = n18290 ^ n18288 ;
  assign n18293 = n18292 ^ n18291 ;
  assign n18294 = ~n18278 & ~n18293 ;
  assign n18295 = ~n18277 & n18294 ;
  assign n18296 = ~n18275 & n18295 ;
  assign n18297 = n17158 ^ n17124 ;
  assign n18298 = ~n17090 & n18297 ;
  assign n18299 = n18296 & ~n18298 ;
  assign n18300 = ~n17201 & n18299 ;
  assign n18301 = ~n17129 & n18300 ;
  assign n18302 = n18301 ^ n15868 ;
  assign n18303 = n18302 ^ x126 ;
  assign n18304 = n18272 & n18303 ;
  assign n18305 = n18304 ^ n18272 ;
  assign n16969 = n16968 ^ x74 ;
  assign n16626 = n15966 ^ x121 ;
  assign n16885 = n16884 ^ n14713 ;
  assign n16865 = ~n16814 & ~n16864 ;
  assign n16857 = n16856 ^ n16833 ;
  assign n16858 = n16815 & ~n16857 ;
  assign n16853 = n16852 ^ n16809 ;
  assign n16854 = ~n16814 & n16853 ;
  assign n16849 = n16821 ^ n16808 ;
  assign n16855 = n16854 ^ n16849 ;
  assign n16859 = n16858 ^ n16855 ;
  assign n16860 = ~n16848 & n16859 ;
  assign n16829 = n16828 ^ n16817 ;
  assign n16837 = n16836 ^ n16829 ;
  assign n16841 = n16840 ^ n16837 ;
  assign n16842 = n16820 & ~n16841 ;
  assign n16843 = n16842 ^ n16817 ;
  assign n16846 = n16845 ^ n16820 ;
  assign n16847 = n16843 & n16846 ;
  assign n16861 = n16860 ^ n16847 ;
  assign n16866 = n16865 ^ n16861 ;
  assign n16818 = n16813 & n16817 ;
  assign n16867 = n16866 ^ n16818 ;
  assign n16876 = n16867 & ~n16875 ;
  assign n16886 = n16885 ^ n16876 ;
  assign n16887 = n16886 ^ x89 ;
  assign n16670 = n15102 & ~n15181 ;
  assign n16671 = n15162 ^ n15159 ;
  assign n16672 = n15207 & n16671 ;
  assign n16716 = n16715 ^ n15205 ;
  assign n16676 = n15092 ^ n15091 ;
  assign n16677 = n16676 ^ n15175 ;
  assign n16697 = n16677 ^ n15179 ;
  assign n16674 = n15181 ^ n15091 ;
  assign n16681 = n16677 ^ n16674 ;
  assign n16678 = n16677 ^ n15141 ;
  assign n16679 = n16678 ^ n15091 ;
  assign n16682 = n16681 ^ n16679 ;
  assign n16683 = n16682 ^ n16681 ;
  assign n16684 = n16681 ^ n16677 ;
  assign n16685 = n16684 ^ n15091 ;
  assign n16686 = ~n16683 & n16685 ;
  assign n16687 = n16686 ^ n16681 ;
  assign n16690 = n16686 ^ n16685 ;
  assign n16691 = n16676 & n16690 ;
  assign n16692 = n16691 ^ n15092 ;
  assign n16693 = n16692 ^ n16676 ;
  assign n16694 = ~n16687 & n16693 ;
  assign n16695 = n16694 ^ n16691 ;
  assign n16696 = n16695 ^ n15091 ;
  assign n16698 = n16697 ^ n16696 ;
  assign n16699 = n16698 ^ n15179 ;
  assign n16700 = n16673 & ~n16699 ;
  assign n16701 = n16700 ^ n15179 ;
  assign n16702 = ~n15207 & n16701 ;
  assign n16703 = n16702 ^ n15179 ;
  assign n16704 = n15178 ^ n15098 ;
  assign n16705 = n16704 ^ n16703 ;
  assign n16707 = n16706 ^ n16673 ;
  assign n16708 = ~n15098 & n16707 ;
  assign n16709 = n16708 ^ n16673 ;
  assign n16710 = n16705 & n16709 ;
  assign n16711 = n16710 ^ n15098 ;
  assign n16712 = ~n16703 & ~n16711 ;
  assign n16717 = n16716 ^ n16712 ;
  assign n16718 = ~n15209 & n16717 ;
  assign n16719 = ~n16672 & n16718 ;
  assign n16720 = ~n16670 & n16719 ;
  assign n16722 = n16721 ^ n15099 ;
  assign n16723 = n16722 ^ n15174 ;
  assign n16724 = n15174 ^ n15141 ;
  assign n16725 = n16724 ^ n15174 ;
  assign n16726 = ~n16723 & n16725 ;
  assign n16727 = n16726 ^ n15174 ;
  assign n16728 = ~n14679 & ~n16727 ;
  assign n16729 = n16720 & ~n16728 ;
  assign n16730 = ~n15216 & n16729 ;
  assign n16731 = n16730 ^ n14746 ;
  assign n16732 = n16731 ^ x98 ;
  assign n16734 = n14640 ^ x99 ;
  assign n16669 = n16668 ^ x80 ;
  assign n16733 = n16732 ^ n16669 ;
  assign n16899 = n16734 ^ n16733 ;
  assign n16919 = ~n16732 & ~n16899 ;
  assign n16920 = n16919 ^ n16733 ;
  assign n16921 = ~n16887 & ~n16920 ;
  assign n16922 = n16921 ^ n16899 ;
  assign n16917 = n16887 ^ n16733 ;
  assign n16893 = n16734 ^ n16669 ;
  assign n16894 = n16887 ^ n16732 ;
  assign n16895 = n16734 & ~n16894 ;
  assign n16896 = n16895 ^ n16732 ;
  assign n16897 = n16893 & n16896 ;
  assign n16918 = n16917 ^ n16897 ;
  assign n16923 = n16922 ^ n16918 ;
  assign n16924 = ~n16626 & ~n16923 ;
  assign n16925 = n16924 ^ n16922 ;
  assign n16914 = n16734 ^ n16732 ;
  assign n16900 = n16887 ^ n16734 ;
  assign n16907 = n16669 & n16732 ;
  assign n16908 = ~n16900 & n16907 ;
  assign n16909 = n16908 ^ n16895 ;
  assign n16910 = n16909 ^ n16897 ;
  assign n16911 = n16910 ^ n16900 ;
  assign n16903 = n16893 & ~n16900 ;
  assign n16904 = n16903 ^ n16669 ;
  assign n16905 = n16899 & ~n16904 ;
  assign n16906 = n16905 ^ n16669 ;
  assign n16912 = n16911 ^ n16906 ;
  assign n16898 = n16897 ^ n16734 ;
  assign n16913 = n16912 ^ n16898 ;
  assign n16915 = n16914 ^ n16913 ;
  assign n16888 = n16734 & n16887 ;
  assign n16889 = n16888 ^ n16732 ;
  assign n16890 = n16733 & ~n16889 ;
  assign n16891 = n16890 ^ n16732 ;
  assign n16892 = n16626 & n16891 ;
  assign n16916 = n16915 ^ n16892 ;
  assign n16971 = n16925 ^ n16916 ;
  assign n16972 = n16969 & ~n16971 ;
  assign n16973 = n16972 ^ n16925 ;
  assign n18306 = n16973 ^ n15833 ;
  assign n18307 = n18306 ^ x86 ;
  assign n18311 = ~n16616 & ~n18310 ;
  assign n18316 = n16571 ^ n16554 ;
  assign n18318 = n18317 ^ n18316 ;
  assign n18319 = n16267 & ~n18318 ;
  assign n18320 = n18319 ^ n16583 ;
  assign n18313 = n18312 ^ n16581 ;
  assign n18337 = n18320 ^ n18313 ;
  assign n16585 = n16584 ^ n16553 ;
  assign n18332 = n16553 ^ n16267 ;
  assign n18333 = n18332 ^ n16553 ;
  assign n18334 = ~n16585 & n18333 ;
  assign n18335 = n18334 ^ n16553 ;
  assign n18336 = n16268 & ~n18335 ;
  assign n18338 = n18337 ^ n18336 ;
  assign n16620 = n16567 & n16604 ;
  assign n18339 = n18338 ^ n16620 ;
  assign n18324 = n16554 ^ n16550 ;
  assign n18325 = n18324 ^ n18322 ;
  assign n18327 = n18326 ^ n18325 ;
  assign n18328 = ~n16267 & n18327 ;
  assign n18323 = n18322 ^ n18320 ;
  assign n18329 = n18328 ^ n18323 ;
  assign n18330 = ~n16237 & ~n18329 ;
  assign n18340 = n18339 ^ n18330 ;
  assign n16555 = n16554 ^ n16538 ;
  assign n16562 = n16561 ^ n16555 ;
  assign n16563 = ~n16267 & n16562 ;
  assign n16564 = n16563 ^ n16554 ;
  assign n18314 = n18313 ^ n16564 ;
  assign n18315 = n16268 & ~n18314 ;
  assign n18341 = n18340 ^ n18315 ;
  assign n18349 = ~n18341 & ~n18348 ;
  assign n18350 = n18311 & n18349 ;
  assign n18351 = n18350 ^ n15830 ;
  assign n18352 = n18351 ^ x76 ;
  assign n18353 = n18307 & n18352 ;
  assign n18354 = n18353 ^ n18307 ;
  assign n18366 = n18305 & n18354 ;
  assign n18355 = n18354 ^ n18352 ;
  assign n18356 = n18355 ^ n18307 ;
  assign n18357 = n18305 & n18356 ;
  assign n18367 = n18366 ^ n18357 ;
  assign n18364 = n18305 & n18353 ;
  assign n18365 = n18364 ^ n18305 ;
  assign n18368 = n18367 ^ n18365 ;
  assign n18363 = n18304 & n18356 ;
  assign n18369 = n18368 ^ n18363 ;
  assign n18360 = n18304 & n18353 ;
  assign n18361 = n18360 ^ n18357 ;
  assign n18359 = n18272 & ~n18355 ;
  assign n18362 = n18361 ^ n18359 ;
  assign n18370 = n18369 ^ n18362 ;
  assign n18358 = n18357 ^ n18304 ;
  assign n18371 = n18370 ^ n18358 ;
  assign n19447 = n18371 ^ n18364 ;
  assign n19448 = n18472 & n19447 ;
  assign n20412 = n19448 ^ n16302 ;
  assign n18473 = n18472 ^ n18470 ;
  assign n18374 = n18305 ^ n18303 ;
  assign n18383 = n18353 & ~n18374 ;
  assign n18379 = n18374 ^ n18272 ;
  assign n18380 = ~n18355 & n18379 ;
  assign n18378 = n18359 ^ n18355 ;
  assign n18381 = n18380 ^ n18378 ;
  assign n18376 = n18356 & ~n18374 ;
  assign n18372 = n18371 ^ n18368 ;
  assign n18373 = n18372 ^ n18360 ;
  assign n18377 = n18376 ^ n18373 ;
  assign n18382 = n18381 ^ n18377 ;
  assign n18384 = n18383 ^ n18382 ;
  assign n18375 = n18374 ^ n18373 ;
  assign n18385 = n18384 ^ n18375 ;
  assign n18407 = n18385 ^ n18380 ;
  assign n18401 = n18356 & n18379 ;
  assign n18408 = n18407 ^ n18401 ;
  assign n18403 = n18381 ^ n18371 ;
  assign n18398 = n18307 ^ n18303 ;
  assign n18399 = n18272 & n18398 ;
  assign n18386 = n18307 ^ n18272 ;
  assign n18387 = n18386 ^ n18303 ;
  assign n18388 = n18387 ^ n18352 ;
  assign n18389 = n18388 ^ n18272 ;
  assign n18390 = n18389 ^ n18303 ;
  assign n18391 = n18303 ^ n18272 ;
  assign n18394 = ~n18352 & ~n18391 ;
  assign n18395 = n18394 ^ n18272 ;
  assign n18396 = n18390 & ~n18395 ;
  assign n18397 = n18396 ^ n18387 ;
  assign n18400 = n18399 ^ n18397 ;
  assign n18402 = n18401 ^ n18400 ;
  assign n18404 = n18403 ^ n18402 ;
  assign n18405 = n18404 ^ n18385 ;
  assign n18406 = n18405 ^ n18379 ;
  assign n18409 = n18408 ^ n18406 ;
  assign n20031 = n18473 ^ n18409 ;
  assign n20032 = n18472 ^ n18471 ;
  assign n18495 = n18401 ^ n18383 ;
  assign n20033 = n20032 ^ n18495 ;
  assign n20034 = n18495 ^ n18409 ;
  assign n20035 = n20034 ^ n18495 ;
  assign n20036 = ~n20033 & n20035 ;
  assign n20037 = n20036 ^ n18495 ;
  assign n20038 = n20031 & ~n20037 ;
  assign n20039 = n20038 ^ n18473 ;
  assign n20394 = n18401 ^ n18361 ;
  assign n20395 = n20394 ^ n18381 ;
  assign n20396 = n20395 ^ n18399 ;
  assign n20397 = ~n18471 & ~n20396 ;
  assign n20398 = n20397 ^ n20394 ;
  assign n18487 = n18404 ^ n18381 ;
  assign n18503 = n18487 ^ n18385 ;
  assign n18504 = n18472 & ~n18503 ;
  assign n20409 = n20398 ^ n18504 ;
  assign n20400 = n18383 ^ n18357 ;
  assign n18488 = n18487 ^ n18363 ;
  assign n18486 = n18366 ^ n18360 ;
  assign n18489 = n18488 ^ n18486 ;
  assign n20401 = n20400 ^ n18489 ;
  assign n20402 = n20401 ^ n20398 ;
  assign n20399 = n20398 ^ n18397 ;
  assign n20403 = n20402 ^ n20399 ;
  assign n20404 = n20402 ^ n18471 ;
  assign n20405 = n20404 ^ n20402 ;
  assign n20406 = ~n20403 & ~n20405 ;
  assign n20407 = n20406 ^ n20402 ;
  assign n20408 = ~n18470 & ~n20407 ;
  assign n20410 = n20409 ^ n20408 ;
  assign n20411 = ~n20039 & ~n20410 ;
  assign n20413 = n20412 ^ n20411 ;
  assign n20692 = n20413 ^ x83 ;
  assign n17975 = n17974 ^ x77 ;
  assign n16970 = n16969 ^ n16925 ;
  assign n16974 = n16973 ^ n16970 ;
  assign n16975 = n16974 ^ n16916 ;
  assign n16976 = n16975 ^ n14805 ;
  assign n18206 = n16976 ^ x91 ;
  assign n18232 = ~n17975 & ~n18206 ;
  assign n18257 = n18232 ^ n17975 ;
  assign n18258 = n18257 ^ n18206 ;
  assign n16597 = n16560 ^ n16539 ;
  assign n16598 = n16597 ^ n16556 ;
  assign n16599 = n16267 & ~n16598 ;
  assign n16600 = n16599 ^ n16560 ;
  assign n16608 = n16607 ^ n16600 ;
  assign n16594 = n16581 ^ n16556 ;
  assign n16596 = n16595 ^ n16594 ;
  assign n16601 = n16600 ^ n16596 ;
  assign n16593 = ~n16267 & ~n16579 ;
  assign n16602 = n16601 ^ n16593 ;
  assign n16603 = ~n16237 & ~n16602 ;
  assign n16609 = n16608 ^ n16603 ;
  assign n16610 = n16609 ^ n16553 ;
  assign n16592 = ~n16267 & n16566 ;
  assign n16611 = n16610 ^ n16592 ;
  assign n16587 = n16553 ^ n16237 ;
  assign n16588 = n16587 ^ n16553 ;
  assign n16589 = n16584 & n16588 ;
  assign n16590 = n16589 ^ n16553 ;
  assign n16591 = n16268 & ~n16590 ;
  assign n16612 = n16611 ^ n16591 ;
  assign n16613 = n16612 ^ n16550 ;
  assign n16574 = n16550 ^ n16237 ;
  assign n16575 = n16574 ^ n16550 ;
  assign n16576 = ~n16571 & ~n16575 ;
  assign n16577 = n16576 ^ n16550 ;
  assign n16578 = ~n16267 & n16577 ;
  assign n16614 = n16613 ^ n16578 ;
  assign n16565 = n16268 & n16564 ;
  assign n16615 = n16614 ^ n16565 ;
  assign n16621 = n16619 & ~n16620 ;
  assign n16622 = n16615 & n16621 ;
  assign n16623 = n16622 ^ n15140 ;
  assign n18143 = n16623 ^ x78 ;
  assign n18192 = n18191 ^ x67 ;
  assign n18193 = n18143 & ~n18192 ;
  assign n18084 = n18064 ^ n18036 ;
  assign n18083 = n18039 ^ n17986 ;
  assign n18085 = n18084 ^ n18083 ;
  assign n18061 = n18060 ^ n18025 ;
  assign n18068 = n18067 ^ n18061 ;
  assign n18086 = n18085 ^ n18068 ;
  assign n18087 = n17977 & n18086 ;
  assign n18077 = n18067 ^ n18063 ;
  assign n18071 = n18067 ^ n18026 ;
  assign n18073 = n18026 ^ n17977 ;
  assign n18074 = n18072 & ~n18073 ;
  assign n18075 = n18074 ^ n17977 ;
  assign n18076 = ~n18071 & ~n18075 ;
  assign n18078 = n18077 ^ n18076 ;
  assign n18082 = n18078 ^ n18046 ;
  assign n18088 = n18087 ^ n18082 ;
  assign n18089 = n17981 & n18088 ;
  assign n18079 = n18064 ^ n18022 ;
  assign n18080 = n17980 & n18079 ;
  assign n18081 = n18080 ^ n18078 ;
  assign n18090 = n18089 ^ n18081 ;
  assign n18091 = n18090 ^ n18038 ;
  assign n18092 = n18091 ^ n15628 ;
  assign n18057 = n18038 ^ n18027 ;
  assign n18069 = n18068 ^ n18057 ;
  assign n18070 = n18056 & ~n18069 ;
  assign n18093 = n18092 ^ n18070 ;
  assign n18048 = n18047 ^ n18042 ;
  assign n18049 = n18048 ^ n18035 ;
  assign n18029 = n18028 ^ n18027 ;
  assign n18050 = n18049 ^ n18029 ;
  assign n18051 = n18029 ^ n17977 ;
  assign n18052 = n18051 ^ n18029 ;
  assign n18053 = ~n18050 & ~n18052 ;
  assign n18054 = n18053 ^ n18029 ;
  assign n18055 = ~n17981 & ~n18054 ;
  assign n18094 = n18093 ^ n18055 ;
  assign n18095 = n18094 ^ x116 ;
  assign n18117 = n17605 ^ n17584 ;
  assign n18115 = n17644 ^ n17618 ;
  assign n18116 = n18115 ^ n18114 ;
  assign n18118 = n18117 ^ n18116 ;
  assign n18119 = n18118 ^ n18114 ;
  assign n18120 = n17493 & n18119 ;
  assign n18121 = n18120 ^ n18116 ;
  assign n18129 = n18128 ^ n18121 ;
  assign n17676 = n17648 & n17675 ;
  assign n18130 = n18129 ^ n17676 ;
  assign n17594 = ~n17494 & n17593 ;
  assign n17595 = n17594 ^ n17584 ;
  assign n17596 = n17595 ^ n17494 ;
  assign n17597 = n17596 ^ n17595 ;
  assign n17598 = n17595 ^ n17586 ;
  assign n17599 = n17598 ^ n17595 ;
  assign n17600 = ~n17597 & n17599 ;
  assign n17601 = n17600 ^ n17595 ;
  assign n17602 = n17493 & n17601 ;
  assign n17603 = n17602 ^ n17595 ;
  assign n18131 = n18130 ^ n17603 ;
  assign n18132 = n18131 ^ n15543 ;
  assign n17617 = n17616 ^ n17587 ;
  assign n18122 = n18121 ^ n17617 ;
  assign n18123 = n18122 ^ n18114 ;
  assign n18107 = n17644 ^ n17634 ;
  assign n18106 = n17616 ^ n17586 ;
  assign n18108 = n18107 ^ n18106 ;
  assign n18109 = n17493 & n18108 ;
  assign n18124 = n18123 ^ n18109 ;
  assign n18125 = n18124 ^ n17663 ;
  assign n18126 = ~n17615 & ~n18125 ;
  assign n18133 = n18132 ^ n18126 ;
  assign n18103 = n17663 ^ n17589 ;
  assign n18104 = n18103 ^ n17636 ;
  assign n18105 = n17675 & ~n18104 ;
  assign n18134 = n18133 ^ n18105 ;
  assign n18100 = n17648 ^ n17617 ;
  assign n18135 = n18134 ^ n18100 ;
  assign n18098 = n17608 ^ n17585 ;
  assign n18099 = n18098 ^ n17584 ;
  assign n18101 = n18100 ^ n18099 ;
  assign n18102 = n17494 & n18101 ;
  assign n18136 = n18135 ^ n18102 ;
  assign n18137 = n18136 ^ n18134 ;
  assign n18096 = n17589 & ~n17615 ;
  assign n18097 = n17663 & n18096 ;
  assign n18138 = n18137 ^ n18097 ;
  assign n18139 = ~n17493 & n18138 ;
  assign n18140 = n18139 ^ n18136 ;
  assign n18141 = n18140 ^ x101 ;
  assign n18142 = ~n18095 & ~n18141 ;
  assign n18196 = n18142 ^ n18095 ;
  assign n18223 = n18193 & ~n18196 ;
  assign n18197 = n18193 ^ n18143 ;
  assign n18217 = n18142 & n18197 ;
  assign n18245 = n18223 ^ n18217 ;
  assign n18201 = n18142 ^ n18141 ;
  assign n18215 = n18197 & ~n18201 ;
  assign n18246 = n18245 ^ n18215 ;
  assign n18244 = n18142 & n18193 ;
  assign n18247 = n18246 ^ n18244 ;
  assign n18248 = n18247 ^ n18193 ;
  assign n18209 = n18196 ^ n18141 ;
  assign n18212 = n18193 & ~n18209 ;
  assign n18216 = n18215 ^ n18212 ;
  assign n18218 = n18217 ^ n18216 ;
  assign n18259 = n18248 ^ n18218 ;
  assign n18214 = ~n18196 & n18197 ;
  assign n18219 = n18218 ^ n18214 ;
  assign n18213 = n18212 ^ n18197 ;
  assign n18220 = n18219 ^ n18213 ;
  assign n18260 = n18259 ^ n18220 ;
  assign n18261 = ~n18258 & n18260 ;
  assign n20738 = n18261 ^ n16331 ;
  assign n18198 = n18197 ^ n18192 ;
  assign n18228 = n18142 & n18198 ;
  assign n18194 = n18193 ^ n18192 ;
  assign n18202 = ~n18194 & ~n18201 ;
  assign n19351 = n18228 ^ n18202 ;
  assign n18210 = ~n18194 & ~n18209 ;
  assign n19352 = n19351 ^ n18210 ;
  assign n18199 = ~n18196 & n18198 ;
  assign n20720 = n19352 ^ n18199 ;
  assign n20721 = ~n18258 & n20720 ;
  assign n18235 = n18206 ^ n17975 ;
  assign n18224 = n18223 ^ n18214 ;
  assign n18225 = n18224 ^ n18196 ;
  assign n18226 = n18225 ^ n18199 ;
  assign n18221 = n18220 ^ n18212 ;
  assign n18211 = n18210 ^ n18209 ;
  assign n18222 = n18221 ^ n18211 ;
  assign n18227 = n18226 ^ n18222 ;
  assign n18229 = n18228 ^ n18227 ;
  assign n18230 = n18229 ^ n18225 ;
  assign n18231 = n18230 ^ n18198 ;
  assign n19396 = n18231 ^ n18210 ;
  assign n20715 = n19396 ^ n18226 ;
  assign n20716 = ~n18257 & n20715 ;
  assign n20703 = n18192 ^ n18143 ;
  assign n20704 = n20703 ^ n18095 ;
  assign n20705 = n20704 ^ n18141 ;
  assign n20709 = n18141 & ~n18192 ;
  assign n20710 = n20709 ^ n18095 ;
  assign n20711 = n20705 & ~n20710 ;
  assign n20712 = ~n18206 & n20711 ;
  assign n18195 = n18142 & ~n18194 ;
  assign n19393 = n18220 ^ n18195 ;
  assign n20714 = n20712 ^ n19393 ;
  assign n20717 = n20716 ^ n20714 ;
  assign n20718 = n18235 & n20717 ;
  assign n18233 = n18232 ^ n18206 ;
  assign n18268 = n18227 & ~n18233 ;
  assign n20713 = n20712 ^ n18268 ;
  assign n20719 = n20718 ^ n20713 ;
  assign n20722 = n20721 ^ n20719 ;
  assign n20701 = n18222 ^ n18202 ;
  assign n20702 = n18232 & ~n20701 ;
  assign n20723 = n20722 ^ n20702 ;
  assign n20724 = n18260 ^ n18217 ;
  assign n20725 = ~n17975 & n20724 ;
  assign n20726 = n20725 ^ n18223 ;
  assign n20727 = n18235 & n20726 ;
  assign n20728 = ~n20723 & n20727 ;
  assign n20729 = n20728 ^ n20723 ;
  assign n20693 = n18259 ^ n18217 ;
  assign n20696 = n18215 ^ n18206 ;
  assign n20697 = n20696 ^ n18215 ;
  assign n20698 = n20693 & ~n20697 ;
  assign n20699 = n20698 ^ n18215 ;
  assign n20700 = n17975 & n20699 ;
  assign n20730 = n20729 ^ n20700 ;
  assign n20731 = n19396 ^ n18244 ;
  assign n20732 = n18244 ^ n17975 ;
  assign n20733 = n20732 ^ n18244 ;
  assign n20734 = ~n20731 & ~n20733 ;
  assign n20735 = n20734 ^ n18244 ;
  assign n20736 = ~n18235 & n20735 ;
  assign n20737 = ~n20730 & ~n20736 ;
  assign n20739 = n20738 ^ n20737 ;
  assign n20740 = n20739 ^ x109 ;
  assign n20741 = n20692 & ~n20740 ;
  assign n20742 = n20741 ^ n20740 ;
  assign n18846 = ~n17129 & ~n18277 ;
  assign n18568 = ~n17127 & n17165 ;
  assign n18569 = n18568 ^ n18278 ;
  assign n18865 = n17178 ^ n17130 ;
  assign n18866 = n17205 & ~n18865 ;
  assign n17206 = n17124 & n17145 ;
  assign n17207 = n17206 ^ n17089 ;
  assign n17208 = n17207 ^ n17178 ;
  assign n17209 = n17208 ^ n17161 ;
  assign n17210 = n17209 ^ n17197 ;
  assign n17211 = n17210 ^ n17207 ;
  assign n17212 = n17124 & ~n17211 ;
  assign n17213 = n17212 ^ n17208 ;
  assign n17214 = ~n17205 & ~n17213 ;
  assign n17215 = n17214 ^ n17207 ;
  assign n17216 = ~n17127 & n17149 ;
  assign n17217 = ~n17215 & n17216 ;
  assign n17218 = n17217 ^ n17215 ;
  assign n17199 = ~n17127 & ~n17198 ;
  assign n17202 = n17201 ^ n17199 ;
  assign n18863 = n17218 ^ n17202 ;
  assign n18856 = n17176 ^ n17156 ;
  assign n18857 = n18856 ^ n17148 ;
  assign n18858 = n17148 ^ n17090 ;
  assign n18859 = n18858 ^ n17148 ;
  assign n18860 = n18857 & ~n18859 ;
  assign n18861 = n18860 ^ n17148 ;
  assign n18862 = n17124 & n18861 ;
  assign n18864 = n18863 ^ n18862 ;
  assign n18867 = n18866 ^ n18864 ;
  assign n18855 = n17126 & n17167 ;
  assign n18868 = n18867 ^ n18855 ;
  assign n18848 = n17135 ^ n17089 ;
  assign n18847 = n17176 ^ n17162 ;
  assign n18849 = n18848 ^ n18847 ;
  assign n18850 = n18848 ^ n17090 ;
  assign n18851 = n18850 ^ n18848 ;
  assign n18852 = ~n18849 & ~n18851 ;
  assign n18853 = n18852 ^ n18848 ;
  assign n18854 = ~n17205 & n18853 ;
  assign n18869 = n18868 ^ n18854 ;
  assign n18870 = ~n18569 & ~n18869 ;
  assign n18871 = n18846 & n18870 ;
  assign n18872 = n18871 ^ n16029 ;
  assign n19453 = n18872 ^ x104 ;
  assign n19481 = n19074 ^ x81 ;
  assign n18835 = n18048 ^ n18036 ;
  assign n18836 = n17976 & n18835 ;
  assign n18723 = n18697 ^ n18060 ;
  assign n18724 = n17978 & n18723 ;
  assign n18837 = n18836 ^ n18724 ;
  assign n18833 = n18697 ^ n18063 ;
  assign n18834 = n18056 & n18833 ;
  assign n18838 = n18837 ^ n18834 ;
  assign n18704 = n18038 ^ n18022 ;
  assign n18716 = n18704 ^ n18044 ;
  assign n18717 = n18716 ^ n18697 ;
  assign n18832 = ~n17979 & ~n18717 ;
  assign n18839 = n18838 ^ n18832 ;
  assign n18825 = n18060 ^ n18038 ;
  assign n18826 = n18825 ^ n18044 ;
  assign n18827 = n18044 ^ n17976 ;
  assign n18828 = n18827 ^ n18044 ;
  assign n18829 = n18826 & n18828 ;
  assign n18830 = n18829 ^ n18044 ;
  assign n18831 = n17977 & n18830 ;
  assign n18840 = n18839 ^ n18831 ;
  assign n18842 = n18841 ^ n18840 ;
  assign n18843 = ~n18080 & ~n18842 ;
  assign n18844 = n18843 ^ n16110 ;
  assign n19455 = n18844 ^ x90 ;
  assign n17460 = n17454 ^ n17422 ;
  assign n17483 = n17413 & n17460 ;
  assign n19473 = ~n17417 & ~n17444 ;
  assign n19471 = n18455 ^ n18411 ;
  assign n19464 = n17467 ^ n17414 ;
  assign n19465 = n18420 ^ n17457 ;
  assign n19468 = ~n17467 & n19465 ;
  assign n19469 = n19468 ^ n17457 ;
  assign n19470 = ~n19464 & ~n19469 ;
  assign n19472 = n19471 ^ n19470 ;
  assign n19474 = n19473 ^ n19472 ;
  assign n19457 = n18422 ^ n17432 ;
  assign n19456 = n17465 ^ n17436 ;
  assign n19458 = n19457 ^ n19456 ;
  assign n19459 = n19456 ^ n17412 ;
  assign n19460 = n19459 ^ n19456 ;
  assign n19461 = ~n19458 & n19460 ;
  assign n19462 = n19461 ^ n19456 ;
  assign n19463 = n17388 & ~n19462 ;
  assign n19475 = n19474 ^ n19463 ;
  assign n19476 = ~n17483 & n19475 ;
  assign n19477 = n19476 ^ n16363 ;
  assign n19478 = n19477 ^ x107 ;
  assign n19479 = ~n19455 & n19478 ;
  assign n19535 = n19479 ^ n19478 ;
  assign n19536 = ~n19481 & n19535 ;
  assign n18596 = n16923 ^ n16896 ;
  assign n18597 = n18596 ^ n16915 ;
  assign n19482 = n18597 ^ n16908 ;
  assign n19483 = n19482 ^ n16626 ;
  assign n19484 = n19483 ^ n19482 ;
  assign n19485 = n19482 ^ n18597 ;
  assign n19486 = n16906 & ~n19485 ;
  assign n19487 = n19486 ^ n19482 ;
  assign n19488 = n19484 & ~n19487 ;
  assign n19489 = n19488 ^ n19482 ;
  assign n19490 = n16969 & ~n19489 ;
  assign n19491 = n19490 ^ n16969 ;
  assign n18593 = n16919 ^ n16734 ;
  assign n18594 = n16887 & n18593 ;
  assign n18595 = n18594 ^ n16899 ;
  assign n19492 = ~n16969 & n18595 ;
  assign n19493 = n19492 ^ n16908 ;
  assign n19494 = n19493 ^ n16969 ;
  assign n19495 = n19494 ^ n19492 ;
  assign n19496 = n19492 ^ n16911 ;
  assign n19497 = n19496 ^ n19492 ;
  assign n19498 = ~n19495 & ~n19497 ;
  assign n19499 = n19498 ^ n19492 ;
  assign n19500 = n16626 & n19499 ;
  assign n19501 = n19500 ^ n19492 ;
  assign n19502 = ~n19491 & ~n19501 ;
  assign n19503 = n19502 ^ n16380 ;
  assign n19504 = n19503 ^ x72 ;
  assign n19505 = ~n19481 & n19504 ;
  assign n19506 = n19505 ^ n19481 ;
  assign n19480 = n19479 ^ n19455 ;
  assign n19509 = n19480 ^ n19478 ;
  assign n19515 = n19509 ^ n19455 ;
  assign n19516 = ~n19506 & n19515 ;
  assign n19537 = n19536 ^ n19516 ;
  assign n19530 = n19479 & n19505 ;
  assign n19518 = n19479 & ~n19506 ;
  assign n19531 = n19530 ^ n19518 ;
  assign n19507 = n19506 ^ n19504 ;
  assign n19524 = n19507 & n19509 ;
  assign n19528 = n19524 ^ n19509 ;
  assign n19514 = ~n19506 & n19509 ;
  assign n19510 = n19505 ^ n19504 ;
  assign n19511 = n19509 & n19510 ;
  assign n19527 = n19514 ^ n19511 ;
  assign n19529 = n19528 ^ n19527 ;
  assign n19532 = n19531 ^ n19529 ;
  assign n19538 = n19537 ^ n19532 ;
  assign n19539 = n19538 ^ n19515 ;
  assign n19533 = n19532 ^ n19516 ;
  assign n19526 = n19510 & n19515 ;
  assign n19534 = n19533 ^ n19526 ;
  assign n19540 = n19539 ^ n19534 ;
  assign n19508 = ~n19480 & n19507 ;
  assign n19541 = n19540 ^ n19508 ;
  assign n19525 = n19524 ^ n19507 ;
  assign n19542 = n19541 ^ n19525 ;
  assign n20280 = n19542 ^ n19537 ;
  assign n19452 = n19171 ^ x114 ;
  assign n20281 = n19537 ^ n19452 ;
  assign n20282 = n20281 ^ n19537 ;
  assign n20283 = n20280 & ~n20282 ;
  assign n20284 = n20283 ^ n19537 ;
  assign n20285 = n19453 & n20284 ;
  assign n19454 = n19453 ^ n19452 ;
  assign n20123 = n19542 ^ n19526 ;
  assign n20124 = n19542 ^ n19452 ;
  assign n20125 = n20124 ^ n19542 ;
  assign n20126 = n20123 & ~n20125 ;
  assign n20127 = n20126 ^ n19542 ;
  assign n20128 = n19454 & n20127 ;
  assign n20781 = n20285 ^ n20128 ;
  assign n19556 = ~n19452 & n19453 ;
  assign n19588 = n19556 ^ n19454 ;
  assign n19589 = n19588 ^ n19453 ;
  assign n19543 = n19542 ^ n19479 ;
  assign n19544 = n19543 ^ n19531 ;
  assign n19549 = n19544 ^ n19527 ;
  assign n19519 = n19518 ^ n19506 ;
  assign n19517 = n19516 ^ n19514 ;
  assign n19520 = n19519 ^ n19517 ;
  assign n19547 = n19530 ^ n19520 ;
  assign n19548 = n19547 ^ n19529 ;
  assign n19550 = n19549 ^ n19548 ;
  assign n19551 = n19550 ^ n19534 ;
  assign n19546 = n19504 ^ n19481 ;
  assign n19552 = n19551 ^ n19546 ;
  assign n19553 = n19552 ^ n19540 ;
  assign n20769 = n19553 ^ n19520 ;
  assign n20770 = ~n19589 & ~n20769 ;
  assign n19512 = n19511 ^ n19508 ;
  assign n19513 = n19452 & n19512 ;
  assign n20766 = n19544 ^ n19513 ;
  assign n20104 = n19519 ^ n19481 ;
  assign n20105 = n20104 ^ n19538 ;
  assign n20106 = n20105 ^ n19537 ;
  assign n20745 = n20106 ^ n19516 ;
  assign n20755 = n20745 ^ n19529 ;
  assign n20743 = n19548 ^ n19526 ;
  assign n20744 = n20743 ^ n19529 ;
  assign n20746 = n20745 ^ n20744 ;
  assign n20749 = n20743 & ~n20746 ;
  assign n20756 = n20755 ^ n20749 ;
  assign n20747 = n20746 ^ n20745 ;
  assign n20751 = n20749 ^ n20747 ;
  assign n20752 = n19452 & ~n20751 ;
  assign n20753 = n20752 ^ n20745 ;
  assign n20754 = ~n19453 & n20753 ;
  assign n20757 = n20756 ^ n20754 ;
  assign n20767 = n20766 ^ n20757 ;
  assign n19572 = n19529 ^ n19518 ;
  assign n20760 = n20106 ^ n19572 ;
  assign n20758 = n19549 ^ n19514 ;
  assign n20759 = n20758 ^ n19541 ;
  assign n20761 = n20760 ^ n20759 ;
  assign n20762 = ~n19452 & n20761 ;
  assign n20763 = n20762 ^ n20759 ;
  assign n20764 = n19453 & n20763 ;
  assign n20765 = ~n20757 & n20764 ;
  assign n20768 = n20767 ^ n20765 ;
  assign n20771 = n20770 ^ n20768 ;
  assign n20782 = n20781 ^ n20771 ;
  assign n20783 = n20782 ^ n16490 ;
  assign n20772 = n20771 ^ n20766 ;
  assign n20774 = n19514 ^ n19508 ;
  assign n20773 = n20105 ^ n19572 ;
  assign n20775 = n20774 ^ n20773 ;
  assign n20776 = ~n19452 & n20775 ;
  assign n20777 = n20776 ^ n20773 ;
  assign n20778 = ~n20772 & n20777 ;
  assign n20779 = n20778 ^ n20766 ;
  assign n20780 = n19453 & n20779 ;
  assign n20784 = n20783 ^ n20780 ;
  assign n20785 = n20784 ^ x108 ;
  assign n18725 = n18724 ^ n18080 ;
  assign n18726 = n18725 ^ n15365 ;
  assign n18705 = n18704 ^ n18039 ;
  assign n18706 = n18705 ^ n18058 ;
  assign n18707 = n18058 ^ n17976 ;
  assign n18708 = n18707 ^ n18058 ;
  assign n18709 = n18706 & ~n18708 ;
  assign n18710 = n18709 ^ n18058 ;
  assign n18711 = n17977 & n18710 ;
  assign n18695 = n18063 ^ n17979 ;
  assign n18696 = n17981 ^ n17980 ;
  assign n18698 = n18697 ^ n18084 ;
  assign n18699 = n18698 ^ n17980 ;
  assign n18700 = ~n18696 & ~n18699 ;
  assign n18701 = n18700 ^ n17980 ;
  assign n18702 = ~n18695 & ~n18701 ;
  assign n18703 = n18702 ^ n18063 ;
  assign n18712 = n18711 ^ n18703 ;
  assign n18714 = n18713 ^ n17976 ;
  assign n18715 = n18714 ^ n18713 ;
  assign n18718 = ~n17977 & ~n18717 ;
  assign n18719 = n18718 ^ n18713 ;
  assign n18720 = n18715 & n18719 ;
  assign n18721 = n18720 ^ n18713 ;
  assign n18722 = ~n18712 & ~n18721 ;
  assign n18727 = n18726 ^ n18722 ;
  assign n18728 = n18727 ^ x121 ;
  assign n18694 = n18693 ^ x99 ;
  assign n18729 = n18728 ^ n18694 ;
  assign n18598 = n18597 ^ n18595 ;
  assign n18599 = n16969 & ~n18598 ;
  assign n18600 = n18599 ^ n18597 ;
  assign n18602 = n18600 ^ n16911 ;
  assign n18601 = n18600 ^ n16906 ;
  assign n18603 = n18602 ^ n18601 ;
  assign n18606 = ~n16969 & ~n18603 ;
  assign n18607 = n18606 ^ n18602 ;
  assign n18608 = n16626 & n18607 ;
  assign n18609 = n18608 ^ n18600 ;
  assign n18610 = ~n16908 & ~n18609 ;
  assign n18611 = n18610 ^ n15323 ;
  assign n18612 = n18611 ^ x97 ;
  assign n18648 = n18647 ^ x66 ;
  assign n18649 = n18612 & n18648 ;
  assign n18550 = n17871 & n17928 ;
  assign n18542 = n17895 ^ n17886 ;
  assign n18543 = n18542 ^ n17896 ;
  assign n18544 = n18543 ^ n17897 ;
  assign n18545 = ~n17879 & n18544 ;
  assign n18546 = n18545 ^ n17897 ;
  assign n18547 = n17880 ^ n17879 ;
  assign n18548 = n18546 & ~n18547 ;
  assign n18537 = n17874 & n17885 ;
  assign n18530 = n17918 ^ n17912 ;
  assign n18531 = n18530 ^ n17918 ;
  assign n18532 = n17918 ^ n17872 ;
  assign n18533 = n18532 ^ n17918 ;
  assign n18534 = n18531 & n18533 ;
  assign n18535 = n18534 ^ n17918 ;
  assign n18536 = ~n18521 & n18535 ;
  assign n18538 = n18537 ^ n18536 ;
  assign n18528 = n17927 ^ n17879 ;
  assign n18527 = n18526 ^ n17964 ;
  assign n18529 = n18528 ^ n18527 ;
  assign n18539 = n18538 ^ n18529 ;
  assign n18540 = n18539 ^ n17955 ;
  assign n18541 = n18540 ^ n15303 ;
  assign n18549 = n18548 ^ n18541 ;
  assign n18551 = n18550 ^ n18549 ;
  assign n18513 = n17933 ^ n17927 ;
  assign n18511 = n17928 ^ n17927 ;
  assign n18514 = n18513 ^ n18511 ;
  assign n18515 = n18511 ^ n17871 ;
  assign n18516 = n18515 ^ n18511 ;
  assign n18517 = n18514 & ~n18516 ;
  assign n18518 = n18517 ^ n18511 ;
  assign n18519 = ~n17872 & n18518 ;
  assign n18552 = n18551 ^ n18519 ;
  assign n18553 = n18552 ^ x106 ;
  assign n18586 = n17125 & ~n17145 ;
  assign n18579 = n17166 ^ n17154 ;
  assign n18580 = n18579 ^ n18276 ;
  assign n18561 = n17170 ^ n17135 ;
  assign n18581 = n18580 ^ n18561 ;
  assign n18582 = n17124 & n18581 ;
  assign n18577 = n18561 ^ n18276 ;
  assign n18571 = n17165 ^ n17053 ;
  assign n18572 = n18571 ^ n17149 ;
  assign n18573 = n17124 & ~n18572 ;
  assign n18574 = n18573 ^ n17169 ;
  assign n18578 = n18577 ^ n18574 ;
  assign n18583 = n18582 ^ n18578 ;
  assign n18584 = ~n17090 & ~n18583 ;
  assign n18570 = n18569 ^ n17215 ;
  assign n18575 = n18574 ^ n18570 ;
  assign n18576 = n18575 ^ n15266 ;
  assign n18585 = n18584 ^ n18576 ;
  assign n18587 = n18586 ^ n18585 ;
  assign n18560 = n17133 ^ n17126 ;
  assign n18562 = n18561 ^ n17128 ;
  assign n18565 = ~n17133 & n18562 ;
  assign n18566 = n18565 ^ n17128 ;
  assign n18567 = n18560 & n18566 ;
  assign n18588 = n18587 ^ n18567 ;
  assign n18554 = n17200 ^ n17161 ;
  assign n18555 = n17200 ^ n17124 ;
  assign n18556 = n18555 ^ n17200 ;
  assign n18557 = ~n18554 & n18556 ;
  assign n18558 = n18557 ^ n17200 ;
  assign n18559 = ~n17090 & n18558 ;
  assign n18589 = n18588 ^ n18559 ;
  assign n18590 = n18589 ^ x80 ;
  assign n18591 = ~n18553 & n18590 ;
  assign n18592 = n18591 ^ n18553 ;
  assign n18735 = n18592 ^ n18590 ;
  assign n18757 = n18649 & n18735 ;
  assign n18730 = n18649 ^ n18648 ;
  assign n18736 = n18730 & n18735 ;
  assign n18746 = n18736 ^ n18730 ;
  assign n18742 = ~n18592 & n18730 ;
  assign n18733 = n18591 & n18730 ;
  assign n18743 = n18742 ^ n18733 ;
  assign n18747 = n18746 ^ n18743 ;
  assign n18788 = n18757 ^ n18747 ;
  assign n18789 = n18757 ^ n18694 ;
  assign n18790 = n18789 ^ n18757 ;
  assign n18791 = n18788 & n18790 ;
  assign n18792 = n18791 ^ n18757 ;
  assign n18793 = n18729 & n18792 ;
  assign n18731 = n18730 ^ n18612 ;
  assign n18741 = ~n18592 & ~n18731 ;
  assign n20788 = n18741 ^ n18736 ;
  assign n18732 = n18591 & ~n18731 ;
  assign n18748 = n18747 ^ n18732 ;
  assign n18745 = ~n18731 & n18735 ;
  assign n18749 = n18748 ^ n18745 ;
  assign n18750 = n18749 ^ n18736 ;
  assign n18751 = n18750 ^ n18612 ;
  assign n18744 = n18743 ^ n18741 ;
  assign n18752 = n18751 ^ n18744 ;
  assign n20789 = n20788 ^ n18752 ;
  assign n18650 = n18649 ^ n18612 ;
  assign n18651 = ~n18592 & n18650 ;
  assign n18760 = n18744 ^ n18651 ;
  assign n18759 = n18733 ^ n18592 ;
  assign n18761 = n18760 ^ n18759 ;
  assign n18753 = n18752 ^ n18747 ;
  assign n18738 = n18735 ^ n18553 ;
  assign n18739 = n18650 & n18738 ;
  assign n18740 = n18739 ^ n18738 ;
  assign n18754 = n18753 ^ n18740 ;
  assign n18762 = n18761 ^ n18754 ;
  assign n18758 = n18757 ^ n18649 ;
  assign n18763 = n18762 ^ n18758 ;
  assign n20044 = n18763 ^ n18651 ;
  assign n18770 = n18650 & n18735 ;
  assign n20045 = n20044 ^ n18770 ;
  assign n20786 = n20045 ^ n18752 ;
  assign n20787 = n18728 & ~n20786 ;
  assign n20790 = n20789 ^ n20787 ;
  assign n20794 = ~n18694 & ~n20790 ;
  assign n20791 = n20790 ^ n18742 ;
  assign n20792 = n20791 ^ n20045 ;
  assign n20793 = n18728 & ~n20792 ;
  assign n20795 = n20794 ^ n20793 ;
  assign n20796 = n20795 ^ n18742 ;
  assign n20803 = n18762 ^ n18739 ;
  assign n18764 = n18763 ^ n18591 ;
  assign n18734 = n18733 ^ n18732 ;
  assign n18765 = n18764 ^ n18734 ;
  assign n18766 = n18765 ^ n18742 ;
  assign n18805 = ~n18728 & n18766 ;
  assign n18806 = n18805 ^ n18742 ;
  assign n18807 = n18806 ^ n18739 ;
  assign n18808 = n18807 ^ n18806 ;
  assign n18811 = n18728 & n18808 ;
  assign n18812 = n18811 ^ n18806 ;
  assign n18813 = n18694 & n18812 ;
  assign n18814 = n18813 ^ n18806 ;
  assign n18771 = n18770 ^ n18761 ;
  assign n18796 = n18694 & ~n18728 ;
  assign n18803 = n18796 ^ n18694 ;
  assign n18804 = ~n18771 & n18803 ;
  assign n18815 = n18814 ^ n18804 ;
  assign n20804 = n20803 ^ n18815 ;
  assign n20799 = n18748 ^ n18741 ;
  assign n20800 = n20799 ^ n18739 ;
  assign n20801 = n20800 ^ n18762 ;
  assign n20802 = n18728 & n20801 ;
  assign n20805 = n20804 ^ n20802 ;
  assign n20075 = n18765 ^ n18757 ;
  assign n20076 = n18757 ^ n18728 ;
  assign n20077 = n20076 ^ n18757 ;
  assign n20078 = n20075 & ~n20077 ;
  assign n20079 = n20078 ^ n18757 ;
  assign n20080 = n18694 & n20079 ;
  assign n20814 = n20805 ^ n20080 ;
  assign n20806 = n20805 ^ n18815 ;
  assign n20807 = n20806 ^ n20045 ;
  assign n20808 = n20807 ^ n20806 ;
  assign n20809 = n20806 ^ n18728 ;
  assign n20810 = n20809 ^ n20806 ;
  assign n20811 = n20808 & ~n20810 ;
  assign n20812 = n20811 ^ n20806 ;
  assign n20813 = n18694 & n20812 ;
  assign n20815 = n20814 ^ n20813 ;
  assign n20230 = n18745 ^ n18739 ;
  assign n20798 = n18796 & n20230 ;
  assign n20816 = n20815 ^ n20798 ;
  assign n20797 = n18734 & n18803 ;
  assign n20817 = n20816 ^ n20797 ;
  assign n20818 = ~n20796 & ~n20817 ;
  assign n20819 = ~n18793 & n20818 ;
  assign n20820 = n20819 ^ n16534 ;
  assign n20821 = n20820 ^ x94 ;
  assign n20822 = ~n20785 & n20821 ;
  assign n20828 = n20822 ^ n20821 ;
  assign n20829 = ~n20742 & n20828 ;
  assign n20823 = n20822 ^ n20785 ;
  assign n20826 = n20741 & ~n20823 ;
  assign n20859 = n20829 ^ n20826 ;
  assign n20840 = n20741 & n20828 ;
  assign n20824 = n20823 ^ n20821 ;
  assign n20825 = ~n20742 & n20824 ;
  assign n20827 = n20826 ^ n20825 ;
  assign n20830 = n20829 ^ n20827 ;
  assign n20854 = n20840 ^ n20830 ;
  assign n20836 = n20742 ^ n20692 ;
  assign n20851 = n20828 & n20836 ;
  assign n20852 = n20851 ^ n20827 ;
  assign n20853 = n20852 ^ n20828 ;
  assign n20855 = n20854 ^ n20853 ;
  assign n20837 = n20822 & n20836 ;
  assign n20856 = n20855 ^ n20837 ;
  assign n20834 = n20741 ^ n20692 ;
  assign n20850 = ~n20823 & n20834 ;
  assign n20857 = n20856 ^ n20850 ;
  assign n20835 = n20822 & n20834 ;
  assign n20838 = n20837 ^ n20835 ;
  assign n20849 = n20838 ^ n20834 ;
  assign n20858 = n20857 ^ n20849 ;
  assign n20860 = n20859 ^ n20858 ;
  assign n16211 = ~n14641 & n16143 ;
  assign n16208 = ~n16146 & n16192 ;
  assign n16209 = n16208 ^ n16207 ;
  assign n16196 = n16168 ^ n16144 ;
  assign n16197 = n16144 ^ n14641 ;
  assign n16198 = n16197 ^ n16144 ;
  assign n16199 = n16196 & ~n16198 ;
  assign n16200 = n16199 ^ n16144 ;
  assign n16201 = n15223 & n16200 ;
  assign n16210 = n16209 ^ n16201 ;
  assign n16212 = n16211 ^ n16210 ;
  assign n16194 = n16152 ^ n16136 ;
  assign n16195 = n16193 & n16194 ;
  assign n16213 = n16212 ^ n16195 ;
  assign n16189 = n16169 ^ n16162 ;
  assign n16190 = n16189 ^ n16151 ;
  assign n16191 = ~n16188 & ~n16190 ;
  assign n16214 = n16213 ^ n16191 ;
  assign n16176 = n16158 ^ n16130 ;
  assign n16182 = n16176 ^ n15223 ;
  assign n16183 = n16182 ^ n16176 ;
  assign n16184 = n16179 & ~n16183 ;
  assign n16185 = n16184 ^ n16176 ;
  assign n16186 = n14641 & n16185 ;
  assign n16215 = n16214 ^ n16186 ;
  assign n16217 = n16216 ^ n16215 ;
  assign n16219 = n16218 ^ n16217 ;
  assign n16220 = n16219 ^ n16175 ;
  assign n16221 = n16220 ^ n14678 ;
  assign n18904 = n16221 ^ x64 ;
  assign n18925 = n16559 ^ n16554 ;
  assign n18926 = n18925 ^ n16556 ;
  assign n18927 = n18926 ^ n18313 ;
  assign n18928 = n16604 & ~n18927 ;
  assign n18923 = n16617 ^ n16556 ;
  assign n18924 = n18923 ^ n18336 ;
  assign n18929 = n18928 ^ n18924 ;
  assign n18910 = n18308 ^ n16569 ;
  assign n18911 = n18910 ^ n16553 ;
  assign n18914 = n18911 ^ n16566 ;
  assign n18909 = n16559 ^ n16548 ;
  assign n18912 = n16605 & ~n18911 ;
  assign n18913 = ~n18909 & n18912 ;
  assign n18915 = n18914 ^ n18913 ;
  assign n18916 = n18915 ^ n16617 ;
  assign n18917 = n16605 ^ n16543 ;
  assign n18920 = ~n18915 & n18917 ;
  assign n18921 = n18920 ^ n16543 ;
  assign n18922 = ~n18916 & ~n18921 ;
  assign n18930 = n18929 ^ n18922 ;
  assign n18931 = n18930 ^ n18675 ;
  assign n18907 = n18322 ^ n16581 ;
  assign n18908 = ~n16267 & ~n18907 ;
  assign n18932 = n18931 ^ n18908 ;
  assign n18906 = ~n16605 & n18322 ;
  assign n18933 = n18932 ^ n18906 ;
  assign n18934 = ~n18683 & ~n18933 ;
  assign n18935 = n18934 ^ n16607 ;
  assign n18936 = ~n16618 & n18935 ;
  assign n18937 = n18936 ^ n16070 ;
  assign n18938 = n18937 ^ x73 ;
  assign n18942 = ~n18904 & n18938 ;
  assign n18973 = n18942 ^ n18904 ;
  assign n18873 = n18872 ^ x112 ;
  assign n18875 = n17923 ^ n17900 ;
  assign n18876 = n18875 ^ n17904 ;
  assign n18874 = n17934 ^ n17918 ;
  assign n18877 = n18876 ^ n18874 ;
  assign n18878 = n17871 & n18877 ;
  assign n18879 = n18878 ^ n18876 ;
  assign n18888 = n18879 ^ n17883 ;
  assign n18895 = n18894 ^ n18888 ;
  assign n18898 = n18897 ^ n18895 ;
  assign n18899 = n18898 ^ n18538 ;
  assign n18900 = n18899 ^ n17955 ;
  assign n18901 = n18900 ^ n15993 ;
  assign n18881 = n18879 ^ n17926 ;
  assign n18880 = n18879 ^ n17911 ;
  assign n18882 = n18881 ^ n18880 ;
  assign n18883 = n18881 ^ n17872 ;
  assign n18884 = n18883 ^ n18881 ;
  assign n18885 = n18882 & ~n18884 ;
  assign n18886 = n18885 ^ n18881 ;
  assign n18887 = ~n18521 & n18886 ;
  assign n18902 = n18901 ^ n18887 ;
  assign n18903 = n18902 ^ x82 ;
  assign n18943 = n18873 & n18903 ;
  assign n18974 = n18943 ^ n18903 ;
  assign n18975 = ~n18973 & n18974 ;
  assign n18944 = n18942 & n18943 ;
  assign n18979 = n18975 ^ n18944 ;
  assign n18845 = n18844 ^ x105 ;
  assign n17677 = n17676 ^ n15030 ;
  assign n17655 = n17619 ^ n17609 ;
  assign n17649 = n17648 ^ n17586 ;
  assign n17650 = n17586 ^ n17494 ;
  assign n17651 = n17650 ^ n17586 ;
  assign n17652 = n17649 & ~n17651 ;
  assign n17653 = n17652 ^ n17586 ;
  assign n17654 = ~n17493 & n17653 ;
  assign n17656 = n17655 ^ n17654 ;
  assign n17645 = n17644 ^ n17589 ;
  assign n17640 = n17639 ^ n17616 ;
  assign n17635 = n17634 ^ n17589 ;
  assign n17638 = n17637 ^ n17635 ;
  assign n17641 = n17640 ^ n17638 ;
  assign n17642 = ~n17494 & n17641 ;
  assign n17646 = n17645 ^ n17642 ;
  assign n17647 = n17493 & n17646 ;
  assign n17657 = n17656 ^ n17647 ;
  assign n17627 = n17609 ^ n17586 ;
  assign n17628 = n17627 ^ n17609 ;
  assign n17629 = n17609 ^ n17493 ;
  assign n17630 = n17629 ^ n17609 ;
  assign n17631 = n17628 & ~n17630 ;
  assign n17632 = n17631 ^ n17609 ;
  assign n17633 = ~n17494 & n17632 ;
  assign n17658 = n17657 ^ n17633 ;
  assign n17620 = n17619 ^ n17617 ;
  assign n17621 = n17620 ^ n17619 ;
  assign n17622 = n17619 ^ n17493 ;
  assign n17623 = n17622 ^ n17619 ;
  assign n17624 = n17621 & ~n17623 ;
  assign n17625 = n17624 ^ n17619 ;
  assign n17626 = n17615 & n17625 ;
  assign n17659 = n17658 ^ n17626 ;
  assign n17660 = ~n17614 & ~n17659 ;
  assign n17672 = n17671 ^ n17660 ;
  assign n17673 = ~n17603 & n17672 ;
  assign n17678 = n17677 ^ n17673 ;
  assign n18824 = n17678 ^ x123 ;
  assign n19945 = n18845 ^ n18824 ;
  assign n18939 = n18938 ^ n18904 ;
  assign n18961 = n18904 ^ n18873 ;
  assign n18962 = ~n18939 & n18961 ;
  assign n18963 = n18962 ^ n18938 ;
  assign n18905 = n18904 ^ n18903 ;
  assign n18970 = n18905 ^ n18873 ;
  assign n18971 = ~n18963 & ~n18970 ;
  assign n18972 = n18971 ^ n18904 ;
  assign n18976 = n18975 ^ n18972 ;
  assign n18950 = n18873 & ~n18938 ;
  assign n18965 = n18950 ^ n18904 ;
  assign n18966 = n18938 ^ n18903 ;
  assign n18967 = n18965 & n18966 ;
  assign n18954 = n18903 ^ n18873 ;
  assign n18968 = n18967 ^ n18954 ;
  assign n18964 = n18963 ^ n18938 ;
  assign n18969 = n18968 ^ n18964 ;
  assign n18977 = n18976 ^ n18969 ;
  assign n18948 = n18938 ^ n18873 ;
  assign n18949 = n18948 ^ n18905 ;
  assign n18951 = n18950 ^ n18873 ;
  assign n18952 = n18951 ^ n18948 ;
  assign n18953 = n18952 ^ n18873 ;
  assign n18955 = n18954 ^ n18873 ;
  assign n18956 = n18955 ^ n18873 ;
  assign n18957 = ~n18953 & n18956 ;
  assign n18958 = n18957 ^ n18873 ;
  assign n18959 = n18949 & n18958 ;
  assign n18960 = n18959 ^ n18950 ;
  assign n18978 = n18977 ^ n18960 ;
  assign n18940 = ~n18905 & n18939 ;
  assign n18941 = n18873 & n18940 ;
  assign n18991 = n18978 ^ n18941 ;
  assign n18988 = n18942 ^ n18873 ;
  assign n18989 = n18970 & n18988 ;
  assign n18990 = n18989 ^ n18948 ;
  assign n18992 = n18991 ^ n18990 ;
  assign n18987 = n18971 ^ n18940 ;
  assign n18993 = n18992 ^ n18987 ;
  assign n20486 = n18993 ^ n18972 ;
  assign n20487 = n18824 & n20486 ;
  assign n20488 = n20487 ^ n18972 ;
  assign n20489 = n20488 ^ n18990 ;
  assign n20490 = n20489 ^ n18992 ;
  assign n20491 = n20490 ^ n20489 ;
  assign n20492 = n20489 ^ n18824 ;
  assign n20493 = n20492 ^ n20489 ;
  assign n20494 = ~n20491 & ~n20493 ;
  assign n20495 = n20494 ^ n20489 ;
  assign n20496 = n19945 & n20495 ;
  assign n20497 = n20496 ^ n20488 ;
  assign n20498 = ~n18979 & ~n20497 ;
  assign n20499 = n20498 ^ n16236 ;
  assign n20864 = n20499 ^ x126 ;
  assign n20865 = n20860 & n20864 ;
  assign n20866 = n20865 ^ n20858 ;
  assign n20861 = n20860 ^ n20824 ;
  assign n20832 = n20741 & n20822 ;
  assign n20833 = n20832 ^ n20822 ;
  assign n20839 = n20838 ^ n20833 ;
  assign n20843 = n20839 ^ n20830 ;
  assign n20842 = n20826 ^ n20742 ;
  assign n20844 = n20843 ^ n20842 ;
  assign n20845 = n20844 ^ n20832 ;
  assign n20841 = n20840 ^ n20839 ;
  assign n20846 = n20845 ^ n20841 ;
  assign n20831 = n20830 ^ n20740 ;
  assign n20847 = n20846 ^ n20831 ;
  assign n20848 = n20847 ^ n20830 ;
  assign n20862 = n20861 ^ n20848 ;
  assign n20863 = n20862 ^ n20856 ;
  assign n20867 = n20866 ^ n20863 ;
  assign n20868 = n20867 ^ n20832 ;
  assign n20869 = n20868 ^ n20856 ;
  assign n20870 = n20869 ^ n20867 ;
  assign n20871 = n20867 ^ n20864 ;
  assign n20872 = n20871 ^ n20867 ;
  assign n20873 = n20870 & n20872 ;
  assign n20874 = n20873 ^ n20867 ;
  assign n20875 = n20691 & n20874 ;
  assign n20876 = n20875 ^ n20866 ;
  assign n20890 = n20864 ^ n20691 ;
  assign n20905 = n20851 ^ n20835 ;
  assign n20906 = ~n20890 & n20905 ;
  assign n20900 = n20691 & ~n20864 ;
  assign n20901 = n20900 ^ n20890 ;
  assign n20902 = n20858 ^ n20839 ;
  assign n20903 = n20901 & n20902 ;
  assign n20877 = n20857 ^ n20846 ;
  assign n20878 = n20691 & ~n20877 ;
  assign n20879 = n20878 ^ n20857 ;
  assign n20892 = n20879 ^ n20826 ;
  assign n20891 = n20879 ^ n20854 ;
  assign n20893 = n20892 ^ n20891 ;
  assign n20896 = ~n20691 & n20893 ;
  assign n20897 = n20896 ^ n20892 ;
  assign n20898 = ~n20890 & n20897 ;
  assign n20880 = ~n20823 & n20836 ;
  assign n20881 = n20880 ^ n20691 ;
  assign n20882 = n20881 ^ n20880 ;
  assign n20883 = n20847 ^ n20844 ;
  assign n20884 = n20883 ^ n20840 ;
  assign n20885 = n20884 ^ n20880 ;
  assign n20886 = n20882 & ~n20885 ;
  assign n20887 = n20886 ^ n20880 ;
  assign n20888 = n20864 & n20887 ;
  assign n20889 = n20888 ^ n20879 ;
  assign n20899 = n20898 ^ n20889 ;
  assign n20904 = n20903 ^ n20899 ;
  assign n20907 = n20906 ^ n20904 ;
  assign n20908 = ~n20876 & ~n20907 ;
  assign n20909 = n20880 ^ n20858 ;
  assign n20910 = n20858 ^ n20691 ;
  assign n20911 = n20910 ^ n20858 ;
  assign n20912 = n20909 & ~n20911 ;
  assign n20913 = n20912 ^ n20858 ;
  assign n20914 = ~n20864 & n20913 ;
  assign n20915 = n20908 & ~n20914 ;
  assign n20916 = n20915 ^ n16623 ;
  assign n20917 = n20916 ^ x83 ;
  assign n18476 = n18471 ^ n18470 ;
  assign n18479 = n18376 ^ n18366 ;
  assign n18480 = n18479 ^ n18376 ;
  assign n18481 = ~n18471 & n18480 ;
  assign n18482 = n18481 ^ n18376 ;
  assign n18483 = n18476 & n18482 ;
  assign n18484 = n18483 ^ n18376 ;
  assign n18474 = n18473 ^ n18471 ;
  assign n18475 = n18409 & ~n18474 ;
  assign n18485 = n18484 ^ n18475 ;
  assign n19406 = n18408 & n18470 ;
  assign n19407 = n19406 ^ n18401 ;
  assign n19408 = n19407 ^ n18363 ;
  assign n19409 = n19408 ^ n18364 ;
  assign n19410 = n19409 ^ n19407 ;
  assign n19411 = n19407 ^ n18470 ;
  assign n19412 = n19411 ^ n19407 ;
  assign n19413 = n19410 & ~n19412 ;
  assign n19414 = n19413 ^ n19407 ;
  assign n19415 = ~n18471 & n19414 ;
  assign n19416 = n19415 ^ n19407 ;
  assign n19417 = ~n18485 & ~n19416 ;
  assign n19424 = n18383 ^ n18371 ;
  assign n19425 = n19424 ^ n18404 ;
  assign n19426 = ~n18470 & n19425 ;
  assign n19427 = n19426 ^ n18487 ;
  assign n19428 = ~n18471 & ~n19427 ;
  assign n19429 = n19428 ^ n18362 ;
  assign n19421 = n18369 & n18471 ;
  assign n19422 = n19421 ^ n18362 ;
  assign n19423 = ~n18476 & n19422 ;
  assign n19430 = n19429 ^ n19423 ;
  assign n19433 = n18405 & n18471 ;
  assign n19434 = n19433 ^ n18401 ;
  assign n19435 = ~n18470 & n19434 ;
  assign n19436 = n19435 ^ n18401 ;
  assign n19437 = ~n19430 & n19436 ;
  assign n19438 = n19437 ^ n19430 ;
  assign n19439 = n18380 ^ n18366 ;
  assign n19442 = ~n18471 & n19439 ;
  assign n19443 = n19442 ^ n18366 ;
  assign n19444 = ~n18470 & n19443 ;
  assign n19445 = ~n19438 & ~n19444 ;
  assign n19446 = n19417 & n19445 ;
  assign n19449 = n19448 ^ n19446 ;
  assign n19450 = n19449 ^ n17082 ;
  assign n19451 = n19450 ^ x104 ;
  assign n19590 = n19541 & ~n19589 ;
  assign n19521 = n19520 ^ n19513 ;
  assign n19522 = ~n19454 & ~n19521 ;
  assign n19523 = n19522 ^ n19520 ;
  assign n19557 = n19542 & n19556 ;
  assign n19558 = n19557 ^ n19526 ;
  assign n19559 = n19453 & n19558 ;
  assign n19554 = n19454 & n19553 ;
  assign n19545 = n19544 ^ n19526 ;
  assign n19555 = n19554 ^ n19545 ;
  assign n19560 = n19559 ^ n19555 ;
  assign n19561 = n19560 ^ n19453 ;
  assign n19564 = n19518 ^ n19514 ;
  assign n19565 = n19564 ^ n19452 ;
  assign n19566 = ~n19560 & n19565 ;
  assign n19567 = n19566 ^ n19452 ;
  assign n19568 = ~n19561 & ~n19567 ;
  assign n19569 = n19568 ^ n19453 ;
  assign n19577 = n19504 ^ n19478 ;
  assign n19574 = n19553 ^ n19511 ;
  assign n19575 = n19574 ^ n19524 ;
  assign n19576 = n19575 ^ n19538 ;
  assign n19578 = n19577 ^ n19576 ;
  assign n19573 = n19572 ^ n19537 ;
  assign n19579 = n19578 ^ n19573 ;
  assign n19580 = n19452 & n19579 ;
  assign n19581 = n19580 ^ n19573 ;
  assign n19582 = n19581 ^ n19529 ;
  assign n19570 = n19530 ^ n19505 ;
  assign n19571 = ~n19452 & n19570 ;
  assign n19583 = n19582 ^ n19571 ;
  assign n19584 = ~n19453 & n19583 ;
  assign n19585 = n19584 ^ n19581 ;
  assign n19586 = n19569 & ~n19585 ;
  assign n19587 = n19523 & n19586 ;
  assign n19591 = n19590 ^ n19587 ;
  assign n19592 = n19591 ^ n17003 ;
  assign n19593 = n19592 ^ x97 ;
  assign n19596 = n18611 ^ x75 ;
  assign n19700 = n18302 ^ x93 ;
  assign n19635 = n18469 ^ x125 ;
  assign n19650 = n18177 ^ n16147 ;
  assign n19649 = n18170 ^ n16136 ;
  assign n19651 = n19650 ^ n19649 ;
  assign n19652 = n19649 ^ n15223 ;
  assign n19653 = n19652 ^ n19649 ;
  assign n19654 = n19651 & ~n19653 ;
  assign n19655 = n19654 ^ n19649 ;
  assign n19656 = ~n14641 & n19655 ;
  assign n19657 = n19656 ^ n16208 ;
  assign n19647 = n16170 ^ n16133 ;
  assign n19648 = n16187 & ~n19647 ;
  assign n19658 = n19657 ^ n19648 ;
  assign n19646 = n16166 & ~n16188 ;
  assign n19659 = n19658 ^ n19646 ;
  assign n19639 = n16177 ^ n16165 ;
  assign n19636 = n18159 ^ n15452 ;
  assign n19637 = n19636 ^ n15741 ;
  assign n19638 = n19637 ^ n16155 ;
  assign n19640 = n19639 ^ n19638 ;
  assign n19641 = n19638 ^ n15223 ;
  assign n19642 = n19641 ^ n19638 ;
  assign n19643 = ~n19640 & ~n19642 ;
  assign n19644 = n19643 ^ n19638 ;
  assign n19645 = n14641 & ~n19644 ;
  assign n19660 = n19659 ^ n19645 ;
  assign n19661 = n19660 ^ n19116 ;
  assign n19662 = ~n16216 & ~n19661 ;
  assign n19663 = n19662 ^ n16218 ;
  assign n19664 = ~n16159 & n19663 ;
  assign n19665 = n19664 ^ n16803 ;
  assign n19666 = n19665 ^ x124 ;
  assign n19667 = ~n19635 & n19666 ;
  assign n19597 = n18727 ^ x68 ;
  assign n19615 = n18107 ^ n17588 ;
  assign n19612 = n17639 ^ n17608 ;
  assign n19613 = n19612 ^ n18103 ;
  assign n19608 = n17605 ^ n17593 ;
  assign n19605 = n17637 ^ n17608 ;
  assign n19606 = n19605 ^ n17593 ;
  assign n19607 = ~n17494 & n19606 ;
  assign n19609 = n19608 ^ n19607 ;
  assign n19610 = n19609 ^ n17640 ;
  assign n19614 = n19613 ^ n19610 ;
  assign n19616 = n19615 ^ n19614 ;
  assign n19617 = n19616 ^ n19610 ;
  assign n19618 = n17493 & ~n19617 ;
  assign n19619 = n19618 ^ n19614 ;
  assign n19620 = n17615 & ~n19619 ;
  assign n19611 = n19610 ^ n17654 ;
  assign n19621 = n19620 ^ n19611 ;
  assign n19622 = n19621 ^ n17654 ;
  assign n19623 = n17663 ^ n17585 ;
  assign n19624 = n19623 ^ n17609 ;
  assign n19625 = n19051 & ~n19624 ;
  assign n19626 = ~n19622 & n19625 ;
  assign n19627 = n19626 ^ n19621 ;
  assign n19604 = n17588 & n17674 ;
  assign n19628 = n19627 ^ n19604 ;
  assign n19598 = n18107 ^ n17618 ;
  assign n19599 = n17618 ^ n17494 ;
  assign n19600 = n19599 ^ n17618 ;
  assign n19601 = n19598 & n19600 ;
  assign n19602 = n19601 ^ n17618 ;
  assign n19603 = ~n17493 & n19602 ;
  assign n19629 = n19628 ^ n19603 ;
  assign n19630 = ~n17676 & ~n19629 ;
  assign n19631 = n19630 ^ n16775 ;
  assign n19632 = n19631 ^ x110 ;
  assign n19633 = ~n19597 & n19632 ;
  assign n19634 = n19633 ^ n19632 ;
  assign n19676 = n19634 ^ n19597 ;
  assign n19682 = n19667 & n19676 ;
  assign n19678 = n19633 & ~n19635 ;
  assign n19670 = n19633 & n19667 ;
  assign n19679 = n19678 ^ n19670 ;
  assign n19668 = n19667 ^ n19635 ;
  assign n19677 = ~n19668 & n19676 ;
  assign n19680 = n19679 ^ n19677 ;
  assign n19683 = n19682 ^ n19680 ;
  assign n19669 = n19634 & ~n19668 ;
  assign n19675 = n19669 ^ n19668 ;
  assign n19681 = n19680 ^ n19675 ;
  assign n19684 = n19683 ^ n19681 ;
  assign n19672 = n19634 & n19667 ;
  assign n19671 = n19670 ^ n19669 ;
  assign n19673 = n19672 ^ n19671 ;
  assign n19674 = n19673 ^ n19635 ;
  assign n19685 = n19684 ^ n19674 ;
  assign n19776 = n19685 ^ n19680 ;
  assign n19779 = n19700 & n19776 ;
  assign n19780 = n19779 ^ n19680 ;
  assign n19781 = n19596 & n19780 ;
  assign n19782 = n19781 ^ n17052 ;
  assign n19687 = n19668 ^ n19666 ;
  assign n19688 = n19633 & n19687 ;
  assign n19725 = n19688 ^ n19687 ;
  assign n19693 = n19633 ^ n19597 ;
  assign n19694 = n19687 & ~n19693 ;
  assign n19692 = n19667 ^ n19666 ;
  assign n19695 = n19694 ^ n19692 ;
  assign n19690 = n19632 & n19687 ;
  assign n19691 = n19690 ^ n19635 ;
  assign n19696 = n19695 ^ n19691 ;
  assign n19726 = n19725 ^ n19696 ;
  assign n19709 = n19694 ^ n19693 ;
  assign n19686 = n19685 ^ n19681 ;
  assign n19710 = n19709 ^ n19686 ;
  assign n19752 = n19726 ^ n19710 ;
  assign n19753 = ~n19700 & n19752 ;
  assign n19756 = n19753 ^ n19710 ;
  assign n19712 = n19634 & n19692 ;
  assign n19757 = n19756 ^ n19712 ;
  assign n19758 = n19757 ^ n19756 ;
  assign n19761 = n19700 & n19758 ;
  assign n19762 = n19761 ^ n19756 ;
  assign n19763 = ~n19596 & n19762 ;
  assign n19764 = n19763 ^ n19756 ;
  assign n19706 = n19677 ^ n19676 ;
  assign n19697 = n19696 ^ n19682 ;
  assign n19707 = n19706 ^ n19697 ;
  assign n19747 = ~n19596 & ~n19700 ;
  assign n19748 = n19747 ^ n19596 ;
  assign n19749 = n19748 ^ n19700 ;
  assign n19750 = n19749 ^ n19596 ;
  assign n19751 = n19707 & ~n19750 ;
  assign n19765 = n19764 ^ n19751 ;
  assign n19708 = n19707 ^ n19694 ;
  assign n19711 = n19710 ^ n19708 ;
  assign n19713 = n19712 ^ n19711 ;
  assign n19714 = n19713 ^ n19695 ;
  assign n19739 = n19714 ^ n19696 ;
  assign n19740 = n19696 ^ n19596 ;
  assign n19741 = n19740 ^ n19696 ;
  assign n19742 = n19739 & ~n19741 ;
  assign n19743 = n19742 ^ n19696 ;
  assign n19744 = n19700 & n19743 ;
  assign n19732 = n19707 ^ n19688 ;
  assign n19733 = n19732 ^ n19672 ;
  assign n19734 = n19672 ^ n19596 ;
  assign n19735 = n19734 ^ n19672 ;
  assign n19736 = n19733 & ~n19735 ;
  assign n19737 = n19736 ^ n19672 ;
  assign n19738 = ~n19700 & n19737 ;
  assign n19745 = n19744 ^ n19738 ;
  assign n19717 = n19690 ^ n19673 ;
  assign n19715 = n19714 ^ n19681 ;
  assign n19689 = n19688 ^ n19686 ;
  assign n19698 = n19697 ^ n19689 ;
  assign n19699 = n19698 ^ n19686 ;
  assign n19703 = n19699 & n19700 ;
  assign n19704 = n19703 ^ n19686 ;
  assign n19705 = ~n19596 & ~n19704 ;
  assign n19716 = n19715 ^ n19705 ;
  assign n19718 = n19717 ^ n19716 ;
  assign n19719 = n19718 ^ n19705 ;
  assign n19720 = n19700 & ~n19719 ;
  assign n19721 = n19720 ^ n19716 ;
  assign n19746 = n19745 ^ n19721 ;
  assign n19766 = n19765 ^ n19746 ;
  assign n19722 = n19721 ^ n19705 ;
  assign n19723 = n19722 ^ n19700 ;
  assign n19724 = n19723 ^ n19722 ;
  assign n19727 = n19726 ^ n19722 ;
  assign n19728 = n19727 ^ n19722 ;
  assign n19729 = ~n19724 & n19728 ;
  assign n19730 = n19729 ^ n19722 ;
  assign n19731 = ~n19596 & ~n19730 ;
  assign n19767 = n19766 ^ n19731 ;
  assign n19772 = n19673 & ~n19700 ;
  assign n19773 = n19772 ^ n19672 ;
  assign n19774 = ~n19596 & n19773 ;
  assign n19775 = n19767 & ~n19774 ;
  assign n19783 = n19782 ^ n19775 ;
  assign n19784 = n19783 ^ x123 ;
  assign n16624 = n16623 ^ x84 ;
  assign n16977 = n16976 ^ x85 ;
  assign n17203 = n17202 ^ n17090 ;
  assign n17174 = n17124 ^ n17090 ;
  assign n17179 = n17178 ^ n17168 ;
  assign n17180 = n17179 ^ n17124 ;
  assign n17181 = ~n17174 & ~n17180 ;
  assign n17182 = n17181 ^ n17124 ;
  assign n17185 = n17179 ^ n17165 ;
  assign n17186 = n17182 & n17185 ;
  assign n17183 = n17165 ^ n17149 ;
  assign n17187 = n17186 ^ n17183 ;
  assign n17204 = n17203 ^ n17187 ;
  assign n17219 = n17218 ^ n17204 ;
  assign n17188 = n17187 ^ n17179 ;
  assign n17189 = n17188 ^ n17176 ;
  assign n17190 = n17189 ^ n17187 ;
  assign n17193 = n17124 & n17190 ;
  assign n17194 = n17193 ^ n17187 ;
  assign n17195 = ~n17174 & ~n17194 ;
  assign n17220 = n17219 ^ n17195 ;
  assign n17172 = n17171 ^ n17145 ;
  assign n17173 = ~n17127 & ~n17172 ;
  assign n17221 = n17220 ^ n17173 ;
  assign n17136 = n17135 ^ n17126 ;
  assign n17138 = n17137 ^ n17128 ;
  assign n17141 = ~n17135 & ~n17138 ;
  assign n17142 = n17141 ^ n17128 ;
  assign n17143 = n17136 & n17142 ;
  assign n17222 = n17221 ^ n17143 ;
  assign n17134 = n17124 & n17133 ;
  assign n17223 = n17222 ^ n17134 ;
  assign n17131 = n17090 & n17130 ;
  assign n17224 = n17223 ^ n17131 ;
  assign n17225 = ~n17129 & ~n17224 ;
  assign n17226 = n17225 ^ n14988 ;
  assign n17227 = n17226 ^ x83 ;
  assign n17228 = ~n16977 & ~n17227 ;
  assign n17685 = n17228 ^ n16977 ;
  assign n17490 = n17388 & n17441 ;
  assign n17484 = n17483 ^ n17412 ;
  assign n17476 = n17475 ^ n17414 ;
  assign n17477 = n17457 ^ n17444 ;
  assign n17478 = n17444 ^ n17414 ;
  assign n17479 = n17478 ^ n17444 ;
  assign n17480 = n17477 & n17479 ;
  assign n17481 = n17480 ^ n17444 ;
  assign n17482 = ~n17476 & ~n17481 ;
  assign n17485 = n17484 ^ n17482 ;
  assign n17452 = n17451 ^ n17428 ;
  assign n17456 = n17455 ^ n17420 ;
  assign n17458 = n17457 ^ n17456 ;
  assign n17459 = n17452 & ~n17458 ;
  assign n17461 = n17460 ^ n17459 ;
  assign n17474 = n17473 ^ n17461 ;
  assign n17486 = n17485 ^ n17474 ;
  assign n17487 = n17486 ^ n15086 ;
  assign n17450 = n17449 ^ n17429 ;
  assign n17462 = n17461 ^ n17450 ;
  assign n17430 = n17429 ^ n17419 ;
  assign n17447 = n17446 ^ n17430 ;
  assign n17448 = ~n17388 & ~n17447 ;
  assign n17463 = n17462 ^ n17448 ;
  assign n17464 = ~n17417 & ~n17463 ;
  assign n17488 = n17487 ^ n17464 ;
  assign n17416 = ~n17360 & ~n17415 ;
  assign n17489 = n17488 ^ n17416 ;
  assign n17491 = n17490 ^ n17489 ;
  assign n17492 = n17491 ^ x102 ;
  assign n17679 = n17678 ^ x108 ;
  assign n17680 = n17492 & ~n17679 ;
  assign n17681 = n17680 ^ n17679 ;
  assign n17703 = n17681 ^ n17492 ;
  assign n17705 = ~n17685 & n17703 ;
  assign n17771 = n16624 & n17705 ;
  assign n16222 = n16221 ^ x70 ;
  assign n17760 = ~n17681 & ~n17685 ;
  assign n17763 = ~n16624 & n17760 ;
  assign n17687 = n17685 ^ n17227 ;
  assign n17712 = n17703 ^ n17679 ;
  assign n17714 = ~n17687 & n17712 ;
  assign n17688 = n17687 ^ n16977 ;
  assign n17704 = ~n17688 & n17703 ;
  assign n17706 = n17705 ^ n17704 ;
  assign n17689 = n17680 & ~n17688 ;
  assign n17686 = n17680 & ~n17685 ;
  assign n17690 = n17689 ^ n17686 ;
  assign n17683 = n17228 & n17680 ;
  assign n17684 = n17683 ^ n17680 ;
  assign n17691 = n17690 ^ n17684 ;
  assign n17707 = n17706 ^ n17691 ;
  assign n17700 = n17492 ^ n17227 ;
  assign n17701 = n17679 & ~n17700 ;
  assign n17693 = n17492 ^ n16977 ;
  assign n17694 = n17679 ^ n17227 ;
  assign n17695 = n17679 ^ n16977 ;
  assign n17696 = n17695 ^ n17679 ;
  assign n17697 = n17694 & n17696 ;
  assign n17698 = n17697 ^ n17679 ;
  assign n17699 = ~n17693 & n17698 ;
  assign n17702 = n17701 ^ n17699 ;
  assign n17708 = n17707 ^ n17702 ;
  assign n17715 = n17714 ^ n17708 ;
  assign n17716 = n17715 ^ n17704 ;
  assign n17717 = n17716 ^ n17701 ;
  assign n17718 = n17717 ^ n17706 ;
  assign n17719 = n17718 ^ n17703 ;
  assign n17713 = n17228 & n17712 ;
  assign n17720 = n17719 ^ n17713 ;
  assign n17721 = n17720 ^ n17715 ;
  assign n17722 = n17721 ^ n17679 ;
  assign n17723 = n17722 ^ n17718 ;
  assign n17724 = n17723 ^ n17689 ;
  assign n17711 = n17704 ^ n17688 ;
  assign n17725 = n17724 ^ n17711 ;
  assign n17755 = n17725 ^ n17723 ;
  assign n17756 = ~n16624 & ~n17755 ;
  assign n17757 = n17756 ^ n17723 ;
  assign n17764 = n17763 ^ n17757 ;
  assign n17765 = ~n16222 & n17764 ;
  assign n17766 = n17765 ^ n17757 ;
  assign n17710 = n17688 ^ n17686 ;
  assign n17726 = n17725 ^ n17710 ;
  assign n17727 = n17726 ^ n17492 ;
  assign n17682 = n17228 & ~n17681 ;
  assign n17692 = n17691 ^ n17682 ;
  assign n17709 = n17708 ^ n17692 ;
  assign n17728 = n17727 ^ n17709 ;
  assign n17729 = n16624 & n17728 ;
  assign n17730 = n17729 ^ n17727 ;
  assign n17767 = n17766 ^ n17730 ;
  assign n16625 = n16624 ^ n16222 ;
  assign n17740 = n17719 ^ n17714 ;
  assign n17748 = n17740 ^ n17720 ;
  assign n17749 = n17748 ^ n17719 ;
  assign n17750 = n17719 ^ n16624 ;
  assign n17751 = n17750 ^ n17719 ;
  assign n17752 = n17749 & n17751 ;
  assign n17753 = n17752 ^ n17719 ;
  assign n17754 = n16625 & n17753 ;
  assign n17768 = n17767 ^ n17754 ;
  assign n17743 = n17714 ^ n16624 ;
  assign n17744 = n17743 ^ n17714 ;
  assign n17745 = n17740 & n17744 ;
  assign n17746 = n17745 ^ n17714 ;
  assign n17747 = n16222 & n17746 ;
  assign n17769 = n17768 ^ n17747 ;
  assign n17733 = n17730 ^ n17717 ;
  assign n17731 = n17725 ^ n17683 ;
  assign n17732 = n17731 ^ n17730 ;
  assign n17734 = n17733 ^ n17732 ;
  assign n17735 = n17733 ^ n16222 ;
  assign n17736 = n17735 ^ n17733 ;
  assign n17737 = ~n17734 & ~n17736 ;
  assign n17738 = n17737 ^ n17733 ;
  assign n17739 = n16625 & n17738 ;
  assign n17770 = n17769 ^ n17739 ;
  assign n17772 = n17771 ^ n17770 ;
  assign n17773 = n17691 ^ n17687 ;
  assign n17774 = n17773 ^ n17740 ;
  assign n17775 = n17774 ^ n17690 ;
  assign n17776 = n17690 ^ n16624 ;
  assign n17777 = n17776 ^ n17690 ;
  assign n17778 = ~n17775 & n17777 ;
  assign n17779 = n17778 ^ n17690 ;
  assign n17780 = n16625 & n17779 ;
  assign n17781 = ~n17772 & ~n17780 ;
  assign n17782 = n17725 ^ n17689 ;
  assign n17783 = n17782 ^ n17774 ;
  assign n17784 = n17774 ^ n16624 ;
  assign n17785 = n17784 ^ n17774 ;
  assign n17786 = n17783 & n17785 ;
  assign n17787 = n17786 ^ n17774 ;
  assign n17788 = n16222 & ~n17787 ;
  assign n17789 = n17760 ^ n17717 ;
  assign n17790 = n17789 ^ n17723 ;
  assign n17791 = n16624 & n17790 ;
  assign n17792 = n17791 ^ n17760 ;
  assign n17793 = n17792 ^ n17774 ;
  assign n17794 = n17793 ^ n17792 ;
  assign n17795 = n17792 ^ n16222 ;
  assign n17796 = n17795 ^ n17792 ;
  assign n17797 = ~n17794 & ~n17796 ;
  assign n17798 = n17797 ^ n17792 ;
  assign n17799 = ~n16625 & n17798 ;
  assign n17800 = n17799 ^ n17792 ;
  assign n17801 = ~n17788 & ~n17800 ;
  assign n17802 = n17781 & n17801 ;
  assign n17803 = n17802 ^ n15222 ;
  assign n19785 = n17803 ^ x114 ;
  assign n19786 = ~n19784 & ~n19785 ;
  assign n19797 = n19593 & n19786 ;
  assign n19807 = n19451 & n19797 ;
  assign n19594 = n19451 & ~n19593 ;
  assign n19803 = n19594 ^ n19451 ;
  assign n19808 = n19807 ^ n19803 ;
  assign n19787 = n19786 ^ n19785 ;
  assign n19805 = ~n19787 & n19803 ;
  assign n19788 = n19787 ^ n19784 ;
  assign n19804 = ~n19788 & n19803 ;
  assign n19806 = n19805 ^ n19804 ;
  assign n19809 = n19808 ^ n19806 ;
  assign n19595 = n19594 ^ n19593 ;
  assign n19792 = n19786 ^ n19784 ;
  assign n19801 = ~n19595 & ~n19792 ;
  assign n19823 = n19809 ^ n19801 ;
  assign n19789 = ~n19595 & ~n19788 ;
  assign n19824 = n19823 ^ n19789 ;
  assign n19795 = ~n19595 & n19786 ;
  assign n19810 = n19809 ^ n19795 ;
  assign n19822 = n19810 ^ n19595 ;
  assign n19825 = n19824 ^ n19822 ;
  assign n19793 = n19595 ^ n19451 ;
  assign n19816 = n19785 & n19793 ;
  assign n19794 = ~n19792 & n19793 ;
  assign n19817 = n19816 ^ n19794 ;
  assign n19826 = n19825 ^ n19817 ;
  assign n19820 = n19816 ^ n19793 ;
  assign n19813 = n19807 ^ n19797 ;
  assign n19821 = n19820 ^ n19813 ;
  assign n19827 = n19826 ^ n19821 ;
  assign n19350 = n18260 ^ n18224 ;
  assign n19360 = n18195 ^ n17975 ;
  assign n19362 = n18218 ^ n18195 ;
  assign n19361 = n18214 ^ n18195 ;
  assign n19363 = n19362 ^ n19361 ;
  assign n19364 = n19362 ^ n18206 ;
  assign n19365 = n19364 ^ n19362 ;
  assign n19366 = n19363 & n19365 ;
  assign n19367 = n19366 ^ n19362 ;
  assign n19368 = n19360 & ~n19367 ;
  assign n19369 = n19368 ^ n17975 ;
  assign n19353 = n19352 ^ n18195 ;
  assign n19354 = n19353 ^ n18247 ;
  assign n19355 = n18247 ^ n18206 ;
  assign n19356 = n19355 ^ n18247 ;
  assign n19357 = n19354 & ~n19356 ;
  assign n19358 = n19357 ^ n18247 ;
  assign n19359 = ~n17975 & n19358 ;
  assign n19370 = n19369 ^ n19359 ;
  assign n19371 = n19370 ^ n18261 ;
  assign n19375 = n18206 & n18229 ;
  assign n19376 = n19375 ^ n18225 ;
  assign n19377 = ~n18235 & ~n19376 ;
  assign n19378 = n19377 ^ n18225 ;
  assign n19379 = ~n19371 & ~n19378 ;
  assign n19380 = n19379 ^ n19371 ;
  assign n19381 = n18232 & ~n19380 ;
  assign n19382 = n19350 & n19381 ;
  assign n19383 = n19382 ^ n19380 ;
  assign n19384 = n18206 & ~n19383 ;
  assign n19385 = n18202 ^ n17975 ;
  assign n19386 = n19385 ^ n18202 ;
  assign n19389 = ~n18231 & ~n19386 ;
  assign n19390 = n19389 ^ n18202 ;
  assign n19391 = n19384 & n19390 ;
  assign n19392 = n19391 ^ n19383 ;
  assign n19394 = n19393 ^ n18202 ;
  assign n19395 = n19394 ^ n18224 ;
  assign n19398 = n19395 ^ n18233 ;
  assign n19399 = n19396 & n19398 ;
  assign n19400 = n19399 ^ n18233 ;
  assign n19397 = n19396 ^ n19395 ;
  assign n19401 = n19400 ^ n19397 ;
  assign n19402 = ~n19392 & n19401 ;
  assign n19403 = n19402 ^ n17123 ;
  assign n19404 = n19403 ^ x99 ;
  assign n18797 = n18796 ^ n18728 ;
  assign n18800 = n18739 & ~n18797 ;
  assign n18798 = n18757 ^ n18741 ;
  assign n18799 = ~n18797 & n18798 ;
  assign n18801 = n18800 ^ n18799 ;
  assign n18781 = n18747 ^ n18694 ;
  assign n18782 = n18781 ^ n18747 ;
  assign n18785 = ~n18753 & ~n18782 ;
  assign n18786 = n18785 ^ n18747 ;
  assign n18787 = n18728 & n18786 ;
  assign n18794 = n18793 ^ n18787 ;
  assign n18767 = n18694 & n18766 ;
  assign n18756 = n18745 ^ n18743 ;
  assign n18768 = n18767 ^ n18756 ;
  assign n18795 = n18794 ^ n18768 ;
  assign n18802 = n18801 ^ n18795 ;
  assign n18816 = n18815 ^ n18802 ;
  assign n18775 = n18754 ^ n18741 ;
  assign n18737 = n18736 ^ n18734 ;
  assign n18776 = n18775 ^ n18737 ;
  assign n18773 = n18763 ^ n18752 ;
  assign n18772 = n18771 ^ n18736 ;
  assign n18774 = n18773 ^ n18772 ;
  assign n18777 = n18776 ^ n18774 ;
  assign n18778 = n18694 & ~n18777 ;
  assign n18755 = n18754 ^ n18737 ;
  assign n18769 = n18768 ^ n18755 ;
  assign n18779 = n18778 ^ n18769 ;
  assign n18780 = n18729 & ~n18779 ;
  assign n18817 = n18816 ^ n18780 ;
  assign n18818 = ~n18651 & ~n18817 ;
  assign n18819 = n18818 ^ n15451 ;
  assign n19405 = n18819 ^ x72 ;
  assign n19859 = n19404 & ~n19405 ;
  assign n19860 = n19859 ^ n19405 ;
  assign n19861 = n19860 ^ n19404 ;
  assign n19864 = n19861 ^ n19405 ;
  assign n19887 = ~n19827 & n19864 ;
  assign n19873 = n19805 & ~n19860 ;
  assign n19845 = n19405 ^ n19404 ;
  assign n19796 = n19795 ^ n19786 ;
  assign n19798 = n19797 ^ n19796 ;
  assign n19799 = n19798 ^ n19794 ;
  assign n19867 = n19813 ^ n19799 ;
  assign n19868 = n19813 ^ n19404 ;
  assign n19869 = n19868 ^ n19813 ;
  assign n19870 = n19867 & ~n19869 ;
  assign n19871 = n19870 ^ n19813 ;
  assign n19872 = n19845 & n19871 ;
  assign n19874 = n19873 ^ n19872 ;
  assign n19875 = n19874 ^ n19801 ;
  assign n19802 = n19801 ^ n19797 ;
  assign n19811 = n19810 ^ n19802 ;
  assign n19800 = n19799 ^ n19784 ;
  assign n19812 = n19811 ^ n19800 ;
  assign n19866 = n19812 ^ n19807 ;
  assign n19876 = n19875 ^ n19866 ;
  assign n19865 = n19798 & n19864 ;
  assign n19877 = n19876 ^ n19865 ;
  assign n19818 = n19817 ^ n19805 ;
  assign n19819 = n19818 ^ n19787 ;
  assign n19828 = n19827 ^ n19819 ;
  assign n19884 = n19877 ^ n19828 ;
  assign n19879 = n19828 ^ n19817 ;
  assign n19880 = n19879 ^ n19804 ;
  assign n19881 = ~n19405 & n19880 ;
  assign n19878 = n19877 ^ n19874 ;
  assign n19882 = n19881 ^ n19878 ;
  assign n19883 = ~n19404 & ~n19882 ;
  assign n19885 = n19884 ^ n19883 ;
  assign n19862 = n19813 ^ n19809 ;
  assign n19863 = n19861 & n19862 ;
  assign n19886 = n19885 ^ n19863 ;
  assign n19888 = n19887 ^ n19886 ;
  assign n19814 = n19813 ^ n19795 ;
  assign n19815 = n19814 ^ n19812 ;
  assign n19829 = n19828 ^ n19815 ;
  assign n19853 = n19829 ^ n19828 ;
  assign n19854 = n19828 ^ n19405 ;
  assign n19855 = n19854 ^ n19828 ;
  assign n19856 = ~n19853 & ~n19855 ;
  assign n19857 = n19856 ^ n19828 ;
  assign n19858 = ~n19845 & n19857 ;
  assign n19889 = n19888 ^ n19858 ;
  assign n19890 = n19889 ^ n19789 ;
  assign n19846 = n19805 ^ n19404 ;
  assign n19847 = n19846 ^ n19805 ;
  assign n19850 = n19806 & ~n19847 ;
  assign n19851 = n19850 ^ n19805 ;
  assign n19852 = n19845 & n19851 ;
  assign n19891 = n19890 ^ n19852 ;
  assign n19839 = n19804 ^ n19801 ;
  assign n19840 = n19804 ^ n19404 ;
  assign n19841 = n19840 ^ n19804 ;
  assign n19842 = n19839 & ~n19841 ;
  assign n19843 = n19842 ^ n19804 ;
  assign n19844 = ~n19405 & n19843 ;
  assign n19892 = n19891 ^ n19844 ;
  assign n19893 = n19892 ^ n17226 ;
  assign n19790 = n19789 ^ n19405 ;
  assign n19791 = n19790 ^ n19789 ;
  assign n19830 = n19814 ^ n19798 ;
  assign n19831 = n19830 ^ n19594 ;
  assign n19832 = n19831 ^ n19829 ;
  assign n19833 = n19832 ^ n19821 ;
  assign n19836 = n19791 & ~n19833 ;
  assign n19837 = n19836 ^ n19789 ;
  assign n19838 = ~n19404 & n19837 ;
  assign n19894 = n19893 ^ n19838 ;
  assign n19895 = n19894 ^ x118 ;
  assign n19896 = n16222 & ~n16624 ;
  assign n19897 = n19896 ^ n16624 ;
  assign n19898 = n17692 & ~n19897 ;
  assign n19899 = n19898 ^ n17780 ;
  assign n19913 = n17705 ^ n17689 ;
  assign n19914 = n19913 ^ n17715 ;
  assign n19915 = n19914 ^ n17720 ;
  assign n19916 = ~n16222 & n19915 ;
  assign n19909 = n17691 ^ n17679 ;
  assign n19910 = ~n16222 & n19909 ;
  assign n19911 = n19910 ^ n17721 ;
  assign n19912 = n19911 ^ n17716 ;
  assign n19917 = n19916 ^ n19912 ;
  assign n19918 = ~n16624 & n19917 ;
  assign n19919 = n19918 ^ n19911 ;
  assign n19907 = n19896 ^ n16222 ;
  assign n19908 = n17760 & n19907 ;
  assign n19920 = n19919 ^ n19908 ;
  assign n19921 = n19920 ^ n17686 ;
  assign n19900 = n17686 ^ n17682 ;
  assign n19901 = n19900 ^ n17686 ;
  assign n19902 = n17686 ^ n16222 ;
  assign n19903 = n19902 ^ n17686 ;
  assign n19904 = n19901 & n19903 ;
  assign n19905 = n19904 ^ n17686 ;
  assign n19906 = ~n16624 & n19905 ;
  assign n19922 = n19921 ^ n19906 ;
  assign n19923 = ~n19899 & ~n19922 ;
  assign n19924 = n16222 & n17720 ;
  assign n19925 = n19924 ^ n17719 ;
  assign n19926 = n19925 ^ n17683 ;
  assign n19927 = n19926 ^ n19925 ;
  assign n19930 = ~n16222 & n19927 ;
  assign n19931 = n19930 ^ n19925 ;
  assign n19932 = ~n16625 & n19931 ;
  assign n19933 = n19932 ^ n19925 ;
  assign n19934 = ~n17788 & ~n19933 ;
  assign n19935 = n19923 & n19934 ;
  assign n19936 = n19935 ^ n17387 ;
  assign n19937 = n19936 ^ x124 ;
  assign n19941 = n18938 ^ n18905 ;
  assign n19942 = n19941 ^ n18969 ;
  assign n19950 = n19942 ^ n18941 ;
  assign n19946 = n18960 ^ n18903 ;
  assign n19947 = n19946 ^ n18873 ;
  assign n19948 = n19947 ^ n18904 ;
  assign n19949 = n19948 ^ n18944 ;
  assign n19951 = n19950 ^ n19949 ;
  assign n19952 = n18845 & ~n19951 ;
  assign n19953 = n19952 ^ n19949 ;
  assign n19954 = n19953 ^ n18968 ;
  assign n19955 = n19954 ^ n19953 ;
  assign n19938 = n18942 ^ n18903 ;
  assign n19939 = ~n18873 & ~n19938 ;
  assign n19940 = n19939 ^ n18939 ;
  assign n19956 = n19955 ^ n19940 ;
  assign n19957 = ~n18845 & n19956 ;
  assign n19958 = n19957 ^ n19954 ;
  assign n18945 = n18944 ^ n18941 ;
  assign n18946 = n18845 & n18945 ;
  assign n18947 = n18946 ^ n18944 ;
  assign n19959 = n19958 ^ n18947 ;
  assign n19960 = n19945 & ~n19959 ;
  assign n19961 = n19960 ^ n19940 ;
  assign n19943 = n19942 ^ n19940 ;
  assign n19944 = n18845 & n19943 ;
  assign n19962 = n19961 ^ n19944 ;
  assign n19964 = n18824 & n18947 ;
  assign n19965 = ~n19962 & n19964 ;
  assign n19963 = n19962 ^ n17411 ;
  assign n19966 = n19965 ^ n19963 ;
  assign n19967 = n19966 ^ x75 ;
  assign n20183 = n19937 & ~n19967 ;
  assign n20185 = n20183 ^ n19967 ;
  assign n20184 = n20183 ^ n19937 ;
  assign n20186 = n20185 ^ n20184 ;
  assign n20017 = n18376 ^ n18359 ;
  assign n20023 = n20017 ^ n18371 ;
  assign n20020 = n18367 ^ n18363 ;
  assign n20021 = n20020 ^ n20017 ;
  assign n20022 = n18471 & n20021 ;
  assign n20024 = n20023 ^ n20022 ;
  assign n20025 = ~n18404 & n18470 ;
  assign n20026 = ~n20024 & n20025 ;
  assign n20027 = n20026 ^ n18470 ;
  assign n20018 = n20017 ^ n18405 ;
  assign n20019 = ~n18474 & n20018 ;
  assign n20028 = n20027 ^ n20019 ;
  assign n20014 = ~n18384 & ~n18470 ;
  assign n20015 = n20014 ^ n18383 ;
  assign n20016 = n18471 & n20015 ;
  assign n20029 = n20028 ^ n20016 ;
  assign n20030 = ~n19416 & ~n20029 ;
  assign n20040 = ~n19444 & ~n20039 ;
  assign n20041 = n20030 & n20040 ;
  assign n20042 = n20041 ^ n17300 ;
  assign n20043 = n20042 ^ x100 ;
  assign n20061 = n18757 ^ n18744 ;
  assign n20062 = n20061 ^ n18771 ;
  assign n20053 = n18752 ^ n18750 ;
  assign n20054 = n20053 ^ n18737 ;
  assign n20055 = n20054 ^ n18750 ;
  assign n20056 = n18750 ^ n18694 ;
  assign n20057 = n20056 ^ n18750 ;
  assign n20058 = ~n20055 & n20057 ;
  assign n20059 = n20058 ^ n18750 ;
  assign n20060 = n18761 & ~n20059 ;
  assign n20063 = n20062 ^ n20060 ;
  assign n20064 = n20063 ^ n18765 ;
  assign n20065 = n20064 ^ n20060 ;
  assign n20066 = n20060 ^ n18694 ;
  assign n20067 = n20066 ^ n20060 ;
  assign n20068 = ~n20065 & ~n20067 ;
  assign n20069 = n20068 ^ n20060 ;
  assign n20070 = n18728 & ~n20069 ;
  assign n20071 = n20070 ^ n20060 ;
  assign n20048 = n18754 ^ n18651 ;
  assign n20046 = n20045 ^ n18742 ;
  assign n20047 = n20046 ^ n18734 ;
  assign n20049 = n20048 ^ n20047 ;
  assign n20050 = n18728 & ~n20049 ;
  assign n20051 = n20050 ^ n20048 ;
  assign n20052 = n18694 & ~n20051 ;
  assign n20072 = n20071 ^ n20052 ;
  assign n20073 = ~n18787 & n20072 ;
  assign n20074 = n20073 ^ n18801 ;
  assign n20081 = n20074 & ~n20080 ;
  assign n20082 = n20081 ^ n17355 ;
  assign n20083 = n20082 ^ x85 ;
  assign n20084 = n20043 & ~n20083 ;
  assign n20085 = n20084 ^ n20043 ;
  assign n20002 = n19679 ^ n19672 ;
  assign n20003 = ~n19749 & n20002 ;
  assign n20001 = n19682 & ~n19749 ;
  assign n20004 = n20003 ^ n20001 ;
  assign n19997 = n19688 & ~n19750 ;
  assign n19998 = n19997 ^ n19744 ;
  assign n19999 = n19998 ^ n19765 ;
  assign n19976 = n19677 ^ n19669 ;
  assign n19977 = n19976 ^ n19714 ;
  assign n19971 = n19632 ^ n19597 ;
  assign n19972 = n19971 ^ n19707 ;
  assign n19970 = n19685 ^ n19679 ;
  assign n19973 = n19972 ^ n19970 ;
  assign n19974 = n19973 ^ n19710 ;
  assign n19975 = ~n19700 & n19974 ;
  assign n19978 = n19977 ^ n19975 ;
  assign n20000 = n19999 ^ n19978 ;
  assign n20005 = n20004 ^ n20000 ;
  assign n19986 = n19712 ^ n19669 ;
  assign n19987 = ~n19596 & n19986 ;
  assign n19988 = n19987 ^ n19669 ;
  assign n19991 = n19988 ^ n19708 ;
  assign n19992 = n19991 ^ n19988 ;
  assign n19993 = ~n19596 & n19992 ;
  assign n19994 = n19993 ^ n19988 ;
  assign n19995 = n19700 & n19994 ;
  assign n19996 = n19995 ^ n19988 ;
  assign n20006 = n20005 ^ n19996 ;
  assign n20007 = n20006 ^ n17262 ;
  assign n19969 = n19700 ^ n19596 ;
  assign n19979 = n19978 ^ n19684 ;
  assign n19980 = n19979 ^ n19686 ;
  assign n19981 = n19980 ^ n19712 ;
  assign n19982 = n19981 ^ n19978 ;
  assign n19983 = ~n19700 & n19982 ;
  assign n19984 = n19983 ^ n19979 ;
  assign n19985 = n19969 & ~n19984 ;
  assign n20008 = n20007 ^ n19985 ;
  assign n20009 = n20008 ^ x125 ;
  assign n20099 = ~n19452 & ~n19551 ;
  assign n20088 = n19558 ^ n19552 ;
  assign n20089 = n20088 ^ n19524 ;
  assign n20090 = n20089 ^ n19588 ;
  assign n20091 = n19556 ^ n19531 ;
  assign n20094 = ~n20089 & ~n20091 ;
  assign n20095 = n20094 ^ n19556 ;
  assign n20096 = n20090 & n20095 ;
  assign n20097 = n20096 ^ n19588 ;
  assign n20098 = n20097 ^ n19534 ;
  assign n20100 = n20099 ^ n20098 ;
  assign n20119 = n20100 ^ n19523 ;
  assign n20112 = n19517 ^ n19516 ;
  assign n20113 = n19516 ^ n19452 ;
  assign n20114 = n20113 ^ n19516 ;
  assign n20115 = n20112 & n20114 ;
  assign n20116 = n20115 ^ n19516 ;
  assign n20117 = ~n19454 & n20116 ;
  assign n20118 = n20117 ^ n19516 ;
  assign n20120 = n20119 ^ n20118 ;
  assign n20101 = n20100 ^ n20097 ;
  assign n20102 = n20101 ^ n19453 ;
  assign n20103 = n20102 ^ n20101 ;
  assign n20109 = n20103 & n20106 ;
  assign n20110 = n20109 ^ n20101 ;
  assign n20111 = n19454 & n20110 ;
  assign n20121 = n20120 ^ n20111 ;
  assign n20122 = n20121 ^ n19590 ;
  assign n20129 = n20122 & ~n20128 ;
  assign n20130 = n20129 ^ n17332 ;
  assign n20131 = n20130 ^ x118 ;
  assign n20132 = n20009 & ~n20131 ;
  assign n20133 = n20132 ^ n20009 ;
  assign n20198 = n20085 & n20133 ;
  assign n20148 = n20084 & n20133 ;
  assign n20199 = n20198 ^ n20148 ;
  assign n20086 = n20085 ^ n20083 ;
  assign n20170 = n20086 & n20133 ;
  assign n20171 = n20170 ^ n20133 ;
  assign n20200 = n20199 ^ n20171 ;
  assign n20134 = n20133 ^ n20131 ;
  assign n20143 = n20084 & n20134 ;
  assign n20215 = n20200 ^ n20143 ;
  assign n20213 = n20083 ^ n20009 ;
  assign n20163 = n20131 ^ n20009 ;
  assign n20164 = n20131 ^ n20043 ;
  assign n20167 = ~n20083 & n20164 ;
  assign n20168 = n20167 ^ n20043 ;
  assign n20169 = ~n20163 & n20168 ;
  assign n20214 = n20213 ^ n20169 ;
  assign n20216 = n20215 ^ n20214 ;
  assign n20140 = n20084 ^ n20083 ;
  assign n20194 = n20132 & ~n20140 ;
  assign n20195 = n20194 ^ n20170 ;
  assign n20187 = n20085 & n20132 ;
  assign n20212 = n20195 ^ n20187 ;
  assign n20217 = n20216 ^ n20212 ;
  assign n20218 = ~n19937 & n20217 ;
  assign n20219 = n20218 ^ n20214 ;
  assign n20220 = n20186 & n20219 ;
  assign n20135 = n20134 ^ n20009 ;
  assign n20146 = n20084 & ~n20135 ;
  assign n20150 = n20146 ^ n20143 ;
  assign n20149 = n20148 ^ n20084 ;
  assign n20151 = n20150 ^ n20149 ;
  assign n20196 = n20195 ^ n20151 ;
  assign n20188 = n20187 ^ n20170 ;
  assign n20193 = n20188 ^ n20132 ;
  assign n20197 = n20196 ^ n20193 ;
  assign n20201 = n20200 ^ n20197 ;
  assign n20172 = n20171 ^ n20169 ;
  assign n20138 = n20086 & n20134 ;
  assign n20173 = n20172 ^ n20138 ;
  assign n20174 = n20173 ^ n20146 ;
  assign n20087 = ~n20009 & n20086 ;
  assign n20136 = n20135 ^ n20087 ;
  assign n20175 = n20174 ^ n20136 ;
  assign n20176 = n20175 ^ n20143 ;
  assign n20202 = n20201 ^ n20176 ;
  assign n20203 = ~n19937 & ~n20202 ;
  assign n20189 = ~n20186 & n20188 ;
  assign n20141 = n20134 & ~n20140 ;
  assign n20177 = n20176 ^ n20141 ;
  assign n20178 = n20141 ^ n19967 ;
  assign n20179 = n20178 ^ n20141 ;
  assign n20180 = ~n20177 & n20179 ;
  assign n20181 = n20180 ^ n20141 ;
  assign n20182 = n19937 & n20181 ;
  assign n20190 = n20189 ^ n20182 ;
  assign n20191 = n20190 ^ n17491 ;
  assign n19968 = n19967 ^ n19937 ;
  assign n20139 = n20138 ^ n20087 ;
  assign n20142 = n20141 ^ n20139 ;
  assign n20144 = n20143 ^ n20142 ;
  assign n20137 = n20136 ^ n20009 ;
  assign n20145 = n20144 ^ n20137 ;
  assign n20147 = n20146 ^ n20145 ;
  assign n20152 = n20151 ^ n20147 ;
  assign n20153 = ~n19937 & n20152 ;
  assign n20154 = n20153 ^ n20151 ;
  assign n20155 = n20154 ^ n20148 ;
  assign n20156 = n20155 ^ n20154 ;
  assign n20159 = n19937 & n20156 ;
  assign n20160 = n20159 ^ n20154 ;
  assign n20161 = n19968 & n20160 ;
  assign n20162 = n20161 ^ n20154 ;
  assign n20192 = n20191 ^ n20162 ;
  assign n20204 = n20203 ^ n20192 ;
  assign n20207 = n20204 ^ n17491 ;
  assign n20208 = n20207 ^ n20162 ;
  assign n20205 = n20172 ^ n20142 ;
  assign n20206 = n20205 ^ n20190 ;
  assign n20209 = n20208 ^ n20206 ;
  assign n20210 = n19967 & n20209 ;
  assign n20211 = n20210 ^ n20204 ;
  assign n20221 = n20220 ^ n20211 ;
  assign n20222 = n20221 ^ x70 ;
  assign n20622 = ~n19895 & ~n20222 ;
  assign n20623 = n20622 ^ n20222 ;
  assign n20624 = n20623 ^ n19895 ;
  assign n20625 = n20624 ^ n20222 ;
  assign n20239 = ~n18729 & ~n18754 ;
  assign n20234 = n18760 ^ n18745 ;
  assign n20225 = n20062 ^ n18747 ;
  assign n20224 = n18770 ^ n18737 ;
  assign n20226 = n20225 ^ n20224 ;
  assign n20227 = n18694 & ~n20226 ;
  assign n20228 = n20227 ^ n20224 ;
  assign n20235 = n20234 ^ n20228 ;
  assign n20231 = n20230 ^ n18744 ;
  assign n20232 = n20231 ^ n18774 ;
  assign n20233 = ~n18694 & n20232 ;
  assign n20236 = n20235 ^ n20233 ;
  assign n20237 = n18728 & n20236 ;
  assign n20229 = n20228 ^ n18799 ;
  assign n20238 = n20237 ^ n20229 ;
  assign n20240 = n20239 ^ n20238 ;
  assign n20241 = ~n18814 & ~n20240 ;
  assign n20242 = ~n20080 & n20241 ;
  assign n20243 = n20242 ^ n16968 ;
  assign n20244 = n20243 ^ x107 ;
  assign n18491 = n18400 & ~n18470 ;
  assign n18492 = n18491 ^ n18399 ;
  assign n18505 = n18504 ^ n18492 ;
  assign n18496 = n18495 ^ n18385 ;
  assign n18494 = n18373 ^ n18363 ;
  assign n18497 = n18496 ^ n18494 ;
  assign n18498 = n18497 ^ n18492 ;
  assign n18490 = n18489 ^ n18368 ;
  assign n18493 = n18492 ^ n18490 ;
  assign n18499 = n18498 ^ n18493 ;
  assign n18500 = ~n18470 & ~n18499 ;
  assign n18501 = n18500 ^ n18498 ;
  assign n18502 = ~n18471 & n18501 ;
  assign n18506 = n18505 ^ n18502 ;
  assign n18507 = ~n18485 & ~n18506 ;
  assign n18508 = n18507 ^ n15966 ;
  assign n20245 = n18508 ^ x89 ;
  assign n20320 = n17723 ^ n17705 ;
  assign n20321 = n20320 ^ n17725 ;
  assign n20322 = ~n16222 & ~n20321 ;
  assign n20333 = n20322 ^ n17766 ;
  assign n20334 = n20333 ^ n17754 ;
  assign n20335 = n20334 ^ n19899 ;
  assign n20331 = n17708 & ~n19897 ;
  assign n20332 = n20331 ^ n19933 ;
  assign n20336 = n20335 ^ n20332 ;
  assign n20337 = n20336 ^ n16731 ;
  assign n20324 = n17731 ^ n17705 ;
  assign n20325 = n20324 ^ n17760 ;
  assign n20326 = n20325 ^ n20322 ;
  assign n20319 = n17690 ^ n17682 ;
  assign n20323 = n20322 ^ n20319 ;
  assign n20327 = n20326 ^ n20323 ;
  assign n20328 = ~n16222 & ~n20327 ;
  assign n20329 = n20328 ^ n20326 ;
  assign n20330 = n16624 & ~n20329 ;
  assign n20338 = n20337 ^ n20330 ;
  assign n20318 = n17707 & n19896 ;
  assign n20339 = n20338 ^ n20318 ;
  assign n20311 = n17717 ^ n16222 ;
  assign n20312 = n20311 ^ n17717 ;
  assign n20315 = n17715 & n20312 ;
  assign n20316 = n20315 ^ n17717 ;
  assign n20317 = n16624 & n20316 ;
  assign n20340 = n20339 ^ n20317 ;
  assign n20341 = n20340 ^ x66 ;
  assign n20250 = n19707 ^ n19690 ;
  assign n20251 = n20250 ^ n19713 ;
  assign n20252 = n19700 & n20251 ;
  assign n20253 = n20252 ^ n19713 ;
  assign n20254 = n20253 ^ n19708 ;
  assign n20255 = n20254 ^ n19671 ;
  assign n20256 = n20255 ^ n20253 ;
  assign n20259 = ~n19700 & n20256 ;
  assign n20260 = n20259 ^ n20253 ;
  assign n20261 = n19596 & n20260 ;
  assign n20262 = n20261 ^ n20253 ;
  assign n20247 = n19677 ^ n19670 ;
  assign n20248 = n20247 ^ n19681 ;
  assign n20249 = ~n19748 & ~n20248 ;
  assign n20263 = n20262 ^ n20249 ;
  assign n20271 = n20263 ^ n20004 ;
  assign n19754 = n19753 ^ n19726 ;
  assign n20269 = n19596 & n19754 ;
  assign n20270 = n20269 ^ n19998 ;
  assign n20272 = n20271 ^ n20270 ;
  assign n20264 = ~n19969 & ~n20263 ;
  assign n20265 = n19712 ^ n19680 ;
  assign n20266 = n19596 & n20265 ;
  assign n20267 = n20266 ^ n19680 ;
  assign n20268 = n20264 & n20267 ;
  assign n20273 = n20272 ^ n20268 ;
  assign n20274 = ~n19781 & ~n20273 ;
  assign n20275 = ~n19774 & n20274 ;
  assign n20276 = n20275 ^ n16886 ;
  assign n20277 = n20276 ^ x122 ;
  assign n20343 = n20341 ^ n20277 ;
  assign n19253 = n19200 ^ n19189 ;
  assign n19254 = ~n19076 & n19253 ;
  assign n19255 = n19254 ^ n19189 ;
  assign n19258 = n19255 ^ n19174 ;
  assign n19259 = n19258 ^ n19255 ;
  assign n19260 = ~n19076 & n19259 ;
  assign n19261 = n19260 ^ n19255 ;
  assign n19262 = ~n19075 & n19261 ;
  assign n19263 = n19262 ^ n19255 ;
  assign n19238 = n19237 ^ n19075 ;
  assign n19252 = ~n19238 & n19246 ;
  assign n19264 = n19263 ^ n19252 ;
  assign n19239 = n19207 ^ n19195 ;
  assign n19240 = ~n19238 & n19239 ;
  assign n19225 = n19224 ^ n19223 ;
  assign n19227 = n19226 ^ n19225 ;
  assign n19229 = n19228 ^ n19227 ;
  assign n19230 = n19229 ^ n19225 ;
  assign n19231 = n19225 ^ n19075 ;
  assign n19232 = n19231 ^ n19225 ;
  assign n19233 = n19230 & ~n19232 ;
  assign n19234 = n19233 ^ n19225 ;
  assign n19235 = n19077 & n19234 ;
  assign n19236 = n19235 ^ n19225 ;
  assign n19241 = n19240 ^ n19236 ;
  assign n19211 = n19210 ^ n19196 ;
  assign n19193 = n19192 ^ n19190 ;
  assign n19188 = n19187 ^ n19140 ;
  assign n19194 = n19193 ^ n19188 ;
  assign n19212 = n19211 ^ n19194 ;
  assign n19215 = n19211 ^ n19076 ;
  assign n19216 = n19215 ^ n19211 ;
  assign n19217 = n19212 & ~n19216 ;
  assign n19218 = n19217 ^ n19211 ;
  assign n19219 = n19075 & n19218 ;
  assign n19242 = n19241 ^ n19219 ;
  assign n19182 = n19181 ^ n19178 ;
  assign n19183 = ~n19075 & n19182 ;
  assign n19184 = n19183 ^ n19181 ;
  assign n19185 = n19077 & n19184 ;
  assign n19243 = n19242 ^ n19185 ;
  assign n19251 = ~n19243 & ~n19250 ;
  assign n19265 = n19264 ^ n19251 ;
  assign n19278 = n19265 & ~n19277 ;
  assign n19279 = n19278 ^ n14640 ;
  assign n20246 = n19279 ^ x96 ;
  assign n20370 = n20246 & ~n20277 ;
  assign n20298 = n19531 ^ n19524 ;
  assign n20299 = n20298 ^ n19576 ;
  assign n20300 = n19452 & n20299 ;
  assign n20287 = n20105 ^ n19527 ;
  assign n20286 = n19529 ^ n19512 ;
  assign n20288 = n20287 ^ n20286 ;
  assign n20289 = n19452 & n20288 ;
  assign n20290 = n20289 ^ n20286 ;
  assign n20296 = n20290 ^ n19524 ;
  assign n20292 = n19544 ^ n19520 ;
  assign n20295 = n20292 ^ n19538 ;
  assign n20297 = n20296 ^ n20295 ;
  assign n20301 = n20300 ^ n20297 ;
  assign n20302 = ~n19454 & ~n20301 ;
  assign n20291 = n20290 ^ n20118 ;
  assign n20293 = n20292 ^ n20291 ;
  assign n20294 = n20293 ^ n20285 ;
  assign n20303 = n20302 ^ n20294 ;
  assign n20304 = n20303 ^ n19590 ;
  assign n20279 = ~n19453 & n19552 ;
  assign n20305 = n20304 ^ n20279 ;
  assign n20306 = ~n20128 & n20305 ;
  assign n20307 = n20306 ^ n16668 ;
  assign n20308 = n20307 ^ x113 ;
  assign n20371 = n20370 ^ n20308 ;
  assign n20372 = ~n20343 & ~n20371 ;
  assign n20349 = n20341 ^ n20246 ;
  assign n20373 = n20372 ^ n20349 ;
  assign n20344 = n20246 & n20343 ;
  assign n20369 = n20344 ^ n20277 ;
  assign n20374 = n20373 ^ n20369 ;
  assign n20375 = n20374 ^ n20349 ;
  assign n20309 = n20308 ^ n20277 ;
  assign n20278 = n20277 ^ n20246 ;
  assign n20310 = n20309 ^ n20278 ;
  assign n20361 = n20308 & ~n20341 ;
  assign n20362 = n20361 ^ n20308 ;
  assign n20363 = n20343 & n20362 ;
  assign n20364 = n20363 ^ n20277 ;
  assign n20365 = ~n20310 & ~n20364 ;
  assign n20366 = n20365 ^ n20361 ;
  assign n20367 = n20366 ^ n20277 ;
  assign n20368 = n20367 ^ n20308 ;
  assign n20376 = n20375 ^ n20368 ;
  assign n20377 = n20376 ^ n20375 ;
  assign n20352 = n20308 ^ n20246 ;
  assign n20378 = n20370 ^ n20352 ;
  assign n20379 = ~n20341 & ~n20378 ;
  assign n20382 = n20377 & ~n20379 ;
  assign n20383 = n20382 ^ n20375 ;
  assign n20384 = n20245 & n20383 ;
  assign n20385 = n20384 ^ n20375 ;
  assign n20353 = n20341 & ~n20352 ;
  assign n20354 = n20353 ^ n20246 ;
  assign n20355 = n20277 & n20354 ;
  assign n20350 = n20349 ^ n20308 ;
  assign n20356 = n20355 ^ n20350 ;
  assign n20351 = n20350 ^ n20344 ;
  assign n20357 = n20356 ^ n20351 ;
  assign n20342 = n20341 ^ n20309 ;
  assign n20345 = n20344 ^ n20342 ;
  assign n20346 = n20345 ^ n20278 ;
  assign n20347 = n20310 & n20346 ;
  assign n20348 = n20347 ^ n20342 ;
  assign n20358 = n20357 ^ n20348 ;
  assign n20359 = ~n20245 & n20358 ;
  assign n20360 = n20359 ^ n20356 ;
  assign n20386 = n20385 ^ n20360 ;
  assign n20387 = n20244 & ~n20386 ;
  assign n20388 = n20387 ^ n20244 ;
  assign n20389 = n20388 ^ n20385 ;
  assign n20390 = n20389 ^ n16976 ;
  assign n20391 = n20390 ^ x116 ;
  assign n20393 = n19783 ^ x112 ;
  assign n20414 = n20413 ^ x105 ;
  assign n20415 = n20393 & ~n20414 ;
  assign n20416 = n20415 ^ n20414 ;
  assign n20439 = n20438 ^ n19177 ;
  assign n20440 = n20439 ^ n19212 ;
  assign n20441 = n19076 & ~n20440 ;
  assign n20442 = n20441 ^ n19228 ;
  assign n20443 = ~n19075 & n20442 ;
  assign n20434 = n19076 & n20433 ;
  assign n20420 = n19199 ^ n19175 ;
  assign n20421 = n20420 ^ n19226 ;
  assign n20422 = n19226 ^ n19076 ;
  assign n20423 = n19077 & n20422 ;
  assign n20424 = n20423 ^ n19076 ;
  assign n20425 = n20421 & n20424 ;
  assign n20426 = n20425 ^ n19226 ;
  assign n20427 = n20426 ^ n19209 ;
  assign n20428 = n20427 ^ n19181 ;
  assign n20431 = n20428 ^ n19263 ;
  assign n20417 = n19221 ^ n19192 ;
  assign n20418 = n20417 ^ n19187 ;
  assign n20419 = n19075 & n20418 ;
  assign n20429 = n20428 ^ n20419 ;
  assign n20430 = n19077 & n20429 ;
  assign n20432 = n20431 ^ n20430 ;
  assign n20435 = n20434 ^ n20432 ;
  assign n20444 = n20443 ^ n20435 ;
  assign n20445 = ~n19252 & ~n20444 ;
  assign n20457 = n20445 & ~n20456 ;
  assign n20458 = n20457 ^ n17549 ;
  assign n20459 = n20458 ^ x64 ;
  assign n20500 = n20499 ^ x81 ;
  assign n20545 = ~n20459 & ~n20500 ;
  assign n20464 = n17715 ^ n17683 ;
  assign n20465 = n20464 ^ n17692 ;
  assign n20462 = n17700 ^ n17699 ;
  assign n20463 = n16222 & ~n20462 ;
  assign n20466 = n20465 ^ n20463 ;
  assign n20478 = n20466 ^ n20332 ;
  assign n20479 = n20478 ^ n17747 ;
  assign n20460 = n17719 ^ n17692 ;
  assign n20461 = n20460 ^ n17724 ;
  assign n20467 = n20466 ^ n20461 ;
  assign n20468 = n20467 ^ n20466 ;
  assign n20469 = n20468 ^ n17718 ;
  assign n20470 = n20469 ^ n20468 ;
  assign n20471 = n20468 ^ n17782 ;
  assign n20472 = n20471 ^ n20468 ;
  assign n20473 = ~n20470 & n20472 ;
  assign n20474 = n20473 ^ n20468 ;
  assign n20475 = ~n16222 & ~n20474 ;
  assign n20476 = n20475 ^ n20467 ;
  assign n20477 = ~n16624 & n20476 ;
  assign n20480 = n20479 ^ n20477 ;
  assign n20481 = ~n17800 & ~n20480 ;
  assign n20482 = n20481 ^ n17579 ;
  assign n20483 = n20482 ^ x90 ;
  assign n20484 = ~n20459 & n20483 ;
  assign n20485 = n20484 ^ n20459 ;
  assign n20501 = n19403 ^ x115 ;
  assign n20502 = ~n20500 & n20501 ;
  assign n20503 = n20502 ^ n20500 ;
  assign n20529 = ~n20485 & ~n20503 ;
  assign n20517 = n20484 & n20502 ;
  assign n20530 = n20529 ^ n20517 ;
  assign n20546 = n20545 ^ n20530 ;
  assign n20513 = n20459 & ~n20501 ;
  assign n20514 = n20483 ^ n20459 ;
  assign n20515 = n20513 & ~n20514 ;
  assign n20526 = n20515 ^ n20514 ;
  assign n20527 = ~n20500 & ~n20526 ;
  assign n20528 = n20527 ^ n20502 ;
  assign n20531 = n20530 ^ n20528 ;
  assign n20504 = n20503 ^ n20501 ;
  assign n20506 = n20485 ^ n20483 ;
  assign n20523 = n20504 & n20506 ;
  assign n20507 = n20504 ^ n20500 ;
  assign n20521 = ~n20485 & n20507 ;
  assign n20524 = n20523 ^ n20521 ;
  assign n20508 = n20506 & n20507 ;
  assign n20525 = n20524 ^ n20508 ;
  assign n20532 = n20531 ^ n20525 ;
  assign n20522 = n20521 ^ n20506 ;
  assign n20533 = n20532 ^ n20522 ;
  assign n20536 = n20533 ^ n20517 ;
  assign n20537 = n20536 ^ n20529 ;
  assign n20511 = n20484 ^ n20483 ;
  assign n20512 = n20504 & n20511 ;
  assign n20516 = n20515 ^ n20512 ;
  assign n20518 = n20517 ^ n20516 ;
  assign n20535 = n20518 ^ n20503 ;
  assign n20538 = n20537 ^ n20535 ;
  assign n20547 = n20546 ^ n20538 ;
  assign n20548 = n20547 ^ n20536 ;
  assign n20534 = n20533 ^ n20531 ;
  assign n20544 = n20534 ^ n20502 ;
  assign n20549 = n20548 ^ n20544 ;
  assign n20550 = n20549 ^ n20538 ;
  assign n20510 = n20484 & n20504 ;
  assign n20551 = n20550 ^ n20510 ;
  assign n20542 = n20483 & n20501 ;
  assign n20543 = n20542 ^ n20484 ;
  assign n20552 = n20551 ^ n20543 ;
  assign n20614 = n20552 ^ n20533 ;
  assign n20615 = ~n20416 & n20614 ;
  assign n20608 = n20549 ^ n20512 ;
  assign n20609 = n20512 ^ n20414 ;
  assign n20610 = n20609 ^ n20512 ;
  assign n20611 = ~n20608 & ~n20610 ;
  assign n20612 = n20611 ^ n20512 ;
  assign n20613 = ~n20393 & n20612 ;
  assign n20616 = n20615 ^ n20613 ;
  assign n20617 = n20616 ^ n17678 ;
  assign n20581 = n20415 ^ n20393 ;
  assign n20582 = n20516 & n20581 ;
  assign n20553 = n20552 ^ n20524 ;
  assign n20554 = n20553 ^ n20512 ;
  assign n20539 = n20538 ^ n20534 ;
  assign n20540 = n20539 ^ n20527 ;
  assign n20519 = n20518 ^ n20510 ;
  assign n20505 = ~n20485 & n20504 ;
  assign n20509 = n20508 ^ n20505 ;
  assign n20520 = n20519 ^ n20509 ;
  assign n20541 = n20540 ^ n20520 ;
  assign n20555 = n20554 ^ n20541 ;
  assign n20567 = n20555 ^ n20523 ;
  assign n20566 = n20552 ^ n20550 ;
  assign n20568 = n20567 ^ n20566 ;
  assign n20569 = n20393 & n20568 ;
  assign n20570 = n20569 ^ n20551 ;
  assign n20558 = n20547 ^ n20512 ;
  assign n20579 = n20570 ^ n20558 ;
  assign n20571 = n20570 ^ n20509 ;
  assign n20572 = n20571 ^ n20552 ;
  assign n20573 = n20572 ^ n20570 ;
  assign n20576 = n20393 & n20573 ;
  assign n20577 = n20576 ^ n20570 ;
  assign n20578 = ~n20414 & n20577 ;
  assign n20580 = n20579 ^ n20578 ;
  assign n20583 = n20582 ^ n20580 ;
  assign n20559 = n20558 ^ n20532 ;
  assign n20560 = n20559 ^ n20558 ;
  assign n20561 = n20558 ^ n20393 ;
  assign n20562 = n20561 ^ n20558 ;
  assign n20563 = n20560 & ~n20562 ;
  assign n20564 = n20563 ^ n20558 ;
  assign n20565 = n20414 & ~n20564 ;
  assign n20584 = n20583 ^ n20565 ;
  assign n20585 = n20414 ^ n20393 ;
  assign n20586 = n20531 ^ n20529 ;
  assign n20587 = n20531 ^ n20414 ;
  assign n20588 = n20587 ^ n20531 ;
  assign n20589 = n20586 & ~n20588 ;
  assign n20590 = n20589 ^ n20531 ;
  assign n20591 = ~n20585 & n20590 ;
  assign n20592 = n20584 & ~n20591 ;
  assign n20556 = n20555 ^ n20505 ;
  assign n20557 = ~n20416 & n20556 ;
  assign n20593 = n20592 ^ n20557 ;
  assign n20596 = n20534 & n20588 ;
  assign n20597 = n20596 ^ n20531 ;
  assign n20598 = n20393 & n20597 ;
  assign n20599 = n20593 & ~n20598 ;
  assign n20600 = n20536 ^ n20414 ;
  assign n20601 = n20600 ^ n20536 ;
  assign n20604 = ~n20548 & n20601 ;
  assign n20605 = n20604 ^ n20536 ;
  assign n20606 = n20393 & n20605 ;
  assign n20607 = n20599 & ~n20606 ;
  assign n20618 = n20617 ^ n20607 ;
  assign n20619 = n20618 ^ x76 ;
  assign n20620 = ~n20391 & n20619 ;
  assign n20621 = n20620 ^ n20391 ;
  assign n20627 = n20621 ^ n20619 ;
  assign n20640 = n20627 ^ n20391 ;
  assign n20650 = ~n20625 & n20640 ;
  assign n20649 = n20620 & n20622 ;
  assign n20651 = n20650 ^ n20649 ;
  assign n20641 = ~n20623 & n20640 ;
  assign n20652 = n20651 ^ n20641 ;
  assign n18509 = n18508 ^ x74 ;
  assign n18997 = n18993 ^ n16126 ;
  assign n18994 = n18993 ^ n18979 ;
  assign n18995 = n18994 ^ n18990 ;
  assign n18996 = ~n18845 & n18995 ;
  assign n18998 = n18997 ^ n18996 ;
  assign n18999 = n18998 ^ n16126 ;
  assign n18980 = n18979 ^ n18978 ;
  assign n18981 = n18980 ^ n18976 ;
  assign n18982 = n18976 ^ n18845 ;
  assign n18983 = n18982 ^ n18976 ;
  assign n18984 = ~n18981 & n18983 ;
  assign n18985 = n18984 ^ n18976 ;
  assign n18986 = ~n18947 & ~n18985 ;
  assign n19000 = n18999 ^ n18986 ;
  assign n19001 = n18824 & n19000 ;
  assign n19002 = n19001 ^ n18998 ;
  assign n19003 = n19002 ^ x121 ;
  assign n19004 = n18509 & ~n19003 ;
  assign n19005 = n19004 ^ n19003 ;
  assign n18263 = n18221 ^ n18209 ;
  assign n18264 = ~n18258 & ~n18263 ;
  assign n18250 = n18141 ^ n18095 ;
  assign n18249 = n18248 ^ n18192 ;
  assign n18251 = n18250 ^ n18249 ;
  assign n18252 = ~n17975 & ~n18251 ;
  assign n18253 = n18252 ^ n18245 ;
  assign n18254 = ~n18206 & n18253 ;
  assign n18255 = n18254 ^ n18245 ;
  assign n18237 = n18228 ^ n18221 ;
  assign n18236 = n18224 ^ n18216 ;
  assign n18238 = n18237 ^ n18236 ;
  assign n18239 = n18237 ^ n17975 ;
  assign n18240 = n18239 ^ n18237 ;
  assign n18241 = n18238 & n18240 ;
  assign n18242 = n18241 ^ n18237 ;
  assign n18243 = n18235 & n18242 ;
  assign n18256 = n18255 ^ n18243 ;
  assign n18262 = n18261 ^ n18256 ;
  assign n18265 = n18264 ^ n18262 ;
  assign n18234 = ~n18231 & ~n18233 ;
  assign n18266 = n18265 ^ n18234 ;
  assign n18200 = n18199 ^ n18195 ;
  assign n18203 = n18202 ^ n18200 ;
  assign n18207 = n18203 & n18206 ;
  assign n18205 = n17975 & n18202 ;
  assign n18208 = n18207 ^ n18205 ;
  assign n18267 = n18266 ^ n18208 ;
  assign n18269 = n18268 ^ n18267 ;
  assign n18270 = n18269 ^ n15740 ;
  assign n18271 = n18270 ^ x120 ;
  assign n18820 = n18819 ^ x65 ;
  assign n19007 = ~n18271 & ~n18820 ;
  assign n19008 = n19007 ^ n18820 ;
  assign n19010 = n19008 ^ n18271 ;
  assign n19030 = ~n19005 & ~n19010 ;
  assign n19011 = n19010 ^ n18820 ;
  assign n19012 = n19004 & ~n19011 ;
  assign n19033 = n19030 ^ n19012 ;
  assign n19021 = n19004 & n19007 ;
  assign n19020 = ~n19005 & n19007 ;
  assign n19022 = n19021 ^ n19020 ;
  assign n19023 = n19022 ^ n19007 ;
  assign n19014 = n19005 ^ n18509 ;
  assign n19018 = n19014 ^ n19003 ;
  assign n19019 = n19007 & n19018 ;
  assign n19024 = n19023 ^ n19019 ;
  assign n19017 = ~n19010 & n19014 ;
  assign n19025 = n19024 ^ n19017 ;
  assign n19015 = ~n19008 & n19014 ;
  assign n19016 = n19015 ^ n19014 ;
  assign n19026 = n19025 ^ n19016 ;
  assign n19034 = n19033 ^ n19026 ;
  assign n19009 = ~n19005 & ~n19008 ;
  assign n19013 = n19012 ^ n19009 ;
  assign n19027 = n19026 ^ n19013 ;
  assign n19028 = n19027 ^ n19025 ;
  assign n18510 = n18509 ^ n18271 ;
  assign n18821 = n18820 ^ n18271 ;
  assign n18822 = ~n18510 & ~n18821 ;
  assign n18823 = n18822 ^ n18820 ;
  assign n19006 = n19005 ^ n18823 ;
  assign n19029 = n19028 ^ n19006 ;
  assign n19031 = n19030 ^ n19029 ;
  assign n19032 = n19031 ^ n19011 ;
  assign n19035 = n19034 ^ n19032 ;
  assign n19036 = n19035 ^ n19029 ;
  assign n19037 = n17803 ^ x98 ;
  assign n19280 = n19279 ^ x88 ;
  assign n19281 = n19037 & ~n19280 ;
  assign n19282 = ~n19036 & n19281 ;
  assign n19283 = n19280 ^ n19037 ;
  assign n19299 = ~n19010 & n19018 ;
  assign n19300 = ~n19283 & n19299 ;
  assign n19293 = n19017 ^ n19015 ;
  assign n19296 = ~n19280 & n19293 ;
  assign n19297 = n19296 ^ n19015 ;
  assign n19298 = ~n19037 & n19297 ;
  assign n19301 = n19300 ^ n19298 ;
  assign n19319 = ~n19008 & n19018 ;
  assign n19310 = n19035 ^ n19019 ;
  assign n19311 = n19310 ^ n19021 ;
  assign n19303 = n19299 ^ n19020 ;
  assign n19304 = n19303 ^ n18822 ;
  assign n19305 = n19304 ^ n19024 ;
  assign n19308 = n19305 ^ n19035 ;
  assign n19309 = n19308 ^ n19019 ;
  assign n19312 = n19311 ^ n19309 ;
  assign n19307 = n19012 ^ n19004 ;
  assign n19313 = n19312 ^ n19307 ;
  assign n19314 = n19313 ^ n19024 ;
  assign n19327 = n19319 ^ n19314 ;
  assign n19321 = n19021 ^ n19009 ;
  assign n19324 = n19281 ^ n19280 ;
  assign n19325 = n19321 & ~n19324 ;
  assign n19326 = n19325 ^ n19015 ;
  assign n19328 = n19327 ^ n19326 ;
  assign n19331 = n19321 ^ n19313 ;
  assign n19332 = ~n19281 & ~n19331 ;
  assign n19333 = n19328 & n19332 ;
  assign n19320 = n19319 ^ n19030 ;
  assign n19322 = n19321 ^ n19320 ;
  assign n19323 = n19037 & n19322 ;
  assign n19329 = n19328 ^ n19323 ;
  assign n19334 = n19333 ^ n19329 ;
  assign n19335 = ~n19280 & n19334 ;
  assign n19336 = n19335 ^ n19323 ;
  assign n19302 = n19036 ^ n19013 ;
  assign n19306 = n19305 ^ n19302 ;
  assign n19315 = n19314 ^ n19306 ;
  assign n19316 = n19280 & ~n19315 ;
  assign n19317 = n19316 ^ n19305 ;
  assign n19318 = ~n19037 & n19317 ;
  assign n19337 = n19336 ^ n19318 ;
  assign n19338 = ~n19301 & ~n19337 ;
  assign n19284 = n19281 ^ n19037 ;
  assign n19287 = n19280 ^ n19020 ;
  assign n19288 = n19287 ^ n19283 ;
  assign n19289 = n19284 & ~n19288 ;
  assign n19290 = n19289 ^ n19283 ;
  assign n19291 = ~n19019 & ~n19290 ;
  assign n19292 = n19291 ^ n19283 ;
  assign n19339 = n19338 ^ n19292 ;
  assign n19340 = ~n19282 & ~n19339 ;
  assign n19341 = n19017 ^ n19012 ;
  assign n19342 = n19341 ^ n19030 ;
  assign n19343 = n19280 & n19342 ;
  assign n19344 = n19343 ^ n19034 ;
  assign n19345 = n19283 & n19344 ;
  assign n19346 = n19345 ^ n19026 ;
  assign n19347 = n19340 & ~n19346 ;
  assign n19348 = n19347 ^ n16221 ;
  assign n19349 = n19348 ^ x101 ;
  assign n20956 = n20641 ^ n19349 ;
  assign n20957 = n20956 ^ n20641 ;
  assign n20958 = n20652 & n20957 ;
  assign n20959 = n20958 ^ n20641 ;
  assign n20960 = n20917 & n20959 ;
  assign n20643 = n20620 & ~n20623 ;
  assign n20644 = n20643 ^ n20623 ;
  assign n20635 = ~n20621 & ~n20624 ;
  assign n20631 = ~n20624 & n20627 ;
  assign n20636 = n20635 ^ n20631 ;
  assign n20628 = n20622 & n20627 ;
  assign n20626 = ~n20621 & ~n20625 ;
  assign n20629 = n20628 ^ n20626 ;
  assign n20637 = n20636 ^ n20629 ;
  assign n20633 = n20391 ^ n20222 ;
  assign n20634 = ~n20619 & ~n20633 ;
  assign n20638 = n20637 ^ n20634 ;
  assign n20632 = n20631 ^ n20619 ;
  assign n20639 = n20638 ^ n20632 ;
  assign n20642 = n20641 ^ n20639 ;
  assign n20645 = n20644 ^ n20642 ;
  assign n20646 = n20645 ^ n20631 ;
  assign n20630 = n20629 ^ n20619 ;
  assign n20647 = n20646 ^ n20630 ;
  assign n20223 = n20222 ^ n19895 ;
  assign n20392 = n20391 ^ n20223 ;
  assign n20648 = n20647 ^ n20392 ;
  assign n20653 = n20652 ^ n20648 ;
  assign n20660 = n20653 ^ n20650 ;
  assign n20661 = n20660 ^ n20643 ;
  assign n20923 = n20661 ^ n20620 ;
  assign n20924 = n20923 ^ n20651 ;
  assign n20654 = n20653 ^ n20624 ;
  assign n20655 = n20654 ^ n20636 ;
  assign n20925 = n20924 ^ n20655 ;
  assign n20936 = n20925 ^ n20653 ;
  assign n20934 = n20655 ^ n20641 ;
  assign n20933 = n20650 ^ n20640 ;
  assign n20935 = n20934 ^ n20933 ;
  assign n20937 = n20936 ^ n20935 ;
  assign n20931 = n20645 ^ n20628 ;
  assign n20930 = n20639 ^ n20635 ;
  assign n20932 = n20931 ^ n20930 ;
  assign n20938 = n20937 ^ n20932 ;
  assign n20939 = ~n19349 & ~n20938 ;
  assign n20940 = n20939 ^ n20937 ;
  assign n20961 = n20960 ^ n20940 ;
  assign n20941 = n20639 ^ n20629 ;
  assign n20944 = n20941 ^ n20621 ;
  assign n20945 = n20944 ^ n20932 ;
  assign n20946 = n20945 ^ n20631 ;
  assign n20657 = n20628 ^ n20621 ;
  assign n20658 = n20657 ^ n20638 ;
  assign n20943 = n20658 ^ n20628 ;
  assign n20947 = n20946 ^ n20943 ;
  assign n20948 = n20947 ^ n20940 ;
  assign n20942 = n20941 ^ n20643 ;
  assign n20949 = n20948 ^ n20942 ;
  assign n20950 = n20949 ^ n20940 ;
  assign n20951 = n19349 & ~n20950 ;
  assign n20952 = n20951 ^ n20948 ;
  assign n20953 = n20917 & n20952 ;
  assign n20962 = n20961 ^ n20953 ;
  assign n20926 = n19349 & n20917 ;
  assign n20928 = n20926 ^ n19349 ;
  assign n20929 = n20646 & n20928 ;
  assign n20963 = n20962 ^ n20929 ;
  assign n20927 = ~n20925 & n20926 ;
  assign n20964 = n20963 ^ n20927 ;
  assign n20656 = n20655 ^ n20649 ;
  assign n20659 = n20658 ^ n20656 ;
  assign n20662 = n20661 ^ n20659 ;
  assign n20920 = n20662 & ~n20917 ;
  assign n20921 = n20920 ^ n20661 ;
  assign n20922 = ~n19349 & n20921 ;
  assign n20965 = n20964 ^ n20922 ;
  assign n20969 = n20626 & n20928 ;
  assign n20966 = ~n20642 & n20957 ;
  assign n20967 = n20966 ^ n20641 ;
  assign n20968 = ~n20917 & n20967 ;
  assign n20970 = n20969 ^ n20968 ;
  assign n20971 = ~n20965 & ~n20970 ;
  assign n20972 = n20971 ^ n17803 ;
  assign n20973 = n20008 ^ x68 ;
  assign n20974 = n20307 ^ x117 ;
  assign n20975 = n20973 & n20974 ;
  assign n20976 = n20975 ^ n20973 ;
  assign n21038 = n20680 ^ n19184 ;
  assign n21039 = n21038 ^ n19223 ;
  assign n21040 = n21039 ^ n19174 ;
  assign n21041 = n21040 ^ n19184 ;
  assign n21042 = n19075 & n21041 ;
  assign n21043 = n21042 ^ n21038 ;
  assign n21044 = ~n19077 & n21043 ;
  assign n21035 = n19177 & n19237 ;
  assign n21029 = n19246 ^ n19221 ;
  assign n21030 = n21029 ^ n19201 ;
  assign n21031 = n19075 & n21030 ;
  assign n21023 = n19226 ^ n19196 ;
  assign n21016 = n19206 ^ n19195 ;
  assign n21017 = n21016 ^ n19196 ;
  assign n21018 = n21016 ^ n19075 ;
  assign n21020 = ~n19076 & n21018 ;
  assign n21021 = n21020 ^ n19075 ;
  assign n21022 = n21017 & ~n21021 ;
  assign n21024 = n21023 ^ n21022 ;
  assign n21027 = n21024 ^ n19201 ;
  assign n21028 = n21027 ^ n19268 ;
  assign n21032 = n21031 ^ n21028 ;
  assign n21033 = ~n19076 & n21032 ;
  assign n21025 = n21024 ^ n19222 ;
  assign n21026 = n21025 ^ n19184 ;
  assign n21034 = n21033 ^ n21026 ;
  assign n21036 = n21035 ^ n21034 ;
  assign n21009 = n19222 ^ n19193 ;
  assign n21010 = n21009 ^ n19222 ;
  assign n21011 = n19222 ^ n19075 ;
  assign n21012 = n21011 ^ n19222 ;
  assign n21013 = n21010 & n21012 ;
  assign n21014 = n21013 ^ n19222 ;
  assign n21015 = n19077 & n21014 ;
  assign n21037 = n21036 ^ n21015 ;
  assign n21045 = n21044 ^ n21037 ;
  assign n21046 = ~n19252 & ~n21045 ;
  assign n21047 = ~n19274 & n21046 ;
  assign n21048 = n21047 ^ n17863 ;
  assign n21049 = n21048 ^ x67 ;
  assign n21050 = n20243 ^ x92 ;
  assign n21051 = n21049 & n21050 ;
  assign n21069 = n21051 ^ n21050 ;
  assign n20977 = n19966 ^ x69 ;
  assign n20997 = n18268 ^ n18206 ;
  assign n20989 = n18227 ^ n18216 ;
  assign n20990 = n20989 ^ n18200 ;
  assign n20988 = n20693 ^ n18221 ;
  assign n20991 = n20990 ^ n20988 ;
  assign n20992 = n20990 ^ n18206 ;
  assign n20993 = n20992 ^ n20990 ;
  assign n20994 = ~n20991 & ~n20993 ;
  assign n20995 = n20994 ^ n20990 ;
  assign n20996 = ~n17975 & ~n20995 ;
  assign n20998 = n20997 ^ n20996 ;
  assign n20986 = n19396 ^ n18258 ;
  assign n20987 = ~n19400 & n20986 ;
  assign n20999 = n20998 ^ n20987 ;
  assign n20985 = ~n18206 & n18228 ;
  assign n21000 = n20999 ^ n20985 ;
  assign n20984 = n18235 & n20693 ;
  assign n21001 = n21000 ^ n20984 ;
  assign n20978 = n18226 ^ n18214 ;
  assign n20979 = n18214 ^ n17975 ;
  assign n20980 = n20979 ^ n18214 ;
  assign n20981 = ~n20978 & ~n20980 ;
  assign n20982 = n20981 ^ n18214 ;
  assign n20983 = ~n18206 & n20982 ;
  assign n21002 = n21001 ^ n20983 ;
  assign n21003 = ~n20736 & ~n21002 ;
  assign n21004 = n21003 ^ n17841 ;
  assign n21005 = n21004 ^ x86 ;
  assign n21006 = ~n20977 & ~n21005 ;
  assign n21076 = n21006 ^ n20977 ;
  assign n21079 = n21069 & ~n21076 ;
  assign n21073 = n21006 & n21069 ;
  assign n21080 = n21079 ^ n21073 ;
  assign n21007 = n21006 ^ n21005 ;
  assign n21070 = ~n21007 & n21069 ;
  assign n21078 = n21070 ^ n21069 ;
  assign n21081 = n21080 ^ n21078 ;
  assign n21082 = n21081 ^ n21079 ;
  assign n21077 = n21051 & ~n21076 ;
  assign n21083 = n21082 ^ n21077 ;
  assign n21008 = n21007 ^ n20977 ;
  assign n21072 = ~n21008 & n21051 ;
  assign n21074 = n21073 ^ n21072 ;
  assign n21068 = n21006 & n21051 ;
  assign n21071 = n21070 ^ n21068 ;
  assign n21075 = n21074 ^ n21071 ;
  assign n21084 = n21083 ^ n21075 ;
  assign n21085 = n21084 ^ n21050 ;
  assign n21089 = n21085 ^ n21068 ;
  assign n21052 = n21051 ^ n21049 ;
  assign n21062 = n21006 & n21052 ;
  assign n21088 = n21079 ^ n21062 ;
  assign n21090 = n21089 ^ n21088 ;
  assign n21086 = n21085 ^ n21080 ;
  assign n21087 = n21086 ^ n21006 ;
  assign n21091 = n21090 ^ n21087 ;
  assign n21060 = ~n21008 & n21052 ;
  assign n21092 = n21091 ^ n21060 ;
  assign n21058 = ~n21007 & n21052 ;
  assign n21093 = n21092 ^ n21058 ;
  assign n21094 = n21093 ^ n21050 ;
  assign n21055 = ~n21007 & ~n21050 ;
  assign n21059 = n21058 ^ n21055 ;
  assign n21061 = n21060 ^ n21059 ;
  assign n21063 = n21062 ^ n21061 ;
  assign n21053 = n21052 ^ n21050 ;
  assign n21056 = n21055 ^ n21053 ;
  assign n21057 = n21056 ^ n21050 ;
  assign n21064 = n21063 ^ n21057 ;
  assign n21054 = ~n21008 & ~n21053 ;
  assign n21065 = n21064 ^ n21054 ;
  assign n21066 = n21065 ^ n21059 ;
  assign n21067 = n21066 ^ n21062 ;
  assign n21095 = n21094 ^ n21067 ;
  assign n21096 = n20976 & ~n21095 ;
  assign n21139 = n20976 & n21081 ;
  assign n21104 = n20976 ^ n20974 ;
  assign n21136 = ~n21056 & ~n21104 ;
  assign n21126 = n20974 ^ n20973 ;
  assign n21131 = n21089 ^ n21074 ;
  assign n21127 = n21088 ^ n20974 ;
  assign n21128 = ~n21126 & ~n21127 ;
  assign n21129 = n21128 ^ n20974 ;
  assign n21130 = n21090 & n21129 ;
  assign n21132 = n21131 ^ n21130 ;
  assign n21114 = n21069 ^ n21006 ;
  assign n21115 = n21114 ^ n21060 ;
  assign n21116 = n20974 & n21115 ;
  assign n21133 = n21132 ^ n21116 ;
  assign n21134 = n21126 & n21133 ;
  assign n21117 = n21070 ^ n21058 ;
  assign n21118 = n21070 ^ n20973 ;
  assign n21119 = n21118 ^ n21070 ;
  assign n21120 = n21117 & n21119 ;
  assign n21121 = n21120 ^ n21070 ;
  assign n21122 = ~n20974 & n21121 ;
  assign n21123 = n21122 ^ n21064 ;
  assign n21124 = n21123 ^ n21116 ;
  assign n21107 = n21085 ^ n21077 ;
  assign n21108 = n21107 ^ n21095 ;
  assign n21109 = n21095 ^ n20974 ;
  assign n21110 = n21109 ^ n21095 ;
  assign n21111 = ~n21108 & ~n21110 ;
  assign n21112 = n21111 ^ n21095 ;
  assign n21113 = ~n20973 & ~n21112 ;
  assign n21125 = n21124 ^ n21113 ;
  assign n21135 = n21134 ^ n21125 ;
  assign n21137 = n21136 ^ n21135 ;
  assign n21105 = n21104 ^ n20973 ;
  assign n21106 = n21066 & n21105 ;
  assign n21138 = n21137 ^ n21106 ;
  assign n21140 = n21139 ^ n21138 ;
  assign n21097 = n21064 ^ n20974 ;
  assign n21098 = n21097 ^ n21064 ;
  assign n21101 = n21073 & ~n21098 ;
  assign n21102 = n21101 ^ n21064 ;
  assign n21103 = ~n20973 & n21102 ;
  assign n21141 = n21140 ^ n21103 ;
  assign n21142 = ~n21096 & ~n21141 ;
  assign n21143 = n21142 ^ n19171 ;
  assign n21144 = n21143 ^ x82 ;
  assign n21172 = n19805 ^ n19789 ;
  assign n21173 = n19861 & n21172 ;
  assign n21158 = ~n19860 & ~n19862 ;
  assign n21168 = n19594 & n19792 ;
  assign n21169 = n21158 & n21168 ;
  assign n21164 = ~n19832 & n19859 ;
  assign n21165 = n21164 ^ n19852 ;
  assign n21160 = n19866 ^ n19795 ;
  assign n21161 = n21160 ^ n19879 ;
  assign n21162 = n19864 & ~n21161 ;
  assign n21155 = n19825 ^ n19804 ;
  assign n21156 = n19864 & ~n21155 ;
  assign n21157 = n21156 ^ n19860 ;
  assign n21159 = n21158 ^ n21157 ;
  assign n21163 = n21162 ^ n21159 ;
  assign n21166 = n21165 ^ n21163 ;
  assign n21167 = n21166 ^ n19872 ;
  assign n21170 = n21169 ^ n21167 ;
  assign n21145 = n19807 ^ n19801 ;
  assign n21146 = n21145 ^ n19821 ;
  assign n21147 = n21146 ^ n19807 ;
  assign n21148 = n21147 ^ n19799 ;
  assign n21149 = n21148 ^ n21146 ;
  assign n21150 = n21146 ^ n19405 ;
  assign n21151 = n21150 ^ n21146 ;
  assign n21152 = n21149 & ~n21151 ;
  assign n21153 = n21152 ^ n21146 ;
  assign n21154 = n19845 & n21153 ;
  assign n21171 = n21170 ^ n21154 ;
  assign n21174 = n21173 ^ n21171 ;
  assign n21175 = ~n19844 & n21174 ;
  assign n21176 = n19825 ^ n19794 ;
  assign n21177 = n21176 ^ n19816 ;
  assign n21178 = n21177 ^ n19794 ;
  assign n21179 = n19794 ^ n19404 ;
  assign n21180 = n21179 ^ n19794 ;
  assign n21181 = ~n21178 & ~n21180 ;
  assign n21182 = n21181 ^ n19794 ;
  assign n21183 = ~n19845 & n21182 ;
  assign n21184 = n21175 & ~n21183 ;
  assign n21185 = n21184 ^ n18872 ;
  assign n21186 = n21185 ^ x72 ;
  assign n21187 = ~n21144 & n21186 ;
  assign n21188 = n21187 ^ n21186 ;
  assign n21190 = n20130 ^ x93 ;
  assign n21191 = n20739 ^ x84 ;
  assign n21285 = ~n21190 & n21191 ;
  assign n21286 = n21285 ^ n21191 ;
  assign n21225 = n20269 ^ n19738 ;
  assign n21204 = n19686 ^ n19671 ;
  assign n21203 = n20248 ^ n19682 ;
  assign n21205 = n21204 ^ n21203 ;
  assign n21206 = n21203 ^ n19700 ;
  assign n21207 = n19969 ^ n19700 ;
  assign n21208 = ~n21206 & n21207 ;
  assign n21209 = n21208 ^ n19700 ;
  assign n21210 = n21205 & n21209 ;
  assign n21211 = n21210 ^ n21203 ;
  assign n21220 = n21211 ^ n19764 ;
  assign n21212 = n21211 ^ n20247 ;
  assign n21213 = n21212 ^ n19707 ;
  assign n21214 = n21213 ^ n21211 ;
  assign n21215 = n21211 ^ n19700 ;
  assign n21216 = n21215 ^ n21211 ;
  assign n21217 = n21214 & n21216 ;
  assign n21218 = n21217 ^ n21211 ;
  assign n21219 = n19596 & ~n21218 ;
  assign n21221 = n21220 ^ n21219 ;
  assign n21202 = n19714 & n19747 ;
  assign n21222 = n21221 ^ n21202 ;
  assign n21197 = n19970 ^ n19696 ;
  assign n21198 = n21197 ^ n19688 ;
  assign n21199 = ~n19700 & n21198 ;
  assign n21200 = n21199 ^ n19688 ;
  assign n21201 = n19969 & n21200 ;
  assign n21223 = n21222 ^ n21201 ;
  assign n21224 = ~n20003 & n21223 ;
  assign n21226 = n21225 ^ n21224 ;
  assign n21227 = ~n19996 & n21226 ;
  assign n21228 = n21227 ^ n18016 ;
  assign n21229 = n21228 ^ x91 ;
  assign n21231 = n18824 & n19958 ;
  assign n21230 = n19953 ^ n17983 ;
  assign n21232 = n21231 ^ n21230 ;
  assign n21233 = n21232 ^ x70 ;
  assign n21234 = ~n21229 & n21233 ;
  assign n21235 = n21234 ^ n21233 ;
  assign n21236 = n21235 ^ n21229 ;
  assign n21237 = n21236 ^ n21233 ;
  assign n21192 = n20690 ^ x110 ;
  assign n21193 = n19936 ^ x116 ;
  assign n21194 = n21192 & n21193 ;
  assign n21239 = n21194 ^ n21192 ;
  assign n21240 = n21239 ^ n21193 ;
  assign n21277 = ~n21237 & ~n21240 ;
  assign n21262 = n21233 ^ n21192 ;
  assign n21263 = n21262 ^ n21193 ;
  assign n21264 = n21239 & n21263 ;
  assign n21267 = n21264 ^ n21239 ;
  assign n21266 = n21234 & n21239 ;
  assign n21268 = n21267 ^ n21266 ;
  assign n21278 = n21277 ^ n21268 ;
  assign n21241 = n21235 & ~n21240 ;
  assign n21290 = n21278 ^ n21241 ;
  assign n21254 = n21240 ^ n21192 ;
  assign n21255 = n21236 & n21254 ;
  assign n21247 = n21233 ^ n21229 ;
  assign n21243 = n21193 ^ n21192 ;
  assign n21250 = n21243 ^ n21193 ;
  assign n21251 = n21233 & ~n21250 ;
  assign n21252 = n21251 ^ n21193 ;
  assign n21253 = n21247 & n21252 ;
  assign n21256 = n21255 ^ n21253 ;
  assign n21257 = n21192 & n21256 ;
  assign n21288 = n21257 ^ n21256 ;
  assign n21289 = n21288 ^ n21268 ;
  assign n21291 = n21290 ^ n21289 ;
  assign n21323 = n21291 ^ n21240 ;
  assign n21324 = n21286 & ~n21323 ;
  assign n21294 = n21290 ^ n21237 ;
  assign n21238 = n21194 & ~n21237 ;
  assign n21246 = n21238 ^ n21194 ;
  assign n21258 = n21257 ^ n21246 ;
  assign n21259 = n21258 ^ n21241 ;
  assign n21260 = n21259 ^ n21255 ;
  assign n21244 = n21229 & ~n21243 ;
  assign n21245 = n21244 ^ n21236 ;
  assign n21261 = n21260 ^ n21245 ;
  assign n21265 = n21264 ^ n21261 ;
  assign n21269 = n21268 ^ n21265 ;
  assign n21242 = n21241 ^ n21238 ;
  assign n21270 = n21269 ^ n21242 ;
  assign n21295 = n21294 ^ n21270 ;
  assign n21322 = n21286 & ~n21295 ;
  assign n21325 = n21324 ^ n21322 ;
  assign n21316 = n21288 ^ n21191 ;
  assign n21317 = n21316 ^ n21288 ;
  assign n21293 = n21277 ^ n21261 ;
  assign n21296 = n21295 ^ n21293 ;
  assign n21297 = n21296 ^ n21268 ;
  assign n21292 = n21260 ^ n21238 ;
  assign n21298 = n21297 ^ n21292 ;
  assign n21273 = n21270 ^ n21263 ;
  assign n21299 = n21298 ^ n21273 ;
  assign n21300 = n21299 ^ n21291 ;
  assign n21301 = n21300 ^ n21257 ;
  assign n21318 = n21301 ^ n21288 ;
  assign n21319 = n21317 & ~n21318 ;
  assign n21320 = n21319 ^ n21288 ;
  assign n21321 = n21190 & n21320 ;
  assign n21326 = n21325 ^ n21321 ;
  assign n21327 = n21326 ^ n18844 ;
  assign n21302 = n21301 ^ n21266 ;
  assign n21287 = n21256 ^ n21234 ;
  assign n21303 = n21302 ^ n21287 ;
  assign n21304 = n21303 ^ n21238 ;
  assign n21305 = n21286 & ~n21304 ;
  assign n21271 = n21270 ^ n21264 ;
  assign n21272 = n21191 & ~n21271 ;
  assign n21274 = n21273 ^ n21272 ;
  assign n21306 = n21305 ^ n21274 ;
  assign n21279 = n21278 ^ n21258 ;
  assign n21275 = n21263 ^ n21253 ;
  assign n21276 = n21275 ^ n21274 ;
  assign n21280 = n21279 ^ n21276 ;
  assign n21281 = n21280 ^ n21274 ;
  assign n21282 = n21191 & n21281 ;
  assign n21283 = n21282 ^ n21276 ;
  assign n21284 = n21190 & ~n21283 ;
  assign n21307 = n21306 ^ n21284 ;
  assign n21308 = n21191 ^ n21190 ;
  assign n21309 = n21303 ^ n21293 ;
  assign n21310 = n21293 ^ n21191 ;
  assign n21311 = n21310 ^ n21293 ;
  assign n21312 = ~n21309 & ~n21311 ;
  assign n21313 = n21312 ^ n21293 ;
  assign n21314 = n21308 & n21313 ;
  assign n21315 = n21307 & ~n21314 ;
  assign n21328 = n21327 ^ n21315 ;
  assign n21329 = n21328 ^ x123 ;
  assign n21330 = n20148 ^ n20142 ;
  assign n21331 = n21330 ^ n20148 ;
  assign n21332 = n20148 ^ n19937 ;
  assign n21333 = n21332 ^ n20148 ;
  assign n21334 = n21331 & ~n21333 ;
  assign n21335 = n21334 ^ n20148 ;
  assign n21336 = n19968 & n21335 ;
  assign n21337 = n21336 ^ n20148 ;
  assign n21360 = n20187 ^ n20147 ;
  assign n21361 = n21360 ^ n20173 ;
  assign n21362 = n21361 ^ n20147 ;
  assign n21363 = n20147 ^ n19937 ;
  assign n21364 = n21363 ^ n20147 ;
  assign n21365 = n21362 & ~n21364 ;
  assign n21366 = n21365 ^ n20147 ;
  assign n21367 = ~n19968 & n21366 ;
  assign n21368 = n21367 ^ n20147 ;
  assign n21353 = n20212 ^ n20175 ;
  assign n21351 = n20198 ^ n20151 ;
  assign n21352 = n21351 ^ n20188 ;
  assign n21354 = n21353 ^ n21352 ;
  assign n21355 = n21352 ^ n19937 ;
  assign n21356 = n21355 ^ n21352 ;
  assign n21357 = ~n21354 & n21356 ;
  assign n21358 = n21357 ^ n21352 ;
  assign n21359 = n20186 & n21358 ;
  assign n21369 = n21368 ^ n21359 ;
  assign n21370 = n21369 ^ n20200 ;
  assign n21345 = n20197 ^ n20194 ;
  assign n21346 = n20194 ^ n19937 ;
  assign n21347 = n21346 ^ n20194 ;
  assign n21348 = n21345 & n21347 ;
  assign n21349 = n21348 ^ n20194 ;
  assign n21350 = ~n20186 & n21349 ;
  assign n21371 = n21370 ^ n21350 ;
  assign n21338 = n20200 ^ n20184 ;
  assign n21339 = n20185 ^ n20087 ;
  assign n21342 = ~n20200 & n21339 ;
  assign n21343 = n21342 ^ n20185 ;
  assign n21344 = n21338 & n21343 ;
  assign n21372 = n21371 ^ n21344 ;
  assign n21373 = ~n21337 & ~n21372 ;
  assign n21374 = ~n20162 & ~n20182 ;
  assign n21375 = n21373 & n21374 ;
  assign n21376 = n21375 ^ n19477 ;
  assign n21377 = n21376 ^ x104 ;
  assign n21378 = n21329 & n21377 ;
  assign n21379 = n21378 ^ n21377 ;
  assign n21391 = n20521 ^ n20508 ;
  assign n21392 = n21391 ^ n20550 ;
  assign n21393 = n20393 & n21392 ;
  assign n21401 = n21393 ^ n20520 ;
  assign n21400 = n20545 ^ n20542 ;
  assign n21402 = n21401 ^ n21400 ;
  assign n21403 = n21402 ^ n21393 ;
  assign n21404 = ~n20393 & n21403 ;
  assign n21405 = n21404 ^ n21401 ;
  assign n21406 = n20414 & n21405 ;
  assign n21395 = n20512 & n20581 ;
  assign n21394 = ~n20416 & n20510 ;
  assign n21396 = n21395 ^ n21394 ;
  assign n21397 = n21396 ^ n21393 ;
  assign n21387 = n20531 ^ n20512 ;
  assign n21388 = n20610 & n21387 ;
  assign n21389 = n21388 ^ n20512 ;
  assign n21390 = n20585 & n21389 ;
  assign n21398 = n21397 ^ n21390 ;
  assign n21399 = n21398 ^ n20606 ;
  assign n21407 = n21406 ^ n21399 ;
  assign n21382 = n20552 ^ n20510 ;
  assign n21383 = n21382 ^ n20508 ;
  assign n21384 = n21383 ^ n20537 ;
  assign n21380 = n20553 ^ n20483 ;
  assign n21381 = n21380 ^ n20519 ;
  assign n21385 = n21384 ^ n21381 ;
  assign n21386 = ~n20416 & ~n21385 ;
  assign n21408 = n21407 ^ n21386 ;
  assign n21409 = n21408 ^ n20523 ;
  assign n21410 = n21409 ^ n20615 ;
  assign n21411 = n21410 ^ n19074 ;
  assign n21412 = n21411 ^ x114 ;
  assign n21426 = n20363 ^ n20354 ;
  assign n21427 = n21426 ^ n20375 ;
  assign n21428 = n21427 ^ n20350 ;
  assign n21429 = n21428 ^ n20348 ;
  assign n21430 = n20245 & n21429 ;
  assign n21431 = n21430 ^ n21428 ;
  assign n21434 = n21431 ^ n19503 ;
  assign n21420 = n20368 ^ n20278 ;
  assign n21421 = n21420 ^ n20373 ;
  assign n21414 = n20379 ^ n20246 ;
  assign n21415 = n21414 ^ n20366 ;
  assign n21413 = n20379 ^ n20370 ;
  assign n21416 = n21415 ^ n21413 ;
  assign n21417 = n21416 ^ n20366 ;
  assign n21418 = ~n20309 & n21417 ;
  assign n21419 = n21418 ^ n21415 ;
  assign n21422 = n21421 ^ n21419 ;
  assign n21423 = n21422 ^ n20373 ;
  assign n21424 = n20245 & n21423 ;
  assign n21425 = n21424 ^ n21422 ;
  assign n21432 = n21431 ^ n21425 ;
  assign n21433 = n20244 & ~n21432 ;
  assign n21435 = n21434 ^ n21433 ;
  assign n21436 = n21435 ^ x105 ;
  assign n21437 = ~n21412 & ~n21436 ;
  assign n21438 = n21437 ^ n21412 ;
  assign n21453 = n21438 ^ n21436 ;
  assign n21454 = n21379 & ~n21453 ;
  assign n21455 = n21454 ^ n21379 ;
  assign n21442 = n21379 ^ n21329 ;
  assign n21445 = ~n21412 & ~n21442 ;
  assign n21444 = ~n21329 & n21437 ;
  assign n21446 = n21445 ^ n21444 ;
  assign n21443 = ~n21438 & ~n21442 ;
  assign n21447 = n21446 ^ n21443 ;
  assign n21440 = n21378 & ~n21438 ;
  assign n21448 = n21447 ^ n21440 ;
  assign n21439 = n21379 & ~n21438 ;
  assign n21441 = n21440 ^ n21439 ;
  assign n21449 = n21448 ^ n21441 ;
  assign n21456 = n21455 ^ n21449 ;
  assign n21457 = n21188 & n21456 ;
  assign n21458 = n21378 & ~n21453 ;
  assign n21459 = n21144 & n21458 ;
  assign n21460 = n21186 ^ n21144 ;
  assign n21489 = n21443 ^ n21438 ;
  assign n21490 = n21489 ^ n21441 ;
  assign n21462 = n21378 ^ n21329 ;
  assign n21463 = ~n21453 & n21462 ;
  assign n21464 = n21463 ^ n21454 ;
  assign n21465 = n21464 ^ n21453 ;
  assign n21466 = n21465 ^ n21458 ;
  assign n21477 = n21466 ^ n21447 ;
  assign n21472 = n21436 ^ n21412 ;
  assign n21474 = n21412 ^ n21377 ;
  assign n21475 = n21474 ^ n21329 ;
  assign n21476 = ~n21472 & ~n21475 ;
  assign n21478 = n21477 ^ n21476 ;
  assign n21473 = n21472 ^ n21458 ;
  assign n21479 = n21478 ^ n21473 ;
  assign n21480 = n21479 ^ n21443 ;
  assign n21481 = n21480 ^ n21412 ;
  assign n21482 = n21481 ^ n21448 ;
  assign n21470 = n21436 ^ n21329 ;
  assign n21471 = n21470 ^ n21377 ;
  assign n21483 = n21482 ^ n21471 ;
  assign n21461 = n21445 ^ n21442 ;
  assign n21467 = n21466 ^ n21461 ;
  assign n21468 = n21467 ^ n21464 ;
  assign n21484 = n21483 ^ n21468 ;
  assign n21502 = n21490 ^ n21484 ;
  assign n21503 = n21502 ^ n21444 ;
  assign n21501 = n21443 ^ n21412 ;
  assign n21504 = n21503 ^ n21501 ;
  assign n21505 = ~n21144 & n21504 ;
  assign n21499 = n21463 ^ n21461 ;
  assign n21485 = n21484 ^ n21456 ;
  assign n21486 = n21485 ^ n21466 ;
  assign n21487 = n21486 ^ n21458 ;
  assign n21469 = n21468 ^ n21412 ;
  assign n21488 = n21487 ^ n21469 ;
  assign n21491 = n21490 ^ n21454 ;
  assign n21492 = n21491 ^ n21485 ;
  assign n21493 = n21490 ^ n21186 ;
  assign n21494 = n21460 & n21493 ;
  assign n21495 = n21494 ^ n21186 ;
  assign n21496 = ~n21492 & ~n21495 ;
  assign n21497 = n21496 ^ n21490 ;
  assign n21498 = n21488 & n21497 ;
  assign n21500 = n21499 ^ n21498 ;
  assign n21506 = n21505 ^ n21500 ;
  assign n21507 = n21460 & n21506 ;
  assign n21508 = n21507 ^ n21498 ;
  assign n21509 = ~n21459 & n21508 ;
  assign n21510 = ~n21457 & n21509 ;
  assign n21189 = n21188 ^ n21144 ;
  assign n21450 = n21449 ^ n21444 ;
  assign n21451 = n21450 ^ n21437 ;
  assign n21452 = n21189 & n21451 ;
  assign n21511 = n21510 ^ n21452 ;
  assign n21512 = n21460 ^ n21445 ;
  assign n21513 = n21448 ^ n21445 ;
  assign n21514 = n21513 ^ n21460 ;
  assign n21515 = n21514 ^ n21186 ;
  assign n21516 = n21515 ^ n21513 ;
  assign n21517 = n21460 ^ n21441 ;
  assign n21518 = n21517 ^ n21513 ;
  assign n21519 = ~n21516 & n21518 ;
  assign n21520 = n21519 ^ n21513 ;
  assign n21521 = ~n21512 & n21520 ;
  assign n21522 = n21521 ^ n21445 ;
  assign n21523 = n21511 & ~n21522 ;
  assign n21524 = n21523 ^ n20307 ;
  assign n21525 = n21524 ^ x93 ;
  assign n21535 = n19404 & n19802 ;
  assign n21543 = n21535 ^ n19833 ;
  assign n21541 = n19799 & ~n19860 ;
  assign n21542 = n21541 ^ n21156 ;
  assign n21544 = n21543 ^ n21542 ;
  assign n21537 = n19817 ^ n19789 ;
  assign n21538 = ~n19404 & n21537 ;
  assign n21533 = n19810 ^ n19789 ;
  assign n21534 = n21533 ^ n19828 ;
  assign n21536 = n21535 ^ n21534 ;
  assign n21539 = n21538 ^ n21536 ;
  assign n21540 = n19845 & n21539 ;
  assign n21545 = n21544 ^ n21540 ;
  assign n21528 = n19833 ^ n19405 ;
  assign n21529 = n21528 ^ n19833 ;
  assign n21530 = ~n19866 & ~n21529 ;
  assign n21531 = n21530 ^ n19833 ;
  assign n21532 = ~n19404 & ~n21531 ;
  assign n21546 = n21545 ^ n21532 ;
  assign n21547 = ~n21173 & n21546 ;
  assign n21548 = ~n21183 & n21547 ;
  assign n21549 = ~n19874 & n21548 ;
  assign n21550 = ~n19844 & n21549 ;
  assign n21551 = n21550 ^ n18302 ;
  assign n21552 = n21551 ^ x124 ;
  assign n21553 = n21424 ^ n21419 ;
  assign n21554 = n21553 ^ n21431 ;
  assign n21555 = n21431 ^ n20244 ;
  assign n21556 = n21555 ^ n21431 ;
  assign n21557 = n21554 & ~n21556 ;
  assign n21558 = n21557 ^ n21431 ;
  assign n21559 = ~n21421 & n21558 ;
  assign n21560 = n21559 ^ n18611 ;
  assign n21561 = n21560 ^ x110 ;
  assign n21710 = n21552 & n21561 ;
  assign n21711 = n21710 ^ n21561 ;
  assign n21712 = n21711 ^ n21552 ;
  assign n21583 = n21350 ^ n20145 ;
  assign n21575 = n20198 ^ n20195 ;
  assign n21576 = n21575 ^ n20197 ;
  assign n21580 = n21576 ^ n20174 ;
  assign n21574 = n20175 ^ n20138 ;
  assign n21577 = n21576 ^ n21574 ;
  assign n21570 = n20143 ^ n20084 ;
  assign n21571 = n21570 ^ n20173 ;
  assign n21572 = n21571 ^ n20169 ;
  assign n21573 = n21572 ^ n20144 ;
  assign n21578 = n21577 ^ n21573 ;
  assign n21579 = ~n19937 & ~n21578 ;
  assign n21581 = n21580 ^ n21579 ;
  assign n21582 = n20186 & n21581 ;
  assign n21584 = n21583 ^ n21582 ;
  assign n21569 = ~n19937 & n20144 ;
  assign n21585 = n21584 ^ n21569 ;
  assign n21562 = n20184 ^ n20145 ;
  assign n21563 = n20194 ^ n20185 ;
  assign n21564 = n20185 ^ n20145 ;
  assign n21565 = n21564 ^ n20185 ;
  assign n21566 = n21563 & ~n21565 ;
  assign n21567 = n21566 ^ n20185 ;
  assign n21568 = n21562 & n21567 ;
  assign n21586 = n21585 ^ n21568 ;
  assign n21587 = ~n20190 & ~n21586 ;
  assign n21588 = ~n21337 & n21587 ;
  assign n21589 = n21588 ^ n18469 ;
  assign n21590 = n21589 ^ x93 ;
  assign n21591 = n19299 ^ n19021 ;
  assign n21592 = n21591 ^ n19308 ;
  assign n21593 = n19308 ^ n19280 ;
  assign n21594 = n21593 ^ n19308 ;
  assign n21595 = n21592 & ~n21594 ;
  assign n21596 = n21595 ^ n19308 ;
  assign n21597 = n19037 & n21596 ;
  assign n21606 = n19031 ^ n19017 ;
  assign n21607 = n21606 ^ n19303 ;
  assign n21608 = n19037 & ~n21607 ;
  assign n21609 = n21608 ^ n19303 ;
  assign n21616 = n21609 ^ n19319 ;
  assign n21617 = n21616 ^ n19292 ;
  assign n21611 = n19313 ^ n19026 ;
  assign n21612 = n21611 ^ n19321 ;
  assign n21613 = n19037 & n21612 ;
  assign n21605 = n19321 ^ n19024 ;
  assign n21610 = n21609 ^ n21605 ;
  assign n21614 = n21613 ^ n21610 ;
  assign n21615 = n19283 & n21614 ;
  assign n21618 = n21617 ^ n21615 ;
  assign n21598 = n19319 ^ n19308 ;
  assign n21599 = n19324 ^ n19284 ;
  assign n21600 = n21599 ^ n19281 ;
  assign n21601 = n19308 ^ n19281 ;
  assign n21602 = n21600 & n21601 ;
  assign n21603 = n21602 ^ n19281 ;
  assign n21604 = n21598 & n21603 ;
  assign n21619 = n21618 ^ n21604 ;
  assign n21620 = n19031 ^ n19012 ;
  assign n21623 = ~n19280 & ~n21620 ;
  assign n21624 = n21623 ^ n19031 ;
  assign n21625 = ~n19037 & ~n21624 ;
  assign n21626 = n21619 & ~n21625 ;
  assign n21627 = ~n21597 & n21626 ;
  assign n21628 = n21627 ^ n19325 ;
  assign n21629 = ~n19030 & n21628 ;
  assign n21630 = n21629 ^ n19665 ;
  assign n21631 = n21630 ^ x92 ;
  assign n21632 = n21590 & ~n21631 ;
  assign n21713 = n21632 ^ n21631 ;
  assign n21714 = n21713 ^ n21590 ;
  assign n21715 = n21714 ^ n21631 ;
  assign n21633 = n21285 ^ n21190 ;
  assign n21652 = n21275 ^ n21244 ;
  assign n21650 = n21268 ^ n21235 ;
  assign n21651 = n21650 ^ n21259 ;
  assign n21653 = n21652 ^ n21651 ;
  assign n21654 = ~n21633 & n21653 ;
  assign n21646 = n21288 ^ n21258 ;
  assign n21643 = n21257 ^ n21243 ;
  assign n21644 = n21643 ^ n21229 ;
  assign n21645 = n21191 & ~n21644 ;
  assign n21647 = n21646 ^ n21645 ;
  assign n21648 = n21308 & n21647 ;
  assign n21649 = n21648 ^ n21646 ;
  assign n21655 = n21654 ^ n21649 ;
  assign n21636 = n21300 ^ n21255 ;
  assign n21637 = n21636 ^ n21273 ;
  assign n21638 = n21273 ^ n21191 ;
  assign n21639 = n21638 ^ n21273 ;
  assign n21640 = n21637 & n21639 ;
  assign n21641 = n21640 ^ n21273 ;
  assign n21642 = n21190 & ~n21641 ;
  assign n21656 = n21655 ^ n21642 ;
  assign n21635 = n21269 & n21286 ;
  assign n21657 = n21656 ^ n21635 ;
  assign n21658 = n21657 ^ n21324 ;
  assign n21659 = n21658 ^ n21322 ;
  assign n21660 = n21659 ^ n18727 ;
  assign n21634 = ~n21301 & ~n21633 ;
  assign n21661 = n21660 ^ n21634 ;
  assign n21662 = n21661 ^ x67 ;
  assign n21680 = ~n20416 & n20508 ;
  assign n21677 = n20524 ^ n20505 ;
  assign n21678 = n20415 & n21677 ;
  assign n21663 = ~n20414 & ~n20540 ;
  assign n21664 = n21663 ^ n20527 ;
  assign n21673 = n21664 ^ n20598 ;
  assign n21666 = n21664 ^ n20553 ;
  assign n21665 = n21664 ^ n20519 ;
  assign n21667 = n21666 ^ n21665 ;
  assign n21668 = n21666 ^ n20393 ;
  assign n21669 = n21668 ^ n21666 ;
  assign n21670 = n21667 & n21669 ;
  assign n21671 = n21670 ^ n21666 ;
  assign n21672 = n20585 & n21671 ;
  assign n21674 = n21673 ^ n21672 ;
  assign n21675 = ~n20613 & ~n21674 ;
  assign n21676 = n21675 ^ n21396 ;
  assign n21679 = n21678 ^ n21676 ;
  assign n21681 = n21680 ^ n21679 ;
  assign n21682 = n21681 ^ n21396 ;
  assign n21685 = n20537 ^ n20393 ;
  assign n21686 = n21685 ^ n20537 ;
  assign n21687 = n21384 & n21686 ;
  assign n21688 = n21687 ^ n20537 ;
  assign n21689 = n20414 & n21688 ;
  assign n21690 = n21682 & n21689 ;
  assign n21691 = n21690 ^ n21681 ;
  assign n21692 = ~n20557 & n21691 ;
  assign n21693 = ~n21390 & n21692 ;
  assign n21694 = n21693 ^ n19631 ;
  assign n21695 = n21694 ^ x78 ;
  assign n21700 = ~n21662 & n21695 ;
  assign n21716 = n21700 ^ n21662 ;
  assign n21717 = n21715 & ~n21716 ;
  assign n21718 = ~n21712 & n21717 ;
  assign n21696 = n21695 ^ n21662 ;
  assign n21697 = n21632 & ~n21696 ;
  assign n21698 = n21697 ^ n21561 ;
  assign n21699 = n21698 ^ n21697 ;
  assign n21701 = n21700 ^ n21695 ;
  assign n21702 = n21701 ^ n21662 ;
  assign n21703 = n21632 & n21702 ;
  assign n21704 = n21703 ^ n21697 ;
  assign n21707 = ~n21699 & n21704 ;
  assign n21708 = n21707 ^ n21697 ;
  assign n21709 = ~n21552 & n21708 ;
  assign n21719 = n21718 ^ n21709 ;
  assign n21720 = n21712 ^ n21561 ;
  assign n21721 = n21717 & n21720 ;
  assign n21726 = n21701 & n21714 ;
  assign n21725 = n21714 & ~n21716 ;
  assign n21727 = n21726 ^ n21725 ;
  assign n21723 = n21700 & n21714 ;
  assign n21724 = n21723 ^ n21714 ;
  assign n21728 = n21727 ^ n21724 ;
  assign n21722 = ~n21713 & ~n21716 ;
  assign n21729 = n21728 ^ n21722 ;
  assign n21730 = n21729 ^ n21726 ;
  assign n21731 = ~n21712 & n21730 ;
  assign n21743 = n21701 & ~n21713 ;
  assign n21744 = n21743 ^ n21728 ;
  assign n21745 = n21744 ^ n21713 ;
  assign n21741 = n21702 & ~n21713 ;
  assign n21742 = n21741 ^ n21729 ;
  assign n21746 = n21745 ^ n21742 ;
  assign n21750 = n21700 & n21715 ;
  assign n21747 = n21632 & ~n21695 ;
  assign n21748 = n21747 ^ n21704 ;
  assign n21751 = n21750 ^ n21748 ;
  assign n21756 = n21751 ^ n21741 ;
  assign n21733 = n21701 & n21715 ;
  assign n21752 = n21751 ^ n21733 ;
  assign n21753 = n21752 ^ n21717 ;
  assign n21749 = n21748 ^ n21715 ;
  assign n21754 = n21753 ^ n21749 ;
  assign n21755 = n21754 ^ n21722 ;
  assign n21757 = n21756 ^ n21755 ;
  assign n21758 = ~n21561 & n21757 ;
  assign n21759 = n21758 ^ n21755 ;
  assign n21760 = n21552 & ~n21759 ;
  assign n21761 = n21746 & n21760 ;
  assign n21762 = n21761 ^ n21552 ;
  assign n21773 = ~n21561 & n21723 ;
  assign n21774 = ~n21762 & n21773 ;
  assign n21763 = n21743 ^ n21711 ;
  assign n21764 = n21750 ^ n21720 ;
  assign n21767 = ~n21743 & ~n21764 ;
  assign n21768 = n21767 ^ n21720 ;
  assign n21769 = n21763 & n21768 ;
  assign n21770 = n21769 ^ n21711 ;
  assign n21771 = n21770 ^ n21762 ;
  assign n21732 = n21704 ^ n21632 ;
  assign n21734 = n21733 ^ n21732 ;
  assign n21735 = n21734 ^ n21717 ;
  assign n21736 = n21717 ^ n21561 ;
  assign n21737 = n21736 ^ n21717 ;
  assign n21738 = n21735 & ~n21737 ;
  assign n21739 = n21738 ^ n21717 ;
  assign n21740 = ~n21552 & n21739 ;
  assign n21772 = n21771 ^ n21740 ;
  assign n21775 = n21774 ^ n21772 ;
  assign n21776 = n21723 ^ n21703 ;
  assign n21777 = n21703 ^ n21552 ;
  assign n21778 = n21777 ^ n21703 ;
  assign n21779 = n21776 & n21778 ;
  assign n21780 = n21779 ^ n21703 ;
  assign n21781 = n21561 & n21780 ;
  assign n21782 = ~n21775 & ~n21781 ;
  assign n21783 = n21754 ^ n21734 ;
  assign n21784 = n21754 ^ n21561 ;
  assign n21785 = n21784 ^ n21754 ;
  assign n21786 = n21783 & n21785 ;
  assign n21787 = n21786 ^ n21754 ;
  assign n21788 = n21552 & n21787 ;
  assign n21789 = n21782 & ~n21788 ;
  assign n21790 = ~n21731 & n21789 ;
  assign n21791 = ~n21721 & n21790 ;
  assign n21792 = ~n21719 & n21791 ;
  assign n21794 = n21741 ^ n21725 ;
  assign n21793 = n21726 ^ n21722 ;
  assign n21795 = n21794 ^ n21793 ;
  assign n21796 = ~n21552 & n21795 ;
  assign n21797 = n21796 ^ n21794 ;
  assign n21798 = n21561 & n21797 ;
  assign n21799 = n21792 & ~n21798 ;
  assign n21800 = n21799 ^ n20008 ;
  assign n21801 = n21800 ^ x75 ;
  assign n22625 = n21525 & n21801 ;
  assign n22626 = n22625 ^ n21801 ;
  assign n22446 = n20618 ^ x120 ;
  assign n22447 = n21328 ^ x73 ;
  assign n22480 = n19348 ^ x97 ;
  assign n21949 = n21081 ^ n21062 ;
  assign n21950 = n21081 ^ n20974 ;
  assign n21951 = n21950 ^ n21081 ;
  assign n21952 = n21949 & n21951 ;
  assign n21953 = n21952 ^ n21081 ;
  assign n21954 = ~n20973 & n21953 ;
  assign n21919 = n20975 & n21073 ;
  assign n22461 = n21081 ^ n21052 ;
  assign n22462 = n22461 ^ n21059 ;
  assign n22463 = n22462 ^ n21054 ;
  assign n22464 = n20974 & n22463 ;
  assign n22465 = n22464 ^ n21063 ;
  assign n22466 = n20973 & n22465 ;
  assign n22467 = n22466 ^ n21096 ;
  assign n22460 = n21071 & ~n21126 ;
  assign n22468 = n22467 ^ n22460 ;
  assign n22457 = n21082 ^ n21064 ;
  assign n21924 = n21091 ^ n21059 ;
  assign n22458 = n22457 ^ n21924 ;
  assign n22459 = n21105 & n22458 ;
  assign n22469 = n22468 ^ n22459 ;
  assign n22470 = n22469 ^ n21072 ;
  assign n21958 = n21107 ^ n21093 ;
  assign n21959 = n21093 ^ n20974 ;
  assign n21960 = n21959 ^ n21093 ;
  assign n21961 = n21958 & n21960 ;
  assign n21962 = n21961 ^ n21093 ;
  assign n21963 = ~n20973 & n21962 ;
  assign n22471 = n22470 ^ n21963 ;
  assign n22456 = n20976 & n21086 ;
  assign n22472 = n22471 ^ n22456 ;
  assign n22449 = n21072 ^ n21065 ;
  assign n22450 = n22449 ^ n21072 ;
  assign n22451 = n21072 ^ n20974 ;
  assign n22452 = n22451 ^ n21072 ;
  assign n22453 = n22450 & ~n22452 ;
  assign n22454 = n22453 ^ n21072 ;
  assign n22455 = ~n20973 & n22454 ;
  assign n22473 = n22472 ^ n22455 ;
  assign n22474 = ~n21919 & ~n22473 ;
  assign n22475 = ~n21954 & n22474 ;
  assign n22476 = n22475 ^ n18902 ;
  assign n22477 = n22476 ^ x115 ;
  assign n22512 = n22480 ^ n22477 ;
  assign n22083 = n20880 & n20900 ;
  assign n22481 = ~n20888 & ~n22083 ;
  assign n22489 = n20838 ^ n20829 ;
  assign n22490 = ~n20858 & ~n20890 ;
  assign n22491 = n20864 & n22490 ;
  assign n22492 = n22489 & n22491 ;
  assign n22493 = n22492 ^ n22490 ;
  assign n22494 = n22493 ^ n20890 ;
  assign n22495 = n22494 ^ n20852 ;
  assign n22483 = n20862 ^ n20855 ;
  assign n22084 = n20847 ^ n20839 ;
  assign n22484 = n22483 ^ n22084 ;
  assign n22482 = n20832 ^ n20825 ;
  assign n22485 = n22484 ^ n22482 ;
  assign n22486 = ~n20864 & n22485 ;
  assign n22487 = n22486 ^ n20852 ;
  assign n22488 = n20691 & n22487 ;
  assign n22496 = n22495 ^ n22488 ;
  assign n22497 = n20850 ^ n20691 ;
  assign n22498 = n22497 ^ n20850 ;
  assign n22501 = ~n20845 & ~n20864 ;
  assign n22502 = n22501 ^ n20850 ;
  assign n22503 = ~n22498 & n22502 ;
  assign n22504 = n22503 ^ n20850 ;
  assign n22505 = n22496 & ~n22504 ;
  assign n22113 = n20856 ^ n20845 ;
  assign n22114 = n22113 ^ n20856 ;
  assign n22115 = n20864 & ~n22114 ;
  assign n22116 = n22115 ^ n20856 ;
  assign n22117 = ~n20691 & n22116 ;
  assign n22506 = n22505 ^ n22117 ;
  assign n22507 = n22481 & n22506 ;
  assign n22508 = n22507 ^ n18937 ;
  assign n22509 = n22508 ^ x106 ;
  assign n22562 = n22512 ^ n22509 ;
  assign n22448 = n21185 ^ x80 ;
  assign n22514 = n22509 ^ n22448 ;
  assign n22550 = n22514 ^ n22477 ;
  assign n22551 = n22550 ^ n22480 ;
  assign n22552 = n22551 ^ n22509 ;
  assign n22556 = n22480 & n22509 ;
  assign n22557 = n22556 ^ n22477 ;
  assign n22558 = n22552 & ~n22557 ;
  assign n22559 = n22558 ^ n22514 ;
  assign n22537 = n22477 ^ n22448 ;
  assign n22540 = n22537 ^ n22480 ;
  assign n22545 = n22480 ^ n22448 ;
  assign n22546 = ~n22514 & n22545 ;
  assign n22547 = n22546 ^ n22448 ;
  assign n22548 = ~n22540 & n22547 ;
  assign n22549 = n22548 ^ n22537 ;
  assign n22560 = n22559 ^ n22549 ;
  assign n22478 = ~n22448 & ~n22477 ;
  assign n22479 = n22478 ^ n22477 ;
  assign n22510 = n22509 ^ n22480 ;
  assign n22513 = n22512 ^ n22510 ;
  assign n22515 = n22510 ^ n22509 ;
  assign n22516 = n22514 & ~n22515 ;
  assign n22517 = n22516 ^ n22509 ;
  assign n22518 = ~n22513 & n22517 ;
  assign n22519 = n22518 ^ n22512 ;
  assign n22520 = n22478 & ~n22519 ;
  assign n22511 = n22480 & n22510 ;
  assign n22521 = n22520 ^ n22511 ;
  assign n22522 = n22521 ^ n22480 ;
  assign n22523 = n22522 ^ n22509 ;
  assign n22524 = n22523 ^ n22521 ;
  assign n22525 = n22479 & ~n22524 ;
  assign n22526 = n22525 ^ n22522 ;
  assign n22542 = n22526 ^ n22448 ;
  assign n22561 = n22560 ^ n22542 ;
  assign n22563 = n22562 ^ n22561 ;
  assign n22541 = n22540 ^ n22521 ;
  assign n22564 = n22563 ^ n22541 ;
  assign n22565 = n22564 ^ n22549 ;
  assign n22566 = ~n22447 & ~n22565 ;
  assign n22567 = n22566 ^ n22563 ;
  assign n22538 = n22537 ^ n22526 ;
  assign n22527 = n22510 ^ n22477 ;
  assign n22528 = n22527 ^ n22526 ;
  assign n22529 = n22528 ^ n22511 ;
  assign n22530 = n22529 ^ n22477 ;
  assign n22531 = n22530 ^ n22528 ;
  assign n22532 = n22528 ^ n22448 ;
  assign n22533 = n22532 ^ n22528 ;
  assign n22534 = ~n22531 & ~n22533 ;
  assign n22535 = n22534 ^ n22528 ;
  assign n22536 = ~n22447 & n22535 ;
  assign n22539 = n22538 ^ n22536 ;
  assign n22568 = n22567 ^ n22539 ;
  assign n22569 = n22446 & ~n22568 ;
  assign n22570 = n22569 ^ n22446 ;
  assign n22571 = n22570 ^ n22539 ;
  assign n22572 = n22571 ^ n19966 ;
  assign n22573 = n22572 ^ x108 ;
  assign n21918 = n20390 ^ x126 ;
  assign n21826 = n20615 ^ n18140 ;
  assign n21827 = n21826 ^ n20613 ;
  assign n21811 = n20567 ^ n20509 ;
  assign n21812 = ~n20414 & n21811 ;
  assign n21813 = ~n20393 & ~n20508 ;
  assign n21814 = n21812 & n21813 ;
  assign n21815 = n21814 ^ n21812 ;
  assign n21816 = n21815 ^ n20581 ;
  assign n21817 = n21816 ^ n21815 ;
  assign n21818 = ~n20530 & ~n20554 ;
  assign n21819 = n21817 & n21818 ;
  assign n21820 = n21819 ^ n21816 ;
  assign n21806 = n20529 ^ n20483 ;
  assign n21807 = n21806 ^ n20553 ;
  assign n21808 = n20414 & ~n21807 ;
  assign n21809 = n21808 ^ n20538 ;
  assign n21810 = n20585 & ~n21809 ;
  assign n21822 = n21820 ^ n21810 ;
  assign n21804 = n20393 & ~n20547 ;
  assign n21803 = ~n20414 & n20518 ;
  assign n21805 = n21804 ^ n21803 ;
  assign n21823 = n21822 ^ n21805 ;
  assign n21824 = n21823 ^ n21394 ;
  assign n21825 = ~n20591 & ~n21824 ;
  assign n21828 = n21827 ^ n21825 ;
  assign n21829 = n21828 ^ x69 ;
  assign n21876 = n21324 ^ n18094 ;
  assign n21858 = n21289 ^ n21265 ;
  assign n21859 = n21858 ^ n21241 ;
  assign n21856 = n21293 ^ n21259 ;
  assign n21857 = n21856 ^ n21636 ;
  assign n21860 = n21859 ^ n21857 ;
  assign n21861 = n21190 & ~n21860 ;
  assign n21862 = n21861 ^ n21859 ;
  assign n21863 = ~n21191 & n21862 ;
  assign n21835 = n21651 ^ n21258 ;
  assign n21836 = n21835 ^ n21303 ;
  assign n21837 = n21303 ^ n21191 ;
  assign n21838 = n21308 ^ n21191 ;
  assign n21839 = ~n21837 & n21838 ;
  assign n21840 = n21839 ^ n21191 ;
  assign n21841 = ~n21836 & n21840 ;
  assign n21842 = n21841 ^ n21303 ;
  assign n21843 = n21842 ^ n21238 ;
  assign n21844 = n21843 ^ n21295 ;
  assign n21853 = n21844 ^ n21305 ;
  assign n21845 = n21844 ^ n21300 ;
  assign n21846 = n21845 ^ n21241 ;
  assign n21847 = n21846 ^ n21844 ;
  assign n21848 = n21844 ^ n21191 ;
  assign n21849 = n21848 ^ n21844 ;
  assign n21850 = ~n21847 & n21849 ;
  assign n21851 = n21850 ^ n21844 ;
  assign n21852 = n21190 & n21851 ;
  assign n21854 = n21853 ^ n21852 ;
  assign n21834 = n21285 & ~n21323 ;
  assign n21855 = n21854 ^ n21834 ;
  assign n21864 = n21863 ^ n21855 ;
  assign n21865 = ~n21314 & ~n21864 ;
  assign n21830 = n21266 ^ n21261 ;
  assign n21831 = n21190 & n21830 ;
  assign n21832 = n21831 ^ n21266 ;
  assign n21833 = n21191 & n21832 ;
  assign n21866 = n21865 ^ n21833 ;
  assign n21867 = ~n21635 & n21866 ;
  assign n21870 = n21266 ^ n21190 ;
  assign n21871 = n21870 ^ n21266 ;
  assign n21872 = ~n21302 & ~n21871 ;
  assign n21873 = n21872 ^ n21266 ;
  assign n21874 = ~n21191 & n21873 ;
  assign n21875 = n21867 & ~n21874 ;
  assign n21877 = n21876 ^ n21875 ;
  assign n21878 = n21877 ^ x84 ;
  assign n21879 = ~n21829 & ~n21878 ;
  assign n21880 = n20916 ^ x109 ;
  assign n21892 = n19020 ^ n19009 ;
  assign n21893 = n19281 & n21892 ;
  assign n21887 = n19346 ^ n19020 ;
  assign n21888 = n21887 ^ n21597 ;
  assign n21889 = n21888 ^ n21625 ;
  assign n21882 = n19003 ^ n18820 ;
  assign n21883 = n21882 ^ n18509 ;
  assign n21884 = n21883 ^ n18271 ;
  assign n21885 = ~n18823 & ~n19283 ;
  assign n21886 = ~n21884 & n21885 ;
  assign n21890 = n21889 ^ n21886 ;
  assign n21881 = ~n19029 & ~n19324 ;
  assign n21891 = n21890 ^ n21881 ;
  assign n21894 = n21893 ^ n21891 ;
  assign n21895 = n19319 ^ n19025 ;
  assign n21896 = n21895 ^ n19028 ;
  assign n21897 = n21896 ^ n21895 ;
  assign n21898 = n21895 ^ n19037 ;
  assign n21899 = n21898 ^ n21895 ;
  assign n21900 = n21897 & ~n21899 ;
  assign n21901 = n21900 ^ n21895 ;
  assign n21902 = n19283 & n21901 ;
  assign n21903 = ~n21894 & ~n21902 ;
  assign n21904 = n21903 ^ n18191 ;
  assign n21905 = n21904 ^ x102 ;
  assign n21906 = n21880 & n21905 ;
  assign n22020 = n21879 & n21906 ;
  assign n21910 = n21879 ^ n21829 ;
  assign n21911 = n21910 ^ n21878 ;
  assign n21975 = n21906 ^ n21905 ;
  assign n21992 = ~n21911 & n21975 ;
  assign n21907 = n21906 ^ n21880 ;
  assign n21908 = n21907 ^ n21905 ;
  assign n21914 = n21911 ^ n21829 ;
  assign n21915 = ~n21908 & ~n21914 ;
  assign n21916 = n21915 ^ n21908 ;
  assign n21912 = ~n21908 & ~n21911 ;
  assign n21909 = n21879 & ~n21908 ;
  assign n21913 = n21912 ^ n21909 ;
  assign n21917 = n21916 ^ n21913 ;
  assign n22018 = n21992 ^ n21917 ;
  assign n22008 = n21907 & ~n21914 ;
  assign n21990 = ~n21914 & n21975 ;
  assign n22017 = n22008 ^ n21990 ;
  assign n22019 = n22018 ^ n22017 ;
  assign n22021 = n22020 ^ n22019 ;
  assign n22022 = n21918 & ~n22021 ;
  assign n22005 = n21906 & ~n21910 ;
  assign n22004 = n21879 & n21907 ;
  assign n22006 = n22005 ^ n22004 ;
  assign n22025 = n22022 ^ n22006 ;
  assign n21921 = n20973 & n21079 ;
  assign n21920 = n20974 & n21070 ;
  assign n21922 = n21921 ^ n21920 ;
  assign n21925 = n21081 ^ n21067 ;
  assign n21926 = n21925 ^ n21924 ;
  assign n21927 = ~n20974 & n21926 ;
  assign n21928 = n21927 ^ n21067 ;
  assign n21945 = n21928 ^ n21096 ;
  assign n21946 = n21945 ^ n21113 ;
  assign n21938 = n21073 ^ n21061 ;
  assign n21936 = n21077 ^ n21072 ;
  assign n21937 = n21936 ^ n21068 ;
  assign n21939 = n21938 ^ n21937 ;
  assign n21940 = n21937 ^ n20974 ;
  assign n21941 = n21940 ^ n21937 ;
  assign n21942 = n21939 & n21941 ;
  assign n21943 = n21942 ^ n21937 ;
  assign n21944 = n21126 & n21943 ;
  assign n21947 = n21946 ^ n21944 ;
  assign n21929 = n21928 ^ n20974 ;
  assign n21930 = n21929 ^ n21928 ;
  assign n21931 = n21928 ^ n21079 ;
  assign n21932 = n21931 ^ n21928 ;
  assign n21933 = ~n21930 & n21932 ;
  assign n21934 = n21933 ^ n21928 ;
  assign n21935 = ~n20973 & n21934 ;
  assign n21948 = n21947 ^ n21935 ;
  assign n21955 = ~n21948 & ~n21954 ;
  assign n21923 = n21062 & ~n21104 ;
  assign n21956 = n21955 ^ n21923 ;
  assign n21957 = ~n21922 & n21956 ;
  assign n21964 = n21957 & ~n21963 ;
  assign n21965 = ~n21919 & n21964 ;
  assign n21967 = n20975 & n21085 ;
  assign n21968 = n21965 & n21967 ;
  assign n21966 = n21965 ^ n17974 ;
  assign n21969 = n21968 ^ n21966 ;
  assign n21970 = n21969 ^ x108 ;
  assign n22015 = n21906 & ~n21911 ;
  assign n21976 = ~n21910 & n21975 ;
  assign n21991 = n21990 ^ n21976 ;
  assign n21993 = n21992 ^ n21991 ;
  assign n21994 = n21993 ^ n21975 ;
  assign n21995 = n21994 ^ n21915 ;
  assign n22016 = n22015 ^ n21995 ;
  assign n22023 = n22022 ^ n22016 ;
  assign n22024 = n21970 & n22023 ;
  assign n22026 = n22025 ^ n22024 ;
  assign n21971 = n21918 & ~n21970 ;
  assign n21986 = n21971 ^ n21970 ;
  assign n21987 = n21986 ^ n21918 ;
  assign n21988 = n21987 ^ n21971 ;
  assign n22012 = n21912 & n21970 ;
  assign n22011 = n22006 ^ n21912 ;
  assign n22013 = n22012 ^ n22011 ;
  assign n22014 = ~n21988 & n22013 ;
  assign n22027 = n22026 ^ n22014 ;
  assign n21978 = n21906 & ~n21914 ;
  assign n22007 = n22006 ^ n21978 ;
  assign n22009 = n22008 ^ n22007 ;
  assign n22010 = ~n21986 & n22009 ;
  assign n22028 = n22027 ^ n22010 ;
  assign n22029 = n22028 ^ n21976 ;
  assign n22002 = n21990 ^ n21912 ;
  assign n22003 = n21987 & n22002 ;
  assign n22030 = n22029 ^ n22003 ;
  assign n21989 = n21907 & ~n21910 ;
  assign n21996 = n21995 ^ n21989 ;
  assign n21997 = n21995 ^ n21970 ;
  assign n21998 = n21997 ^ n21995 ;
  assign n21999 = n21996 & n21998 ;
  assign n22000 = n21999 ^ n21995 ;
  assign n22001 = ~n21988 & n22000 ;
  assign n22031 = n22030 ^ n22001 ;
  assign n21974 = n21907 & ~n21911 ;
  assign n21977 = n21976 ^ n21974 ;
  assign n21979 = n21978 ^ n21977 ;
  assign n21980 = n21979 ^ n21976 ;
  assign n21981 = n21976 ^ n21970 ;
  assign n21982 = n21981 ^ n21976 ;
  assign n21983 = n21980 & n21982 ;
  assign n21984 = n21983 ^ n21976 ;
  assign n21985 = n21918 & n21984 ;
  assign n22032 = n22031 ^ n21985 ;
  assign n21972 = n21971 ^ n21918 ;
  assign n21973 = ~n21917 & n21972 ;
  assign n22033 = n22032 ^ n21973 ;
  assign n22038 = n21913 & n21970 ;
  assign n22039 = n22038 ^ n21912 ;
  assign n22040 = n21918 & n22039 ;
  assign n22041 = ~n22033 & ~n22040 ;
  assign n22042 = n22041 ^ n21004 ;
  assign n22043 = n22042 ^ x125 ;
  assign n22277 = n21661 ^ x89 ;
  assign n22099 = n20843 & ~n20864 ;
  assign n22100 = n22099 ^ n20850 ;
  assign n22101 = n22100 ^ n20862 ;
  assign n22102 = ~n20890 & n22101 ;
  assign n22089 = n20835 ^ n20691 ;
  assign n22092 = n20848 ^ n20835 ;
  assign n22090 = n20841 ^ n20827 ;
  assign n22091 = ~n20864 & n22090 ;
  assign n22093 = n22092 ^ n22091 ;
  assign n22094 = n22089 & ~n22093 ;
  assign n22095 = n22094 ^ n20691 ;
  assign n22096 = n22095 ^ n20862 ;
  assign n22085 = n22084 ^ n20880 ;
  assign n22086 = ~n20882 & n22085 ;
  assign n22087 = n22086 ^ n20880 ;
  assign n22088 = n20864 & n22087 ;
  assign n22097 = n22096 ^ n22088 ;
  assign n22103 = n22102 ^ n22097 ;
  assign n22104 = n20851 ^ n20850 ;
  assign n22105 = n20851 ^ n20691 ;
  assign n22106 = n22105 ^ n20851 ;
  assign n22107 = n22104 & ~n22106 ;
  assign n22108 = n22107 ^ n20851 ;
  assign n22109 = n20864 & n22108 ;
  assign n22110 = ~n22103 & ~n22109 ;
  assign n22118 = n22110 & ~n22117 ;
  assign n22119 = ~n22083 & n22118 ;
  assign n22120 = ~n20914 & n22119 ;
  assign n22121 = n22120 ^ n18693 ;
  assign n22278 = n22121 ^ x96 ;
  assign n22426 = ~n22277 & n22278 ;
  assign n22427 = n22426 ^ n22277 ;
  assign n22428 = n22427 ^ n22278 ;
  assign n22291 = n19784 ^ n19451 ;
  assign n22292 = n22291 ^ n19785 ;
  assign n22293 = n22292 ^ n19816 ;
  assign n22294 = n19404 & ~n22293 ;
  assign n22289 = n19828 ^ n19795 ;
  assign n22290 = n22289 ^ n21172 ;
  assign n22295 = n22294 ^ n22290 ;
  assign n22296 = n22295 ^ n19801 ;
  assign n22297 = n22296 ^ n19830 ;
  assign n22298 = n22297 ^ n22295 ;
  assign n22301 = n19404 & n22298 ;
  assign n22302 = n22301 ^ n22295 ;
  assign n22303 = n19405 & n22302 ;
  assign n22304 = n22303 ^ n22295 ;
  assign n22286 = n19812 ^ n19794 ;
  assign n22287 = n22286 ^ n19797 ;
  assign n22288 = n19861 & ~n22287 ;
  assign n22305 = n22304 ^ n22288 ;
  assign n22306 = n22305 ^ n19789 ;
  assign n22307 = n22306 ^ n21165 ;
  assign n22308 = n22307 ^ n21542 ;
  assign n22309 = n22308 ^ n18589 ;
  assign n22285 = n19818 & n19864 ;
  assign n22310 = n22309 ^ n22285 ;
  assign n22313 = n22310 ^ n19825 ;
  assign n22311 = n22310 ^ n19789 ;
  assign n22284 = ~n19404 & n19823 ;
  assign n22312 = n22311 ^ n22284 ;
  assign n22314 = n22313 ^ n22312 ;
  assign n22315 = n22314 ^ n22289 ;
  assign n22316 = n22315 ^ n19825 ;
  assign n22317 = n22316 ^ n22314 ;
  assign n22320 = n19405 & ~n22317 ;
  assign n22321 = n22320 ^ n22314 ;
  assign n22322 = n19845 & ~n22321 ;
  assign n22323 = n22322 ^ n22312 ;
  assign n22324 = n22323 ^ x113 ;
  assign n22342 = n21079 ^ n21060 ;
  assign n22343 = n20976 & n22342 ;
  assign n22336 = n21064 ^ n21058 ;
  assign n22339 = n22336 ^ n21919 ;
  assign n22332 = n21086 ^ n21068 ;
  assign n22333 = n22332 ^ n21092 ;
  assign n22334 = n22333 ^ n21054 ;
  assign n22335 = n20974 & n22334 ;
  assign n22337 = n22336 ^ n22335 ;
  assign n22338 = n21126 & n22337 ;
  assign n22340 = n22339 ^ n22338 ;
  assign n22327 = n21083 ^ n20974 ;
  assign n22328 = n22327 ^ n21083 ;
  assign n22329 = n21084 & ~n22328 ;
  assign n22330 = n22329 ^ n21083 ;
  assign n22331 = n20973 & n22330 ;
  assign n22341 = n22340 ^ n22331 ;
  assign n22344 = n22343 ^ n22341 ;
  assign n22345 = n21091 & ~n22344 ;
  assign n22346 = n20973 & n22345 ;
  assign n22347 = n22346 ^ n21126 ;
  assign n22348 = n21062 ^ n21059 ;
  assign n22349 = n22348 ^ n21095 ;
  assign n22350 = n22349 ^ n21936 ;
  assign n22351 = ~n20974 & ~n22350 ;
  assign n22352 = n22351 ^ n21059 ;
  assign n22353 = n22346 ^ n22344 ;
  assign n22354 = ~n21122 & ~n22353 ;
  assign n22355 = n22352 & n22354 ;
  assign n22356 = ~n22347 & n22355 ;
  assign n22357 = n22356 ^ n22354 ;
  assign n22358 = ~n21954 & n22357 ;
  assign n22359 = n22358 ^ n18552 ;
  assign n22360 = n22359 ^ x74 ;
  assign n22361 = n22324 & ~n22360 ;
  assign n22362 = n22361 ^ n22360 ;
  assign n22363 = n22362 ^ n22324 ;
  assign n22067 = n20150 & ~n20186 ;
  assign n22048 = n20200 ^ n20145 ;
  assign n22049 = n22048 ^ n19937 ;
  assign n22050 = n19968 & ~n22049 ;
  assign n22051 = n22050 ^ n19937 ;
  assign n22054 = n22048 ^ n20199 ;
  assign n22055 = n22051 & n22054 ;
  assign n22052 = n20199 ^ n20187 ;
  assign n22056 = n22055 ^ n22052 ;
  assign n22057 = n22056 ^ n20197 ;
  assign n22064 = n22057 ^ n18647 ;
  assign n22059 = n20141 ^ n19937 ;
  assign n22060 = n22059 ^ n20173 ;
  assign n22061 = n19967 & n22060 ;
  assign n22047 = n20196 ^ n20145 ;
  assign n22058 = n22057 ^ n22047 ;
  assign n22062 = n22061 ^ n22058 ;
  assign n22063 = n20186 & n22062 ;
  assign n22065 = n22064 ^ n22063 ;
  assign n22045 = n20176 ^ n20173 ;
  assign n22046 = n20183 & ~n22045 ;
  assign n22066 = n22065 ^ n22046 ;
  assign n22068 = n22067 ^ n22066 ;
  assign n22044 = n20142 & n20184 ;
  assign n22069 = n22068 ^ n22044 ;
  assign n22070 = n22069 ^ n18647 ;
  assign n22071 = n20148 ^ n20087 ;
  assign n22072 = n20148 ^ n19967 ;
  assign n22073 = n22072 ^ n20148 ;
  assign n22074 = n22071 & ~n22073 ;
  assign n22075 = n22074 ^ n20148 ;
  assign n22076 = ~n19937 & n22075 ;
  assign n22077 = ~n22070 & n22076 ;
  assign n22078 = n22077 ^ n22069 ;
  assign n22280 = n22078 ^ x99 ;
  assign n22281 = n21560 ^ x65 ;
  assign n22282 = n22280 & ~n22281 ;
  assign n22283 = n22282 ^ n22281 ;
  assign n22369 = n22283 ^ n22280 ;
  assign n22431 = n22363 & n22369 ;
  assign n22365 = n22361 ^ n22324 ;
  assign n22383 = n22369 ^ n22281 ;
  assign n22384 = n22365 & n22383 ;
  assign n22385 = n22384 ^ n22365 ;
  assign n22381 = ~n22283 & n22365 ;
  assign n22366 = n22282 & n22365 ;
  assign n22382 = n22381 ^ n22366 ;
  assign n22386 = n22385 ^ n22382 ;
  assign n22372 = n22361 ^ n22280 ;
  assign n22373 = n22281 & n22372 ;
  assign n22374 = n22373 ^ n22281 ;
  assign n22370 = n22361 & n22369 ;
  assign n22371 = n22370 ^ n22369 ;
  assign n22375 = n22374 ^ n22371 ;
  assign n22387 = n22386 ^ n22375 ;
  assign n22435 = n22431 ^ n22387 ;
  assign n22436 = n22435 ^ n22374 ;
  assign n22377 = n22282 & n22363 ;
  assign n22378 = n22377 ^ n22370 ;
  assign n22424 = n22378 ^ n22375 ;
  assign n22406 = n22360 ^ n22324 ;
  assign n22407 = n22281 ^ n22280 ;
  assign n22410 = ~n22360 & n22407 ;
  assign n22411 = n22410 ^ n22280 ;
  assign n22412 = n22406 & n22411 ;
  assign n22425 = n22424 ^ n22412 ;
  assign n22437 = n22436 ^ n22425 ;
  assign n22438 = n22428 & n22437 ;
  assign n22364 = ~n22283 & n22363 ;
  assign n22434 = n22364 & n22426 ;
  assign n22439 = n22438 ^ n22434 ;
  assign n22432 = n22431 ^ n22384 ;
  assign n22433 = ~n22427 & n22432 ;
  assign n22440 = n22439 ^ n22433 ;
  assign n22403 = n22324 ^ n22280 ;
  assign n22367 = ~n22283 & n22361 ;
  assign n22390 = n22367 ^ n22283 ;
  assign n22401 = n22390 ^ n22366 ;
  assign n22393 = n22361 ^ n22282 ;
  assign n22368 = n22367 ^ n22366 ;
  assign n22376 = n22375 ^ n22368 ;
  assign n22379 = n22378 ^ n22376 ;
  assign n22394 = n22393 ^ n22379 ;
  assign n22395 = n22394 ^ n22367 ;
  assign n22396 = n22395 ^ n22363 ;
  assign n22389 = n22381 ^ n22364 ;
  assign n22391 = n22390 ^ n22389 ;
  assign n22392 = n22391 ^ n22370 ;
  assign n22397 = n22396 ^ n22392 ;
  assign n22398 = ~n22277 & n22397 ;
  assign n22388 = n22387 ^ n22370 ;
  assign n22399 = n22398 ^ n22388 ;
  assign n22400 = n22278 & n22399 ;
  assign n22402 = n22401 ^ n22400 ;
  assign n22404 = n22403 ^ n22402 ;
  assign n22405 = n22404 ^ n22400 ;
  assign n22413 = n22412 ^ n22405 ;
  assign n22414 = ~n22278 & ~n22413 ;
  assign n22415 = n22414 ^ n22402 ;
  assign n22441 = n22440 ^ n22415 ;
  assign n22429 = n22428 ^ n22277 ;
  assign n22430 = n22425 & n22429 ;
  assign n22442 = n22441 ^ n22430 ;
  assign n22443 = n22442 ^ n20243 ;
  assign n22279 = n22278 ^ n22277 ;
  assign n22416 = n22415 ^ n22400 ;
  assign n22380 = n22379 ^ n22364 ;
  assign n22417 = n22416 ^ n22380 ;
  assign n22418 = n22417 ^ n22416 ;
  assign n22419 = n22416 ^ n22277 ;
  assign n22420 = n22419 ^ n22416 ;
  assign n22421 = n22418 & n22420 ;
  assign n22422 = n22421 ^ n22416 ;
  assign n22423 = n22279 & ~n22422 ;
  assign n22444 = n22443 ^ n22423 ;
  assign n22445 = n22444 ^ x68 ;
  assign n22590 = n22043 & ~n22445 ;
  assign n22591 = ~n22573 & n22590 ;
  assign n22640 = n22591 ^ n22590 ;
  assign n22574 = n22445 & ~n22573 ;
  assign n22608 = n22574 ^ n22445 ;
  assign n22080 = n21411 ^ x121 ;
  assign n22079 = n22078 ^ x112 ;
  assign n22081 = n22080 ^ n22079 ;
  assign n22082 = n21143 ^ x98 ;
  assign n22122 = n22121 ^ x107 ;
  assign n22123 = ~n22082 & n22122 ;
  assign n22138 = n19022 & ~n19280 ;
  assign n22135 = n19314 ^ n19031 ;
  assign n22136 = ~n19283 & ~n22135 ;
  assign n22132 = n19301 ^ n19282 ;
  assign n22133 = n22132 ^ n21902 ;
  assign n22134 = n22133 ^ n19139 ;
  assign n22137 = n22136 ^ n22134 ;
  assign n22139 = n22138 ^ n22137 ;
  assign n22131 = n19281 & n19305 ;
  assign n22140 = n22139 ^ n22131 ;
  assign n22126 = n19311 ^ n19037 ;
  assign n22127 = n22126 ^ n19311 ;
  assign n22128 = n19312 & ~n22127 ;
  assign n22129 = n22128 ^ n19311 ;
  assign n22130 = n19280 & n22129 ;
  assign n22141 = n22140 ^ n22130 ;
  assign n22142 = n22141 ^ x81 ;
  assign n22143 = n21651 ^ n21303 ;
  assign n22144 = n22143 ^ n21300 ;
  assign n22168 = n22144 ^ n21322 ;
  assign n22157 = ~n21190 & ~n21298 ;
  assign n22158 = n22157 ^ n21292 ;
  assign n22169 = n22168 ^ n22158 ;
  assign n22170 = n22169 ^ n21321 ;
  assign n22171 = n22170 ^ n21874 ;
  assign n22172 = n22171 ^ n19112 ;
  assign n22156 = n21832 ^ n21290 ;
  assign n22159 = n22158 ^ n22156 ;
  assign n22160 = n22159 ^ n21289 ;
  assign n22161 = n22160 ^ n21290 ;
  assign n22162 = n22161 ^ n22159 ;
  assign n22165 = n21190 & n22162 ;
  assign n22166 = n22165 ^ n22159 ;
  assign n22167 = n21191 & n22166 ;
  assign n22173 = n22172 ^ n22167 ;
  assign n22153 = n21292 ^ n21241 ;
  assign n22154 = n22153 ^ n21303 ;
  assign n22155 = n21285 & ~n22154 ;
  assign n22174 = n22173 ^ n22155 ;
  assign n22145 = n22144 ^ n21323 ;
  assign n22146 = n22145 ^ n21265 ;
  assign n22147 = n22146 ^ n22144 ;
  assign n22148 = n22144 ^ n21191 ;
  assign n22149 = n22148 ^ n22144 ;
  assign n22150 = ~n22147 & ~n22149 ;
  assign n22151 = n22150 ^ n22144 ;
  assign n22152 = n21308 & n22151 ;
  assign n22175 = n22174 ^ n22152 ;
  assign n22176 = n22175 ^ x88 ;
  assign n22177 = n22142 & n22176 ;
  assign n22178 = n22177 ^ n22142 ;
  assign n22194 = n22123 & n22178 ;
  assign n22179 = n22178 ^ n22176 ;
  assign n22180 = n22179 ^ n22142 ;
  assign n22184 = n22123 ^ n22122 ;
  assign n22186 = n22184 ^ n22082 ;
  assign n22190 = n22180 & n22186 ;
  assign n22189 = n22177 & n22186 ;
  assign n22191 = n22190 ^ n22189 ;
  assign n22187 = ~n22179 & n22186 ;
  assign n22188 = n22187 ^ n22186 ;
  assign n22192 = n22191 ^ n22188 ;
  assign n22185 = ~n22179 & n22184 ;
  assign n22193 = n22192 ^ n22185 ;
  assign n22195 = n22194 ^ n22193 ;
  assign n22196 = ~n22079 & n22195 ;
  assign n22197 = n22196 ^ n22192 ;
  assign n22181 = n22123 & n22180 ;
  assign n22182 = n22079 & n22181 ;
  assign n22183 = n22182 ^ n22181 ;
  assign n22198 = n22197 ^ n22183 ;
  assign n22199 = ~n22081 & n22198 ;
  assign n22200 = n22199 ^ n22197 ;
  assign n22201 = n22186 ^ n22122 ;
  assign n22205 = ~n22179 & ~n22201 ;
  assign n22236 = n22205 ^ n22181 ;
  assign n22237 = n22236 ^ n22180 ;
  assign n22206 = n22180 & ~n22201 ;
  assign n22207 = n22206 ^ n22189 ;
  assign n22208 = n22207 ^ n22205 ;
  assign n22209 = n22208 ^ n22191 ;
  assign n22238 = n22237 ^ n22209 ;
  assign n22202 = n22178 & ~n22201 ;
  assign n22245 = n22238 ^ n22202 ;
  assign n22211 = n22178 & n22184 ;
  assign n22243 = n22211 ^ n22189 ;
  assign n22244 = n22243 ^ n22205 ;
  assign n22246 = n22245 ^ n22244 ;
  assign n22247 = n22079 & n22246 ;
  assign n22248 = n22247 ^ n22211 ;
  assign n22249 = n22081 & n22248 ;
  assign n22235 = n22123 & n22177 ;
  assign n22239 = n22238 ^ n22235 ;
  assign n22240 = ~n22081 & n22239 ;
  assign n22250 = n22249 ^ n22240 ;
  assign n22234 = n22207 ^ n22192 ;
  assign n22241 = ~n22079 & ~n22240 ;
  assign n22242 = n22234 & n22241 ;
  assign n22251 = n22250 ^ n22242 ;
  assign n22221 = n22205 ^ n22185 ;
  assign n22222 = n22221 ^ n22179 ;
  assign n22223 = n22222 ^ n22187 ;
  assign n22252 = n22251 ^ n22223 ;
  assign n22218 = ~n22079 & ~n22080 ;
  assign n22219 = n22218 ^ n22079 ;
  assign n22220 = n22219 ^ n22080 ;
  assign n22224 = n22223 ^ n22220 ;
  assign n22226 = n22205 ^ n22190 ;
  assign n22225 = n22177 & n22184 ;
  assign n22227 = n22226 ^ n22225 ;
  assign n22228 = n22227 ^ n22219 ;
  assign n22231 = n22223 & n22228 ;
  assign n22232 = n22231 ^ n22219 ;
  assign n22233 = n22224 & n22232 ;
  assign n22253 = n22252 ^ n22233 ;
  assign n22203 = n22202 ^ n22190 ;
  assign n22204 = n22203 ^ n22201 ;
  assign n22210 = n22209 ^ n22204 ;
  assign n22212 = n22211 ^ n22210 ;
  assign n22213 = n22211 ^ n22080 ;
  assign n22214 = n22213 ^ n22211 ;
  assign n22215 = ~n22212 & n22214 ;
  assign n22216 = n22215 ^ n22211 ;
  assign n22217 = ~n22079 & n22216 ;
  assign n22254 = n22253 ^ n22217 ;
  assign n22255 = ~n22200 & n22254 ;
  assign n22263 = n22079 & ~n22080 ;
  assign n22264 = n22235 & n22263 ;
  assign n22258 = n22185 ^ n22079 ;
  assign n22259 = n22258 ^ n22185 ;
  assign n22260 = n22221 & ~n22259 ;
  assign n22261 = n22260 ^ n22185 ;
  assign n22262 = ~n22080 & n22261 ;
  assign n22265 = n22264 ^ n22262 ;
  assign n22266 = n22210 ^ n22187 ;
  assign n22267 = n22266 ^ n22181 ;
  assign n22268 = n22181 ^ n22080 ;
  assign n22269 = n22268 ^ n22181 ;
  assign n22270 = ~n22267 & n22269 ;
  assign n22271 = n22270 ^ n22181 ;
  assign n22272 = n22079 & n22271 ;
  assign n22273 = ~n22265 & ~n22272 ;
  assign n22274 = n22255 & n22273 ;
  assign n22275 = n22274 ^ n21048 ;
  assign n22276 = n22275 ^ x110 ;
  assign n22579 = n22276 & n22573 ;
  assign n22580 = n22445 & n22579 ;
  assign n22609 = n22608 ^ n22580 ;
  assign n22607 = n22579 ^ n22573 ;
  assign n22610 = n22609 ^ n22607 ;
  assign n22618 = n22610 ^ n22445 ;
  assign n22595 = n22276 & n22591 ;
  assign n22596 = n22595 ^ n22591 ;
  assign n22593 = n22590 ^ n22445 ;
  assign n22594 = n22579 & ~n22593 ;
  assign n22597 = n22596 ^ n22594 ;
  assign n22598 = n22597 ^ n22595 ;
  assign n22589 = n22574 ^ n22573 ;
  assign n22592 = n22591 ^ n22589 ;
  assign n22599 = n22598 ^ n22592 ;
  assign n22619 = n22618 ^ n22599 ;
  assign n22641 = n22640 ^ n22619 ;
  assign n22642 = n22641 ^ n22596 ;
  assign n22643 = n22642 ^ n22619 ;
  assign n22636 = n22276 ^ n22043 ;
  assign n22637 = n22636 ^ n22573 ;
  assign n22638 = ~n22445 & ~n22637 ;
  assign n22639 = n22638 ^ n22618 ;
  assign n22644 = n22643 ^ n22639 ;
  assign n22681 = n22626 & ~n22644 ;
  assign n22575 = n22276 & n22574 ;
  assign n22576 = n22575 ^ n22574 ;
  assign n22577 = ~n22043 & n22576 ;
  assign n22578 = n22577 ^ n22576 ;
  assign n22627 = n22626 ^ n21525 ;
  assign n22680 = n22578 & ~n22627 ;
  assign n22682 = n22681 ^ n22680 ;
  assign n22613 = n22043 & n22575 ;
  assign n22668 = n22619 ^ n22613 ;
  assign n22669 = n22619 ^ n21801 ;
  assign n22670 = n22669 ^ n22619 ;
  assign n22671 = n22668 & n22670 ;
  assign n22672 = n22671 ^ n22619 ;
  assign n22673 = n21525 & n22672 ;
  assign n22614 = n22613 ^ n22575 ;
  assign n22581 = ~n22043 & n22580 ;
  assign n22615 = n22614 ^ n22581 ;
  assign n22616 = n22615 ^ n22577 ;
  assign n22612 = n22593 ^ n22043 ;
  assign n22617 = n22616 ^ n22612 ;
  assign n22631 = n22617 ^ n22609 ;
  assign n22655 = n22631 ^ n22613 ;
  assign n22652 = n22641 ^ n22610 ;
  assign n22653 = n22652 ^ n22596 ;
  assign n21802 = n21801 ^ n21525 ;
  assign n22645 = n22644 ^ n22592 ;
  assign n22635 = n22617 ^ n22577 ;
  assign n22646 = n22645 ^ n22635 ;
  assign n22647 = n22635 ^ n21525 ;
  assign n22648 = n22647 ^ n22635 ;
  assign n22649 = n22646 & n22648 ;
  assign n22650 = n22649 ^ n22635 ;
  assign n22651 = n21802 & n22650 ;
  assign n22654 = n22653 ^ n22651 ;
  assign n22656 = n22655 ^ n22654 ;
  assign n22657 = n22656 ^ n22651 ;
  assign n22658 = ~n21525 & n22657 ;
  assign n22659 = n22658 ^ n22654 ;
  assign n22674 = n22673 ^ n22659 ;
  assign n22660 = n22659 ^ n22651 ;
  assign n22629 = n22581 ^ n22580 ;
  assign n22661 = n22660 ^ n22629 ;
  assign n22662 = n22661 ^ n22660 ;
  assign n22663 = n22660 ^ n21801 ;
  assign n22664 = n22663 ^ n22660 ;
  assign n22665 = n22662 & n22664 ;
  assign n22666 = n22665 ^ n22660 ;
  assign n22667 = ~n21802 & n22666 ;
  assign n22675 = n22674 ^ n22667 ;
  assign n22628 = n22627 ^ n21801 ;
  assign n22632 = n22631 ^ n22578 ;
  assign n22630 = n22629 ^ n22614 ;
  assign n22633 = n22632 ^ n22630 ;
  assign n22634 = n22628 & n22633 ;
  assign n22676 = n22675 ^ n22634 ;
  assign n22620 = n22619 ^ n22617 ;
  assign n22606 = n22595 ^ n22581 ;
  assign n22611 = n22610 ^ n22606 ;
  assign n22621 = n22620 ^ n22611 ;
  assign n22622 = ~n21525 & n22621 ;
  assign n22623 = n22622 ^ n22620 ;
  assign n22624 = ~n21802 & n22623 ;
  assign n22677 = n22676 ^ n22624 ;
  assign n22678 = n22677 ^ n22592 ;
  assign n22601 = n22592 ^ n21525 ;
  assign n22602 = n22601 ^ n22592 ;
  assign n22603 = n22598 & ~n22602 ;
  assign n22604 = n22603 ^ n22592 ;
  assign n22605 = n21802 & ~n22604 ;
  assign n22679 = n22678 ^ n22605 ;
  assign n22683 = n22682 ^ n22679 ;
  assign n22582 = n22581 ^ n22578 ;
  assign n22583 = n22582 ^ n22577 ;
  assign n22584 = n22577 ^ n21525 ;
  assign n22585 = n22584 ^ n22577 ;
  assign n22586 = n22583 & n22585 ;
  assign n22587 = n22586 ^ n22577 ;
  assign n22588 = ~n21802 & n22587 ;
  assign n22684 = n22683 ^ n22588 ;
  assign n22685 = n22684 ^ n21143 ;
  assign n22972 = n20972 ^ x74 ;
  assign n22930 = n22436 ^ n22381 ;
  assign n22931 = ~n22427 & n22930 ;
  assign n22927 = n22429 & n22435 ;
  assign n22924 = ~n22384 & ~n22428 ;
  assign n22925 = n22373 & ~n22924 ;
  assign n22918 = n22395 ^ n22364 ;
  assign n22919 = n22918 ^ n22377 ;
  assign n22920 = ~n22427 & n22919 ;
  assign n22916 = n22394 & n22429 ;
  assign n22917 = n22916 ^ n22434 ;
  assign n22921 = n22920 ^ n22917 ;
  assign n22911 = n22370 ^ n22278 ;
  assign n22912 = n22911 ^ n22370 ;
  assign n22913 = ~n22392 & n22912 ;
  assign n22914 = n22913 ^ n22370 ;
  assign n22915 = ~n22279 & n22914 ;
  assign n22922 = n22921 ^ n22915 ;
  assign n22923 = n22922 ^ n18819 ;
  assign n22926 = n22925 ^ n22923 ;
  assign n22928 = n22927 ^ n22926 ;
  assign n22901 = n22425 ^ n22387 ;
  assign n22903 = n22901 ^ n22394 ;
  assign n22890 = n22382 ^ n22364 ;
  assign n22904 = n22903 ^ n22890 ;
  assign n22905 = n22904 ^ n22403 ;
  assign n22906 = n22905 ^ n22380 ;
  assign n22902 = n22901 ^ n22391 ;
  assign n22907 = n22906 ^ n22902 ;
  assign n22908 = n22426 & ~n22907 ;
  assign n22929 = n22928 ^ n22908 ;
  assign n22932 = n22931 ^ n22929 ;
  assign n22900 = n22368 & n22429 ;
  assign n22933 = n22932 ^ n22900 ;
  assign n22891 = n22390 ^ n22372 ;
  assign n22892 = n22891 ^ n22374 ;
  assign n22893 = n22892 ^ n22890 ;
  assign n22894 = n22893 ^ n22892 ;
  assign n22895 = n22892 ^ n22277 ;
  assign n22896 = n22895 ^ n22892 ;
  assign n22897 = n22894 & n22896 ;
  assign n22898 = n22897 ^ n22892 ;
  assign n22899 = n22279 & n22898 ;
  assign n22934 = n22933 ^ n22899 ;
  assign n22935 = n22934 ^ x106 ;
  assign n22553 = n22509 ^ n22477 ;
  assign n22941 = n22537 ^ n22477 ;
  assign n22942 = ~n22553 & n22941 ;
  assign n22943 = n22942 ^ n22477 ;
  assign n22944 = n22510 & n22943 ;
  assign n22945 = n22944 ^ n22537 ;
  assign n22947 = n22446 & ~n22945 ;
  assign n22946 = n22945 ^ n22446 ;
  assign n22948 = n22947 ^ n22946 ;
  assign n22949 = n22948 ^ n22519 ;
  assign n22957 = n22949 ^ n19002 ;
  assign n22936 = n22521 ^ n22519 ;
  assign n22937 = n22936 ^ n22561 ;
  assign n22940 = n22937 ^ n22559 ;
  assign n22950 = n22949 ^ n22940 ;
  assign n22939 = n22549 ^ n22519 ;
  assign n22951 = n22950 ^ n22939 ;
  assign n22954 = n22446 & ~n22951 ;
  assign n22955 = n22954 ^ n22950 ;
  assign n22956 = ~n22447 & n22955 ;
  assign n22958 = n22957 ^ n22956 ;
  assign n22938 = n22446 & ~n22937 ;
  assign n22959 = n22958 ^ n22938 ;
  assign n22960 = n22959 ^ x97 ;
  assign n22961 = n22935 & n22960 ;
  assign n22982 = n22961 ^ n22935 ;
  assign n22983 = n22982 ^ n22960 ;
  assign n22775 = n21904 ^ x77 ;
  assign n22776 = n21589 ^ x68 ;
  assign n22779 = n22775 & ~n22776 ;
  assign n22780 = n22779 ^ n22775 ;
  assign n22721 = n20387 ^ n20360 ;
  assign n22722 = n22721 ^ n18306 ;
  assign n22723 = n22722 ^ x117 ;
  assign n22724 = n21551 ^ x94 ;
  assign n22725 = n22723 & n22724 ;
  assign n22726 = n22725 ^ n22724 ;
  assign n22727 = n22726 ^ n22723 ;
  assign n22728 = n21969 ^ x100 ;
  assign n22729 = ~n20691 & n20866 ;
  assign n22744 = n20883 ^ n20837 ;
  assign n22745 = n22744 ^ n20905 ;
  assign n22746 = n20864 & ~n22745 ;
  assign n22747 = n22746 ^ n20856 ;
  assign n22748 = ~n20691 & n22747 ;
  assign n22749 = n22748 ^ n20856 ;
  assign n22740 = n22483 ^ n20850 ;
  assign n22741 = ~n20864 & n22740 ;
  assign n22742 = n22741 ^ n20850 ;
  assign n22743 = ~n20890 & n22742 ;
  assign n22750 = n22749 ^ n22743 ;
  assign n22751 = n22750 ^ n20843 ;
  assign n22731 = n22482 ^ n20841 ;
  assign n22730 = n22482 ^ n20883 ;
  assign n22732 = n22731 ^ n22730 ;
  assign n22733 = n22730 ^ n20864 ;
  assign n22734 = n22733 ^ n22730 ;
  assign n22735 = ~n22732 & ~n22734 ;
  assign n22736 = n22735 ^ n22730 ;
  assign n22737 = ~n20890 & ~n22736 ;
  assign n22738 = n22737 ^ n20843 ;
  assign n22739 = ~n20900 & n22738 ;
  assign n22752 = n22751 ^ n22739 ;
  assign n22753 = ~n22109 & ~n22752 ;
  assign n22754 = ~n22729 & n22753 ;
  assign n22755 = n22754 ^ n22083 ;
  assign n22756 = ~n20914 & n22755 ;
  assign n22757 = n22756 ^ n18351 ;
  assign n22758 = n22757 ^ x75 ;
  assign n22759 = n22728 & n22758 ;
  assign n22760 = n22759 ^ n22758 ;
  assign n22771 = n22760 ^ n22728 ;
  assign n22794 = ~n22727 & ~n22771 ;
  assign n22787 = n22725 & n22760 ;
  assign n22786 = n22724 & n22760 ;
  assign n22788 = n22787 ^ n22786 ;
  assign n22838 = n22794 ^ n22788 ;
  assign n22839 = n22780 & n22838 ;
  assign n22770 = n22725 ^ n22723 ;
  assign n22807 = n22770 & ~n22771 ;
  assign n22837 = n22780 & n22807 ;
  assign n22840 = n22839 ^ n22837 ;
  assign n22841 = n22840 ^ n18508 ;
  assign n22777 = n22727 ^ n22725 ;
  assign n22798 = n22777 ^ n22728 ;
  assign n22764 = n22758 ^ n22723 ;
  assign n22765 = n22758 ^ n22724 ;
  assign n22766 = ~n22758 & ~n22765 ;
  assign n22767 = n22766 ^ n22759 ;
  assign n22768 = ~n22764 & ~n22767 ;
  assign n22799 = n22798 ^ n22768 ;
  assign n22796 = n22725 & n22759 ;
  assign n22772 = n22771 ^ n22758 ;
  assign n22773 = n22770 & n22772 ;
  assign n22782 = n22773 ^ n22772 ;
  assign n22781 = n22724 & n22772 ;
  assign n22783 = n22782 ^ n22781 ;
  assign n22797 = n22796 ^ n22783 ;
  assign n22800 = n22799 ^ n22797 ;
  assign n22793 = n22765 ^ n22728 ;
  assign n22795 = n22794 ^ n22793 ;
  assign n22801 = n22800 ^ n22795 ;
  assign n22804 = n22801 ^ n22788 ;
  assign n22761 = ~n22727 & n22760 ;
  assign n22762 = n22761 ^ n22760 ;
  assign n22763 = n22762 ^ n22726 ;
  assign n22769 = n22768 ^ n22763 ;
  assign n22805 = n22804 ^ n22769 ;
  assign n22791 = n22725 & n22772 ;
  assign n22792 = n22791 ^ n22781 ;
  assign n22802 = n22801 ^ n22792 ;
  assign n22803 = n22802 ^ n22726 ;
  assign n22806 = n22805 ^ n22803 ;
  assign n22808 = n22807 ^ n22806 ;
  assign n22790 = n22786 ^ n22762 ;
  assign n22809 = n22808 ^ n22790 ;
  assign n22778 = n22728 & ~n22777 ;
  assign n22784 = ~n22780 & ~n22783 ;
  assign n22785 = n22778 & ~n22784 ;
  assign n22789 = n22788 ^ n22785 ;
  assign n22810 = n22809 ^ n22789 ;
  assign n22811 = n22810 ^ n22785 ;
  assign n22812 = n22785 ^ n22775 ;
  assign n22813 = n22812 ^ n22785 ;
  assign n22814 = n22811 & ~n22813 ;
  assign n22815 = n22814 ^ n22785 ;
  assign n22816 = ~n22776 & n22815 ;
  assign n22817 = n22816 ^ n22785 ;
  assign n22821 = n22796 ^ n22761 ;
  assign n22819 = n22794 ^ n22787 ;
  assign n22818 = n22792 ^ n22790 ;
  assign n22820 = n22819 ^ n22818 ;
  assign n22822 = n22821 ^ n22820 ;
  assign n22823 = ~n22775 & n22822 ;
  assign n22824 = n22823 ^ n22790 ;
  assign n22825 = n22824 ^ n22799 ;
  assign n22826 = n22825 ^ n22800 ;
  assign n22827 = n22826 ^ n22825 ;
  assign n22830 = ~n22775 & ~n22827 ;
  assign n22831 = n22830 ^ n22825 ;
  assign n22832 = ~n22776 & ~n22831 ;
  assign n22833 = n22832 ^ n22824 ;
  assign n22834 = ~n22817 & ~n22833 ;
  assign n22842 = n22841 ^ n22834 ;
  assign n22774 = n22773 ^ n22769 ;
  assign n22835 = ~n22775 & n22834 ;
  assign n22836 = n22774 & n22835 ;
  assign n22843 = n22842 ^ n22836 ;
  assign n22844 = n22843 ^ x115 ;
  assign n22882 = n22005 ^ n21974 ;
  assign n22883 = n21971 & n22882 ;
  assign n22881 = ~n21986 & n22015 ;
  assign n22884 = n22883 ^ n22881 ;
  assign n22845 = ~n21986 & n21989 ;
  assign n22846 = n22845 ^ n22003 ;
  assign n22874 = n22018 ^ n21995 ;
  assign n22875 = n22874 ^ n22006 ;
  assign n22876 = ~n21986 & ~n22875 ;
  assign n22864 = n22015 ^ n21974 ;
  assign n22862 = n21879 & ~n21880 ;
  assign n22863 = n22862 ^ n22020 ;
  assign n22865 = n22864 ^ n22863 ;
  assign n22866 = n22865 ^ n21971 ;
  assign n22867 = n21987 & ~n22866 ;
  assign n22868 = n22867 ^ n21971 ;
  assign n22853 = n21992 ^ n21915 ;
  assign n22854 = ~n21971 & ~n22853 ;
  assign n22855 = n22854 ^ n21990 ;
  assign n22856 = n21918 & ~n22855 ;
  assign n22870 = n22856 ^ n21987 ;
  assign n22869 = n22856 ^ n22008 ;
  assign n22871 = n22870 ^ n22869 ;
  assign n22872 = n22868 & n22871 ;
  assign n22873 = n22872 ^ n22870 ;
  assign n22877 = n22876 ^ n22873 ;
  assign n22849 = n21976 ^ n21909 ;
  assign n22850 = n22849 ^ n21978 ;
  assign n22851 = n22850 ^ n22018 ;
  assign n22852 = n22851 ^ n21978 ;
  assign n22859 = n22852 & n22856 ;
  assign n22860 = n22859 ^ n21978 ;
  assign n22861 = n21971 & n22860 ;
  assign n22878 = n22877 ^ n22861 ;
  assign n22847 = n22007 ^ n21974 ;
  assign n22848 = n21972 & n22847 ;
  assign n22879 = n22878 ^ n22848 ;
  assign n22880 = ~n22846 & ~n22879 ;
  assign n22885 = n22884 ^ n22880 ;
  assign n22886 = n22885 ^ n21973 ;
  assign n22887 = n22886 ^ n18270 ;
  assign n22888 = n22887 ^ x96 ;
  assign n22889 = n22844 & n22888 ;
  assign n22965 = n22889 ^ n22888 ;
  assign n22987 = n22965 ^ n22844 ;
  assign n22988 = ~n22983 & ~n22987 ;
  assign n23046 = n22972 & n22988 ;
  assign n23011 = n22961 & ~n22987 ;
  assign n23010 = n22889 & n22961 ;
  assign n23012 = n23011 ^ n23010 ;
  assign n23008 = n22961 & n22965 ;
  assign n23009 = n23008 ^ n22961 ;
  assign n23013 = n23012 ^ n23009 ;
  assign n22714 = n22218 & n22225 ;
  assign n22687 = n22238 ^ n22223 ;
  assign n22711 = n22218 & ~n22687 ;
  assign n22702 = n22194 ^ n22181 ;
  assign n22703 = n22702 ^ n22187 ;
  assign n22704 = n22187 ^ n22079 ;
  assign n22705 = n22704 ^ n22187 ;
  assign n22706 = n22703 & n22705 ;
  assign n22707 = n22706 ^ n22187 ;
  assign n22708 = n22081 & n22707 ;
  assign n22709 = n22708 ^ n22182 ;
  assign n22697 = n22235 ^ n22207 ;
  assign n22698 = n22697 ^ n22245 ;
  assign n22699 = ~n22079 & n22698 ;
  assign n22710 = n22709 ^ n22699 ;
  assign n22712 = n22711 ^ n22710 ;
  assign n22713 = n22712 ^ n22265 ;
  assign n22715 = n22714 ^ n22713 ;
  assign n22696 = n22266 ^ n22192 ;
  assign n22700 = n22699 ^ n22696 ;
  assign n22701 = ~n22081 & ~n22700 ;
  assign n22716 = n22715 ^ n22701 ;
  assign n22688 = n22687 ^ n22206 ;
  assign n22689 = n22688 ^ n22211 ;
  assign n22686 = n22227 ^ n22210 ;
  assign n22690 = n22689 ^ n22686 ;
  assign n22691 = n22686 ^ n22080 ;
  assign n22692 = n22691 ^ n22686 ;
  assign n22693 = n22690 & n22692 ;
  assign n22694 = n22693 ^ n22686 ;
  assign n22695 = n22079 & ~n22694 ;
  assign n22717 = n22716 ^ n22695 ;
  assign n22718 = ~n22200 & ~n22717 ;
  assign n22719 = n22718 ^ n19279 ;
  assign n22720 = n22719 ^ x64 ;
  assign n22978 = n22972 ^ n22720 ;
  assign n22979 = ~n22972 & n22978 ;
  assign n23042 = n23013 ^ n22979 ;
  assign n22967 = n22889 ^ n22844 ;
  assign n22995 = n22967 & n22982 ;
  assign n22980 = n22979 ^ n22720 ;
  assign n22981 = n22980 ^ n22972 ;
  assign n23043 = n22995 ^ n22981 ;
  assign n23044 = n23042 & n23043 ;
  assign n22994 = n22965 & n22982 ;
  assign n22996 = n22995 ^ n22994 ;
  assign n23024 = n22979 ^ n22972 ;
  assign n23038 = n22996 & ~n23024 ;
  assign n23034 = n22980 & n22994 ;
  assign n22997 = n22982 & ~n22987 ;
  assign n22998 = n22997 ^ n22982 ;
  assign n22999 = n22998 ^ n22996 ;
  assign n23032 = n23008 ^ n22999 ;
  assign n23033 = n22979 & n23032 ;
  assign n23035 = n23034 ^ n23033 ;
  assign n22986 = n22965 & ~n22983 ;
  assign n22989 = n22988 ^ n22986 ;
  assign n22984 = n22889 & ~n22983 ;
  assign n22985 = n22984 ^ n22983 ;
  assign n22990 = n22989 ^ n22985 ;
  assign n23029 = n22979 & ~n22990 ;
  assign n23028 = n22978 & n22986 ;
  assign n23030 = n23029 ^ n23028 ;
  assign n22962 = n22961 ^ n22960 ;
  assign n22968 = n22962 & n22967 ;
  assign n22966 = n22962 & n22965 ;
  assign n22969 = n22968 ^ n22966 ;
  assign n22963 = n22889 & n22962 ;
  assign n22964 = n22963 ^ n22962 ;
  assign n22970 = n22969 ^ n22964 ;
  assign n22971 = n22970 ^ n22966 ;
  assign n23025 = n22971 & ~n23024 ;
  assign n23014 = n23013 ^ n22997 ;
  assign n23015 = n23014 ^ n23012 ;
  assign n23018 = n23015 ^ n22720 ;
  assign n23019 = n23018 ^ n23015 ;
  assign n23020 = n23011 & n23019 ;
  assign n23021 = n23020 ^ n23015 ;
  assign n23022 = ~n22978 & n23021 ;
  assign n23023 = n23022 ^ n23012 ;
  assign n23026 = n23025 ^ n23023 ;
  assign n22993 = n22984 ^ n22963 ;
  assign n23027 = n23026 ^ n22993 ;
  assign n23031 = n23030 ^ n23027 ;
  assign n23036 = n23035 ^ n23031 ;
  assign n23000 = n22999 ^ n22968 ;
  assign n23003 = n22993 ^ n22720 ;
  assign n23004 = n23003 ^ n22993 ;
  assign n23005 = n23000 & ~n23004 ;
  assign n23006 = n23005 ^ n22993 ;
  assign n23007 = n22978 & n23006 ;
  assign n23037 = n23036 ^ n23007 ;
  assign n23039 = n23038 ^ n23037 ;
  assign n22991 = n22981 & ~n22990 ;
  assign n22975 = n22971 & ~n22972 ;
  assign n22976 = n22975 ^ n22966 ;
  assign n22977 = n22720 & n22976 ;
  assign n22992 = n22991 ^ n22977 ;
  assign n23040 = n23039 ^ n22992 ;
  assign n23041 = n23040 ^ n19348 ;
  assign n23045 = n23044 ^ n23041 ;
  assign n23047 = n23046 ^ n23045 ;
  assign n23066 = n21461 ^ n21458 ;
  assign n23067 = n23066 ^ n21502 ;
  assign n23068 = n21187 & n23067 ;
  assign n23063 = ~n21460 & ~n21482 ;
  assign n23056 = n21453 ^ n21412 ;
  assign n23057 = n23056 ^ n21456 ;
  assign n23058 = n23057 ^ n21458 ;
  assign n23059 = ~n21144 & ~n23058 ;
  assign n23060 = n23059 ^ n21487 ;
  assign n23061 = ~n21186 & ~n23060 ;
  assign n23053 = n21187 & ~n21488 ;
  assign n23052 = n21189 & n21480 ;
  assign n23054 = n23053 ^ n23052 ;
  assign n23051 = n21457 ^ n20130 ;
  assign n23055 = n23054 ^ n23051 ;
  assign n23062 = n23061 ^ n23055 ;
  assign n23064 = n23063 ^ n23062 ;
  assign n23049 = n21488 ^ n21464 ;
  assign n23050 = n21188 & ~n23049 ;
  assign n23065 = n23064 ^ n23050 ;
  assign n23069 = n23068 ^ n23065 ;
  assign n23048 = n21448 & n21460 ;
  assign n23070 = n23069 ^ n23048 ;
  assign n23099 = ~n22990 & ~n23024 ;
  assign n23097 = n23011 ^ n22995 ;
  assign n23098 = n22980 & n23097 ;
  assign n23100 = n23099 ^ n23098 ;
  assign n23101 = n23100 ^ n23030 ;
  assign n23096 = n22981 & n23032 ;
  assign n23102 = n23101 ^ n23096 ;
  assign n23103 = n23102 ^ n23014 ;
  assign n23094 = n23033 ^ n22991 ;
  assign n23084 = n22720 & n22989 ;
  assign n23085 = n23084 ^ n22988 ;
  assign n23086 = n23085 ^ n22966 ;
  assign n23087 = n23086 ^ n23085 ;
  assign n23090 = n22720 & n23087 ;
  assign n23091 = n23090 ^ n23085 ;
  assign n23092 = n22978 & n23091 ;
  assign n23093 = n23092 ^ n23085 ;
  assign n23095 = n23094 ^ n23093 ;
  assign n23104 = n23103 ^ n23095 ;
  assign n23077 = n23008 ^ n22988 ;
  assign n23078 = n23077 ^ n22968 ;
  assign n23081 = n22972 & n23078 ;
  assign n23082 = n23081 ^ n22968 ;
  assign n23083 = n22720 & n23082 ;
  assign n23105 = n23104 ^ n23083 ;
  assign n23073 = n23012 ^ n22963 ;
  assign n23074 = ~n22720 & n23073 ;
  assign n23072 = n23014 ^ n22970 ;
  assign n23075 = n23074 ^ n23072 ;
  assign n23076 = ~n22978 & n23075 ;
  assign n23106 = n23105 ^ n23076 ;
  assign n23107 = n23106 ^ n23038 ;
  assign n23108 = n23107 ^ n21904 ;
  assign n23071 = n22972 & n22993 ;
  assign n23109 = n23108 ^ n23071 ;
  assign n23139 = n22779 ^ n22776 ;
  assign n23140 = n23139 ^ n22775 ;
  assign n23144 = n22806 & n23140 ;
  assign n23141 = n22807 ^ n22787 ;
  assign n23142 = n23141 ^ n22783 ;
  assign n23143 = n23140 & n23142 ;
  assign n23145 = n23144 ^ n23143 ;
  assign n23121 = ~n22727 & n22759 ;
  assign n23114 = n22787 ^ n22769 ;
  assign n23110 = n22786 ^ n22783 ;
  assign n23111 = n23110 ^ n22801 ;
  assign n23112 = n23111 ^ n22808 ;
  assign n23113 = ~n22776 & ~n23112 ;
  assign n23115 = n23114 ^ n23113 ;
  assign n23116 = n22776 ^ n22775 ;
  assign n23117 = n22821 & n23116 ;
  assign n23118 = n22775 & ~n23117 ;
  assign n23119 = n23115 & n23118 ;
  assign n23120 = n23119 ^ n23117 ;
  assign n23122 = n23121 ^ n23120 ;
  assign n23146 = n23145 ^ n23122 ;
  assign n23131 = n22801 ^ n22791 ;
  assign n23132 = n23131 ^ n22781 ;
  assign n23133 = n23132 ^ n22791 ;
  assign n23134 = n22791 ^ n22775 ;
  assign n23135 = n23134 ^ n22791 ;
  assign n23136 = ~n23133 & n23135 ;
  assign n23137 = n23136 ^ n22791 ;
  assign n23138 = n22776 & n23137 ;
  assign n23147 = n23146 ^ n23138 ;
  assign n23148 = n23147 ^ n22840 ;
  assign n23149 = n23148 ^ n20413 ;
  assign n23124 = n23121 ^ n22775 ;
  assign n23125 = n23124 ^ n23121 ;
  assign n23126 = n23121 ^ n22799 ;
  assign n23127 = n23126 ^ n23121 ;
  assign n23128 = ~n23125 & ~n23127 ;
  assign n23129 = n23128 ^ n23121 ;
  assign n23130 = ~n22776 & n23129 ;
  assign n23150 = n23149 ^ n23130 ;
  assign n23151 = n23070 ^ x69 ;
  assign n23152 = ~n22881 & ~n22883 ;
  assign n23175 = n21970 & n22020 ;
  assign n23156 = n22854 ^ n21976 ;
  assign n23159 = n21995 ^ n21917 ;
  assign n23160 = ~n21972 & n23159 ;
  assign n23161 = ~n23156 & n23160 ;
  assign n23155 = n22004 ^ n21978 ;
  assign n23157 = n23156 ^ n23155 ;
  assign n23162 = n23161 ^ n23157 ;
  assign n23171 = n23162 ^ n22846 ;
  assign n23172 = n23171 ^ n22001 ;
  assign n23163 = n23162 ^ n22849 ;
  assign n23164 = n23163 ^ n22017 ;
  assign n23165 = n23164 ^ n23162 ;
  assign n23166 = n23162 ^ n21970 ;
  assign n23167 = n23166 ^ n23162 ;
  assign n23168 = n23165 & ~n23167 ;
  assign n23169 = n23168 ^ n23162 ;
  assign n23170 = ~n21918 & ~n23169 ;
  assign n23173 = n23172 ^ n23170 ;
  assign n23153 = n22847 ^ n21917 ;
  assign n23154 = n21987 & ~n23153 ;
  assign n23174 = n23173 ^ n23154 ;
  assign n23176 = n23175 ^ n23174 ;
  assign n23177 = ~n22040 & n23176 ;
  assign n23178 = n23152 & n23177 ;
  assign n23179 = n23178 ^ n20739 ;
  assign n23180 = n23179 ^ x91 ;
  assign n23181 = ~n23151 & ~n23180 ;
  assign n23182 = n23181 ^ n23180 ;
  assign n23183 = n23182 ^ n23151 ;
  assign n23230 = n20935 ^ n20643 ;
  assign n23242 = n23230 ^ n20641 ;
  assign n23243 = n23242 ^ n20924 ;
  assign n23236 = n20391 ^ n19895 ;
  assign n23237 = ~n20619 & n23236 ;
  assign n23235 = n20937 ^ n20647 ;
  assign n23238 = n23237 ^ n23235 ;
  assign n23239 = ~n20917 & ~n23238 ;
  assign n23240 = n23239 ^ n23237 ;
  assign n23241 = n23240 ^ n20658 ;
  assign n23244 = n23243 ^ n23241 ;
  assign n23245 = n23244 ^ n23240 ;
  assign n23248 = ~n20917 & n23245 ;
  assign n23249 = n23248 ^ n23240 ;
  assign n23250 = n19349 & n23249 ;
  assign n23251 = n23250 ^ n23240 ;
  assign n23228 = n20639 ^ n20624 ;
  assign n23229 = n23228 ^ n20924 ;
  assign n23231 = n23230 ^ n23229 ;
  assign n23232 = n19349 & ~n23231 ;
  assign n23233 = n23232 ^ n20936 ;
  assign n23234 = n20917 & ~n23233 ;
  assign n23252 = n23251 ^ n23234 ;
  assign n23253 = ~n20960 & ~n23252 ;
  assign n23226 = n20928 & ~n20946 ;
  assign n23225 = n20641 & n20926 ;
  assign n23227 = n23226 ^ n23225 ;
  assign n23254 = n23253 ^ n23227 ;
  assign n23255 = ~n20969 & n23254 ;
  assign n23256 = n23255 ^ n19936 ;
  assign n23257 = n23256 ^ x92 ;
  assign n23258 = n21750 ^ n21703 ;
  assign n23259 = ~n21552 & n23258 ;
  assign n23260 = n23259 ^ n21703 ;
  assign n23263 = n23260 ^ n21794 ;
  assign n23264 = n23263 ^ n23260 ;
  assign n23265 = ~n21552 & n23264 ;
  assign n23266 = n23265 ^ n23260 ;
  assign n23267 = n21561 & n23266 ;
  assign n23268 = n23267 ^ n23260 ;
  assign n23269 = ~n21719 & ~n23268 ;
  assign n23285 = n21754 ^ n21746 ;
  assign n23277 = n21751 ^ n21717 ;
  assign n23279 = n21733 ^ n21721 ;
  assign n23278 = n21750 ^ n21697 ;
  assign n23280 = n23279 ^ n23278 ;
  assign n23281 = ~n21710 & n23280 ;
  assign n23282 = ~n23277 & n23281 ;
  assign n23283 = n23282 ^ n23280 ;
  assign n23284 = n23283 ^ n21723 ;
  assign n23286 = n23285 ^ n23284 ;
  assign n23287 = n23286 ^ n23283 ;
  assign n23288 = n23283 ^ n21561 ;
  assign n23289 = n23288 ^ n23283 ;
  assign n23290 = ~n23287 & ~n23289 ;
  assign n23291 = n23290 ^ n23283 ;
  assign n23292 = ~n21552 & n23291 ;
  assign n23293 = n23292 ^ n23283 ;
  assign n23270 = n21746 ^ n21728 ;
  assign n23271 = n23270 ^ n21734 ;
  assign n23272 = n21734 ^ n21552 ;
  assign n23273 = n23272 ^ n21734 ;
  assign n23274 = ~n23271 & n23273 ;
  assign n23275 = n23274 ^ n21734 ;
  assign n23276 = n21561 & n23275 ;
  assign n23294 = n23293 ^ n23276 ;
  assign n23295 = n21793 ^ n21744 ;
  assign n23296 = n23295 ^ n21794 ;
  assign n23297 = n23296 ^ n23295 ;
  assign n23298 = n23295 ^ n21552 ;
  assign n23299 = n23298 ^ n23295 ;
  assign n23300 = n23297 & n23299 ;
  assign n23301 = n23300 ^ n23295 ;
  assign n23302 = ~n21561 & n23301 ;
  assign n23303 = n23302 ^ n21797 ;
  assign n23304 = ~n23294 & ~n23303 ;
  assign n23305 = n23269 & n23304 ;
  assign n23306 = n23305 ^ n21228 ;
  assign n23307 = n23306 ^ x67 ;
  assign n23308 = n23257 & ~n23307 ;
  assign n23311 = n23308 ^ n23257 ;
  assign n23314 = n23311 ^ n23307 ;
  assign n23217 = n22714 ^ n20690 ;
  assign n23204 = ~n22081 & n22203 ;
  assign n23187 = n22235 ^ n22211 ;
  assign n23185 = n22205 ^ n22194 ;
  assign n23184 = n22688 ^ n22225 ;
  assign n23186 = n23185 ^ n23184 ;
  assign n23188 = n23187 ^ n23186 ;
  assign n23189 = n22080 & ~n23188 ;
  assign n23190 = n23189 ^ n23187 ;
  assign n23199 = n23190 ^ n22262 ;
  assign n23200 = n23199 ^ n22272 ;
  assign n23201 = n23200 ^ n22709 ;
  assign n23202 = n23201 ^ n22711 ;
  assign n23192 = n23190 ^ n22185 ;
  assign n23191 = n23190 ^ n22234 ;
  assign n23193 = n23192 ^ n23191 ;
  assign n23196 = ~n22080 & n23193 ;
  assign n23197 = n23196 ^ n23192 ;
  assign n23198 = n22079 & n23197 ;
  assign n23203 = n23202 ^ n23198 ;
  assign n23205 = n23204 ^ n23203 ;
  assign n23206 = n22079 & ~n22696 ;
  assign n23207 = n23206 ^ n22192 ;
  assign n23208 = n23207 ^ n23187 ;
  assign n23209 = n23208 ^ n23207 ;
  assign n23212 = n22079 & n23209 ;
  assign n23213 = n23212 ^ n23207 ;
  assign n23214 = ~n22081 & n23213 ;
  assign n23215 = n23214 ^ n23207 ;
  assign n23216 = ~n23205 & ~n23215 ;
  assign n23218 = n23217 ^ n23216 ;
  assign n23219 = n23218 ^ x86 ;
  assign n23220 = n22569 ^ n22567 ;
  assign n23221 = n23220 ^ n21232 ;
  assign n23222 = n23221 ^ x109 ;
  assign n23223 = ~n23219 & ~n23222 ;
  assign n23224 = n23223 ^ n23222 ;
  assign n23319 = n23224 ^ n23219 ;
  assign n23324 = n23314 & ~n23319 ;
  assign n23309 = n23308 ^ n23307 ;
  assign n23320 = ~n23309 & ~n23319 ;
  assign n23316 = n23223 & n23308 ;
  assign n23315 = n23223 & n23314 ;
  assign n23317 = n23316 ^ n23315 ;
  assign n23312 = n23223 & n23311 ;
  assign n23313 = n23312 ^ n23223 ;
  assign n23318 = n23317 ^ n23313 ;
  assign n23321 = n23320 ^ n23318 ;
  assign n23322 = n23321 ^ n23309 ;
  assign n23310 = ~n23224 & ~n23309 ;
  assign n23323 = n23322 ^ n23310 ;
  assign n23325 = n23324 ^ n23323 ;
  assign n23326 = n23325 ^ n23318 ;
  assign n23327 = ~n23183 & ~n23326 ;
  assign n23334 = n23311 & ~n23319 ;
  assign n23346 = n23334 ^ n23316 ;
  assign n23339 = n23319 ^ n23222 ;
  assign n23340 = n23308 & ~n23339 ;
  assign n23347 = n23346 ^ n23340 ;
  assign n23336 = n23324 ^ n23320 ;
  assign n23335 = n23334 ^ n23319 ;
  assign n23337 = n23336 ^ n23335 ;
  assign n23348 = n23347 ^ n23337 ;
  assign n23345 = n23334 ^ n23308 ;
  assign n23349 = n23348 ^ n23345 ;
  assign n23350 = n23349 ^ n23346 ;
  assign n23351 = n23350 ^ n23312 ;
  assign n23343 = n23311 & ~n23339 ;
  assign n23344 = n23343 ^ n23337 ;
  assign n23352 = n23351 ^ n23344 ;
  assign n23342 = n23340 ^ n23257 ;
  assign n23353 = n23352 ^ n23342 ;
  assign n23375 = n23353 ^ n23321 ;
  assign n23376 = n23375 ^ n23340 ;
  assign n23377 = n23376 ^ n23181 ;
  assign n23378 = n23377 ^ n23151 ;
  assign n23354 = n23349 ^ n23343 ;
  assign n23379 = n23354 ^ n23182 ;
  assign n23380 = n23354 ^ n23151 ;
  assign n23381 = n23380 ^ n23181 ;
  assign n23382 = n23381 ^ n23354 ;
  assign n23383 = ~n23379 & n23382 ;
  assign n23384 = n23383 ^ n23354 ;
  assign n23385 = ~n23378 & n23384 ;
  assign n23386 = n23385 ^ n23181 ;
  assign n23330 = ~n23224 & n23314 ;
  assign n23368 = n23344 ^ n23330 ;
  assign n23366 = n23315 ^ n23314 ;
  assign n23367 = n23366 ^ n23330 ;
  assign n23369 = n23368 ^ n23367 ;
  assign n23370 = n23368 ^ n23180 ;
  assign n23371 = n23370 ^ n23368 ;
  assign n23372 = ~n23369 & ~n23371 ;
  assign n23373 = n23372 ^ n23368 ;
  assign n23374 = n23151 & n23373 ;
  assign n23387 = n23386 ^ n23374 ;
  assign n23358 = n23334 ^ n23312 ;
  assign n23388 = n23387 ^ n23358 ;
  assign n23355 = n23354 ^ n23353 ;
  assign n23331 = n23330 ^ n23324 ;
  assign n23332 = n23331 ^ n23318 ;
  assign n23328 = n23307 ^ n23257 ;
  assign n23329 = n23328 ^ n23219 ;
  assign n23333 = n23332 ^ n23329 ;
  assign n23338 = n23337 ^ n23333 ;
  assign n23341 = n23340 ^ n23338 ;
  assign n23356 = n23355 ^ n23341 ;
  assign n23357 = n23356 ^ n23329 ;
  assign n23359 = n23358 ^ n23357 ;
  assign n23360 = n23359 ^ n23358 ;
  assign n23361 = n23358 ^ n23180 ;
  assign n23362 = n23361 ^ n23358 ;
  assign n23363 = ~n23360 & ~n23362 ;
  assign n23364 = n23363 ^ n23358 ;
  assign n23365 = ~n23151 & n23364 ;
  assign n23389 = n23388 ^ n23365 ;
  assign n23390 = n23181 ^ n23151 ;
  assign n23391 = n23366 ^ n23324 ;
  assign n23392 = ~n23390 & n23391 ;
  assign n23393 = n23389 & ~n23392 ;
  assign n23394 = ~n23327 & n23393 ;
  assign n23395 = n23394 ^ n21661 ;
  assign n23421 = n23141 ^ n22766 ;
  assign n23397 = n22805 ^ n22791 ;
  assign n23422 = n23421 ^ n23397 ;
  assign n23423 = ~n23139 & n23422 ;
  assign n23416 = n23397 ^ n23143 ;
  assign n23408 = n22779 ^ n22773 ;
  assign n23409 = n23140 ^ n22783 ;
  assign n23412 = n22773 & ~n23409 ;
  assign n23413 = n23412 ^ n22783 ;
  assign n23414 = n23408 & ~n23413 ;
  assign n23415 = n23414 ^ n22779 ;
  assign n23417 = n23416 ^ n23415 ;
  assign n23418 = n23417 ^ n19450 ;
  assign n23399 = n22777 ^ n22758 ;
  assign n23400 = n23399 ^ n22728 ;
  assign n23398 = n23397 ^ n22786 ;
  assign n23401 = n23400 ^ n23398 ;
  assign n23402 = n23401 ^ n23397 ;
  assign n23403 = n23397 ^ n22776 ;
  assign n23404 = n23403 ^ n23397 ;
  assign n23405 = ~n23402 & n23404 ;
  assign n23406 = n23405 ^ n23397 ;
  assign n23407 = ~n23116 & ~n23406 ;
  assign n23419 = n23418 ^ n23407 ;
  assign n23396 = n22779 & n22819 ;
  assign n23420 = n23419 ^ n23396 ;
  assign n23424 = n23423 ^ n23420 ;
  assign n23426 = ~n23183 & n23310 ;
  assign n23440 = n23366 ^ n23331 ;
  assign n23441 = ~n23180 & n23440 ;
  assign n23445 = n23441 ^ n23180 ;
  assign n23439 = n23330 ^ n23325 ;
  assign n23442 = n23441 ^ n23439 ;
  assign n23437 = n23324 ^ n23317 ;
  assign n23438 = n23180 & ~n23437 ;
  assign n23443 = n23442 ^ n23438 ;
  assign n23444 = n23151 & ~n23443 ;
  assign n23446 = n23445 ^ n23444 ;
  assign n23430 = n23390 ^ n23340 ;
  assign n23431 = n23332 ^ n23182 ;
  assign n23434 = n23390 & n23431 ;
  assign n23435 = n23434 ^ n23332 ;
  assign n23436 = ~n23430 & ~n23435 ;
  assign n23447 = n23446 ^ n23436 ;
  assign n23448 = n23447 ^ n23344 ;
  assign n23429 = n23181 & n23310 ;
  assign n23449 = n23448 ^ n23429 ;
  assign n23427 = n23180 ^ n23151 ;
  assign n23428 = n23352 & n23427 ;
  assign n23450 = n23449 ^ n23428 ;
  assign n23451 = ~n23426 & n23450 ;
  assign n23425 = n23181 & n23375 ;
  assign n23452 = n23451 ^ n23425 ;
  assign n23453 = n23353 ^ n23315 ;
  assign n23454 = n23353 ^ n23180 ;
  assign n23455 = n23454 ^ n23353 ;
  assign n23456 = n23453 & ~n23455 ;
  assign n23457 = n23456 ^ n23353 ;
  assign n23458 = ~n23427 & n23457 ;
  assign n23459 = n23452 & ~n23458 ;
  assign n23460 = n23459 ^ n22175 ;
  assign n23494 = n21794 ^ n21726 ;
  assign n23495 = n21710 & n23494 ;
  assign n23477 = n21750 ^ n21747 ;
  assign n23478 = n23477 ^ n21754 ;
  assign n23479 = n23478 ^ n21745 ;
  assign n23480 = n21552 & ~n23479 ;
  assign n23481 = n23480 ^ n21745 ;
  assign n23491 = n23481 ^ n20276 ;
  assign n23492 = n23491 ^ n21781 ;
  assign n23475 = n21561 ^ n21552 ;
  assign n23482 = n21732 ^ n21717 ;
  assign n23483 = n23482 ^ n21697 ;
  assign n23484 = n23483 ^ n23481 ;
  assign n23476 = n21753 ^ n21745 ;
  assign n23485 = n23484 ^ n23476 ;
  assign n23486 = n23484 ^ n21552 ;
  assign n23487 = n23486 ^ n23484 ;
  assign n23488 = n23485 & ~n23487 ;
  assign n23489 = n23488 ^ n23484 ;
  assign n23490 = ~n23475 & ~n23489 ;
  assign n23493 = n23492 ^ n23490 ;
  assign n23496 = n23495 ^ n23493 ;
  assign n23467 = n21746 ^ n21744 ;
  assign n23468 = n23467 ^ n21725 ;
  assign n23469 = n23468 ^ n21746 ;
  assign n23470 = n21746 ^ n21552 ;
  assign n23471 = n23470 ^ n21746 ;
  assign n23472 = n23469 & n23471 ;
  assign n23473 = n23472 ^ n21746 ;
  assign n23474 = ~n21561 & ~n23473 ;
  assign n23497 = n23496 ^ n23474 ;
  assign n23461 = n21752 ^ n21742 ;
  assign n23462 = n21752 ^ n21561 ;
  assign n23463 = n23462 ^ n21752 ;
  assign n23464 = n23461 & ~n23463 ;
  assign n23465 = n23464 ^ n21752 ;
  assign n23466 = ~n21552 & n23465 ;
  assign n23498 = n23497 ^ n23466 ;
  assign n23516 = n23179 ^ x85 ;
  assign n23517 = ~n22430 & ~n22915 ;
  assign n23540 = n22382 ^ n22375 ;
  assign n23539 = n22391 ^ n22377 ;
  assign n23541 = n23540 ^ n23539 ;
  assign n23542 = ~n22278 & ~n23541 ;
  assign n23524 = n22906 ^ n22892 ;
  assign n23525 = n23524 ^ n22381 ;
  assign n23526 = n22395 ^ n22382 ;
  assign n23527 = n23526 ^ n23524 ;
  assign n23528 = n23527 ^ n23526 ;
  assign n23529 = n23526 ^ n22278 ;
  assign n23530 = n23529 ^ n23526 ;
  assign n23531 = n23528 & n23530 ;
  assign n23532 = n23531 ^ n23526 ;
  assign n23533 = n22277 & n23532 ;
  assign n23534 = n22278 & n23533 ;
  assign n23535 = ~n23525 & n23534 ;
  assign n23538 = n23535 ^ n23533 ;
  assign n23543 = n23542 ^ n23538 ;
  assign n23536 = n22906 ^ n22386 ;
  assign n23537 = n23536 ^ n23535 ;
  assign n23544 = n23543 ^ n23537 ;
  assign n23545 = n23544 ^ n23533 ;
  assign n23546 = n22279 & n23545 ;
  assign n23547 = n23546 ^ n23543 ;
  assign n23550 = n23547 ^ n22440 ;
  assign n23518 = n22432 ^ n22375 ;
  assign n23519 = n23518 ^ n22379 ;
  assign n23520 = n22379 ^ n22277 ;
  assign n23521 = n23520 ^ n22379 ;
  assign n23522 = n23519 & n23521 ;
  assign n23523 = n23522 ^ n22379 ;
  assign n23548 = n22278 & ~n23547 ;
  assign n23549 = n23523 & n23548 ;
  assign n23551 = n23550 ^ n23549 ;
  assign n23552 = n23517 & ~n23551 ;
  assign n23553 = n23552 ^ n20820 ;
  assign n23554 = n23553 ^ x70 ;
  assign n23555 = n23516 & ~n23554 ;
  assign n23556 = n23555 ^ n23516 ;
  assign n23557 = n23150 ^ x126 ;
  assign n23571 = n21189 ^ n21186 ;
  assign n23572 = n21458 ^ n21456 ;
  assign n23573 = ~n23571 & n23572 ;
  assign n23574 = n23573 ^ n21459 ;
  assign n23564 = n23049 ^ n21480 ;
  assign n23565 = n21144 & ~n23564 ;
  assign n23566 = n23565 ^ n21480 ;
  assign n23575 = n23574 ^ n23566 ;
  assign n23570 = n21187 & n21448 ;
  assign n23576 = n23575 ^ n23570 ;
  assign n23567 = n23566 ^ n21468 ;
  assign n23561 = n21490 ^ n21464 ;
  assign n23562 = n23561 ^ n21461 ;
  assign n23563 = ~n21144 & n23562 ;
  assign n23568 = n23567 ^ n23563 ;
  assign n23569 = ~n21460 & n23568 ;
  assign n23577 = n23576 ^ n23569 ;
  assign n23559 = n21461 ^ n21453 ;
  assign n23560 = n21187 & n23559 ;
  assign n23578 = n23577 ^ n23560 ;
  assign n23558 = n21188 & ~n21503 ;
  assign n23579 = n23578 ^ n23558 ;
  assign n23580 = n21456 ^ n21439 ;
  assign n23581 = n23580 ^ n21513 ;
  assign n23582 = n21144 & n23581 ;
  assign n23583 = n23582 ^ n21513 ;
  assign n23584 = ~n21186 & n23583 ;
  assign n23585 = ~n23579 & n23584 ;
  assign n23586 = n23585 ^ n23579 ;
  assign n23587 = ~n23052 & ~n23586 ;
  assign n23588 = n23587 ^ n20784 ;
  assign n23589 = n23588 ^ x84 ;
  assign n23590 = n23557 & ~n23589 ;
  assign n23596 = n23556 & n23590 ;
  assign n23591 = n23590 ^ n23557 ;
  assign n23594 = n23591 ^ n23589 ;
  assign n23660 = n23596 ^ n23594 ;
  assign n23499 = n22947 ^ n22519 ;
  assign n23503 = n23499 ^ n22549 ;
  assign n23500 = n23499 ^ n22559 ;
  assign n23504 = n23503 ^ n23500 ;
  assign n23505 = ~n22446 & ~n23504 ;
  assign n23506 = n23505 ^ n23500 ;
  assign n23507 = ~n22447 & n23506 ;
  assign n23508 = n23507 ^ n23499 ;
  assign n23509 = n22937 & n23508 ;
  assign n23510 = n23509 ^ n20499 ;
  assign n23511 = n23510 ^ x102 ;
  assign n23512 = n23218 ^ x116 ;
  assign n23513 = n23511 & ~n23512 ;
  assign n23665 = ~n23513 & n23554 ;
  assign n23514 = n23513 ^ n23512 ;
  assign n23515 = n23514 ^ n23511 ;
  assign n23666 = n23665 ^ n23515 ;
  assign n23667 = n23516 & n23666 ;
  assign n23668 = n23660 & ~n23667 ;
  assign n23632 = n23515 ^ n23512 ;
  assign n23599 = n23555 ^ n23554 ;
  assign n23600 = n23590 & ~n23599 ;
  assign n23595 = n23556 & n23594 ;
  assign n23597 = n23596 ^ n23595 ;
  assign n23592 = n23556 & n23591 ;
  assign n23593 = n23592 ^ n23556 ;
  assign n23598 = n23597 ^ n23593 ;
  assign n23601 = n23600 ^ n23598 ;
  assign n23648 = n23601 ^ n23596 ;
  assign n23615 = n23555 & n23594 ;
  assign n23610 = n23555 & n23590 ;
  assign n23616 = n23615 ^ n23610 ;
  assign n23649 = n23648 ^ n23616 ;
  assign n23602 = n23556 ^ n23554 ;
  assign n23605 = ~n23589 & n23602 ;
  assign n23650 = n23649 ^ n23605 ;
  assign n23646 = n23615 ^ n23590 ;
  assign n23647 = n23646 ^ n23598 ;
  assign n23651 = n23650 ^ n23647 ;
  assign n23652 = n23651 ^ n23602 ;
  assign n23606 = n23594 & n23602 ;
  assign n23607 = n23606 ^ n23602 ;
  assign n23608 = n23607 ^ n23605 ;
  assign n23653 = n23652 ^ n23608 ;
  assign n23654 = n23632 & n23653 ;
  assign n23612 = n23594 ^ n23557 ;
  assign n23613 = n23555 & ~n23612 ;
  assign n23614 = n23613 ^ n23555 ;
  assign n23617 = n23616 ^ n23614 ;
  assign n23643 = ~n23514 & n23617 ;
  assign n23642 = n23613 & n23632 ;
  assign n23644 = n23643 ^ n23642 ;
  assign n23637 = n23594 & ~n23599 ;
  assign n23636 = n23591 & ~n23599 ;
  assign n23638 = n23637 ^ n23636 ;
  assign n23633 = n23605 ^ n23599 ;
  assign n23634 = n23633 ^ n23600 ;
  assign n23635 = ~n23632 & ~n23634 ;
  assign n23639 = n23638 ^ n23635 ;
  assign n23624 = n23616 ^ n23511 ;
  assign n23625 = n23624 ^ n23616 ;
  assign n23626 = n23616 ^ n23592 ;
  assign n23627 = n23626 ^ n23616 ;
  assign n23628 = ~n23625 & n23627 ;
  assign n23629 = n23628 ^ n23616 ;
  assign n23630 = n23512 & n23629 ;
  assign n23631 = n23630 ^ n23616 ;
  assign n23640 = n23639 ^ n23631 ;
  assign n23611 = n23610 ^ n23598 ;
  assign n23618 = n23617 ^ n23611 ;
  assign n23619 = n23617 ^ n23512 ;
  assign n23620 = n23619 ^ n23617 ;
  assign n23621 = n23618 & n23620 ;
  assign n23622 = n23621 ^ n23617 ;
  assign n23623 = n23511 & n23622 ;
  assign n23641 = n23640 ^ n23623 ;
  assign n23645 = n23644 ^ n23641 ;
  assign n23655 = n23654 ^ n23645 ;
  assign n23656 = n23655 ^ n22508 ;
  assign n23657 = n23656 ^ n23594 ;
  assign n23609 = ~n23512 & n23608 ;
  assign n23658 = n23657 ^ n23609 ;
  assign n23603 = n23602 ^ n23601 ;
  assign n23604 = n23515 & n23603 ;
  assign n23659 = n23658 ^ n23604 ;
  assign n23669 = n23668 ^ n23659 ;
  assign n23697 = n22917 ^ n22430 ;
  assign n23683 = ~n22386 & n22924 ;
  assign n23684 = n23683 ^ n22436 ;
  assign n23685 = ~n22429 & ~n23684 ;
  assign n23686 = n23536 ^ n22366 ;
  assign n23687 = n23686 ^ n22370 ;
  assign n23688 = n23685 & ~n23687 ;
  assign n23689 = n23688 ^ n23684 ;
  assign n23698 = n23697 ^ n23689 ;
  assign n23690 = n23689 ^ n22904 ;
  assign n23691 = n23690 ^ n22370 ;
  assign n23692 = n23691 ^ n23518 ;
  assign n23693 = n23692 ^ n23689 ;
  assign n23694 = n22278 & n23693 ;
  assign n23695 = n23694 ^ n23690 ;
  assign n23696 = ~n22277 & ~n23695 ;
  assign n23699 = n23698 ^ n23696 ;
  assign n23682 = n22279 & ~n23539 ;
  assign n23700 = n23699 ^ n23682 ;
  assign n23677 = n22381 ^ n22277 ;
  assign n23678 = n23677 ^ n22381 ;
  assign n23679 = n22389 & n23678 ;
  assign n23680 = n23679 ^ n22381 ;
  assign n23681 = n22278 & n23680 ;
  assign n23701 = n23700 ^ n23681 ;
  assign n23670 = n22892 ^ n22278 ;
  assign n23671 = n23670 ^ n22892 ;
  assign n23674 = n22367 & ~n23671 ;
  assign n23675 = n23674 ^ n22892 ;
  assign n23676 = n22277 & n23675 ;
  assign n23702 = n23701 ^ n23676 ;
  assign n23703 = ~n22915 & n23702 ;
  assign n23704 = n23703 ^ n20082 ;
  assign n23705 = n23150 ^ x81 ;
  assign n23733 = n21731 ^ n19783 ;
  assign n23734 = n23733 ^ n21788 ;
  assign n23729 = n23268 ^ n21770 ;
  assign n23716 = n21747 ^ n21729 ;
  assign n23714 = n21743 ^ n21697 ;
  assign n23706 = n21727 ^ n21723 ;
  assign n23707 = n23706 ^ n23482 ;
  assign n23708 = n23707 ^ n21727 ;
  assign n23709 = n21727 ^ n21561 ;
  assign n23710 = n23709 ^ n21727 ;
  assign n23711 = n23708 & ~n23710 ;
  assign n23712 = n23711 ^ n21727 ;
  assign n23713 = n21552 & n23712 ;
  assign n23715 = n23714 ^ n23713 ;
  assign n23717 = n23716 ^ n23715 ;
  assign n23718 = n23717 ^ n23713 ;
  assign n23719 = n21552 & n23718 ;
  assign n23720 = n23719 ^ n23715 ;
  assign n23730 = n23729 ^ n23720 ;
  assign n23721 = n23720 ^ n23713 ;
  assign n23722 = n23721 ^ n23285 ;
  assign n23723 = n23722 ^ n23721 ;
  assign n23726 = ~n21552 & ~n23723 ;
  assign n23727 = n23726 ^ n23721 ;
  assign n23728 = n23475 & n23727 ;
  assign n23731 = n23730 ^ n23728 ;
  assign n23732 = ~n21709 & ~n23731 ;
  assign n23735 = n23734 ^ n23732 ;
  assign n23736 = n23735 ^ x88 ;
  assign n23844 = n23705 & ~n23736 ;
  assign n23792 = n23510 ^ x122 ;
  assign n23809 = n22020 ^ n21989 ;
  assign n23805 = n21989 ^ n21917 ;
  assign n23806 = n23805 ^ n22008 ;
  assign n23807 = n23806 ^ n22005 ;
  assign n23808 = n21970 & ~n23807 ;
  assign n23810 = n23809 ^ n23808 ;
  assign n23811 = n21988 & n23810 ;
  assign n23800 = ~n21829 & ~n21880 ;
  assign n23801 = ~n21970 & n23800 ;
  assign n23795 = n22862 ^ n22015 ;
  assign n23796 = n23795 ^ n23155 ;
  assign n23797 = n21970 & n23796 ;
  assign n23798 = n23797 ^ n22862 ;
  assign n23799 = n23798 ^ n21995 ;
  assign n23802 = n23801 ^ n23799 ;
  assign n23803 = ~n21918 & n23802 ;
  assign n23804 = n23803 ^ n23798 ;
  assign n23812 = n23811 ^ n23804 ;
  assign n23813 = n23812 ^ n21973 ;
  assign n23814 = n23813 ^ n22883 ;
  assign n23793 = n23155 ^ n21974 ;
  assign n23794 = ~n21986 & n23793 ;
  assign n23815 = n23814 ^ n23794 ;
  assign n23816 = ~n22012 & ~n23815 ;
  assign n23817 = n21970 ^ n21918 ;
  assign n23818 = n21993 ^ n21992 ;
  assign n23819 = n21992 ^ n21970 ;
  assign n23820 = n23819 ^ n21992 ;
  assign n23821 = n23818 & n23820 ;
  assign n23822 = n23821 ^ n21992 ;
  assign n23823 = ~n23817 & n23822 ;
  assign n23824 = n23823 ^ n21992 ;
  assign n23825 = n23816 & ~n23824 ;
  assign n23826 = ~n22881 & n23825 ;
  assign n23827 = ~n22040 & n23826 ;
  assign n23828 = n23827 ^ n19403 ;
  assign n23829 = n23828 ^ x120 ;
  assign n23830 = n23792 & ~n23829 ;
  assign n23831 = n23830 ^ n23792 ;
  assign n23752 = n22245 ^ n22217 ;
  assign n23753 = n23752 ^ n23215 ;
  assign n23745 = n23185 ^ n22209 ;
  assign n23746 = n23745 ^ n22236 ;
  assign n23747 = n22236 ^ n22080 ;
  assign n23748 = n23747 ^ n22236 ;
  assign n23749 = n23746 & ~n23748 ;
  assign n23750 = n23749 ^ n22236 ;
  assign n23751 = ~n22079 & n23750 ;
  assign n23754 = n23753 ^ n23751 ;
  assign n23755 = n23754 ^ n22714 ;
  assign n23756 = n23755 ^ n22200 ;
  assign n23757 = n23756 ^ n20458 ;
  assign n23743 = n22208 ^ n22187 ;
  assign n23744 = ~n22081 & n23743 ;
  assign n23758 = n23757 ^ n23744 ;
  assign n23738 = n22203 ^ n22181 ;
  assign n23739 = n23738 ^ n23187 ;
  assign n23740 = n22079 & n23739 ;
  assign n23741 = n23740 ^ n22245 ;
  assign n23742 = ~n22080 & n23741 ;
  assign n23759 = n23758 ^ n23742 ;
  assign n23760 = n23759 ^ x105 ;
  assign n23788 = n20970 ^ n20482 ;
  assign n23761 = n20917 ^ n19349 ;
  assign n23777 = n20925 ^ n20650 ;
  assign n23774 = n20660 ^ n20626 ;
  assign n23775 = n23774 ^ n20656 ;
  assign n23776 = n23775 ^ n20946 ;
  assign n23778 = n23777 ^ n23776 ;
  assign n23779 = n23776 ^ n20917 ;
  assign n23780 = n23779 ^ n23776 ;
  assign n23781 = ~n23778 & ~n23780 ;
  assign n23782 = n23781 ^ n23776 ;
  assign n23783 = ~n23761 & n23782 ;
  assign n23767 = n20934 ^ n20637 ;
  assign n23768 = n23767 ^ n20634 ;
  assign n23771 = n20917 & ~n23768 ;
  assign n23772 = n23771 ^ n20634 ;
  assign n23773 = ~n19349 & n23772 ;
  assign n23784 = n23783 ^ n23773 ;
  assign n23763 = n20943 ^ n20653 ;
  assign n23764 = n23763 ^ n20649 ;
  assign n23765 = n20928 & ~n23764 ;
  assign n23785 = n23784 ^ n23765 ;
  assign n23762 = ~n23230 & n23761 ;
  assign n23786 = n23785 ^ n23762 ;
  assign n23787 = ~n23225 & ~n23786 ;
  assign n23789 = n23788 ^ n23787 ;
  assign n23790 = n23789 ^ x66 ;
  assign n23791 = ~n23760 & n23790 ;
  assign n23835 = n23791 ^ n23790 ;
  assign n23845 = n23835 ^ n23760 ;
  assign n23862 = n23845 ^ n23790 ;
  assign n23864 = n23831 & ~n23862 ;
  assign n23913 = n23844 & n23864 ;
  assign n23832 = n23831 ^ n23829 ;
  assign n23846 = n23832 ^ n23792 ;
  assign n23847 = n23845 & ~n23846 ;
  assign n23836 = n23830 & n23835 ;
  assign n23834 = n23791 & n23831 ;
  assign n23837 = n23836 ^ n23834 ;
  assign n23906 = n23847 ^ n23837 ;
  assign n23907 = ~n23736 & n23906 ;
  assign n23854 = n23836 ^ n23835 ;
  assign n23852 = n23835 & ~n23846 ;
  assign n23851 = n23831 & n23835 ;
  assign n23853 = n23852 ^ n23851 ;
  assign n23855 = n23854 ^ n23853 ;
  assign n23833 = n23791 & n23832 ;
  assign n23856 = n23855 ^ n23833 ;
  assign n23848 = ~n23792 & n23845 ;
  assign n23849 = n23848 ^ n23847 ;
  assign n23850 = n23849 ^ n23832 ;
  assign n23857 = n23856 ^ n23850 ;
  assign n23866 = n23862 ^ n23857 ;
  assign n23863 = n23830 & ~n23862 ;
  assign n23865 = n23864 ^ n23863 ;
  assign n23867 = n23866 ^ n23865 ;
  assign n23858 = n23857 ^ n23852 ;
  assign n23859 = n23844 & n23858 ;
  assign n23860 = n23859 ^ n23855 ;
  assign n23861 = n23860 ^ n23848 ;
  assign n23868 = n23867 ^ n23861 ;
  assign n23869 = n23868 ^ n23867 ;
  assign n23870 = n23858 ^ n23849 ;
  assign n23871 = n23844 ^ n23705 ;
  assign n23872 = ~n23870 & ~n23871 ;
  assign n23873 = n23869 & n23872 ;
  assign n23874 = n23873 ^ n23868 ;
  assign n23908 = n23907 ^ n23874 ;
  assign n23910 = n23908 ^ n23855 ;
  assign n23911 = ~n23705 & ~n23910 ;
  assign n23893 = n23791 & ~n23846 ;
  assign n23875 = n23830 & n23845 ;
  assign n23876 = n23875 ^ n23834 ;
  assign n23901 = n23893 ^ n23876 ;
  assign n23902 = n23844 & n23901 ;
  assign n23894 = n23893 ^ n23865 ;
  assign n23895 = n23894 ^ n23865 ;
  assign n23896 = n23865 ^ n23736 ;
  assign n23897 = n23896 ^ n23865 ;
  assign n23898 = n23895 & ~n23897 ;
  assign n23899 = n23898 ^ n23865 ;
  assign n23900 = ~n23705 & n23899 ;
  assign n23903 = n23902 ^ n23900 ;
  assign n23877 = n23876 ^ n23863 ;
  assign n23878 = n23877 ^ n23830 ;
  assign n23879 = n23878 ^ n23837 ;
  assign n23880 = n23879 ^ n23736 ;
  assign n23881 = n23875 ^ n23845 ;
  assign n23882 = n23881 ^ n23848 ;
  assign n23887 = n23882 ^ n23879 ;
  assign n23884 = n23849 ^ n23833 ;
  assign n23883 = n23882 ^ n23853 ;
  assign n23885 = n23884 ^ n23883 ;
  assign n23886 = ~n23705 & n23885 ;
  assign n23888 = n23887 ^ n23886 ;
  assign n23889 = n23880 & ~n23888 ;
  assign n23890 = n23889 ^ n23736 ;
  assign n23891 = n23890 ^ n23874 ;
  assign n23737 = n23736 ^ n23705 ;
  assign n23838 = n23837 ^ n23833 ;
  assign n23839 = n23837 ^ n23705 ;
  assign n23840 = n23839 ^ n23837 ;
  assign n23841 = n23838 & ~n23840 ;
  assign n23842 = n23841 ^ n23837 ;
  assign n23843 = ~n23737 & n23842 ;
  assign n23892 = n23891 ^ n23843 ;
  assign n23904 = n23903 ^ n23892 ;
  assign n23905 = n23904 ^ n21828 ;
  assign n23912 = n23911 ^ n23905 ;
  assign n23914 = n23913 ^ n23912 ;
  assign n23952 = n23882 ^ n23836 ;
  assign n23953 = n23844 & n23952 ;
  assign n23954 = n23953 ^ n23903 ;
  assign n23955 = n23954 ^ n21694 ;
  assign n23915 = n23879 ^ n23851 ;
  assign n23916 = n23915 ^ n23884 ;
  assign n23917 = n23884 ^ n23705 ;
  assign n23918 = n23917 ^ n23884 ;
  assign n23919 = n23916 & ~n23918 ;
  assign n23920 = n23919 ^ n23884 ;
  assign n23921 = ~n23737 & n23920 ;
  assign n23934 = n23855 ^ n23705 ;
  assign n23935 = n23934 ^ n23855 ;
  assign n23938 = n23856 & n23935 ;
  assign n23939 = n23938 ^ n23855 ;
  assign n23940 = n23737 & n23939 ;
  assign n23927 = n23857 ^ n23847 ;
  assign n23928 = n23927 ^ n23884 ;
  assign n23929 = n23705 & n23928 ;
  assign n23930 = n23929 ^ n23884 ;
  assign n23941 = n23940 ^ n23930 ;
  assign n23926 = n23901 ^ n23858 ;
  assign n23931 = n23930 ^ n23926 ;
  assign n23922 = n23867 ^ n23830 ;
  assign n23923 = n23922 ^ n23858 ;
  assign n23924 = n23923 ^ n23901 ;
  assign n23925 = n23705 & ~n23924 ;
  assign n23932 = n23931 ^ n23925 ;
  assign n23933 = n23736 & n23932 ;
  assign n23942 = n23941 ^ n23933 ;
  assign n23943 = n23852 ^ n23705 ;
  assign n23944 = n23943 ^ n23852 ;
  assign n23947 = n23853 & n23944 ;
  assign n23948 = n23947 ^ n23852 ;
  assign n23949 = ~n23737 & n23948 ;
  assign n23950 = ~n23942 & ~n23949 ;
  assign n23951 = ~n23921 & n23950 ;
  assign n23956 = n23955 ^ n23951 ;
  assign n23957 = ~n21457 & ~n23573 ;
  assign n23990 = n21188 & n21458 ;
  assign n23987 = ~n21186 & ~n21490 ;
  assign n23969 = n21467 ^ n21186 ;
  assign n23972 = n21144 & ~n21464 ;
  assign n23973 = n23972 ^ n21484 ;
  assign n23976 = n23969 ^ n21467 ;
  assign n23977 = ~n23973 & ~n23976 ;
  assign n23978 = n23977 ^ n21144 ;
  assign n23979 = ~n23969 & n23978 ;
  assign n23980 = n23979 ^ n21186 ;
  assign n23968 = n21443 & ~n23571 ;
  assign n23981 = n23980 ^ n23968 ;
  assign n23984 = n23981 ^ n23054 ;
  assign n23967 = n21479 ^ n21439 ;
  assign n23982 = ~n21460 & n23981 ;
  assign n23983 = n23967 & n23982 ;
  assign n23985 = n23984 ^ n23983 ;
  assign n23965 = n21463 ^ n21445 ;
  assign n23966 = n21188 & n23965 ;
  assign n23986 = n23985 ^ n23966 ;
  assign n23988 = n23987 ^ n23986 ;
  assign n23960 = n21447 ^ n21186 ;
  assign n23961 = n23960 ^ n21447 ;
  assign n23962 = ~n21478 & n23961 ;
  assign n23963 = n23962 ^ n21447 ;
  assign n23964 = n21460 & n23963 ;
  assign n23989 = n23988 ^ n23964 ;
  assign n23991 = n23990 ^ n23989 ;
  assign n23992 = ~n23570 & n23991 ;
  assign n23993 = n23957 & n23992 ;
  assign n23994 = n23993 ^ n19592 ;
  assign n24016 = n22997 ^ n22963 ;
  assign n24017 = n24016 ^ n23000 ;
  assign n24018 = n22720 & n24017 ;
  assign n24006 = n23010 ^ n23008 ;
  assign n23997 = n23013 ^ n22994 ;
  assign n23998 = n23997 ^ n23010 ;
  assign n24005 = n23998 ^ n22999 ;
  assign n24007 = n24006 ^ n24005 ;
  assign n24004 = n22984 ^ n22969 ;
  assign n24008 = n24007 ^ n24004 ;
  assign n24009 = ~n22720 & n24008 ;
  assign n24010 = n24009 ^ n24005 ;
  assign n24019 = n24018 ^ n24010 ;
  assign n24020 = n22972 & n24019 ;
  assign n23995 = n22979 ^ n22970 ;
  assign n23996 = n23995 ^ n23077 ;
  assign n23999 = n23998 ^ n23996 ;
  assign n24000 = ~n22984 & ~n23999 ;
  assign n24001 = n24000 ^ n22979 ;
  assign n24003 = n23098 ^ n22981 ;
  assign n24011 = n24010 ^ n24003 ;
  assign n24002 = n23098 ^ n22984 ;
  assign n24012 = n24011 ^ n24002 ;
  assign n24013 = n24012 ^ n24010 ;
  assign n24014 = n24001 & n24013 ;
  assign n24015 = n24014 ^ n24011 ;
  assign n24021 = n24020 ^ n24015 ;
  assign n24022 = n24021 ^ n23029 ;
  assign n24023 = n24022 ^ n23093 ;
  assign n24024 = ~n23038 & ~n24023 ;
  assign n24025 = ~n22992 & n24024 ;
  assign n24026 = n24025 ^ n22141 ;
  assign n24046 = ~n20647 & n20926 ;
  assign n24039 = n20656 ^ n20626 ;
  assign n24040 = ~n19349 & ~n24039 ;
  assign n24036 = n20931 ^ n20660 ;
  assign n24030 = n20925 ^ n20649 ;
  assign n24028 = n20943 ^ n20636 ;
  assign n24029 = n24028 ^ n23243 ;
  assign n24031 = n24030 ^ n24029 ;
  assign n24032 = ~n20917 & ~n24031 ;
  assign n24033 = n24032 ^ n24030 ;
  assign n24037 = n24036 ^ n24033 ;
  assign n24034 = n24033 ^ n23227 ;
  assign n24038 = n24037 ^ n24034 ;
  assign n24041 = n24040 ^ n24038 ;
  assign n24042 = ~n20643 & ~n24041 ;
  assign n24043 = n24042 ^ n24034 ;
  assign n24044 = n23761 & n24043 ;
  assign n24027 = n20969 ^ n20340 ;
  assign n24035 = n24034 ^ n24027 ;
  assign n24045 = n24044 ^ n24035 ;
  assign n24047 = n24046 ^ n24045 ;
  assign n24074 = n22629 ^ n22577 ;
  assign n24075 = n22625 & n24074 ;
  assign n24059 = n22681 ^ n22627 ;
  assign n24060 = n22644 ^ n22595 ;
  assign n24061 = n24060 ^ n22642 ;
  assign n24062 = ~n24059 & ~n24061 ;
  assign n24057 = n22644 ^ n22597 ;
  assign n24058 = n22628 & ~n24057 ;
  assign n24063 = n24062 ^ n24058 ;
  assign n24055 = n22652 ^ n22619 ;
  assign n24054 = n22613 ^ n22609 ;
  assign n24056 = n24055 ^ n24054 ;
  assign n24064 = n24063 ^ n24056 ;
  assign n24065 = n24064 ^ n24063 ;
  assign n24066 = n24065 ^ n22638 ;
  assign n24067 = n24066 ^ n24065 ;
  assign n24070 = n21525 & n24067 ;
  assign n24071 = n24070 ^ n24065 ;
  assign n24072 = ~n21802 & n24071 ;
  assign n24073 = n24072 ^ n24064 ;
  assign n24076 = n24075 ^ n24073 ;
  assign n24048 = n22617 ^ n22581 ;
  assign n24049 = n22581 ^ n21801 ;
  assign n24050 = n24049 ^ n22581 ;
  assign n24051 = n24048 & ~n24050 ;
  assign n24052 = n24051 ^ n22581 ;
  assign n24053 = ~n21525 & n24052 ;
  assign n24077 = n24076 ^ n24053 ;
  assign n24078 = ~n22588 & ~n24077 ;
  assign n24081 = n22632 ^ n21801 ;
  assign n24082 = n24081 ^ n22632 ;
  assign n24083 = n22633 & ~n24082 ;
  assign n24084 = n24083 ^ n22632 ;
  assign n24085 = ~n21525 & n24084 ;
  assign n24086 = n24078 & ~n24085 ;
  assign n24087 = n24086 ^ n22476 ;
  assign n24120 = n22769 & n22779 ;
  assign n24117 = n23400 ^ n22781 ;
  assign n24118 = ~n23139 & ~n24117 ;
  assign n24113 = n22839 ^ n22775 ;
  assign n24103 = n22788 ^ n22761 ;
  assign n24104 = n24103 ^ n22809 ;
  assign n24105 = n22809 ^ n22776 ;
  assign n24106 = ~n23116 & n24105 ;
  assign n24107 = n24106 ^ n22776 ;
  assign n24108 = n24104 & n24107 ;
  assign n24109 = n24108 ^ n22809 ;
  assign n24110 = n24109 ^ n22787 ;
  assign n24114 = n24113 ^ n24110 ;
  assign n24115 = n24114 ^ n23144 ;
  assign n24095 = n22758 ^ n22725 ;
  assign n24096 = n24095 ^ n22728 ;
  assign n24097 = n24096 ^ n22725 ;
  assign n24100 = ~n22777 & n24097 ;
  assign n24101 = n24100 ^ n22725 ;
  assign n24102 = n22776 & ~n24101 ;
  assign n24111 = n24110 ^ n24102 ;
  assign n24112 = ~n23116 & ~n24111 ;
  assign n24116 = n24115 ^ n24112 ;
  assign n24119 = n24118 ^ n24116 ;
  assign n24121 = n24120 ^ n24119 ;
  assign n24088 = n23140 ^ n22792 ;
  assign n24089 = n22790 ^ n22779 ;
  assign n24092 = n23140 & ~n24089 ;
  assign n24093 = n24092 ^ n22779 ;
  assign n24094 = n24088 & n24093 ;
  assign n24122 = n24121 ^ n24094 ;
  assign n24123 = ~n23138 & n24122 ;
  assign n24124 = ~n23415 & n24123 ;
  assign n24125 = n24124 ^ n20042 ;
  assign n24134 = n23355 ^ n23316 ;
  assign n24126 = n23307 ^ n23222 ;
  assign n24127 = n24126 ^ n23219 ;
  assign n24128 = n24127 ^ n23222 ;
  assign n24129 = n23328 ^ n23222 ;
  assign n24130 = n24129 ^ n23222 ;
  assign n24131 = n24128 & ~n24130 ;
  assign n24132 = n24131 ^ n23222 ;
  assign n24133 = n23151 & ~n24132 ;
  assign n24135 = n24134 ^ n24133 ;
  assign n24136 = ~n23180 & ~n24135 ;
  assign n24137 = n23440 ^ n23325 ;
  assign n24138 = ~n23183 & ~n24137 ;
  assign n24154 = n23336 & ~n23390 ;
  assign n24145 = n23337 ^ n23180 ;
  assign n24147 = n23340 ^ n23312 ;
  assign n24150 = n24147 ^ n23337 ;
  assign n24146 = n23349 ^ n23317 ;
  assign n24148 = n24147 ^ n24146 ;
  assign n24149 = ~n23151 & ~n24148 ;
  assign n24151 = n24150 ^ n24149 ;
  assign n24152 = ~n24145 & n24151 ;
  assign n24153 = n24152 ^ n23180 ;
  assign n24155 = n24154 ^ n24153 ;
  assign n24139 = n23348 ^ n23325 ;
  assign n24140 = n23348 ^ n23151 ;
  assign n24141 = n24140 ^ n23348 ;
  assign n24142 = n24139 & ~n24141 ;
  assign n24143 = n24142 ^ n23348 ;
  assign n24144 = ~n23180 & ~n24143 ;
  assign n24156 = n24155 ^ n24144 ;
  assign n24157 = ~n23429 & ~n24156 ;
  assign n24158 = ~n23458 & n24157 ;
  assign n24159 = ~n24138 & n24158 ;
  assign n24160 = ~n24136 & n24159 ;
  assign n24161 = ~n23426 & n24160 ;
  assign n24162 = ~n23392 & n24161 ;
  assign n24163 = n24162 ^ n21877 ;
  assign n24172 = n24004 ^ n22988 ;
  assign n24173 = n24172 ^ n22981 ;
  assign n24175 = ~n22995 & ~n24173 ;
  assign n24176 = n24175 ^ n22981 ;
  assign n24178 = n23074 ^ n22979 ;
  assign n24177 = n23074 ^ n22995 ;
  assign n24179 = n24178 ^ n24177 ;
  assign n24180 = n24176 & n24179 ;
  assign n24181 = n24180 ^ n24178 ;
  assign n24182 = n24181 ^ n23025 ;
  assign n24168 = n23074 ^ n22968 ;
  assign n24165 = n23010 ^ n22984 ;
  assign n24169 = n24168 ^ n24165 ;
  assign n24164 = n23998 ^ n22986 ;
  assign n24166 = n24165 ^ n24164 ;
  assign n24167 = ~n22720 & n24166 ;
  assign n24170 = n24169 ^ n24167 ;
  assign n24171 = ~n22978 & n24170 ;
  assign n24183 = n24182 ^ n24171 ;
  assign n24184 = n24183 ^ n23096 ;
  assign n24185 = n24184 ^ n23035 ;
  assign n24186 = n24185 ^ n23100 ;
  assign n24187 = n24186 ^ n22992 ;
  assign n24188 = ~n22970 & ~n24187 ;
  assign n24189 = n24188 ^ n21630 ;
  assign n24190 = n23617 & n23632 ;
  assign n24199 = n23651 ^ n23636 ;
  assign n24200 = n24199 ^ n23608 ;
  assign n24224 = n24200 ^ n23600 ;
  assign n24225 = ~n23514 & n24224 ;
  assign n24223 = ~n23612 & n23667 ;
  assign n24226 = n24225 ^ n24223 ;
  assign n24191 = n23512 ^ n23511 ;
  assign n24221 = n23596 & ~n24191 ;
  assign n24198 = n23638 ^ n23600 ;
  assign n24210 = n24198 ^ n23599 ;
  assign n24211 = n24210 ^ n23592 ;
  assign n24212 = n24211 ^ n23600 ;
  assign n24207 = n24200 ^ n23606 ;
  assign n24201 = n24200 ^ n24198 ;
  assign n24202 = n24198 ^ n23511 ;
  assign n24204 = ~n23512 & n24202 ;
  assign n24205 = n24204 ^ n23511 ;
  assign n24206 = n24201 & ~n24205 ;
  assign n24208 = n24207 ^ n24206 ;
  assign n24209 = n24208 ^ n23598 ;
  assign n24213 = n24212 ^ n24209 ;
  assign n24214 = n24213 ^ n24208 ;
  assign n24215 = n24208 ^ n23511 ;
  assign n24216 = n24215 ^ n24208 ;
  assign n24217 = ~n24214 & n24216 ;
  assign n24218 = n24217 ^ n24208 ;
  assign n24219 = ~n23512 & n24218 ;
  assign n24220 = n24219 ^ n24208 ;
  assign n24222 = n24221 ^ n24220 ;
  assign n24227 = n24226 ^ n24222 ;
  assign n24228 = n24227 ^ n23642 ;
  assign n24229 = n24228 ^ n23631 ;
  assign n24192 = n23653 ^ n23597 ;
  assign n24193 = n23597 ^ n23512 ;
  assign n24194 = n24193 ^ n23597 ;
  assign n24195 = n24192 & ~n24194 ;
  assign n24196 = n24195 ^ n23597 ;
  assign n24197 = n24191 & n24196 ;
  assign n24230 = n24229 ^ n24197 ;
  assign n24231 = ~n24190 & ~n24230 ;
  assign n24232 = n24231 ^ n22121 ;
  assign n24233 = n22934 ^ x113 ;
  assign n24234 = n23828 ^ x104 ;
  assign n24235 = n24233 & ~n24234 ;
  assign n24236 = n24235 ^ n24233 ;
  assign n24237 = n24236 ^ n24234 ;
  assign n24238 = n24237 ^ n24233 ;
  assign n24239 = n23424 ^ x80 ;
  assign n24240 = n20972 ^ x90 ;
  assign n24241 = ~n24239 & ~n24240 ;
  assign n24242 = n24241 ^ n24240 ;
  assign n24248 = n24242 ^ n24239 ;
  assign n24249 = n24248 ^ n24240 ;
  assign n24243 = n23735 ^ x99 ;
  assign n24244 = n23994 ^ x73 ;
  assign n24245 = n24243 & ~n24244 ;
  assign n24252 = n24245 ^ n24244 ;
  assign n24263 = ~n24249 & ~n24252 ;
  assign n24253 = n24252 ^ n24243 ;
  assign n24254 = ~n24242 & n24253 ;
  assign n24267 = n24263 ^ n24254 ;
  assign n24266 = n24241 & n24253 ;
  assign n24268 = n24267 ^ n24266 ;
  assign n24265 = ~n24249 & n24253 ;
  assign n24269 = n24268 ^ n24265 ;
  assign n24264 = n24263 ^ n24253 ;
  assign n24270 = n24269 ^ n24264 ;
  assign n24271 = n24270 ^ n24248 ;
  assign n24261 = ~n24248 & ~n24252 ;
  assign n24260 = n24245 & ~n24248 ;
  assign n24262 = n24261 ^ n24260 ;
  assign n24272 = n24271 ^ n24262 ;
  assign n24257 = n24239 & n24243 ;
  assign n24250 = n24245 & ~n24249 ;
  assign n24246 = n24245 ^ n24243 ;
  assign n24247 = ~n24242 & n24246 ;
  assign n24251 = n24250 ^ n24247 ;
  assign n24258 = n24257 ^ n24251 ;
  assign n24259 = n24258 ^ n24245 ;
  assign n24273 = n24272 ^ n24259 ;
  assign n24274 = n24273 ^ n24260 ;
  assign n24256 = n24250 ^ n24245 ;
  assign n24275 = n24274 ^ n24256 ;
  assign n24276 = n24275 ^ n24250 ;
  assign n24277 = n24276 ^ n24242 ;
  assign n24255 = n24254 ^ n24251 ;
  assign n24278 = n24277 ^ n24255 ;
  assign n24279 = n24278 ^ n24265 ;
  assign n24280 = ~n24238 & n24279 ;
  assign n24297 = n24261 ^ n24252 ;
  assign n24285 = n24278 ^ n24263 ;
  assign n24298 = n24297 ^ n24285 ;
  assign n24299 = n24298 ^ n24270 ;
  assign n24300 = n24299 ^ n24255 ;
  assign n24294 = n24273 ^ n24247 ;
  assign n24293 = n24246 & ~n24249 ;
  assign n24295 = n24294 ^ n24293 ;
  assign n24296 = n24295 ^ n24270 ;
  assign n24301 = n24300 ^ n24296 ;
  assign n24292 = n24269 ^ n24239 ;
  assign n24302 = n24301 ^ n24292 ;
  assign n24303 = n24236 & ~n24302 ;
  assign n24313 = ~n24238 & ~n24294 ;
  assign n24311 = n24260 ^ n24254 ;
  assign n24312 = n24311 ^ n24250 ;
  assign n24314 = n24313 ^ n24312 ;
  assign n24315 = n24314 ^ n24236 ;
  assign n24316 = n24279 ^ n24273 ;
  assign n24317 = n24316 ^ n24238 ;
  assign n24318 = n24314 ^ n24238 ;
  assign n24319 = n24318 ^ n24238 ;
  assign n24320 = ~n24317 & ~n24319 ;
  assign n24321 = n24320 ^ n24238 ;
  assign n24322 = n24315 & ~n24321 ;
  assign n24323 = n24322 ^ n24236 ;
  assign n24309 = n24293 ^ n24266 ;
  assign n24310 = n24237 & n24309 ;
  assign n24324 = n24323 ^ n24310 ;
  assign n24305 = n24261 ^ n24254 ;
  assign n24306 = n24305 ^ n24265 ;
  assign n24304 = n24302 ^ n24298 ;
  assign n24307 = n24306 ^ n24304 ;
  assign n24308 = n24235 & n24307 ;
  assign n24325 = n24324 ^ n24308 ;
  assign n24326 = ~n24303 & ~n24325 ;
  assign n24284 = n24234 ^ n24233 ;
  assign n24327 = n24263 ^ n24261 ;
  assign n24328 = n24263 ^ n24234 ;
  assign n24329 = n24328 ^ n24263 ;
  assign n24330 = n24327 & n24329 ;
  assign n24331 = n24330 ^ n24263 ;
  assign n24332 = ~n24284 & n24331 ;
  assign n24333 = n24293 ^ n24270 ;
  assign n24334 = n24270 ^ n24234 ;
  assign n24335 = n24334 ^ n24270 ;
  assign n24336 = n24333 & ~n24335 ;
  assign n24337 = n24336 ^ n24270 ;
  assign n24338 = n24284 & n24337 ;
  assign n24339 = ~n24332 & ~n24338 ;
  assign n24340 = n24326 & n24339 ;
  assign n24281 = n24275 ^ n24272 ;
  assign n24286 = n24285 ^ n24281 ;
  assign n24287 = n24285 ^ n24234 ;
  assign n24288 = n24287 ^ n24285 ;
  assign n24289 = n24286 & ~n24288 ;
  assign n24290 = n24289 ^ n24285 ;
  assign n24291 = n24284 & n24290 ;
  assign n24341 = n24340 ^ n24291 ;
  assign n24282 = n24281 ^ n24273 ;
  assign n24283 = n24237 & ~n24282 ;
  assign n24342 = n24341 ^ n24283 ;
  assign n24343 = ~n24280 & n24342 ;
  assign n24344 = n24343 ^ n21185 ;
  assign n24366 = n23514 & n23612 ;
  assign n24367 = n24200 & n24366 ;
  assign n24363 = n23637 ^ n23595 ;
  assign n24364 = n24363 ^ n24200 ;
  assign n24354 = n24212 ^ n23637 ;
  assign n24355 = n24354 ^ n23647 ;
  assign n24356 = n23512 & ~n24355 ;
  assign n24357 = n24356 ^ n23649 ;
  assign n24362 = n24357 ^ n23592 ;
  assign n24365 = n24364 ^ n24362 ;
  assign n24368 = n24367 ^ n24365 ;
  assign n24360 = n23613 ^ n23592 ;
  assign n24361 = ~n23512 & n24360 ;
  assign n24369 = n24368 ^ n24361 ;
  assign n24370 = ~n24191 & n24369 ;
  assign n24353 = n23644 ^ n23595 ;
  assign n24358 = n24357 ^ n24353 ;
  assign n24349 = n23616 ^ n23597 ;
  assign n24350 = n24194 & n24349 ;
  assign n24351 = n24350 ^ n23597 ;
  assign n24352 = ~n23511 & n24351 ;
  assign n24359 = n24358 ^ n24352 ;
  assign n24371 = n24370 ^ n24359 ;
  assign n24372 = n24371 ^ n24190 ;
  assign n24373 = n24372 ^ n23654 ;
  assign n24374 = n24373 ^ n20916 ;
  assign n24345 = n24210 ^ n24199 ;
  assign n24346 = n23512 & ~n24345 ;
  assign n24347 = n24346 ^ n24199 ;
  assign n24348 = n23511 & n24347 ;
  assign n24375 = n24374 ^ n24348 ;
  assign n24376 = n23256 ^ x100 ;
  assign n24377 = n22572 ^ x118 ;
  assign n24380 = n21800 ^ x101 ;
  assign n24383 = n23704 ^ x124 ;
  assign n24402 = ~n24380 & n24383 ;
  assign n24379 = n23070 ^ x94 ;
  assign n24381 = ~n24379 & n24380 ;
  assign n24382 = n24381 ^ n24379 ;
  assign n24384 = n24125 ^ x76 ;
  assign n24385 = ~n24383 & n24384 ;
  assign n24400 = ~n24382 & n24385 ;
  assign n24420 = n24402 ^ n24400 ;
  assign n24389 = n24382 ^ n24380 ;
  assign n24404 = n24385 ^ n24383 ;
  assign n24405 = n24389 & ~n24404 ;
  assign n24386 = n24385 ^ n24384 ;
  assign n24387 = n24386 ^ n24383 ;
  assign n24388 = ~n24382 & n24387 ;
  assign n24406 = n24405 ^ n24388 ;
  assign n24390 = n24385 & n24389 ;
  assign n24407 = n24406 ^ n24390 ;
  assign n24403 = n24402 ^ n24389 ;
  assign n24408 = n24407 ^ n24403 ;
  assign n24398 = n24386 & n24389 ;
  assign n24401 = n24400 ^ n24398 ;
  assign n24409 = n24408 ^ n24401 ;
  assign n24410 = n24409 ^ n24388 ;
  assign n24421 = n24420 ^ n24410 ;
  assign n24422 = n24421 ^ n24408 ;
  assign n24475 = n24422 ^ n24400 ;
  assign n24412 = n24389 ^ n24379 ;
  assign n24416 = n24386 & n24412 ;
  assign n24415 = n24385 & n24412 ;
  assign n24417 = n24416 ^ n24415 ;
  assign n24413 = n24387 & n24412 ;
  assign n24414 = n24413 ^ n24412 ;
  assign n24418 = n24417 ^ n24414 ;
  assign n24476 = n24475 ^ n24418 ;
  assign n24477 = n24476 ^ n24385 ;
  assign n24441 = n24381 & n24387 ;
  assign n24473 = n24441 ^ n24418 ;
  assign n24474 = n24473 ^ n24415 ;
  assign n24478 = n24477 ^ n24474 ;
  assign n24479 = n24377 & n24478 ;
  assign n24435 = ~n24376 & ~n24377 ;
  assign n24436 = n24435 ^ n24377 ;
  assign n24437 = n24436 ^ n24376 ;
  assign n24432 = n24408 ^ n24398 ;
  assign n24431 = n24416 ^ n24386 ;
  assign n24433 = n24432 ^ n24431 ;
  assign n24438 = n24433 ^ n24415 ;
  assign n24439 = ~n24436 & n24438 ;
  assign n24440 = n24439 ^ n24416 ;
  assign n24442 = n24441 ^ n24440 ;
  assign n24443 = n24437 & ~n24442 ;
  assign n24444 = n24443 ^ n24377 ;
  assign n24445 = n24444 ^ n24443 ;
  assign n24434 = n24433 ^ n24413 ;
  assign n24446 = n24445 ^ n24434 ;
  assign n24447 = n24446 ^ n24445 ;
  assign n24378 = n24377 ^ n24376 ;
  assign n24448 = n24381 & ~n24404 ;
  assign n24449 = n24448 ^ n24438 ;
  assign n24450 = n24376 & ~n24449 ;
  assign n24451 = n24450 ^ n24449 ;
  assign n24452 = n24451 ^ n24443 ;
  assign n24453 = n24452 ^ n24451 ;
  assign n24456 = n24451 ^ n24416 ;
  assign n24457 = n24456 ^ n24451 ;
  assign n24458 = n24450 & ~n24457 ;
  assign n24459 = ~n24453 & n24458 ;
  assign n24460 = n24459 ^ n24453 ;
  assign n24461 = n24460 ^ n24452 ;
  assign n24462 = ~n24378 & ~n24461 ;
  assign n24463 = ~n24447 & n24462 ;
  assign n24464 = n24463 ^ n24377 ;
  assign n24399 = n24398 ^ n24382 ;
  assign n24411 = n24410 ^ n24399 ;
  assign n24423 = n24422 ^ n24411 ;
  assign n24419 = n24418 ^ n24411 ;
  assign n24424 = n24423 ^ n24419 ;
  assign n24425 = n24423 ^ n24376 ;
  assign n24426 = n24425 ^ n24423 ;
  assign n24427 = n24424 & ~n24426 ;
  assign n24428 = n24427 ^ n24423 ;
  assign n24429 = n24378 & ~n24428 ;
  assign n24430 = n24429 ^ n24411 ;
  assign n24465 = n24464 ^ n24430 ;
  assign n24466 = n24465 ^ n21589 ;
  assign n24471 = n24466 ^ n24401 ;
  assign n24468 = n24405 ^ n24400 ;
  assign n24469 = ~n24436 & n24468 ;
  assign n24472 = n24471 ^ n24469 ;
  assign n24480 = n24479 ^ n24472 ;
  assign n24467 = n24466 ^ n24444 ;
  assign n24470 = n24469 ^ n24467 ;
  assign n24481 = n24480 ^ n24470 ;
  assign n24482 = n24376 & n24481 ;
  assign n24483 = n24482 ^ n24480 ;
  assign n24393 = n24388 ^ n24376 ;
  assign n24394 = n24393 ^ n24388 ;
  assign n24395 = n24390 & n24394 ;
  assign n24396 = n24395 ^ n24388 ;
  assign n24397 = ~n24378 & n24396 ;
  assign n24484 = n24483 ^ n24397 ;
  assign n24497 = n24448 ^ n24443 ;
  assign n24498 = n24439 ^ n24378 ;
  assign n24499 = ~n24413 & ~n24498 ;
  assign n24500 = n24497 & n24499 ;
  assign n24501 = n24500 ^ n24498 ;
  assign n24517 = n24501 ^ n24432 ;
  assign n24509 = n24418 ^ n24388 ;
  assign n24510 = n24509 ^ n24476 ;
  assign n24511 = n24510 ^ n24509 ;
  assign n24512 = n24509 ^ n24376 ;
  assign n24513 = n24512 ^ n24509 ;
  assign n24514 = n24511 & ~n24513 ;
  assign n24515 = n24514 ^ n24509 ;
  assign n24516 = n24378 & n24515 ;
  assign n24518 = n24517 ^ n24516 ;
  assign n24504 = n24440 ^ n24388 ;
  assign n24502 = n24381 & n24385 ;
  assign n24503 = n24502 ^ n24413 ;
  assign n24505 = n24504 ^ n24503 ;
  assign n24506 = ~n24501 & ~n24505 ;
  assign n24507 = n24506 ^ n24432 ;
  assign n24508 = ~n24435 & n24507 ;
  assign n24519 = n24518 ^ n24508 ;
  assign n24496 = n24400 & ~n24437 ;
  assign n24520 = n24519 ^ n24496 ;
  assign n24521 = n24520 ^ n24405 ;
  assign n24522 = n24521 ^ n24430 ;
  assign n24488 = n24411 ^ n24390 ;
  assign n24486 = n24449 ^ n24405 ;
  assign n24487 = n24486 ^ n24449 ;
  assign n24489 = n24488 ^ n24487 ;
  assign n24490 = n24489 ^ n24486 ;
  assign n24491 = n24486 ^ n24376 ;
  assign n24492 = n24491 ^ n24486 ;
  assign n24493 = ~n24490 & n24492 ;
  assign n24494 = n24493 ^ n24486 ;
  assign n24495 = n24378 & n24494 ;
  assign n24523 = n24522 ^ n24495 ;
  assign n24485 = n24398 & ~n24437 ;
  assign n24524 = n24523 ^ n24485 ;
  assign n24525 = n24524 ^ n22078 ;
  assign n24536 = n23354 ^ n23315 ;
  assign n24534 = n23346 ^ n23324 ;
  assign n24537 = n24536 ^ n24534 ;
  assign n24538 = n23180 & ~n24537 ;
  assign n24527 = n23354 ^ n23352 ;
  assign n24528 = n24527 ^ n23329 ;
  assign n24529 = n23180 & ~n24528 ;
  assign n24530 = n24529 ^ n23357 ;
  assign n24533 = n24530 ^ n23340 ;
  assign n24535 = n24534 ^ n24533 ;
  assign n24539 = n24538 ^ n24535 ;
  assign n24540 = ~n23427 & ~n24539 ;
  assign n24526 = n23425 ^ n23327 ;
  assign n24531 = n24530 ^ n24526 ;
  assign n24532 = n24531 ^ n23392 ;
  assign n24541 = n24540 ^ n24532 ;
  assign n24542 = ~n23458 & n24541 ;
  assign n24543 = n24542 ^ n21328 ;
  assign n24584 = n22444 ^ x112 ;
  assign n24544 = n22843 ^ x65 ;
  assign n24548 = n22719 ^ x72 ;
  assign n24546 = n21524 ^ x89 ;
  assign n24586 = n24548 ^ n24546 ;
  assign n24545 = n23498 ^ x98 ;
  assign n24553 = n24545 & ~n24548 ;
  assign n24560 = n24553 ^ n24545 ;
  assign n24558 = n24047 ^ x107 ;
  assign n24562 = n24558 ^ n24548 ;
  assign n24563 = ~n24560 & ~n24562 ;
  assign n24575 = ~n24546 & n24563 ;
  assign n24597 = n24575 ^ n24546 ;
  assign n24551 = ~n24545 & ~n24546 ;
  assign n24552 = n24548 & ~n24551 ;
  assign n24554 = n24553 ^ n24552 ;
  assign n24555 = n24554 ^ n24551 ;
  assign n24549 = n24548 ^ n24545 ;
  assign n24550 = n24546 & ~n24549 ;
  assign n24556 = n24555 ^ n24550 ;
  assign n24571 = n24560 ^ n24556 ;
  assign n24572 = n24558 & ~n24571 ;
  assign n24596 = n24572 ^ n24551 ;
  assign n24598 = n24597 ^ n24596 ;
  assign n24589 = n24558 & n24586 ;
  assign n24590 = n24589 ^ n24546 ;
  assign n24591 = ~n24545 & n24590 ;
  assign n24588 = n24562 ^ n24546 ;
  assign n24592 = n24591 ^ n24588 ;
  assign n24587 = n24558 ^ n24549 ;
  assign n24593 = n24592 ^ n24587 ;
  assign n24594 = n24593 ^ n24549 ;
  assign n24595 = n24594 ^ n24592 ;
  assign n24599 = n24598 ^ n24595 ;
  assign n24600 = n24586 & ~n24599 ;
  assign n24601 = n24600 ^ n24593 ;
  assign n24602 = ~n24544 & ~n24601 ;
  assign n24603 = n24602 ^ n24592 ;
  assign n24567 = n24555 ^ n24546 ;
  assign n24576 = n24575 ^ n24567 ;
  assign n24573 = n24572 ^ n24556 ;
  assign n24564 = n24563 ^ n24562 ;
  assign n24574 = n24573 ^ n24564 ;
  assign n24577 = n24576 ^ n24574 ;
  assign n24559 = n24548 & ~n24558 ;
  assign n24561 = n24560 ^ n24559 ;
  assign n24565 = n24564 ^ n24561 ;
  assign n24566 = n24565 ^ n24563 ;
  assign n24568 = n24567 ^ n24566 ;
  assign n24578 = n24577 ^ n24568 ;
  assign n24579 = n24578 ^ n24567 ;
  assign n24580 = n24579 ^ n24549 ;
  assign n24557 = n24556 ^ n24552 ;
  assign n24569 = n24568 ^ n24557 ;
  assign n24547 = n24546 ^ n24545 ;
  assign n24570 = n24569 ^ n24547 ;
  assign n24581 = n24580 ^ n24570 ;
  assign n24582 = n24544 & ~n24581 ;
  assign n24583 = n24582 ^ n24580 ;
  assign n24604 = n24603 ^ n24583 ;
  assign n24605 = n24584 & n24604 ;
  assign n24606 = n24605 ^ n24603 ;
  assign n24585 = n24584 ^ n24583 ;
  assign n24607 = n24606 ^ n24585 ;
  assign n24608 = n24607 ^ n24603 ;
  assign n24609 = n24608 ^ n20390 ;
  assign n24635 = n24272 ^ n24254 ;
  assign n24636 = n24635 ^ n24273 ;
  assign n24637 = n24636 ^ n24302 ;
  assign n24638 = ~n24233 & ~n24637 ;
  assign n24639 = n24638 ^ n24262 ;
  assign n24640 = n24234 & n24639 ;
  assign n24622 = n24293 ^ n24236 ;
  assign n24623 = n24273 ^ n24238 ;
  assign n24626 = ~n24293 & ~n24623 ;
  assign n24627 = n24626 ^ n24238 ;
  assign n24628 = n24622 & ~n24627 ;
  assign n24629 = n24628 ^ n24236 ;
  assign n24611 = n24299 ^ n24247 ;
  assign n24630 = n24629 ^ n24611 ;
  assign n24631 = n24630 ^ n24291 ;
  assign n24620 = n24235 & n24279 ;
  assign n24621 = n24620 ^ n24303 ;
  assign n24632 = n24631 ^ n24621 ;
  assign n24612 = n24611 ^ n24250 ;
  assign n24613 = n24612 ^ n24268 ;
  assign n24614 = n24613 ^ n24611 ;
  assign n24615 = n24611 ^ n24234 ;
  assign n24616 = n24615 ^ n24611 ;
  assign n24617 = n24614 & ~n24616 ;
  assign n24618 = n24617 ^ n24611 ;
  assign n24619 = n24284 & ~n24618 ;
  assign n24633 = n24632 ^ n24619 ;
  assign n24610 = ~n24238 & ~n24276 ;
  assign n24634 = n24633 ^ n24610 ;
  assign n24641 = n24640 ^ n24634 ;
  assign n24642 = n24641 ^ n24280 ;
  assign n24643 = n24642 ^ n21551 ;
  assign n24672 = n24060 ^ n22619 ;
  assign n24673 = n22628 & ~n24672 ;
  assign n24654 = n22597 ^ n22577 ;
  assign n24655 = n24654 ^ n22619 ;
  assign n24653 = n22652 ^ n22598 ;
  assign n24656 = n24655 ^ n24653 ;
  assign n24657 = ~n21525 & n24656 ;
  assign n24658 = n24657 ^ n24655 ;
  assign n24666 = n24658 ^ n22682 ;
  assign n24667 = n24666 ^ n22651 ;
  assign n24668 = n24667 ^ n22588 ;
  assign n24669 = n24668 ^ n22359 ;
  assign n24659 = n24658 ^ n22643 ;
  assign n24660 = n24659 ^ n22609 ;
  assign n24661 = n24660 ^ n22615 ;
  assign n24662 = n24661 ^ n24658 ;
  assign n24663 = n21525 & n24662 ;
  assign n24664 = n24663 ^ n24659 ;
  assign n24665 = n21802 & n24664 ;
  assign n24670 = n24669 ^ n24665 ;
  assign n24652 = ~n22627 & n22629 ;
  assign n24671 = n24670 ^ n24652 ;
  assign n24674 = n24673 ^ n24671 ;
  assign n24651 = ~n21802 & n22613 ;
  assign n24675 = n24674 ^ n24651 ;
  assign n24644 = n22614 ^ n22578 ;
  assign n24645 = n24644 ^ n22631 ;
  assign n24646 = n22631 ^ n21525 ;
  assign n24647 = n24646 ^ n22631 ;
  assign n24648 = n24645 & ~n24647 ;
  assign n24649 = n24648 ^ n22631 ;
  assign n24650 = n21801 & n24649 ;
  assign n24676 = n24675 ^ n24650 ;
  assign n24693 = n24502 ^ n24408 ;
  assign n24691 = n24421 ^ n24406 ;
  assign n24692 = n24435 & n24691 ;
  assign n24694 = n24693 ^ n24692 ;
  assign n24695 = n24694 ^ n24448 ;
  assign n24690 = ~n24437 & ~n24488 ;
  assign n24696 = n24695 ^ n24690 ;
  assign n24700 = n24696 ^ n24485 ;
  assign n24679 = n24416 ^ n24376 ;
  assign n24680 = n24679 ^ n24416 ;
  assign n24681 = n24417 & ~n24680 ;
  assign n24682 = n24681 ^ n24416 ;
  assign n24683 = ~n24378 & n24682 ;
  assign n24701 = n24700 ^ n24683 ;
  assign n24689 = n24473 ^ n24434 ;
  assign n24697 = n24696 ^ n24689 ;
  assign n24685 = n24407 ^ n24400 ;
  assign n24686 = n24685 ^ n24473 ;
  assign n24687 = n24686 ^ n24434 ;
  assign n24688 = n24376 & n24687 ;
  assign n24698 = n24697 ^ n24688 ;
  assign n24699 = n24378 & n24698 ;
  assign n24702 = n24701 ^ n24699 ;
  assign n24684 = ~n24377 & n24413 ;
  assign n24703 = n24702 ^ n24684 ;
  assign n24704 = n24703 ^ n24683 ;
  assign n24705 = n24437 ^ n24377 ;
  assign n24706 = n24406 & ~n24705 ;
  assign n24707 = ~n24704 & n24706 ;
  assign n24708 = n24707 ^ n24703 ;
  assign n24709 = n24418 ^ n24401 ;
  assign n24710 = n24376 & n24709 ;
  assign n24711 = n24710 ^ n24401 ;
  assign n24714 = n24711 ^ n24448 ;
  assign n24715 = n24714 ^ n24711 ;
  assign n24716 = n24376 & n24715 ;
  assign n24717 = n24716 ^ n24711 ;
  assign n24718 = ~n24377 & n24717 ;
  assign n24719 = n24718 ^ n24711 ;
  assign n24720 = ~n24439 & ~n24719 ;
  assign n24721 = ~n24708 & n24720 ;
  assign n24722 = n24721 ^ n21376 ;
  assign n24726 = n24438 ^ n24410 ;
  assign n24727 = n24726 ^ n24503 ;
  assign n24728 = ~n24376 & n24727 ;
  assign n24729 = n24728 ^ n24410 ;
  assign n24737 = n24729 ^ n24485 ;
  assign n24733 = n24502 ^ n24416 ;
  assign n24734 = ~n24376 & n24733 ;
  assign n24731 = n24406 & n24435 ;
  assign n24725 = n24496 ^ n24488 ;
  assign n24730 = n24729 ^ n24725 ;
  assign n24732 = n24731 ^ n24730 ;
  assign n24735 = n24734 ^ n24732 ;
  assign n24736 = ~n24378 & ~n24735 ;
  assign n24738 = n24737 ^ n24736 ;
  assign n24724 = ~n24436 & n24474 ;
  assign n24739 = n24738 ^ n24724 ;
  assign n24740 = n24377 & ~n24739 ;
  assign n24741 = n24421 ^ n24376 ;
  assign n24742 = n24741 ^ n24421 ;
  assign n24743 = n24421 ^ n24411 ;
  assign n24744 = n24743 ^ n24421 ;
  assign n24745 = ~n24742 & ~n24744 ;
  assign n24746 = n24745 ^ n24421 ;
  assign n24747 = n24740 & n24746 ;
  assign n24748 = n24747 ^ n24739 ;
  assign n24749 = ~n24719 & ~n24748 ;
  assign n24750 = n24749 ^ n20221 ;
  assign n24723 = ~n24378 & n24434 ;
  assign n24753 = n24750 ^ n24723 ;
  assign n24754 = n23615 ^ n23608 ;
  assign n24771 = n24754 ^ n23623 ;
  assign n24772 = n24771 ^ n24347 ;
  assign n24773 = n24772 ^ n24197 ;
  assign n24774 = n24773 ^ n24352 ;
  assign n24764 = n24347 ^ n24224 ;
  assign n24763 = n24354 ^ n24347 ;
  assign n24765 = n24764 ^ n24763 ;
  assign n24768 = ~n23512 & ~n24765 ;
  assign n24769 = n24768 ^ n24764 ;
  assign n24770 = ~n23511 & n24769 ;
  assign n24775 = n24774 ^ n24770 ;
  assign n24755 = n24754 ^ n23611 ;
  assign n24756 = n24755 ^ n23613 ;
  assign n24757 = n24756 ^ n24754 ;
  assign n24758 = n24754 ^ n23512 ;
  assign n24759 = n24758 ^ n24754 ;
  assign n24760 = n24757 & ~n24759 ;
  assign n24761 = n24760 ^ n24754 ;
  assign n24762 = n24191 & n24761 ;
  assign n24776 = n24775 ^ n24762 ;
  assign n24777 = n24776 ^ n24190 ;
  assign n24778 = n24777 ^ n23654 ;
  assign n24779 = n24778 ^ n22757 ;
  assign n24793 = n24283 ^ n24266 ;
  assign n24794 = n24793 ^ n24283 ;
  assign n24795 = n24794 ^ n24250 ;
  assign n24796 = n24795 ^ n24794 ;
  assign n24797 = n24794 ^ n24234 ;
  assign n24798 = n24797 ^ n24794 ;
  assign n24799 = n24796 & n24798 ;
  assign n24800 = n24799 ^ n24794 ;
  assign n24801 = n24284 & n24800 ;
  assign n24802 = n24801 ^ n24793 ;
  assign n24803 = n24802 ^ n24621 ;
  assign n24790 = n24272 ^ n24251 ;
  assign n24791 = n24790 ^ n24298 ;
  assign n24792 = n24236 & n24791 ;
  assign n24804 = n24803 ^ n24792 ;
  assign n24789 = n24278 & ~n24284 ;
  assign n24805 = n24804 ^ n24789 ;
  assign n24784 = n24296 ^ n24233 ;
  assign n24785 = n24784 ^ n24296 ;
  assign n24786 = n24301 & n24785 ;
  assign n24787 = n24786 ^ n24296 ;
  assign n24788 = ~n24234 & ~n24787 ;
  assign n24806 = n24805 ^ n24788 ;
  assign n24781 = n24237 & n24306 ;
  assign n24807 = n24806 ^ n24781 ;
  assign n24808 = ~n24332 & ~n24807 ;
  assign n24809 = ~n24338 & n24808 ;
  assign n24810 = n24809 ^ n22323 ;
  assign n24780 = ~n24238 & n24261 ;
  assign n24813 = n24810 ^ n24780 ;
  assign n24823 = n24551 & n24559 ;
  assign n24821 = n24565 ^ n24554 ;
  assign n24820 = n24590 ^ n24574 ;
  assign n24822 = n24821 ^ n24820 ;
  assign n24824 = n24823 ^ n24822 ;
  assign n24814 = n24551 ^ n24546 ;
  assign n24817 = ~n24562 & n24814 ;
  assign n24818 = n24817 ^ n24551 ;
  assign n24819 = n24573 & ~n24818 ;
  assign n24825 = n24824 ^ n24819 ;
  assign n24826 = ~n24544 & n24825 ;
  assign n24827 = n24826 ^ n24824 ;
  assign n24836 = n24827 ^ n21435 ;
  assign n24829 = n24827 ^ n24577 ;
  assign n24828 = n24827 ^ n24568 ;
  assign n24830 = n24829 ^ n24828 ;
  assign n24833 = ~n24544 & n24830 ;
  assign n24834 = n24833 ^ n24829 ;
  assign n24835 = n24584 & n24834 ;
  assign n24837 = n24836 ^ n24835 ;
  assign n24847 = n24298 ^ n24234 ;
  assign n24848 = n24284 & ~n24847 ;
  assign n24849 = n24848 ^ n24234 ;
  assign n24852 = n24298 ^ n24268 ;
  assign n24853 = ~n24849 & ~n24852 ;
  assign n24850 = n24268 ^ n24261 ;
  assign n24854 = n24853 ^ n24850 ;
  assign n24865 = n24854 ^ n24629 ;
  assign n24859 = n24244 ^ n24239 ;
  assign n24860 = n24240 & n24859 ;
  assign n24857 = n24854 ^ n24269 ;
  assign n24855 = n24244 ^ n24243 ;
  assign n24856 = n24855 ^ n24854 ;
  assign n24858 = n24857 ^ n24856 ;
  assign n24861 = n24860 ^ n24858 ;
  assign n24862 = ~n24234 & n24861 ;
  assign n24863 = n24862 ^ n24857 ;
  assign n24864 = n24284 & n24863 ;
  assign n24866 = n24865 ^ n24864 ;
  assign n24845 = n24302 ^ n24274 ;
  assign n24846 = ~n24238 & n24845 ;
  assign n24867 = n24866 ^ n24846 ;
  assign n24840 = n24251 ^ n24233 ;
  assign n24841 = n24840 ^ n24251 ;
  assign n24842 = n24258 & ~n24841 ;
  assign n24843 = n24842 ^ n24251 ;
  assign n24844 = n24234 & n24843 ;
  assign n24868 = n24867 ^ n24844 ;
  assign n24869 = ~n24280 & ~n24868 ;
  assign n24870 = n24869 ^ n19894 ;
  assign n24871 = n24606 ^ n22722 ;
  assign n24873 = n24577 ^ n24549 ;
  assign n24874 = n24873 ^ n24601 ;
  assign n24876 = ~n24544 & ~n24584 ;
  assign n24877 = ~n24874 & n24876 ;
  assign n24872 = n24574 ^ n24568 ;
  assign n24875 = n24874 ^ n24872 ;
  assign n24878 = n24877 ^ n24875 ;
  assign n24879 = n24819 ^ n24576 ;
  assign n24880 = ~n24544 & ~n24879 ;
  assign n24881 = n24880 ^ n24576 ;
  assign n24882 = n24881 ^ n24584 ;
  assign n24883 = n24882 ^ n24544 ;
  assign n24884 = n24883 ^ n24881 ;
  assign n24885 = n24544 & ~n24824 ;
  assign n24886 = n24885 ^ n24881 ;
  assign n24887 = ~n24884 & n24886 ;
  assign n24888 = n24887 ^ n24881 ;
  assign n24889 = n24878 & n24888 ;
  assign n24890 = n24889 ^ n24878 ;
  assign n24891 = ~n24574 & n24890 ;
  assign n24892 = n24891 ^ n21560 ;
  assign n24933 = n23736 & n23849 ;
  assign n24926 = n23893 ^ n23834 ;
  assign n24927 = n24926 ^ n23927 ;
  assign n24921 = n23875 ^ n23836 ;
  assign n24922 = n24921 ^ n23867 ;
  assign n24923 = n24922 ^ n23864 ;
  assign n24928 = n24927 ^ n24923 ;
  assign n24929 = n23736 & ~n24928 ;
  assign n24910 = n23864 ^ n23833 ;
  assign n24911 = n24910 ^ n23882 ;
  assign n24912 = n24911 ^ n23855 ;
  assign n24909 = n23863 ^ n23837 ;
  assign n24913 = n24912 ^ n24909 ;
  assign n24914 = n23736 & n24913 ;
  assign n24915 = n24914 ^ n24912 ;
  assign n24924 = n24923 ^ n24915 ;
  assign n24930 = n24929 ^ n24924 ;
  assign n24931 = n23705 & ~n24930 ;
  assign n24916 = n24915 ^ n23940 ;
  assign n24905 = n23867 ^ n23855 ;
  assign n24906 = ~n23935 & ~n24905 ;
  assign n24907 = n24906 ^ n23855 ;
  assign n24908 = n23737 & n24907 ;
  assign n24917 = n24916 ^ n24908 ;
  assign n24918 = n24917 ^ n23949 ;
  assign n24899 = n23893 ^ n23875 ;
  assign n24900 = n23875 ^ n23705 ;
  assign n24901 = n24900 ^ n23875 ;
  assign n24902 = n24899 & n24901 ;
  assign n24903 = n24902 ^ n23875 ;
  assign n24904 = n23737 & n24903 ;
  assign n24919 = n24918 ^ n24904 ;
  assign n24893 = n23927 ^ n23863 ;
  assign n24894 = n23863 ^ n23705 ;
  assign n24895 = n24894 ^ n23863 ;
  assign n24896 = n24893 & ~n24895 ;
  assign n24897 = n24896 ^ n23863 ;
  assign n24898 = ~n23737 & n24897 ;
  assign n24920 = n24919 ^ n24898 ;
  assign n24932 = n24931 ^ n24920 ;
  assign n24934 = n24933 ^ n24932 ;
  assign n24935 = ~n23879 & ~n24934 ;
  assign n24936 = n24935 ^ n21411 ;
  assign n24962 = ~n23879 & n23921 ;
  assign n24957 = n23877 ^ n23855 ;
  assign n24958 = n24957 ^ n23893 ;
  assign n24959 = n24958 ^ n24911 ;
  assign n24960 = n23736 & n24959 ;
  assign n24954 = n24911 ^ n23876 ;
  assign n24955 = n23844 & n24954 ;
  assign n24946 = n23879 ^ n23863 ;
  assign n24947 = n24946 ^ n24904 ;
  assign n24943 = n24908 ^ n23864 ;
  assign n24942 = n24898 ^ n23843 ;
  assign n24944 = n24943 ^ n24942 ;
  assign n24941 = n24911 ^ n23877 ;
  assign n24945 = n24944 ^ n24941 ;
  assign n24948 = n24947 ^ n24945 ;
  assign n24949 = n24948 ^ n23953 ;
  assign n24950 = n24949 ^ n23859 ;
  assign n24951 = n24950 ^ n20618 ;
  assign n24939 = n23887 ^ n23833 ;
  assign n24940 = n23705 & n24939 ;
  assign n24952 = n24951 ^ n24940 ;
  assign n24937 = n24911 ^ n23863 ;
  assign n24938 = ~n23864 & n24937 ;
  assign n24953 = n24952 ^ n24938 ;
  assign n24956 = n24955 ^ n24953 ;
  assign n24961 = n24960 ^ n24956 ;
  assign n24963 = n24962 ^ n24961 ;
  assign n24979 = n24060 ^ n22610 ;
  assign n24976 = n22617 ^ n22598 ;
  assign n24977 = n21525 & n24976 ;
  assign n24978 = n24977 ^ n22638 ;
  assign n24980 = n24979 ^ n24978 ;
  assign n24972 = n22635 ^ n22610 ;
  assign n24973 = n24972 ^ n22630 ;
  assign n24974 = n24973 ^ n24060 ;
  assign n24975 = n21525 & ~n24974 ;
  assign n24981 = n24980 ^ n24975 ;
  assign n24982 = n21802 & ~n24981 ;
  assign n24983 = n24982 ^ n24978 ;
  assign n24971 = n22616 & n22625 ;
  assign n24984 = n24983 ^ n24971 ;
  assign n24970 = n22626 & n24074 ;
  assign n24985 = n24984 ^ n24970 ;
  assign n24964 = n22632 ^ n22598 ;
  assign n24965 = n22598 ^ n21525 ;
  assign n24966 = n24965 ^ n22598 ;
  assign n24967 = n24964 & ~n24966 ;
  assign n24968 = n24967 ^ n22598 ;
  assign n24969 = ~n21801 & n24968 ;
  assign n24986 = n24985 ^ n24969 ;
  assign n24987 = ~n22673 & ~n24986 ;
  assign n24988 = ~n24085 & n24987 ;
  assign n24989 = n24988 ^ n21969 ;
  assign y0 = ~n20972 ;
  assign y1 = ~n22685 ;
  assign y2 = ~n21524 ;
  assign y3 = ~n23047 ;
  assign y4 = n23070 ;
  assign y5 = ~n23109 ;
  assign y6 = n23150 ;
  assign y7 = n23395 ;
  assign y8 = ~n23424 ;
  assign y9 = ~n23460 ;
  assign y10 = n23498 ;
  assign y11 = ~n23669 ;
  assign y12 = ~n23704 ;
  assign y13 = n23914 ;
  assign y14 = ~n23553 ;
  assign y15 = ~n23956 ;
  assign y16 = ~n23994 ;
  assign y17 = n24026 ;
  assign y18 = ~n24047 ;
  assign y19 = n24087 ;
  assign y20 = n24125 ;
  assign y21 = n24163 ;
  assign y22 = ~n23588 ;
  assign y23 = ~n24189 ;
  assign y24 = ~n23735 ;
  assign y25 = ~n24232 ;
  assign y26 = n22719 ;
  assign y27 = n24344 ;
  assign y28 = ~n21800 ;
  assign y29 = n24375 ;
  assign y30 = n23179 ;
  assign y31 = ~n24484 ;
  assign y32 = n23828 ;
  assign y33 = n24525 ;
  assign y34 = n22843 ;
  assign y35 = ~n24543 ;
  assign y36 = ~n22572 ;
  assign y37 = ~n24609 ;
  assign y38 = n23218 ;
  assign y39 = n24643 ;
  assign y40 = n23789 ;
  assign y41 = n24676 ;
  assign y42 = ~n22887 ;
  assign y43 = ~n24722 ;
  assign y44 = n22042 ;
  assign y45 = ~n24753 ;
  assign y46 = ~n23306 ;
  assign y47 = n24779 ;
  assign y48 = ~n23759 ;
  assign y49 = n24813 ;
  assign y50 = ~n22959 ;
  assign y51 = ~n24837 ;
  assign y52 = n22275 ;
  assign y53 = ~n24870 ;
  assign y54 = n23221 ;
  assign y55 = n24871 ;
  assign y56 = n23510 ;
  assign y57 = n24892 ;
  assign y58 = n22934 ;
  assign y59 = ~n24936 ;
  assign y60 = n22444 ;
  assign y61 = ~n24963 ;
  assign y62 = ~n23256 ;
  assign y63 = ~n24989 ;
endmodule
