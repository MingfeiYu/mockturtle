module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n200 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n221 , n222 , n223 , n224 , n225 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n536 , n537 , n538 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n613 , n614 , n615 , n616 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1052 , n1053 , n1054 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1302 , n1303 , n1304 , n1305 , n1306 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1374 , n1375 , n1376 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2373 , n2374 , n2375 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3538 , n3539 , n3540 , n3541 , n3542 , n3547 , n3548 , n3550 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4217 , n4218 , n4219 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4939 , n4940 , n4941 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5526 , n5527 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5796 , n5797 , n5798 , n5801 , n5802 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6372 , n6373 , n6374 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6836 , n6837 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7472 , n7477 , n7478 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7497 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8175 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8469 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9577 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10139 , n10140 , n10143 , n10144 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10169 , n10170 , n10171 , n10172 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10184 , n10185 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10200 , n10201 , n10202 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10567 , n10568 , n10569 , n10570 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10757 , n10758 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11176 , n11177 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11548 , n11549 , n11550 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12998 , n12999 , n13000 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13901 , n13902 , n13903 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14104 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14355 , n14356 , n14357 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 ;
  assign n129 = ~x126 & ~x127 ;
  assign n130 = ~x125 & n129 ;
  assign n131 = ~x124 & n130 ;
  assign n9923 = x12 & x65 ;
  assign n9920 = x65 ^ x11 ;
  assign n9916 = x64 ^ x12 ;
  assign n9917 = n9916 ^ x65 ;
  assign n132 = ~x123 & n131 ;
  assign n133 = ~x122 & n132 ;
  assign n134 = ~x121 & n133 ;
  assign n135 = ~x120 & n134 ;
  assign n136 = ~x119 & n135 ;
  assign n137 = ~x118 & n136 ;
  assign n138 = ~x117 & n137 ;
  assign n139 = ~x116 & n138 ;
  assign n7828 = ~x17 & x64 ;
  assign n7829 = n7828 ^ x65 ;
  assign n142 = ~x111 & ~x112 ;
  assign n140 = ~x115 & n139 ;
  assign n143 = ~x113 & ~x114 ;
  assign n144 = n140 & n143 ;
  assign n145 = n142 & n144 ;
  assign n147 = ~x110 & n145 ;
  assign n148 = ~x109 & n147 ;
  assign n5813 = ~x108 & n148 ;
  assign n149 = ~x104 & ~x105 ;
  assign n150 = ~x106 & ~x107 ;
  assign n151 = ~x108 & n150 ;
  assign n152 = n149 & n151 ;
  assign n153 = n148 & n152 ;
  assign n154 = ~x103 & n153 ;
  assign n155 = ~x102 & n154 ;
  assign n156 = ~x101 & n155 ;
  assign n157 = ~x100 & n156 ;
  assign n158 = ~x99 & n157 ;
  assign n159 = ~x98 & n158 ;
  assign n160 = ~x97 & n159 ;
  assign n161 = ~x96 & n160 ;
  assign n162 = ~x95 & n161 ;
  assign n163 = ~x94 & n162 ;
  assign n164 = ~x93 & n163 ;
  assign n165 = ~x92 & n164 ;
  assign n166 = ~x91 & n165 ;
  assign n167 = ~x90 & n166 ;
  assign n168 = ~x89 & n167 ;
  assign n169 = ~x88 & n168 ;
  assign n170 = ~x85 & ~x86 ;
  assign n271 = ~x87 & n169 ;
  assign n272 = n170 & n271 ;
  assign n146 = ~x84 & ~x87 ;
  assign n171 = n169 & n170 ;
  assign n172 = n146 & n171 ;
  assign n173 = ~x83 & n172 ;
  assign n174 = ~x82 & n173 ;
  assign n175 = ~x81 & n174 ;
  assign n176 = ~x80 & n175 ;
  assign n177 = ~x79 & n176 ;
  assign n178 = ~x78 & n177 ;
  assign n179 = ~x77 & n178 ;
  assign n180 = ~x76 & n179 ;
  assign n181 = ~x75 & n180 ;
  assign n182 = ~x74 & n181 ;
  assign n183 = ~x73 & n182 ;
  assign n184 = ~x72 & n183 ;
  assign n185 = ~x71 & n184 ;
  assign n186 = ~x70 & n185 ;
  assign n187 = ~x69 & n186 ;
  assign n188 = ~x68 & n187 ;
  assign n189 = ~x67 & n188 ;
  assign n190 = x63 & n189 ;
  assign n247 = x65 ^ x61 ;
  assign n200 = n247 ^ x62 ;
  assign n203 = x64 & ~n200 ;
  assign n204 = n203 ^ x62 ;
  assign n205 = ~x66 & n189 ;
  assign n206 = ~x63 & x65 ;
  assign n207 = n205 & n206 ;
  assign n208 = n207 ^ n205 ;
  assign n211 = n203 ^ x64 ;
  assign n212 = ~n208 & n211 ;
  assign n191 = x65 ^ x64 ;
  assign n209 = n208 ^ n191 ;
  assign n213 = n212 ^ n209 ;
  assign n214 = n213 ^ n208 ;
  assign n215 = ~n204 & n214 ;
  assign n216 = n215 ^ n212 ;
  assign n217 = n216 ^ x65 ;
  assign n218 = n217 ^ n191 ;
  assign n221 = ~x66 & ~n191 ;
  assign n222 = x65 & n221 ;
  assign n223 = x62 & n222 ;
  assign n224 = n223 ^ n221 ;
  assign n225 = n224 ^ x66 ;
  assign n230 = ~n218 & n225 ;
  assign n231 = n230 ^ x66 ;
  assign n232 = n190 & ~n231 ;
  assign n233 = n232 ^ x63 ;
  assign n250 = x64 & n208 ;
  assign n253 = n250 ^ x62 ;
  assign n248 = x61 & ~x65 ;
  assign n249 = n248 ^ n247 ;
  assign n251 = ~x62 & n250 ;
  assign n252 = n249 & n251 ;
  assign n254 = n253 ^ n252 ;
  assign n263 = n254 ^ n251 ;
  assign n235 = x63 & n225 ;
  assign n236 = n235 ^ x66 ;
  assign n237 = n218 ^ x63 ;
  assign n238 = n237 ^ n189 ;
  assign n239 = ~n236 & n238 ;
  assign n240 = n239 ^ x63 ;
  assign n241 = n189 & n240 ;
  assign n259 = n248 ^ x65 ;
  assign n260 = x64 & ~n259 ;
  assign n261 = n260 ^ x65 ;
  assign n262 = n241 & n261 ;
  assign n264 = n263 ^ n262 ;
  assign n234 = x65 ^ x60 ;
  assign n242 = n241 ^ x61 ;
  assign n243 = n242 ^ x60 ;
  assign n244 = ~n234 & n243 ;
  assign n245 = n244 ^ x60 ;
  assign n246 = x64 & ~n245 ;
  assign n255 = n254 ^ n249 ;
  assign n256 = n255 ^ n253 ;
  assign n257 = ~n246 & ~n256 ;
  assign n265 = n264 ^ n257 ;
  assign n266 = n264 ^ x66 ;
  assign n267 = ~n265 & ~n266 ;
  assign n268 = n267 ^ x66 ;
  assign n273 = n268 ^ x67 ;
  assign n274 = n188 & n273 ;
  assign n275 = n233 & n274 ;
  assign n276 = n275 ^ n233 ;
  assign n277 = n187 & n276 ;
  assign n317 = x68 ^ x67 ;
  assign n280 = ~x67 & ~n232 ;
  assign n281 = n280 ^ x63 ;
  assign n282 = n273 ^ n188 ;
  assign n283 = n281 & ~n282 ;
  assign n284 = n283 ^ x67 ;
  assign n285 = n188 & ~n284 ;
  assign n293 = ~x60 & n285 ;
  assign n294 = n293 ^ n241 ;
  assign n295 = x64 & n294 ;
  assign n296 = n295 ^ x61 ;
  assign n288 = x65 & n285 ;
  assign n297 = n296 ^ n288 ;
  assign n298 = n297 ^ x66 ;
  assign n304 = x60 & x65 ;
  assign n299 = x65 ^ x59 ;
  assign n300 = x64 ^ x60 ;
  assign n301 = n300 ^ x65 ;
  assign n302 = n301 ^ n285 ;
  assign n303 = ~n299 & n302 ;
  assign n305 = n304 ^ n303 ;
  assign n308 = x64 & n305 ;
  assign n309 = n308 ^ n304 ;
  assign n310 = n309 ^ x65 ;
  assign n311 = n310 ^ n297 ;
  assign n312 = ~n298 & n311 ;
  assign n313 = n312 ^ x66 ;
  assign n278 = n257 ^ x66 ;
  assign n286 = ~n278 & n285 ;
  assign n287 = n286 ^ n264 ;
  assign n314 = n313 ^ n287 ;
  assign n315 = n313 ^ x67 ;
  assign n316 = n314 & n315 ;
  assign n318 = n317 ^ n316 ;
  assign n319 = n277 & n318 ;
  assign n320 = n319 ^ n276 ;
  assign n321 = x69 & ~n276 ;
  assign n322 = n186 & ~n321 ;
  assign n323 = n321 ^ x69 ;
  assign n324 = n323 ^ n320 ;
  assign n325 = n276 ^ x68 ;
  assign n328 = n318 & ~n325 ;
  assign n329 = n328 ^ x68 ;
  assign n330 = n187 & ~n329 ;
  assign n331 = n315 & n330 ;
  assign n332 = n331 ^ n287 ;
  assign n333 = n332 ^ x68 ;
  assign n342 = ~x59 & n330 ;
  assign n343 = n342 ^ n285 ;
  assign n344 = x64 & n343 ;
  assign n345 = n344 ^ x60 ;
  assign n337 = x65 & n330 ;
  assign n346 = n345 ^ n337 ;
  assign n347 = n346 ^ x66 ;
  assign n355 = x59 & x65 ;
  assign n352 = x65 ^ x58 ;
  assign n348 = x64 ^ x59 ;
  assign n349 = n348 ^ x65 ;
  assign n353 = n349 ^ n330 ;
  assign n354 = ~n352 & n353 ;
  assign n356 = n355 ^ n354 ;
  assign n357 = x64 & n356 ;
  assign n358 = n357 ^ n355 ;
  assign n359 = n358 ^ x65 ;
  assign n360 = n359 ^ n346 ;
  assign n361 = ~n347 & n360 ;
  assign n362 = n361 ^ x66 ;
  assign n334 = n310 ^ x66 ;
  assign n335 = n330 & n334 ;
  assign n336 = n335 ^ n297 ;
  assign n363 = n362 ^ n336 ;
  assign n364 = n362 ^ x67 ;
  assign n365 = n363 & n364 ;
  assign n366 = n365 ^ n317 ;
  assign n369 = ~n333 & n366 ;
  assign n370 = n369 ^ x68 ;
  assign n371 = ~n324 & n370 ;
  assign n372 = n322 & ~n371 ;
  assign n373 = n320 & ~n372 ;
  assign n269 = n189 & ~n268 ;
  assign n270 = n233 & n269 ;
  assign n374 = n373 ^ n270 ;
  assign n375 = ~n184 & n374 ;
  assign n414 = n374 ^ x70 ;
  assign n387 = x64 & n330 ;
  assign n383 = ~x58 & x64 ;
  assign n384 = n383 ^ x65 ;
  assign n385 = n372 & n384 ;
  assign n386 = n385 ^ x59 ;
  assign n388 = n387 ^ n386 ;
  assign n389 = n388 ^ x66 ;
  assign n395 = x58 & x65 ;
  assign n390 = x65 ^ x57 ;
  assign n391 = x64 ^ x58 ;
  assign n392 = n391 ^ x65 ;
  assign n393 = n392 ^ n372 ;
  assign n394 = ~n390 & n393 ;
  assign n396 = n395 ^ n394 ;
  assign n399 = x64 & n396 ;
  assign n400 = n399 ^ n395 ;
  assign n401 = n400 ^ x65 ;
  assign n402 = n401 ^ n388 ;
  assign n403 = ~n389 & n402 ;
  assign n404 = n403 ^ x66 ;
  assign n379 = n359 ^ x66 ;
  assign n380 = n372 & n379 ;
  assign n381 = n380 ^ n346 ;
  assign n405 = n404 ^ n381 ;
  assign n406 = n404 ^ x67 ;
  assign n407 = n405 & n406 ;
  assign n408 = n407 ^ x67 ;
  assign n377 = n364 & n372 ;
  assign n378 = n377 ^ n336 ;
  assign n409 = n408 ^ n378 ;
  assign n410 = n408 ^ x68 ;
  assign n411 = n409 & n410 ;
  assign n412 = n411 ^ x68 ;
  assign n413 = n412 ^ x69 ;
  assign n415 = n366 & n372 ;
  assign n416 = n415 ^ n332 ;
  assign n417 = n416 ^ n412 ;
  assign n418 = n413 & n417 ;
  assign n419 = n418 ^ x69 ;
  assign n420 = n419 ^ x70 ;
  assign n421 = ~n414 & n420 ;
  assign n422 = n421 ^ x70 ;
  assign n423 = n185 & ~n422 ;
  assign n376 = n374 ^ x71 ;
  assign n474 = x70 & n419 ;
  assign n447 = x57 & x65 ;
  assign n444 = x65 ^ x56 ;
  assign n440 = x64 ^ x57 ;
  assign n441 = n440 ^ x65 ;
  assign n445 = n441 ^ n423 ;
  assign n446 = ~n444 & n445 ;
  assign n448 = n447 ^ n446 ;
  assign n449 = x64 & n448 ;
  assign n450 = n449 ^ n447 ;
  assign n451 = n450 ^ x65 ;
  assign n437 = x64 & n423 ;
  assign n438 = ~x57 & n437 ;
  assign n434 = x65 & n423 ;
  assign n433 = x64 & n372 ;
  assign n435 = n434 ^ n433 ;
  assign n436 = n435 ^ x58 ;
  assign n439 = n438 ^ n436 ;
  assign n452 = n451 ^ n439 ;
  assign n453 = n451 ^ x66 ;
  assign n454 = n452 & n453 ;
  assign n455 = n454 ^ x66 ;
  assign n430 = n401 ^ x66 ;
  assign n431 = n423 & n430 ;
  assign n432 = n431 ^ n388 ;
  assign n456 = n455 ^ n432 ;
  assign n457 = n455 ^ x67 ;
  assign n458 = n456 & n457 ;
  assign n459 = n458 ^ x67 ;
  assign n428 = n406 & n423 ;
  assign n429 = n428 ^ n381 ;
  assign n460 = n459 ^ n429 ;
  assign n461 = n459 ^ x68 ;
  assign n462 = n460 & n461 ;
  assign n463 = n462 ^ x68 ;
  assign n426 = n410 & n423 ;
  assign n427 = n426 ^ n378 ;
  assign n464 = n463 ^ n427 ;
  assign n465 = n463 ^ x69 ;
  assign n466 = n464 & n465 ;
  assign n467 = n466 ^ x69 ;
  assign n424 = n413 & n423 ;
  assign n425 = n424 ^ n416 ;
  assign n468 = n467 ^ n425 ;
  assign n469 = n467 ^ x70 ;
  assign n470 = n468 & n469 ;
  assign n471 = n470 ^ x70 ;
  assign n475 = n474 ^ n471 ;
  assign n476 = n374 & ~n475 ;
  assign n477 = n476 ^ n471 ;
  assign n478 = n376 & ~n477 ;
  assign n479 = n478 ^ n471 ;
  assign n480 = n184 & ~n479 ;
  assign n481 = n374 & ~n480 ;
  assign n482 = ~n423 & n481 ;
  assign n483 = n482 ^ n270 ;
  assign n484 = n483 ^ x72 ;
  assign n485 = n183 & ~n484 ;
  assign n486 = n469 & n480 ;
  assign n487 = n486 ^ n425 ;
  assign n488 = n487 ^ x71 ;
  assign n510 = x56 & x65 ;
  assign n505 = x65 ^ x55 ;
  assign n506 = x64 ^ x56 ;
  assign n507 = n506 ^ x65 ;
  assign n508 = n507 ^ n480 ;
  assign n509 = ~n505 & n508 ;
  assign n511 = n510 ^ n509 ;
  assign n514 = x64 & n511 ;
  assign n515 = n514 ^ n510 ;
  assign n516 = n515 ^ x65 ;
  assign n503 = n437 ^ x57 ;
  assign n500 = ~x56 & x64 ;
  assign n501 = n500 ^ x65 ;
  assign n502 = n480 & n501 ;
  assign n504 = n503 ^ n502 ;
  assign n517 = n516 ^ n504 ;
  assign n518 = n516 ^ x66 ;
  assign n519 = n517 & n518 ;
  assign n520 = n519 ^ x66 ;
  assign n495 = n453 & n480 ;
  assign n496 = n495 ^ n439 ;
  assign n521 = n520 ^ n496 ;
  assign n522 = n520 ^ x67 ;
  assign n523 = n521 & n522 ;
  assign n524 = n523 ^ x67 ;
  assign n493 = n457 & n480 ;
  assign n494 = n493 ^ n432 ;
  assign n525 = n524 ^ n494 ;
  assign n526 = n524 ^ x68 ;
  assign n527 = n525 & n526 ;
  assign n528 = n527 ^ x68 ;
  assign n491 = n461 & n480 ;
  assign n492 = n491 ^ n429 ;
  assign n529 = n528 ^ n492 ;
  assign n530 = n528 ^ x69 ;
  assign n531 = n529 & n530 ;
  assign n532 = n531 ^ x69 ;
  assign n489 = n465 & n480 ;
  assign n490 = n489 ^ n427 ;
  assign n533 = n532 ^ n490 ;
  assign n536 = n490 ^ x70 ;
  assign n537 = n533 & ~n536 ;
  assign n534 = x71 ^ x70 ;
  assign n538 = n537 ^ n534 ;
  assign n541 = ~n488 & n538 ;
  assign n542 = n541 ^ x71 ;
  assign n543 = n485 & ~n542 ;
  assign n544 = n375 & ~n543 ;
  assign n545 = n184 & n483 ;
  assign n546 = n545 ^ n543 ;
  assign n603 = n538 & n546 ;
  assign n604 = n603 ^ n487 ;
  assign n547 = n532 ^ x70 ;
  assign n548 = n546 & n547 ;
  assign n549 = n548 ^ n490 ;
  assign n550 = n549 ^ x71 ;
  assign n554 = n549 ^ x70 ;
  assign n551 = n530 & n546 ;
  assign n552 = n551 ^ n492 ;
  assign n553 = n552 ^ n549 ;
  assign n555 = n554 ^ n553 ;
  assign n566 = x64 & n546 ;
  assign n567 = ~x55 & n566 ;
  assign n563 = x64 & n480 ;
  assign n562 = x65 & n546 ;
  assign n564 = n563 ^ n562 ;
  assign n565 = n564 ^ x56 ;
  assign n568 = n567 ^ n565 ;
  assign n569 = n568 ^ x66 ;
  assign n577 = x55 & x65 ;
  assign n574 = x65 ^ x54 ;
  assign n570 = x64 ^ x55 ;
  assign n571 = n570 ^ x65 ;
  assign n575 = n571 ^ n546 ;
  assign n576 = ~n574 & n575 ;
  assign n578 = n577 ^ n576 ;
  assign n579 = x64 & n578 ;
  assign n580 = n579 ^ n577 ;
  assign n581 = n580 ^ x65 ;
  assign n582 = n581 ^ n568 ;
  assign n583 = ~n569 & n582 ;
  assign n584 = n583 ^ x66 ;
  assign n560 = n518 & n546 ;
  assign n561 = n560 ^ n504 ;
  assign n585 = n584 ^ n561 ;
  assign n586 = n584 ^ x67 ;
  assign n587 = n585 & n586 ;
  assign n588 = n587 ^ x67 ;
  assign n558 = n522 & n546 ;
  assign n559 = n558 ^ n496 ;
  assign n589 = n588 ^ n559 ;
  assign n590 = n588 ^ x68 ;
  assign n591 = n589 & n590 ;
  assign n592 = n591 ^ x68 ;
  assign n556 = n526 & n546 ;
  assign n557 = n556 ^ n494 ;
  assign n593 = n592 ^ n557 ;
  assign n594 = n592 ^ x69 ;
  assign n595 = n593 & n594 ;
  assign n596 = n595 ^ x69 ;
  assign n647 = n596 ^ x70 ;
  assign n599 = ~n555 & n647 ;
  assign n600 = n599 ^ n554 ;
  assign n601 = ~n550 & n600 ;
  assign n602 = n601 ^ x71 ;
  assign n605 = n604 ^ n602 ;
  assign n606 = x73 ^ x72 ;
  assign n607 = n606 ^ n544 ;
  assign n608 = n607 ^ n604 ;
  assign n609 = n605 & ~n608 ;
  assign n613 = n608 ^ x73 ;
  assign n614 = n613 ^ n605 ;
  assign n615 = n614 ^ n602 ;
  assign n616 = ~n606 & n615 ;
  assign n619 = n607 & n616 ;
  assign n620 = n619 ^ n615 ;
  assign n621 = n620 ^ n606 ;
  assign n622 = n609 & ~n621 ;
  assign n623 = n622 ^ n619 ;
  assign n624 = n623 ^ n616 ;
  assign n625 = n624 ^ n607 ;
  assign n626 = n182 & ~n625 ;
  assign n627 = n544 & ~n626 ;
  assign n628 = n627 ^ n270 ;
  assign n629 = n628 ^ x74 ;
  assign n634 = n628 ^ x73 ;
  assign n630 = n602 ^ x72 ;
  assign n631 = n626 & n630 ;
  assign n632 = n631 ^ n604 ;
  assign n633 = n632 ^ n628 ;
  assign n635 = n634 ^ n633 ;
  assign n666 = x54 & x65 ;
  assign n663 = x65 ^ x53 ;
  assign n659 = x64 ^ x54 ;
  assign n660 = n659 ^ x65 ;
  assign n664 = n660 ^ n626 ;
  assign n665 = ~n663 & n664 ;
  assign n667 = n666 ^ n665 ;
  assign n668 = x64 & n667 ;
  assign n669 = n668 ^ n666 ;
  assign n670 = n669 ^ x65 ;
  assign n671 = n670 ^ x66 ;
  assign n676 = n566 ^ x55 ;
  assign n673 = ~x54 & x64 ;
  assign n674 = n673 ^ x65 ;
  assign n675 = n626 & n674 ;
  assign n677 = n676 ^ n675 ;
  assign n678 = n677 ^ n670 ;
  assign n679 = n671 & n678 ;
  assign n680 = n679 ^ x66 ;
  assign n656 = n581 ^ x66 ;
  assign n657 = n626 & n656 ;
  assign n658 = n657 ^ n568 ;
  assign n681 = n680 ^ n658 ;
  assign n682 = n680 ^ x67 ;
  assign n683 = n681 & n682 ;
  assign n684 = n683 ^ x67 ;
  assign n654 = n586 & n626 ;
  assign n655 = n654 ^ n561 ;
  assign n685 = n684 ^ n655 ;
  assign n686 = n684 ^ x68 ;
  assign n687 = n685 & n686 ;
  assign n688 = n687 ^ x68 ;
  assign n652 = n590 & n626 ;
  assign n653 = n652 ^ n559 ;
  assign n689 = n688 ^ n653 ;
  assign n690 = n688 ^ x69 ;
  assign n691 = n689 & n690 ;
  assign n692 = n691 ^ x69 ;
  assign n650 = n594 & n626 ;
  assign n651 = n650 ^ n557 ;
  assign n693 = n692 ^ n651 ;
  assign n694 = n692 ^ x70 ;
  assign n695 = n693 & n694 ;
  assign n696 = n695 ^ x70 ;
  assign n648 = n626 & n647 ;
  assign n649 = n648 ^ n552 ;
  assign n697 = n696 ^ n649 ;
  assign n698 = n696 ^ x71 ;
  assign n699 = n697 & n698 ;
  assign n700 = n699 ^ x71 ;
  assign n641 = n596 ^ x71 ;
  assign n636 = n552 ^ x71 ;
  assign n642 = n641 ^ n636 ;
  assign n643 = ~n642 & ~n647 ;
  assign n644 = n643 ^ n636 ;
  assign n645 = n626 & ~n644 ;
  assign n646 = n645 ^ n549 ;
  assign n701 = n700 ^ n646 ;
  assign n702 = n700 ^ x72 ;
  assign n703 = n701 & n702 ;
  assign n704 = n703 ^ x72 ;
  assign n716 = n704 ^ x73 ;
  assign n707 = ~n635 & n716 ;
  assign n708 = n707 ^ n634 ;
  assign n709 = ~n629 & n708 ;
  assign n710 = n709 ^ x74 ;
  assign n711 = n181 & ~n710 ;
  assign n712 = n711 ^ n270 ;
  assign n713 = n628 & ~n712 ;
  assign n714 = n180 & n713 ;
  assign n715 = x75 & n714 ;
  assign n733 = ~x52 & x64 ;
  assign n738 = n711 ^ x53 ;
  assign n739 = n733 & ~n738 ;
  assign n735 = x64 & n711 ;
  assign n734 = n733 ^ x53 ;
  assign n736 = n735 ^ n734 ;
  assign n737 = x65 & ~n736 ;
  assign n740 = n739 ^ n737 ;
  assign n741 = n740 ^ x66 ;
  assign n747 = x64 & n626 ;
  assign n743 = ~x53 & x64 ;
  assign n744 = n743 ^ x65 ;
  assign n745 = n711 & n744 ;
  assign n746 = n745 ^ x54 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = n748 ^ n740 ;
  assign n750 = n741 & n749 ;
  assign n751 = n750 ^ x66 ;
  assign n731 = n671 & n711 ;
  assign n732 = n731 ^ n677 ;
  assign n752 = n751 ^ n732 ;
  assign n753 = n751 ^ x67 ;
  assign n754 = n752 & n753 ;
  assign n755 = n754 ^ x67 ;
  assign n729 = n682 & n711 ;
  assign n730 = n729 ^ n658 ;
  assign n756 = n755 ^ n730 ;
  assign n757 = n755 ^ x68 ;
  assign n758 = n756 & n757 ;
  assign n759 = n758 ^ x68 ;
  assign n727 = n686 & n711 ;
  assign n728 = n727 ^ n655 ;
  assign n760 = n759 ^ n728 ;
  assign n761 = n759 ^ x69 ;
  assign n762 = n760 & n761 ;
  assign n763 = n762 ^ x69 ;
  assign n725 = n690 & n711 ;
  assign n726 = n725 ^ n653 ;
  assign n764 = n763 ^ n726 ;
  assign n765 = n763 ^ x70 ;
  assign n766 = n764 & n765 ;
  assign n767 = n766 ^ x70 ;
  assign n723 = n694 & n711 ;
  assign n724 = n723 ^ n651 ;
  assign n768 = n767 ^ n724 ;
  assign n769 = n767 ^ x71 ;
  assign n770 = n768 & n769 ;
  assign n771 = n770 ^ x71 ;
  assign n721 = n698 & n711 ;
  assign n722 = n721 ^ n649 ;
  assign n772 = n771 ^ n722 ;
  assign n773 = n771 ^ x72 ;
  assign n774 = n772 & n773 ;
  assign n775 = n774 ^ x72 ;
  assign n719 = n702 & n711 ;
  assign n720 = n719 ^ n646 ;
  assign n776 = n775 ^ n720 ;
  assign n777 = n775 ^ x73 ;
  assign n778 = n776 & n777 ;
  assign n779 = n778 ^ x73 ;
  assign n717 = n711 & n716 ;
  assign n718 = n717 ^ n632 ;
  assign n780 = n779 ^ n718 ;
  assign n781 = n779 ^ x74 ;
  assign n782 = n780 & n781 ;
  assign n783 = n782 ^ x74 ;
  assign n784 = n715 & n783 ;
  assign n785 = n784 ^ n714 ;
  assign n786 = n785 ^ n713 ;
  assign n787 = ~n178 & n786 ;
  assign n811 = ~x51 & x64 ;
  assign n812 = n811 ^ x65 ;
  assign n814 = n811 ^ x52 ;
  assign n788 = n713 ^ x75 ;
  assign n789 = n783 ^ x75 ;
  assign n790 = ~n788 & n789 ;
  assign n791 = n790 ^ x75 ;
  assign n792 = n180 & ~n791 ;
  assign n813 = x64 & n792 ;
  assign n815 = n814 ^ n813 ;
  assign n816 = n812 & n815 ;
  assign n817 = n816 ^ x65 ;
  assign n818 = n817 ^ x66 ;
  assign n821 = n735 ^ x53 ;
  assign n819 = n733 ^ x65 ;
  assign n820 = n792 & n819 ;
  assign n822 = n821 ^ n820 ;
  assign n823 = n822 ^ n817 ;
  assign n824 = n818 & n823 ;
  assign n825 = n824 ^ x66 ;
  assign n809 = n741 & n792 ;
  assign n810 = n809 ^ n748 ;
  assign n826 = n825 ^ n810 ;
  assign n827 = n825 ^ x67 ;
  assign n828 = n826 & n827 ;
  assign n829 = n828 ^ x67 ;
  assign n807 = n753 & n792 ;
  assign n808 = n807 ^ n732 ;
  assign n830 = n829 ^ n808 ;
  assign n831 = n829 ^ x68 ;
  assign n832 = n830 & n831 ;
  assign n833 = n832 ^ x68 ;
  assign n805 = n757 & n792 ;
  assign n806 = n805 ^ n730 ;
  assign n834 = n833 ^ n806 ;
  assign n835 = n833 ^ x69 ;
  assign n836 = n834 & n835 ;
  assign n837 = n836 ^ x69 ;
  assign n803 = n761 & n792 ;
  assign n804 = n803 ^ n728 ;
  assign n838 = n837 ^ n804 ;
  assign n839 = n837 ^ x70 ;
  assign n840 = n838 & n839 ;
  assign n841 = n840 ^ x70 ;
  assign n801 = n765 & n792 ;
  assign n802 = n801 ^ n726 ;
  assign n842 = n841 ^ n802 ;
  assign n843 = n841 ^ x71 ;
  assign n844 = n842 & n843 ;
  assign n845 = n844 ^ x71 ;
  assign n799 = n769 & n792 ;
  assign n800 = n799 ^ n724 ;
  assign n846 = n845 ^ n800 ;
  assign n847 = n845 ^ x72 ;
  assign n848 = n846 & n847 ;
  assign n849 = n848 ^ x72 ;
  assign n797 = n773 & n792 ;
  assign n798 = n797 ^ n722 ;
  assign n850 = n849 ^ n798 ;
  assign n851 = n849 ^ x73 ;
  assign n852 = n850 & n851 ;
  assign n853 = n852 ^ x73 ;
  assign n795 = n777 & n792 ;
  assign n796 = n795 ^ n720 ;
  assign n854 = n853 ^ n796 ;
  assign n855 = n853 ^ x74 ;
  assign n856 = n854 & n855 ;
  assign n857 = n856 ^ x74 ;
  assign n793 = n781 & n792 ;
  assign n794 = n793 ^ n718 ;
  assign n858 = n857 ^ n794 ;
  assign n859 = x76 ^ x75 ;
  assign n860 = n859 ^ n786 ;
  assign n861 = n860 ^ n857 ;
  assign n862 = n858 & n861 ;
  assign n868 = n861 ^ x76 ;
  assign n869 = n868 ^ n858 ;
  assign n870 = n869 ^ n794 ;
  assign n871 = ~n859 & n870 ;
  assign n872 = n860 & n871 ;
  assign n873 = n872 ^ n870 ;
  assign n874 = n873 ^ n859 ;
  assign n875 = n862 & ~n874 ;
  assign n876 = n875 ^ n872 ;
  assign n877 = n876 ^ n871 ;
  assign n878 = n877 ^ n860 ;
  assign n879 = n179 & ~n878 ;
  assign n880 = n786 & ~n879 ;
  assign n881 = n880 ^ n270 ;
  assign n882 = n881 ^ x77 ;
  assign n887 = n881 ^ x76 ;
  assign n883 = n857 ^ x75 ;
  assign n884 = n879 & n883 ;
  assign n885 = n884 ^ n794 ;
  assign n886 = n885 ^ n881 ;
  assign n888 = n887 ^ n886 ;
  assign n908 = n813 ^ x52 ;
  assign n907 = n812 & n879 ;
  assign n909 = n908 ^ n907 ;
  assign n910 = n909 ^ x66 ;
  assign n914 = x64 ^ x51 ;
  assign n915 = n914 ^ x65 ;
  assign n912 = x64 & n879 ;
  assign n911 = ~x64 & x65 ;
  assign n913 = n912 ^ n911 ;
  assign n916 = n915 ^ n913 ;
  assign n917 = ~x50 & x64 ;
  assign n918 = n917 ^ x65 ;
  assign n919 = n916 & n918 ;
  assign n920 = n919 ^ x65 ;
  assign n921 = n920 ^ n909 ;
  assign n922 = ~n910 & n921 ;
  assign n923 = n922 ^ x66 ;
  assign n905 = n818 & n879 ;
  assign n906 = n905 ^ n822 ;
  assign n924 = n923 ^ n906 ;
  assign n925 = n923 ^ x67 ;
  assign n926 = n924 & n925 ;
  assign n927 = n926 ^ x67 ;
  assign n903 = n827 & n879 ;
  assign n904 = n903 ^ n810 ;
  assign n928 = n927 ^ n904 ;
  assign n929 = n927 ^ x68 ;
  assign n930 = n928 & n929 ;
  assign n931 = n930 ^ x68 ;
  assign n901 = n831 & n879 ;
  assign n902 = n901 ^ n808 ;
  assign n932 = n931 ^ n902 ;
  assign n933 = n931 ^ x69 ;
  assign n934 = n932 & n933 ;
  assign n935 = n934 ^ x69 ;
  assign n899 = n835 & n879 ;
  assign n900 = n899 ^ n806 ;
  assign n936 = n935 ^ n900 ;
  assign n937 = n935 ^ x70 ;
  assign n938 = n936 & n937 ;
  assign n939 = n938 ^ x70 ;
  assign n897 = n839 & n879 ;
  assign n898 = n897 ^ n804 ;
  assign n940 = n939 ^ n898 ;
  assign n941 = n939 ^ x71 ;
  assign n942 = n940 & n941 ;
  assign n943 = n942 ^ x71 ;
  assign n895 = n843 & n879 ;
  assign n896 = n895 ^ n802 ;
  assign n944 = n943 ^ n896 ;
  assign n945 = n943 ^ x72 ;
  assign n946 = n944 & n945 ;
  assign n947 = n946 ^ x72 ;
  assign n893 = n847 & n879 ;
  assign n894 = n893 ^ n800 ;
  assign n948 = n947 ^ n894 ;
  assign n949 = n947 ^ x73 ;
  assign n950 = n948 & n949 ;
  assign n951 = n950 ^ x73 ;
  assign n891 = n851 & n879 ;
  assign n892 = n891 ^ n798 ;
  assign n952 = n951 ^ n892 ;
  assign n953 = n951 ^ x74 ;
  assign n954 = n952 & n953 ;
  assign n955 = n954 ^ x74 ;
  assign n889 = n855 & n879 ;
  assign n890 = n889 ^ n796 ;
  assign n956 = n955 ^ n890 ;
  assign n957 = n955 ^ x75 ;
  assign n958 = n956 & n957 ;
  assign n959 = n958 ^ x75 ;
  assign n971 = n959 ^ x76 ;
  assign n962 = ~n888 & n971 ;
  assign n963 = n962 ^ n887 ;
  assign n964 = ~n882 & n963 ;
  assign n965 = n964 ^ x77 ;
  assign n966 = n178 & ~n965 ;
  assign n967 = n880 & ~n966 ;
  assign n968 = n967 ^ n270 ;
  assign n969 = n968 ^ x78 ;
  assign n970 = n177 & ~n969 ;
  assign n972 = n966 & n971 ;
  assign n973 = n972 ^ n885 ;
  assign n974 = n973 ^ x77 ;
  assign n1007 = n918 & n966 ;
  assign n1006 = n912 ^ x51 ;
  assign n1008 = n1007 ^ n1006 ;
  assign n996 = ~x49 & x64 ;
  assign n997 = n996 ^ n966 ;
  assign n998 = n997 ^ x50 ;
  assign n1002 = n996 ^ x65 ;
  assign n1003 = ~n998 & ~n1002 ;
  assign n1001 = ~n911 & n966 ;
  assign n1004 = n1003 ^ n1001 ;
  assign n1005 = n1004 ^ x50 ;
  assign n1009 = n1008 ^ n1005 ;
  assign n1010 = n1008 ^ x66 ;
  assign n1011 = ~n1009 & ~n1010 ;
  assign n1012 = n1011 ^ x66 ;
  assign n993 = n920 ^ x66 ;
  assign n994 = n966 & n993 ;
  assign n995 = n994 ^ n909 ;
  assign n1013 = n1012 ^ n995 ;
  assign n1014 = n1012 ^ x67 ;
  assign n1015 = n1013 & n1014 ;
  assign n1016 = n1015 ^ x67 ;
  assign n991 = n925 & n966 ;
  assign n992 = n991 ^ n906 ;
  assign n1017 = n1016 ^ n992 ;
  assign n1018 = n1016 ^ x68 ;
  assign n1019 = n1017 & n1018 ;
  assign n1020 = n1019 ^ x68 ;
  assign n989 = n929 & n966 ;
  assign n990 = n989 ^ n904 ;
  assign n1021 = n1020 ^ n990 ;
  assign n1022 = n1020 ^ x69 ;
  assign n1023 = n1021 & n1022 ;
  assign n1024 = n1023 ^ x69 ;
  assign n987 = n933 & n966 ;
  assign n988 = n987 ^ n902 ;
  assign n1025 = n1024 ^ n988 ;
  assign n1026 = n1024 ^ x70 ;
  assign n1027 = n1025 & n1026 ;
  assign n1028 = n1027 ^ x70 ;
  assign n985 = n937 & n966 ;
  assign n986 = n985 ^ n900 ;
  assign n1029 = n1028 ^ n986 ;
  assign n1030 = n1028 ^ x71 ;
  assign n1031 = n1029 & n1030 ;
  assign n1032 = n1031 ^ x71 ;
  assign n983 = n941 & n966 ;
  assign n984 = n983 ^ n898 ;
  assign n1033 = n1032 ^ n984 ;
  assign n1034 = n1032 ^ x72 ;
  assign n1035 = n1033 & n1034 ;
  assign n1036 = n1035 ^ x72 ;
  assign n981 = n945 & n966 ;
  assign n982 = n981 ^ n896 ;
  assign n1037 = n1036 ^ n982 ;
  assign n1038 = n1036 ^ x73 ;
  assign n1039 = n1037 & n1038 ;
  assign n1040 = n1039 ^ x73 ;
  assign n979 = n949 & n966 ;
  assign n980 = n979 ^ n894 ;
  assign n1041 = n1040 ^ n980 ;
  assign n1042 = n1040 ^ x74 ;
  assign n1043 = n1041 & n1042 ;
  assign n1044 = n1043 ^ x74 ;
  assign n977 = n953 & n966 ;
  assign n978 = n977 ^ n892 ;
  assign n1045 = n1044 ^ n978 ;
  assign n1046 = n1044 ^ x75 ;
  assign n1047 = n1045 & n1046 ;
  assign n1048 = n1047 ^ x75 ;
  assign n975 = n957 & n966 ;
  assign n976 = n975 ^ n890 ;
  assign n1049 = n1048 ^ n976 ;
  assign n1052 = n976 ^ x76 ;
  assign n1053 = n1049 & ~n1052 ;
  assign n1050 = x77 ^ x76 ;
  assign n1054 = n1053 ^ n1050 ;
  assign n1057 = ~n974 & n1054 ;
  assign n1058 = n1057 ^ x77 ;
  assign n1059 = n970 & ~n1058 ;
  assign n1060 = n787 & ~n1059 ;
  assign n1061 = ~n175 & n1060 ;
  assign n1062 = n1060 ^ n270 ;
  assign n1063 = n1062 ^ x79 ;
  assign n1096 = ~x48 & x64 ;
  assign n1097 = n1096 ^ x65 ;
  assign n1099 = n1096 ^ x49 ;
  assign n1064 = n178 & n968 ;
  assign n1065 = n1064 ^ n1059 ;
  assign n1098 = x64 & n1065 ;
  assign n1100 = n1099 ^ n1098 ;
  assign n1101 = n1097 & n1100 ;
  assign n1102 = n1101 ^ x65 ;
  assign n1093 = n1002 & n1065 ;
  assign n1092 = x64 & n966 ;
  assign n1094 = n1093 ^ n1092 ;
  assign n1095 = n1094 ^ x50 ;
  assign n1103 = n1102 ^ n1095 ;
  assign n1104 = n1102 ^ x66 ;
  assign n1105 = n1103 & n1104 ;
  assign n1106 = n1105 ^ x66 ;
  assign n1089 = n1005 ^ x66 ;
  assign n1090 = n1065 & ~n1089 ;
  assign n1091 = n1090 ^ n1008 ;
  assign n1107 = n1106 ^ n1091 ;
  assign n1108 = n1106 ^ x67 ;
  assign n1109 = n1107 & n1108 ;
  assign n1110 = n1109 ^ x67 ;
  assign n1087 = n1014 & n1065 ;
  assign n1088 = n1087 ^ n995 ;
  assign n1111 = n1110 ^ n1088 ;
  assign n1112 = n1110 ^ x68 ;
  assign n1113 = n1111 & n1112 ;
  assign n1114 = n1113 ^ x68 ;
  assign n1085 = n1018 & n1065 ;
  assign n1086 = n1085 ^ n992 ;
  assign n1115 = n1114 ^ n1086 ;
  assign n1116 = n1114 ^ x69 ;
  assign n1117 = n1115 & n1116 ;
  assign n1118 = n1117 ^ x69 ;
  assign n1083 = n1022 & n1065 ;
  assign n1084 = n1083 ^ n990 ;
  assign n1119 = n1118 ^ n1084 ;
  assign n1120 = n1118 ^ x70 ;
  assign n1121 = n1119 & n1120 ;
  assign n1122 = n1121 ^ x70 ;
  assign n1081 = n1026 & n1065 ;
  assign n1082 = n1081 ^ n988 ;
  assign n1123 = n1122 ^ n1082 ;
  assign n1124 = n1122 ^ x71 ;
  assign n1125 = n1123 & n1124 ;
  assign n1126 = n1125 ^ x71 ;
  assign n1079 = n1030 & n1065 ;
  assign n1080 = n1079 ^ n986 ;
  assign n1127 = n1126 ^ n1080 ;
  assign n1128 = n1126 ^ x72 ;
  assign n1129 = n1127 & n1128 ;
  assign n1130 = n1129 ^ x72 ;
  assign n1077 = n1034 & n1065 ;
  assign n1078 = n1077 ^ n984 ;
  assign n1131 = n1130 ^ n1078 ;
  assign n1132 = n1130 ^ x73 ;
  assign n1133 = n1131 & n1132 ;
  assign n1134 = n1133 ^ x73 ;
  assign n1075 = n1038 & n1065 ;
  assign n1076 = n1075 ^ n982 ;
  assign n1135 = n1134 ^ n1076 ;
  assign n1136 = n1134 ^ x74 ;
  assign n1137 = n1135 & n1136 ;
  assign n1138 = n1137 ^ x74 ;
  assign n1073 = n1042 & n1065 ;
  assign n1074 = n1073 ^ n980 ;
  assign n1139 = n1138 ^ n1074 ;
  assign n1140 = n1138 ^ x75 ;
  assign n1141 = n1139 & n1140 ;
  assign n1142 = n1141 ^ x75 ;
  assign n1071 = n1046 & n1065 ;
  assign n1072 = n1071 ^ n978 ;
  assign n1143 = n1142 ^ n1072 ;
  assign n1144 = n1142 ^ x76 ;
  assign n1145 = n1143 & n1144 ;
  assign n1146 = n1145 ^ x76 ;
  assign n1068 = n1048 ^ x76 ;
  assign n1069 = n1065 & n1068 ;
  assign n1070 = n1069 ^ n976 ;
  assign n1147 = n1146 ^ n1070 ;
  assign n1148 = n1146 ^ x77 ;
  assign n1149 = n1147 & n1148 ;
  assign n1150 = n1149 ^ x77 ;
  assign n1066 = n1054 & n1065 ;
  assign n1067 = n1066 ^ n973 ;
  assign n1151 = n1150 ^ n1067 ;
  assign n1154 = n1067 ^ x78 ;
  assign n1155 = n1151 & ~n1154 ;
  assign n1152 = x79 ^ x78 ;
  assign n1156 = n1155 ^ n1152 ;
  assign n1157 = ~n1063 & n1156 ;
  assign n1158 = n1157 ^ x79 ;
  assign n1159 = n176 & ~n1158 ;
  assign n1160 = n1060 & ~n1159 ;
  assign n1161 = n1160 ^ n270 ;
  assign n1162 = n1161 ^ x80 ;
  assign n1167 = n1161 ^ x79 ;
  assign n1163 = n1150 ^ x78 ;
  assign n1164 = n1159 & n1163 ;
  assign n1165 = n1164 ^ n1067 ;
  assign n1166 = n1165 ^ n1161 ;
  assign n1168 = n1167 ^ n1166 ;
  assign n1191 = n1104 & n1159 ;
  assign n1192 = n1191 ^ n1095 ;
  assign n1193 = n1192 ^ x67 ;
  assign n1204 = x48 & x65 ;
  assign n1201 = x65 ^ x47 ;
  assign n1197 = x64 ^ x48 ;
  assign n1198 = n1197 ^ x65 ;
  assign n1202 = n1198 ^ n1159 ;
  assign n1203 = ~n1201 & n1202 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1206 = x64 & n1205 ;
  assign n1207 = n1206 ^ n1204 ;
  assign n1208 = n1207 ^ x65 ;
  assign n1195 = n1097 & n1159 ;
  assign n1194 = n1098 ^ x49 ;
  assign n1196 = n1195 ^ n1194 ;
  assign n1209 = n1208 ^ n1196 ;
  assign n1210 = n1208 ^ x66 ;
  assign n1211 = n1209 & n1210 ;
  assign n1212 = n1211 ^ x66 ;
  assign n1213 = n1212 ^ n1192 ;
  assign n1214 = ~n1193 & n1213 ;
  assign n1215 = n1214 ^ x67 ;
  assign n1189 = n1108 & n1159 ;
  assign n1190 = n1189 ^ n1091 ;
  assign n1216 = n1215 ^ n1190 ;
  assign n1217 = n1215 ^ x68 ;
  assign n1218 = n1216 & n1217 ;
  assign n1219 = n1218 ^ x68 ;
  assign n1187 = n1112 & n1159 ;
  assign n1188 = n1187 ^ n1088 ;
  assign n1220 = n1219 ^ n1188 ;
  assign n1221 = n1219 ^ x69 ;
  assign n1222 = n1220 & n1221 ;
  assign n1223 = n1222 ^ x69 ;
  assign n1185 = n1116 & n1159 ;
  assign n1186 = n1185 ^ n1086 ;
  assign n1224 = n1223 ^ n1186 ;
  assign n1225 = n1223 ^ x70 ;
  assign n1226 = n1224 & n1225 ;
  assign n1227 = n1226 ^ x70 ;
  assign n1183 = n1120 & n1159 ;
  assign n1184 = n1183 ^ n1084 ;
  assign n1228 = n1227 ^ n1184 ;
  assign n1229 = n1227 ^ x71 ;
  assign n1230 = n1228 & n1229 ;
  assign n1231 = n1230 ^ x71 ;
  assign n1181 = n1124 & n1159 ;
  assign n1182 = n1181 ^ n1082 ;
  assign n1232 = n1231 ^ n1182 ;
  assign n1233 = n1231 ^ x72 ;
  assign n1234 = n1232 & n1233 ;
  assign n1235 = n1234 ^ x72 ;
  assign n1179 = n1128 & n1159 ;
  assign n1180 = n1179 ^ n1080 ;
  assign n1236 = n1235 ^ n1180 ;
  assign n1237 = n1235 ^ x73 ;
  assign n1238 = n1236 & n1237 ;
  assign n1239 = n1238 ^ x73 ;
  assign n1177 = n1132 & n1159 ;
  assign n1178 = n1177 ^ n1078 ;
  assign n1240 = n1239 ^ n1178 ;
  assign n1241 = n1239 ^ x74 ;
  assign n1242 = n1240 & n1241 ;
  assign n1243 = n1242 ^ x74 ;
  assign n1175 = n1136 & n1159 ;
  assign n1176 = n1175 ^ n1076 ;
  assign n1244 = n1243 ^ n1176 ;
  assign n1245 = n1243 ^ x75 ;
  assign n1246 = n1244 & n1245 ;
  assign n1247 = n1246 ^ x75 ;
  assign n1173 = n1140 & n1159 ;
  assign n1174 = n1173 ^ n1074 ;
  assign n1248 = n1247 ^ n1174 ;
  assign n1249 = n1247 ^ x76 ;
  assign n1250 = n1248 & n1249 ;
  assign n1251 = n1250 ^ x76 ;
  assign n1171 = n1144 & n1159 ;
  assign n1172 = n1171 ^ n1072 ;
  assign n1252 = n1251 ^ n1172 ;
  assign n1253 = n1251 ^ x77 ;
  assign n1254 = n1252 & n1253 ;
  assign n1255 = n1254 ^ x77 ;
  assign n1169 = n1148 & n1159 ;
  assign n1170 = n1169 ^ n1070 ;
  assign n1256 = n1255 ^ n1170 ;
  assign n1257 = n1255 ^ x78 ;
  assign n1258 = n1256 & n1257 ;
  assign n1259 = n1258 ^ x78 ;
  assign n1260 = n1259 ^ n1161 ;
  assign n1261 = n1260 ^ n1167 ;
  assign n1262 = ~n1168 & n1261 ;
  assign n1263 = n1262 ^ n1167 ;
  assign n1264 = ~n1162 & n1263 ;
  assign n1265 = n1264 ^ x80 ;
  assign n1266 = n175 & ~n1265 ;
  assign n1267 = n1266 ^ n270 ;
  assign n1268 = n1161 & ~n1267 ;
  assign n1269 = n1268 ^ x81 ;
  assign n1270 = n174 & ~n1269 ;
  assign n1271 = n1259 ^ x79 ;
  assign n1272 = n1266 & n1271 ;
  assign n1273 = n1272 ^ n1165 ;
  assign n1274 = n1273 ^ x80 ;
  assign n1324 = n1212 ^ x67 ;
  assign n1325 = n1266 & n1324 ;
  assign n1326 = n1325 ^ n1192 ;
  assign n1318 = n1210 & n1266 ;
  assign n1319 = n1318 ^ n1196 ;
  assign n1312 = x64 & n1159 ;
  assign n1308 = ~x47 & x64 ;
  assign n1309 = n1308 ^ x65 ;
  assign n1310 = n1266 & n1309 ;
  assign n1311 = n1310 ^ x48 ;
  assign n1313 = n1312 ^ n1311 ;
  assign n1299 = x65 ^ x46 ;
  assign n1303 = x64 & n1266 ;
  assign n1304 = ~n1299 & ~n1303 ;
  assign n1297 = ~x46 & x64 ;
  assign n1298 = n1297 ^ x65 ;
  assign n1302 = ~n1201 & n1298 ;
  assign n1305 = n1304 ^ n1302 ;
  assign n1306 = n1305 ^ x46 ;
  assign n1314 = n1313 ^ n1306 ;
  assign n1315 = n1313 ^ x66 ;
  assign n1316 = ~n1314 & ~n1315 ;
  assign n1317 = n1316 ^ x66 ;
  assign n1320 = n1319 ^ n1317 ;
  assign n1321 = n1319 ^ x67 ;
  assign n1322 = n1320 & ~n1321 ;
  assign n1323 = n1322 ^ x67 ;
  assign n1327 = n1326 ^ n1323 ;
  assign n1328 = n1326 ^ x68 ;
  assign n1329 = n1327 & ~n1328 ;
  assign n1330 = n1329 ^ x68 ;
  assign n1295 = n1217 & n1266 ;
  assign n1296 = n1295 ^ n1190 ;
  assign n1331 = n1330 ^ n1296 ;
  assign n1332 = n1330 ^ x69 ;
  assign n1333 = n1331 & n1332 ;
  assign n1334 = n1333 ^ x69 ;
  assign n1293 = n1221 & n1266 ;
  assign n1294 = n1293 ^ n1188 ;
  assign n1335 = n1334 ^ n1294 ;
  assign n1336 = n1334 ^ x70 ;
  assign n1337 = n1335 & n1336 ;
  assign n1338 = n1337 ^ x70 ;
  assign n1291 = n1225 & n1266 ;
  assign n1292 = n1291 ^ n1186 ;
  assign n1339 = n1338 ^ n1292 ;
  assign n1340 = n1338 ^ x71 ;
  assign n1341 = n1339 & n1340 ;
  assign n1342 = n1341 ^ x71 ;
  assign n1289 = n1229 & n1266 ;
  assign n1290 = n1289 ^ n1184 ;
  assign n1343 = n1342 ^ n1290 ;
  assign n1344 = n1342 ^ x72 ;
  assign n1345 = n1343 & n1344 ;
  assign n1346 = n1345 ^ x72 ;
  assign n1287 = n1233 & n1266 ;
  assign n1288 = n1287 ^ n1182 ;
  assign n1347 = n1346 ^ n1288 ;
  assign n1348 = n1346 ^ x73 ;
  assign n1349 = n1347 & n1348 ;
  assign n1350 = n1349 ^ x73 ;
  assign n1285 = n1237 & n1266 ;
  assign n1286 = n1285 ^ n1180 ;
  assign n1351 = n1350 ^ n1286 ;
  assign n1352 = n1350 ^ x74 ;
  assign n1353 = n1351 & n1352 ;
  assign n1354 = n1353 ^ x74 ;
  assign n1283 = n1241 & n1266 ;
  assign n1284 = n1283 ^ n1178 ;
  assign n1355 = n1354 ^ n1284 ;
  assign n1356 = n1354 ^ x75 ;
  assign n1357 = n1355 & n1356 ;
  assign n1358 = n1357 ^ x75 ;
  assign n1281 = n1245 & n1266 ;
  assign n1282 = n1281 ^ n1176 ;
  assign n1359 = n1358 ^ n1282 ;
  assign n1360 = n1358 ^ x76 ;
  assign n1361 = n1359 & n1360 ;
  assign n1362 = n1361 ^ x76 ;
  assign n1279 = n1249 & n1266 ;
  assign n1280 = n1279 ^ n1174 ;
  assign n1363 = n1362 ^ n1280 ;
  assign n1364 = n1362 ^ x77 ;
  assign n1365 = n1363 & n1364 ;
  assign n1366 = n1365 ^ x77 ;
  assign n1277 = n1253 & n1266 ;
  assign n1278 = n1277 ^ n1172 ;
  assign n1367 = n1366 ^ n1278 ;
  assign n1368 = n1366 ^ x78 ;
  assign n1369 = n1367 & n1368 ;
  assign n1370 = n1369 ^ x78 ;
  assign n1275 = n1257 & n1266 ;
  assign n1276 = n1275 ^ n1170 ;
  assign n1371 = n1370 ^ n1276 ;
  assign n1374 = n1276 ^ x79 ;
  assign n1375 = n1371 & ~n1374 ;
  assign n1372 = x80 ^ x79 ;
  assign n1376 = n1375 ^ n1372 ;
  assign n1379 = ~n1274 & n1376 ;
  assign n1380 = n1379 ^ x80 ;
  assign n1381 = n1270 & ~n1380 ;
  assign n1382 = n1061 & ~n1381 ;
  assign n1383 = n1382 ^ n270 ;
  assign n1384 = n1383 ^ x82 ;
  assign n1390 = n1383 ^ x81 ;
  assign n1385 = n175 & n1268 ;
  assign n1386 = n1385 ^ n1381 ;
  assign n1387 = n1376 & n1386 ;
  assign n1388 = n1387 ^ n1273 ;
  assign n1389 = n1388 ^ n1383 ;
  assign n1391 = n1390 ^ n1389 ;
  assign n1450 = n1332 & n1386 ;
  assign n1451 = n1450 ^ n1296 ;
  assign n1413 = n1323 ^ x68 ;
  assign n1414 = n1386 & n1413 ;
  assign n1415 = n1414 ^ n1326 ;
  assign n1416 = n1415 ^ x69 ;
  assign n1421 = n1415 ^ x68 ;
  assign n1417 = n1317 ^ x67 ;
  assign n1418 = n1386 & n1417 ;
  assign n1419 = n1418 ^ n1319 ;
  assign n1420 = n1419 ^ n1415 ;
  assign n1422 = n1421 ^ n1420 ;
  assign n1437 = n1306 ^ x66 ;
  assign n1438 = n1386 & ~n1437 ;
  assign n1439 = n1438 ^ n1313 ;
  assign n1431 = n1303 ^ x47 ;
  assign n1430 = n1298 & n1386 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1423 = ~x45 & x64 ;
  assign n1424 = n1423 ^ x65 ;
  assign n1425 = x64 & n1386 ;
  assign n1426 = n1425 ^ x46 ;
  assign n1427 = n1426 ^ n1423 ;
  assign n1428 = n1424 & n1427 ;
  assign n1429 = n1428 ^ x65 ;
  assign n1433 = n1432 ^ n1429 ;
  assign n1434 = n1432 ^ x66 ;
  assign n1435 = n1433 & ~n1434 ;
  assign n1436 = n1435 ^ x66 ;
  assign n1440 = n1439 ^ n1436 ;
  assign n1441 = n1439 ^ x67 ;
  assign n1442 = n1440 & ~n1441 ;
  assign n1443 = n1442 ^ x67 ;
  assign n1444 = n1443 ^ n1415 ;
  assign n1445 = n1444 ^ n1421 ;
  assign n1446 = ~n1422 & n1445 ;
  assign n1447 = n1446 ^ n1421 ;
  assign n1448 = ~n1416 & n1447 ;
  assign n1449 = n1448 ^ x69 ;
  assign n1452 = n1451 ^ n1449 ;
  assign n1453 = n1451 ^ x70 ;
  assign n1454 = n1452 & ~n1453 ;
  assign n1455 = n1454 ^ x70 ;
  assign n1411 = n1336 & n1386 ;
  assign n1412 = n1411 ^ n1294 ;
  assign n1456 = n1455 ^ n1412 ;
  assign n1457 = n1455 ^ x71 ;
  assign n1458 = n1456 & n1457 ;
  assign n1459 = n1458 ^ x71 ;
  assign n1409 = n1340 & n1386 ;
  assign n1410 = n1409 ^ n1292 ;
  assign n1460 = n1459 ^ n1410 ;
  assign n1461 = n1459 ^ x72 ;
  assign n1462 = n1460 & n1461 ;
  assign n1463 = n1462 ^ x72 ;
  assign n1407 = n1344 & n1386 ;
  assign n1408 = n1407 ^ n1290 ;
  assign n1464 = n1463 ^ n1408 ;
  assign n1465 = n1463 ^ x73 ;
  assign n1466 = n1464 & n1465 ;
  assign n1467 = n1466 ^ x73 ;
  assign n1405 = n1348 & n1386 ;
  assign n1406 = n1405 ^ n1288 ;
  assign n1468 = n1467 ^ n1406 ;
  assign n1469 = n1467 ^ x74 ;
  assign n1470 = n1468 & n1469 ;
  assign n1471 = n1470 ^ x74 ;
  assign n1403 = n1352 & n1386 ;
  assign n1404 = n1403 ^ n1286 ;
  assign n1472 = n1471 ^ n1404 ;
  assign n1473 = n1471 ^ x75 ;
  assign n1474 = n1472 & n1473 ;
  assign n1475 = n1474 ^ x75 ;
  assign n1401 = n1356 & n1386 ;
  assign n1402 = n1401 ^ n1284 ;
  assign n1476 = n1475 ^ n1402 ;
  assign n1477 = n1475 ^ x76 ;
  assign n1478 = n1476 & n1477 ;
  assign n1479 = n1478 ^ x76 ;
  assign n1399 = n1360 & n1386 ;
  assign n1400 = n1399 ^ n1282 ;
  assign n1480 = n1479 ^ n1400 ;
  assign n1481 = n1479 ^ x77 ;
  assign n1482 = n1480 & n1481 ;
  assign n1483 = n1482 ^ x77 ;
  assign n1397 = n1364 & n1386 ;
  assign n1398 = n1397 ^ n1280 ;
  assign n1484 = n1483 ^ n1398 ;
  assign n1485 = n1483 ^ x78 ;
  assign n1486 = n1484 & n1485 ;
  assign n1487 = n1486 ^ x78 ;
  assign n1395 = n1368 & n1386 ;
  assign n1396 = n1395 ^ n1278 ;
  assign n1488 = n1487 ^ n1396 ;
  assign n1489 = n1487 ^ x79 ;
  assign n1490 = n1488 & n1489 ;
  assign n1491 = n1490 ^ x79 ;
  assign n1392 = n1370 ^ x79 ;
  assign n1393 = n1386 & n1392 ;
  assign n1394 = n1393 ^ n1276 ;
  assign n1492 = n1491 ^ n1394 ;
  assign n1493 = n1491 ^ x80 ;
  assign n1494 = n1492 & n1493 ;
  assign n1495 = n1494 ^ x80 ;
  assign n1496 = n1495 ^ n1383 ;
  assign n1497 = n1496 ^ n1390 ;
  assign n1498 = ~n1391 & n1497 ;
  assign n1499 = n1498 ^ n1390 ;
  assign n1500 = ~n1384 & n1499 ;
  assign n1501 = n1500 ^ x82 ;
  assign n1502 = n173 & ~n1501 ;
  assign n1503 = n1382 & ~n1502 ;
  assign n1504 = n1503 ^ n270 ;
  assign n1505 = n1504 ^ x83 ;
  assign n1510 = n1504 ^ x82 ;
  assign n1506 = n1495 ^ x81 ;
  assign n1507 = n1502 & n1506 ;
  assign n1508 = n1507 ^ n1388 ;
  assign n1509 = n1508 ^ n1504 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1555 = n1424 & n1502 ;
  assign n1556 = n1555 ^ n1426 ;
  assign n1557 = n1556 ^ x66 ;
  assign n1563 = x45 & x65 ;
  assign n1558 = x65 ^ x44 ;
  assign n1559 = x64 ^ x45 ;
  assign n1560 = n1559 ^ x65 ;
  assign n1561 = n1560 ^ n1502 ;
  assign n1562 = ~n1558 & n1561 ;
  assign n1564 = n1563 ^ n1562 ;
  assign n1567 = x64 & n1564 ;
  assign n1568 = n1567 ^ n1563 ;
  assign n1569 = n1568 ^ x65 ;
  assign n1570 = n1569 ^ n1556 ;
  assign n1571 = ~n1557 & n1570 ;
  assign n1572 = n1571 ^ x66 ;
  assign n1552 = n1429 ^ x66 ;
  assign n1553 = n1502 & n1552 ;
  assign n1554 = n1553 ^ n1432 ;
  assign n1573 = n1572 ^ n1554 ;
  assign n1574 = n1572 ^ x67 ;
  assign n1575 = n1573 & n1574 ;
  assign n1576 = n1575 ^ x67 ;
  assign n1549 = n1436 ^ x67 ;
  assign n1550 = n1502 & n1549 ;
  assign n1551 = n1550 ^ n1439 ;
  assign n1577 = n1576 ^ n1551 ;
  assign n1578 = n1576 ^ x68 ;
  assign n1579 = n1577 & n1578 ;
  assign n1580 = n1579 ^ x68 ;
  assign n1546 = n1443 ^ x68 ;
  assign n1547 = n1502 & n1546 ;
  assign n1548 = n1547 ^ n1419 ;
  assign n1581 = n1580 ^ n1548 ;
  assign n1582 = n1580 ^ x69 ;
  assign n1583 = n1581 & n1582 ;
  assign n1584 = n1583 ^ x69 ;
  assign n1535 = n1419 ^ x69 ;
  assign n1536 = n1535 ^ x68 ;
  assign n1537 = n1536 ^ n1443 ;
  assign n1538 = n1537 ^ n1535 ;
  assign n1540 = x69 ^ x68 ;
  assign n1541 = n1540 ^ n1535 ;
  assign n1542 = ~n1538 & ~n1541 ;
  assign n1543 = n1542 ^ n1535 ;
  assign n1544 = n1502 & ~n1543 ;
  assign n1545 = n1544 ^ n1415 ;
  assign n1585 = n1584 ^ n1545 ;
  assign n1586 = n1584 ^ x70 ;
  assign n1587 = n1585 & n1586 ;
  assign n1588 = n1587 ^ x70 ;
  assign n1532 = n1449 ^ x70 ;
  assign n1533 = n1502 & n1532 ;
  assign n1534 = n1533 ^ n1451 ;
  assign n1589 = n1588 ^ n1534 ;
  assign n1590 = n1588 ^ x71 ;
  assign n1591 = n1589 & n1590 ;
  assign n1592 = n1591 ^ x71 ;
  assign n1530 = n1457 & n1502 ;
  assign n1531 = n1530 ^ n1412 ;
  assign n1593 = n1592 ^ n1531 ;
  assign n1594 = n1592 ^ x72 ;
  assign n1595 = n1593 & n1594 ;
  assign n1596 = n1595 ^ x72 ;
  assign n1528 = n1461 & n1502 ;
  assign n1529 = n1528 ^ n1410 ;
  assign n1597 = n1596 ^ n1529 ;
  assign n1598 = n1596 ^ x73 ;
  assign n1599 = n1597 & n1598 ;
  assign n1600 = n1599 ^ x73 ;
  assign n1526 = n1465 & n1502 ;
  assign n1527 = n1526 ^ n1408 ;
  assign n1601 = n1600 ^ n1527 ;
  assign n1602 = n1600 ^ x74 ;
  assign n1603 = n1601 & n1602 ;
  assign n1604 = n1603 ^ x74 ;
  assign n1524 = n1469 & n1502 ;
  assign n1525 = n1524 ^ n1406 ;
  assign n1605 = n1604 ^ n1525 ;
  assign n1606 = n1604 ^ x75 ;
  assign n1607 = n1605 & n1606 ;
  assign n1608 = n1607 ^ x75 ;
  assign n1522 = n1473 & n1502 ;
  assign n1523 = n1522 ^ n1404 ;
  assign n1609 = n1608 ^ n1523 ;
  assign n1610 = n1608 ^ x76 ;
  assign n1611 = n1609 & n1610 ;
  assign n1612 = n1611 ^ x76 ;
  assign n1520 = n1477 & n1502 ;
  assign n1521 = n1520 ^ n1402 ;
  assign n1613 = n1612 ^ n1521 ;
  assign n1614 = n1612 ^ x77 ;
  assign n1615 = n1613 & n1614 ;
  assign n1616 = n1615 ^ x77 ;
  assign n1518 = n1481 & n1502 ;
  assign n1519 = n1518 ^ n1400 ;
  assign n1617 = n1616 ^ n1519 ;
  assign n1618 = n1616 ^ x78 ;
  assign n1619 = n1617 & n1618 ;
  assign n1620 = n1619 ^ x78 ;
  assign n1516 = n1485 & n1502 ;
  assign n1517 = n1516 ^ n1398 ;
  assign n1621 = n1620 ^ n1517 ;
  assign n1622 = n1620 ^ x79 ;
  assign n1623 = n1621 & n1622 ;
  assign n1624 = n1623 ^ x79 ;
  assign n1514 = n1489 & n1502 ;
  assign n1515 = n1514 ^ n1396 ;
  assign n1625 = n1624 ^ n1515 ;
  assign n1626 = n1624 ^ x80 ;
  assign n1627 = n1625 & n1626 ;
  assign n1628 = n1627 ^ x80 ;
  assign n1512 = n1493 & n1502 ;
  assign n1513 = n1512 ^ n1394 ;
  assign n1629 = n1628 ^ n1513 ;
  assign n1630 = n1628 ^ x81 ;
  assign n1631 = n1629 & n1630 ;
  assign n1632 = n1631 ^ x81 ;
  assign n1633 = n1632 ^ n1504 ;
  assign n1634 = n1633 ^ n1510 ;
  assign n1635 = ~n1511 & n1634 ;
  assign n1636 = n1635 ^ n1510 ;
  assign n1637 = ~n1505 & n1636 ;
  assign n1638 = n1637 ^ x83 ;
  assign n1639 = n172 & ~n1638 ;
  assign n1640 = n1639 ^ n270 ;
  assign n1641 = n1504 & ~n1640 ;
  assign n1642 = n272 & n1641 ;
  assign n1643 = x84 & n1642 ;
  assign n1677 = n1569 ^ x66 ;
  assign n1678 = n1639 & n1677 ;
  assign n1679 = n1678 ^ n1556 ;
  assign n1680 = n1679 ^ x67 ;
  assign n1684 = x64 & n1639 ;
  assign n1685 = n1684 ^ x44 ;
  assign n1681 = ~x43 & x64 ;
  assign n1686 = n1685 ^ n1681 ;
  assign n1687 = x65 & ~n1686 ;
  assign n1682 = n1639 ^ x44 ;
  assign n1683 = n1681 & ~n1682 ;
  assign n1688 = n1687 ^ n1683 ;
  assign n1689 = n1688 ^ x66 ;
  assign n1693 = n1502 ^ x44 ;
  assign n1694 = n1693 ^ n1502 ;
  assign n1695 = n1639 & ~n1694 ;
  assign n1696 = n1695 ^ n1502 ;
  assign n1697 = x64 & n1696 ;
  assign n1698 = n1697 ^ x45 ;
  assign n1690 = x65 & n1639 ;
  assign n1699 = n1698 ^ n1690 ;
  assign n1700 = n1699 ^ n1688 ;
  assign n1701 = n1689 & n1700 ;
  assign n1702 = n1701 ^ x66 ;
  assign n1703 = n1702 ^ n1679 ;
  assign n1704 = ~n1680 & n1703 ;
  assign n1705 = n1704 ^ x67 ;
  assign n1675 = n1574 & n1639 ;
  assign n1676 = n1675 ^ n1554 ;
  assign n1706 = n1705 ^ n1676 ;
  assign n1707 = n1705 ^ x68 ;
  assign n1708 = n1706 & n1707 ;
  assign n1709 = n1708 ^ x68 ;
  assign n1673 = n1578 & n1639 ;
  assign n1674 = n1673 ^ n1551 ;
  assign n1710 = n1709 ^ n1674 ;
  assign n1711 = n1709 ^ x69 ;
  assign n1712 = n1710 & n1711 ;
  assign n1713 = n1712 ^ x69 ;
  assign n1671 = n1582 & n1639 ;
  assign n1672 = n1671 ^ n1548 ;
  assign n1714 = n1713 ^ n1672 ;
  assign n1715 = n1713 ^ x70 ;
  assign n1716 = n1714 & n1715 ;
  assign n1717 = n1716 ^ x70 ;
  assign n1669 = n1586 & n1639 ;
  assign n1670 = n1669 ^ n1545 ;
  assign n1718 = n1717 ^ n1670 ;
  assign n1719 = n1717 ^ x71 ;
  assign n1720 = n1718 & n1719 ;
  assign n1721 = n1720 ^ x71 ;
  assign n1667 = n1590 & n1639 ;
  assign n1668 = n1667 ^ n1534 ;
  assign n1722 = n1721 ^ n1668 ;
  assign n1723 = n1721 ^ x72 ;
  assign n1724 = n1722 & n1723 ;
  assign n1725 = n1724 ^ x72 ;
  assign n1665 = n1594 & n1639 ;
  assign n1666 = n1665 ^ n1531 ;
  assign n1726 = n1725 ^ n1666 ;
  assign n1727 = n1725 ^ x73 ;
  assign n1728 = n1726 & n1727 ;
  assign n1729 = n1728 ^ x73 ;
  assign n1663 = n1598 & n1639 ;
  assign n1664 = n1663 ^ n1529 ;
  assign n1730 = n1729 ^ n1664 ;
  assign n1731 = n1729 ^ x74 ;
  assign n1732 = n1730 & n1731 ;
  assign n1733 = n1732 ^ x74 ;
  assign n1661 = n1602 & n1639 ;
  assign n1662 = n1661 ^ n1527 ;
  assign n1734 = n1733 ^ n1662 ;
  assign n1735 = n1733 ^ x75 ;
  assign n1736 = n1734 & n1735 ;
  assign n1737 = n1736 ^ x75 ;
  assign n1659 = n1606 & n1639 ;
  assign n1660 = n1659 ^ n1525 ;
  assign n1738 = n1737 ^ n1660 ;
  assign n1739 = n1737 ^ x76 ;
  assign n1740 = n1738 & n1739 ;
  assign n1741 = n1740 ^ x76 ;
  assign n1657 = n1610 & n1639 ;
  assign n1658 = n1657 ^ n1523 ;
  assign n1742 = n1741 ^ n1658 ;
  assign n1743 = n1741 ^ x77 ;
  assign n1744 = n1742 & n1743 ;
  assign n1745 = n1744 ^ x77 ;
  assign n1655 = n1614 & n1639 ;
  assign n1656 = n1655 ^ n1521 ;
  assign n1746 = n1745 ^ n1656 ;
  assign n1747 = n1745 ^ x78 ;
  assign n1748 = n1746 & n1747 ;
  assign n1749 = n1748 ^ x78 ;
  assign n1653 = n1618 & n1639 ;
  assign n1654 = n1653 ^ n1519 ;
  assign n1750 = n1749 ^ n1654 ;
  assign n1751 = n1749 ^ x79 ;
  assign n1752 = n1750 & n1751 ;
  assign n1753 = n1752 ^ x79 ;
  assign n1651 = n1622 & n1639 ;
  assign n1652 = n1651 ^ n1517 ;
  assign n1754 = n1753 ^ n1652 ;
  assign n1755 = n1753 ^ x80 ;
  assign n1756 = n1754 & n1755 ;
  assign n1757 = n1756 ^ x80 ;
  assign n1649 = n1626 & n1639 ;
  assign n1650 = n1649 ^ n1515 ;
  assign n1758 = n1757 ^ n1650 ;
  assign n1759 = n1757 ^ x81 ;
  assign n1760 = n1758 & n1759 ;
  assign n1761 = n1760 ^ x81 ;
  assign n1647 = n1630 & n1639 ;
  assign n1648 = n1647 ^ n1513 ;
  assign n1762 = n1761 ^ n1648 ;
  assign n1763 = n1761 ^ x82 ;
  assign n1764 = n1762 & n1763 ;
  assign n1765 = n1764 ^ x82 ;
  assign n1644 = n1632 ^ x82 ;
  assign n1645 = n1639 & n1644 ;
  assign n1646 = n1645 ^ n1508 ;
  assign n1766 = n1765 ^ n1646 ;
  assign n1767 = n1765 ^ x83 ;
  assign n1768 = n1766 & n1767 ;
  assign n1769 = n1768 ^ x83 ;
  assign n1770 = n1643 & n1769 ;
  assign n1771 = n1770 ^ n1642 ;
  assign n1772 = n1771 ^ n1641 ;
  assign n1773 = ~x86 & n271 ;
  assign n1774 = n1772 ^ x85 ;
  assign n1783 = n1772 ^ x84 ;
  assign n1775 = n1641 ^ x84 ;
  assign n1776 = n1769 ^ x84 ;
  assign n1777 = ~n1775 & n1776 ;
  assign n1778 = n1777 ^ x84 ;
  assign n1779 = n272 & ~n1778 ;
  assign n1780 = n1767 & n1779 ;
  assign n1781 = n1780 ^ n1646 ;
  assign n1782 = n1781 ^ n1772 ;
  assign n1784 = n1783 ^ n1782 ;
  assign n1799 = n1735 & n1779 ;
  assign n1800 = n1799 ^ n1662 ;
  assign n1801 = n1800 ^ x76 ;
  assign n1802 = n1731 & n1779 ;
  assign n1803 = n1802 ^ n1664 ;
  assign n1804 = n1803 ^ x75 ;
  assign n1822 = n1681 ^ x65 ;
  assign n1823 = n1779 & n1822 ;
  assign n1824 = n1823 ^ n1685 ;
  assign n1825 = n1824 ^ x66 ;
  assign n1826 = ~x42 & x64 ;
  assign n1827 = n1826 ^ x43 ;
  assign n1834 = x65 & n1827 ;
  assign n1831 = n1826 ^ x65 ;
  assign n1832 = n1827 ^ n1779 ;
  assign n1833 = n1831 & n1832 ;
  assign n1835 = n1834 ^ n1833 ;
  assign n1836 = x64 & n1835 ;
  assign n1837 = n1836 ^ n1834 ;
  assign n1838 = n1837 ^ x65 ;
  assign n1839 = n1838 ^ n1824 ;
  assign n1840 = ~n1825 & n1839 ;
  assign n1841 = n1840 ^ x66 ;
  assign n1820 = n1689 & n1779 ;
  assign n1821 = n1820 ^ n1699 ;
  assign n1842 = n1841 ^ n1821 ;
  assign n1843 = n1841 ^ x67 ;
  assign n1844 = n1842 & n1843 ;
  assign n1845 = n1844 ^ x67 ;
  assign n1817 = n1702 ^ x67 ;
  assign n1818 = n1779 & n1817 ;
  assign n1819 = n1818 ^ n1679 ;
  assign n1846 = n1845 ^ n1819 ;
  assign n1847 = n1845 ^ x68 ;
  assign n1848 = n1846 & n1847 ;
  assign n1849 = n1848 ^ x68 ;
  assign n1815 = n1707 & n1779 ;
  assign n1816 = n1815 ^ n1676 ;
  assign n1850 = n1849 ^ n1816 ;
  assign n1851 = n1849 ^ x69 ;
  assign n1852 = n1850 & n1851 ;
  assign n1853 = n1852 ^ x69 ;
  assign n1813 = n1711 & n1779 ;
  assign n1814 = n1813 ^ n1674 ;
  assign n1854 = n1853 ^ n1814 ;
  assign n1855 = n1853 ^ x70 ;
  assign n1856 = n1854 & n1855 ;
  assign n1857 = n1856 ^ x70 ;
  assign n1811 = n1715 & n1779 ;
  assign n1812 = n1811 ^ n1672 ;
  assign n1858 = n1857 ^ n1812 ;
  assign n1859 = n1857 ^ x71 ;
  assign n1860 = n1858 & n1859 ;
  assign n1861 = n1860 ^ x71 ;
  assign n1809 = n1719 & n1779 ;
  assign n1810 = n1809 ^ n1670 ;
  assign n1862 = n1861 ^ n1810 ;
  assign n1863 = n1861 ^ x72 ;
  assign n1864 = n1862 & n1863 ;
  assign n1865 = n1864 ^ x72 ;
  assign n1807 = n1723 & n1779 ;
  assign n1808 = n1807 ^ n1668 ;
  assign n1866 = n1865 ^ n1808 ;
  assign n1867 = n1865 ^ x73 ;
  assign n1868 = n1866 & n1867 ;
  assign n1869 = n1868 ^ x73 ;
  assign n1805 = n1727 & n1779 ;
  assign n1806 = n1805 ^ n1666 ;
  assign n1870 = n1869 ^ n1806 ;
  assign n1871 = n1869 ^ x74 ;
  assign n1872 = n1870 & n1871 ;
  assign n1873 = n1872 ^ x74 ;
  assign n1874 = n1873 ^ n1803 ;
  assign n1875 = ~n1804 & n1874 ;
  assign n1876 = n1875 ^ x75 ;
  assign n1877 = n1876 ^ n1800 ;
  assign n1878 = ~n1801 & n1877 ;
  assign n1879 = n1878 ^ x76 ;
  assign n1797 = n1739 & n1779 ;
  assign n1798 = n1797 ^ n1660 ;
  assign n1880 = n1879 ^ n1798 ;
  assign n1881 = n1879 ^ x77 ;
  assign n1882 = n1880 & n1881 ;
  assign n1883 = n1882 ^ x77 ;
  assign n1795 = n1743 & n1779 ;
  assign n1796 = n1795 ^ n1658 ;
  assign n1884 = n1883 ^ n1796 ;
  assign n1885 = n1883 ^ x78 ;
  assign n1886 = n1884 & n1885 ;
  assign n1887 = n1886 ^ x78 ;
  assign n1793 = n1747 & n1779 ;
  assign n1794 = n1793 ^ n1656 ;
  assign n1888 = n1887 ^ n1794 ;
  assign n1889 = n1887 ^ x79 ;
  assign n1890 = n1888 & n1889 ;
  assign n1891 = n1890 ^ x79 ;
  assign n1791 = n1751 & n1779 ;
  assign n1792 = n1791 ^ n1654 ;
  assign n1892 = n1891 ^ n1792 ;
  assign n1893 = n1891 ^ x80 ;
  assign n1894 = n1892 & n1893 ;
  assign n1895 = n1894 ^ x80 ;
  assign n1789 = n1755 & n1779 ;
  assign n1790 = n1789 ^ n1652 ;
  assign n1896 = n1895 ^ n1790 ;
  assign n1897 = n1895 ^ x81 ;
  assign n1898 = n1896 & n1897 ;
  assign n1899 = n1898 ^ x81 ;
  assign n1787 = n1759 & n1779 ;
  assign n1788 = n1787 ^ n1650 ;
  assign n1900 = n1899 ^ n1788 ;
  assign n1901 = n1899 ^ x82 ;
  assign n1902 = n1900 & n1901 ;
  assign n1903 = n1902 ^ x82 ;
  assign n1785 = n1763 & n1779 ;
  assign n1786 = n1785 ^ n1648 ;
  assign n1904 = n1903 ^ n1786 ;
  assign n1905 = n1903 ^ x83 ;
  assign n1906 = n1904 & n1905 ;
  assign n1907 = n1906 ^ x83 ;
  assign n1908 = n1907 ^ n1772 ;
  assign n1909 = n1908 ^ n1783 ;
  assign n1910 = ~n1784 & n1909 ;
  assign n1911 = n1910 ^ n1783 ;
  assign n1912 = ~n1774 & n1911 ;
  assign n1913 = n1912 ^ x85 ;
  assign n1914 = n1773 & ~n1913 ;
  assign n1915 = n1772 & ~n1914 ;
  assign n1916 = n1915 ^ n270 ;
  assign n1917 = n1916 ^ x86 ;
  assign n2049 = n1907 ^ x84 ;
  assign n2050 = n1914 & n2049 ;
  assign n2051 = n2050 ^ n1781 ;
  assign n1918 = n1905 & n1914 ;
  assign n1919 = n1918 ^ n1786 ;
  assign n1921 = ~x84 & n1919 ;
  assign n1920 = n1919 ^ x84 ;
  assign n1922 = n1921 ^ n1920 ;
  assign n1927 = n1893 & n1914 ;
  assign n1928 = n1927 ^ n1792 ;
  assign n1929 = n1928 ^ x81 ;
  assign n1930 = n1889 & n1914 ;
  assign n1931 = n1930 ^ n1794 ;
  assign n1932 = n1931 ^ x80 ;
  assign n1973 = x42 & x65 ;
  assign n1970 = x65 ^ x41 ;
  assign n1966 = x64 ^ x42 ;
  assign n1967 = n1966 ^ x65 ;
  assign n1971 = n1967 ^ n1914 ;
  assign n1972 = ~n1970 & n1971 ;
  assign n1974 = n1973 ^ n1972 ;
  assign n1975 = x64 & n1974 ;
  assign n1976 = n1975 ^ n1973 ;
  assign n1977 = n1976 ^ x65 ;
  assign n1963 = n1831 & n1914 ;
  assign n1962 = x64 & n1779 ;
  assign n1964 = n1963 ^ n1962 ;
  assign n1965 = n1964 ^ x43 ;
  assign n1978 = n1977 ^ n1965 ;
  assign n1979 = n1977 ^ x66 ;
  assign n1980 = n1978 & n1979 ;
  assign n1981 = n1980 ^ x66 ;
  assign n1959 = n1838 ^ x66 ;
  assign n1960 = n1914 & n1959 ;
  assign n1961 = n1960 ^ n1824 ;
  assign n1982 = n1981 ^ n1961 ;
  assign n1983 = n1981 ^ x67 ;
  assign n1984 = n1982 & n1983 ;
  assign n1985 = n1984 ^ x67 ;
  assign n1957 = n1843 & n1914 ;
  assign n1958 = n1957 ^ n1821 ;
  assign n1986 = n1985 ^ n1958 ;
  assign n1987 = n1985 ^ x68 ;
  assign n1988 = n1986 & n1987 ;
  assign n1989 = n1988 ^ x68 ;
  assign n1955 = n1847 & n1914 ;
  assign n1956 = n1955 ^ n1819 ;
  assign n1990 = n1989 ^ n1956 ;
  assign n1991 = n1989 ^ x69 ;
  assign n1992 = n1990 & n1991 ;
  assign n1993 = n1992 ^ x69 ;
  assign n1953 = n1851 & n1914 ;
  assign n1954 = n1953 ^ n1816 ;
  assign n1994 = n1993 ^ n1954 ;
  assign n1995 = n1993 ^ x70 ;
  assign n1996 = n1994 & n1995 ;
  assign n1997 = n1996 ^ x70 ;
  assign n1951 = n1855 & n1914 ;
  assign n1952 = n1951 ^ n1814 ;
  assign n1998 = n1997 ^ n1952 ;
  assign n1999 = n1997 ^ x71 ;
  assign n2000 = n1998 & n1999 ;
  assign n2001 = n2000 ^ x71 ;
  assign n1949 = n1859 & n1914 ;
  assign n1950 = n1949 ^ n1812 ;
  assign n2002 = n2001 ^ n1950 ;
  assign n2003 = n2001 ^ x72 ;
  assign n2004 = n2002 & n2003 ;
  assign n2005 = n2004 ^ x72 ;
  assign n1947 = n1863 & n1914 ;
  assign n1948 = n1947 ^ n1810 ;
  assign n2006 = n2005 ^ n1948 ;
  assign n2007 = n2005 ^ x73 ;
  assign n2008 = n2006 & n2007 ;
  assign n2009 = n2008 ^ x73 ;
  assign n1945 = n1867 & n1914 ;
  assign n1946 = n1945 ^ n1808 ;
  assign n2010 = n2009 ^ n1946 ;
  assign n2011 = n2009 ^ x74 ;
  assign n2012 = n2010 & n2011 ;
  assign n2013 = n2012 ^ x74 ;
  assign n1943 = n1871 & n1914 ;
  assign n1944 = n1943 ^ n1806 ;
  assign n2014 = n2013 ^ n1944 ;
  assign n2015 = n2013 ^ x75 ;
  assign n2016 = n2014 & n2015 ;
  assign n2017 = n2016 ^ x75 ;
  assign n1940 = n1873 ^ x75 ;
  assign n1941 = n1914 & n1940 ;
  assign n1942 = n1941 ^ n1803 ;
  assign n2018 = n2017 ^ n1942 ;
  assign n2019 = n2017 ^ x76 ;
  assign n2020 = n2018 & n2019 ;
  assign n2021 = n2020 ^ x76 ;
  assign n1937 = n1876 ^ x76 ;
  assign n1938 = n1914 & n1937 ;
  assign n1939 = n1938 ^ n1800 ;
  assign n2022 = n2021 ^ n1939 ;
  assign n2023 = n2021 ^ x77 ;
  assign n2024 = n2022 & n2023 ;
  assign n2025 = n2024 ^ x77 ;
  assign n1935 = n1881 & n1914 ;
  assign n1936 = n1935 ^ n1798 ;
  assign n2026 = n2025 ^ n1936 ;
  assign n2027 = n2025 ^ x78 ;
  assign n2028 = n2026 & n2027 ;
  assign n2029 = n2028 ^ x78 ;
  assign n1933 = n1885 & n1914 ;
  assign n1934 = n1933 ^ n1796 ;
  assign n2030 = n2029 ^ n1934 ;
  assign n2031 = n2029 ^ x79 ;
  assign n2032 = n2030 & n2031 ;
  assign n2033 = n2032 ^ x79 ;
  assign n2034 = n2033 ^ n1931 ;
  assign n2035 = ~n1932 & n2034 ;
  assign n2036 = n2035 ^ x80 ;
  assign n2037 = n2036 ^ n1928 ;
  assign n2038 = ~n1929 & n2037 ;
  assign n2039 = n2038 ^ x81 ;
  assign n1925 = n1897 & n1914 ;
  assign n1926 = n1925 ^ n1790 ;
  assign n2040 = n2039 ^ n1926 ;
  assign n2041 = n2039 ^ x82 ;
  assign n2042 = n2040 & n2041 ;
  assign n2043 = n2042 ^ x82 ;
  assign n1923 = n1901 & n1914 ;
  assign n1924 = n1923 ^ n1788 ;
  assign n2044 = n2043 ^ n1924 ;
  assign n2045 = n2043 ^ x83 ;
  assign n2046 = n2044 & n2045 ;
  assign n2047 = n2046 ^ x83 ;
  assign n2048 = ~n1922 & ~n2047 ;
  assign n2052 = n2051 ^ n2048 ;
  assign n2053 = n2052 ^ n2051 ;
  assign n2054 = n2051 ^ n1921 ;
  assign n2055 = n2054 ^ n2051 ;
  assign n2056 = ~n2053 & ~n2055 ;
  assign n2057 = n2056 ^ n2051 ;
  assign n2060 = n2051 ^ x85 ;
  assign n2061 = n2057 & ~n2060 ;
  assign n2058 = x86 ^ x85 ;
  assign n2062 = n2061 ^ n2058 ;
  assign n2063 = ~n1917 & n2062 ;
  assign n2064 = n2063 ^ x86 ;
  assign n2065 = n271 & ~n2064 ;
  assign n2066 = n2065 ^ n270 ;
  assign n2067 = n1916 & ~n2066 ;
  assign n2068 = n169 & n2067 ;
  assign n2069 = x87 & n2068 ;
  assign n2113 = n1987 & n2065 ;
  assign n2114 = n2113 ^ n1958 ;
  assign n2115 = n2114 ^ x69 ;
  assign n2116 = n1983 & n2065 ;
  assign n2117 = n2116 ^ n1961 ;
  assign n2118 = n2117 ^ x68 ;
  assign n2133 = ~x40 & x64 ;
  assign n2134 = n2133 ^ x65 ;
  assign n2135 = x64 & n2065 ;
  assign n2136 = n2135 ^ n1970 ;
  assign n2137 = n2134 & ~n2136 ;
  assign n2138 = n2137 ^ x65 ;
  assign n2131 = ~x41 & x65 ;
  assign n2129 = x64 & n1914 ;
  assign n2127 = x65 ^ x42 ;
  assign n2121 = n2065 ^ x41 ;
  assign n2125 = n2135 ^ x65 ;
  assign n2126 = n2121 & n2125 ;
  assign n2128 = n2127 ^ n2126 ;
  assign n2130 = n2129 ^ n2128 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2139 = n2138 ^ n2132 ;
  assign n2140 = n2138 ^ x66 ;
  assign n2141 = n2139 & n2140 ;
  assign n2142 = n2141 ^ x66 ;
  assign n2119 = n1979 & n2065 ;
  assign n2120 = n2119 ^ n1965 ;
  assign n2143 = n2142 ^ n2120 ;
  assign n2144 = n2142 ^ x67 ;
  assign n2145 = n2143 & n2144 ;
  assign n2146 = n2145 ^ x67 ;
  assign n2147 = n2146 ^ n2117 ;
  assign n2148 = ~n2118 & n2147 ;
  assign n2149 = n2148 ^ x68 ;
  assign n2150 = n2149 ^ n2114 ;
  assign n2151 = ~n2115 & n2150 ;
  assign n2152 = n2151 ^ x69 ;
  assign n2111 = n1991 & n2065 ;
  assign n2112 = n2111 ^ n1956 ;
  assign n2153 = n2152 ^ n2112 ;
  assign n2154 = n2152 ^ x70 ;
  assign n2155 = n2153 & n2154 ;
  assign n2156 = n2155 ^ x70 ;
  assign n2109 = n1995 & n2065 ;
  assign n2110 = n2109 ^ n1954 ;
  assign n2157 = n2156 ^ n2110 ;
  assign n2158 = n2156 ^ x71 ;
  assign n2159 = n2157 & n2158 ;
  assign n2160 = n2159 ^ x71 ;
  assign n2107 = n1999 & n2065 ;
  assign n2108 = n2107 ^ n1952 ;
  assign n2161 = n2160 ^ n2108 ;
  assign n2162 = n2160 ^ x72 ;
  assign n2163 = n2161 & n2162 ;
  assign n2164 = n2163 ^ x72 ;
  assign n2105 = n2003 & n2065 ;
  assign n2106 = n2105 ^ n1950 ;
  assign n2165 = n2164 ^ n2106 ;
  assign n2166 = n2164 ^ x73 ;
  assign n2167 = n2165 & n2166 ;
  assign n2168 = n2167 ^ x73 ;
  assign n2103 = n2007 & n2065 ;
  assign n2104 = n2103 ^ n1948 ;
  assign n2169 = n2168 ^ n2104 ;
  assign n2170 = n2168 ^ x74 ;
  assign n2171 = n2169 & n2170 ;
  assign n2172 = n2171 ^ x74 ;
  assign n2101 = n2011 & n2065 ;
  assign n2102 = n2101 ^ n1946 ;
  assign n2173 = n2172 ^ n2102 ;
  assign n2174 = n2172 ^ x75 ;
  assign n2175 = n2173 & n2174 ;
  assign n2176 = n2175 ^ x75 ;
  assign n2099 = n2015 & n2065 ;
  assign n2100 = n2099 ^ n1944 ;
  assign n2177 = n2176 ^ n2100 ;
  assign n2178 = n2176 ^ x76 ;
  assign n2179 = n2177 & n2178 ;
  assign n2180 = n2179 ^ x76 ;
  assign n2097 = n2019 & n2065 ;
  assign n2098 = n2097 ^ n1942 ;
  assign n2181 = n2180 ^ n2098 ;
  assign n2182 = n2180 ^ x77 ;
  assign n2183 = n2181 & n2182 ;
  assign n2184 = n2183 ^ x77 ;
  assign n2095 = n2023 & n2065 ;
  assign n2096 = n2095 ^ n1939 ;
  assign n2185 = n2184 ^ n2096 ;
  assign n2186 = n2184 ^ x78 ;
  assign n2187 = n2185 & n2186 ;
  assign n2188 = n2187 ^ x78 ;
  assign n2093 = n2027 & n2065 ;
  assign n2094 = n2093 ^ n1936 ;
  assign n2189 = n2188 ^ n2094 ;
  assign n2190 = n2188 ^ x79 ;
  assign n2191 = n2189 & n2190 ;
  assign n2192 = n2191 ^ x79 ;
  assign n2091 = n2031 & n2065 ;
  assign n2092 = n2091 ^ n1934 ;
  assign n2193 = n2192 ^ n2092 ;
  assign n2194 = n2192 ^ x80 ;
  assign n2195 = n2193 & n2194 ;
  assign n2196 = n2195 ^ x80 ;
  assign n2088 = n2033 ^ x80 ;
  assign n2089 = n2065 & n2088 ;
  assign n2090 = n2089 ^ n1931 ;
  assign n2197 = n2196 ^ n2090 ;
  assign n2198 = n2196 ^ x81 ;
  assign n2199 = n2197 & n2198 ;
  assign n2200 = n2199 ^ x81 ;
  assign n2085 = n2036 ^ x81 ;
  assign n2086 = n2065 & n2085 ;
  assign n2087 = n2086 ^ n1928 ;
  assign n2201 = n2200 ^ n2087 ;
  assign n2202 = n2200 ^ x82 ;
  assign n2203 = n2201 & n2202 ;
  assign n2204 = n2203 ^ x82 ;
  assign n2083 = n2041 & n2065 ;
  assign n2084 = n2083 ^ n1926 ;
  assign n2205 = n2204 ^ n2084 ;
  assign n2206 = n2204 ^ x83 ;
  assign n2207 = n2205 & n2206 ;
  assign n2208 = n2207 ^ x83 ;
  assign n2081 = n2045 & n2065 ;
  assign n2082 = n2081 ^ n1924 ;
  assign n2209 = n2208 ^ n2082 ;
  assign n2210 = n2208 ^ x84 ;
  assign n2211 = n2209 & n2210 ;
  assign n2212 = n2211 ^ x84 ;
  assign n2078 = n2047 ^ x84 ;
  assign n2079 = n2065 & n2078 ;
  assign n2080 = n2079 ^ n1919 ;
  assign n2213 = n2212 ^ n2080 ;
  assign n2214 = n2212 ^ x85 ;
  assign n2215 = n2213 & n2214 ;
  assign n2216 = n2215 ^ x85 ;
  assign n2074 = ~n1921 & ~n2048 ;
  assign n2075 = n2074 ^ x85 ;
  assign n2076 = n2065 & n2075 ;
  assign n2077 = n2076 ^ n2051 ;
  assign n2217 = n2216 ^ n2077 ;
  assign n2218 = n2216 ^ x86 ;
  assign n2219 = n2217 & n2218 ;
  assign n2220 = n2219 ^ x86 ;
  assign n2221 = n2069 & n2220 ;
  assign n2222 = n2221 ^ n2068 ;
  assign n2223 = n2222 ^ n2067 ;
  assign n2224 = n2223 ^ x88 ;
  assign n2225 = n2067 ^ x87 ;
  assign n2226 = n2220 ^ x87 ;
  assign n2227 = ~n2225 & n2226 ;
  assign n2228 = n2227 ^ x87 ;
  assign n2229 = n169 & ~n2228 ;
  assign n2230 = n2218 & n2229 ;
  assign n2231 = n2230 ^ n2077 ;
  assign n2232 = n2231 ^ x87 ;
  assign n2257 = n2166 & n2229 ;
  assign n2258 = n2257 ^ n2106 ;
  assign n2259 = n2258 ^ x74 ;
  assign n2260 = n2162 & n2229 ;
  assign n2261 = n2260 ^ n2108 ;
  assign n2262 = n2261 ^ x73 ;
  assign n2278 = n2135 ^ x41 ;
  assign n2277 = n2134 & n2229 ;
  assign n2279 = n2278 ^ n2277 ;
  assign n2280 = n2279 ^ x66 ;
  assign n2286 = x40 & x65 ;
  assign n2281 = x65 ^ x39 ;
  assign n2282 = x64 ^ x40 ;
  assign n2283 = n2282 ^ x65 ;
  assign n2284 = n2283 ^ n2229 ;
  assign n2285 = ~n2281 & n2284 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2290 = x64 & n2287 ;
  assign n2291 = n2290 ^ n2286 ;
  assign n2292 = n2291 ^ x65 ;
  assign n2293 = n2292 ^ n2279 ;
  assign n2294 = ~n2280 & n2293 ;
  assign n2295 = n2294 ^ x66 ;
  assign n2275 = n2140 & n2229 ;
  assign n2276 = n2275 ^ n2132 ;
  assign n2296 = n2295 ^ n2276 ;
  assign n2297 = n2295 ^ x67 ;
  assign n2298 = n2296 & n2297 ;
  assign n2299 = n2298 ^ x67 ;
  assign n2273 = n2144 & n2229 ;
  assign n2274 = n2273 ^ n2120 ;
  assign n2300 = n2299 ^ n2274 ;
  assign n2301 = n2299 ^ x68 ;
  assign n2302 = n2300 & n2301 ;
  assign n2303 = n2302 ^ x68 ;
  assign n2270 = n2146 ^ x68 ;
  assign n2271 = n2229 & n2270 ;
  assign n2272 = n2271 ^ n2117 ;
  assign n2304 = n2303 ^ n2272 ;
  assign n2305 = n2303 ^ x69 ;
  assign n2306 = n2304 & n2305 ;
  assign n2307 = n2306 ^ x69 ;
  assign n2267 = n2149 ^ x69 ;
  assign n2268 = n2229 & n2267 ;
  assign n2269 = n2268 ^ n2114 ;
  assign n2308 = n2307 ^ n2269 ;
  assign n2309 = n2307 ^ x70 ;
  assign n2310 = n2308 & n2309 ;
  assign n2311 = n2310 ^ x70 ;
  assign n2265 = n2154 & n2229 ;
  assign n2266 = n2265 ^ n2112 ;
  assign n2312 = n2311 ^ n2266 ;
  assign n2313 = n2311 ^ x71 ;
  assign n2314 = n2312 & n2313 ;
  assign n2315 = n2314 ^ x71 ;
  assign n2263 = n2158 & n2229 ;
  assign n2264 = n2263 ^ n2110 ;
  assign n2316 = n2315 ^ n2264 ;
  assign n2317 = n2315 ^ x72 ;
  assign n2318 = n2316 & n2317 ;
  assign n2319 = n2318 ^ x72 ;
  assign n2320 = n2319 ^ n2261 ;
  assign n2321 = ~n2262 & n2320 ;
  assign n2322 = n2321 ^ x73 ;
  assign n2323 = n2322 ^ n2258 ;
  assign n2324 = ~n2259 & n2323 ;
  assign n2325 = n2324 ^ x74 ;
  assign n2255 = n2170 & n2229 ;
  assign n2256 = n2255 ^ n2104 ;
  assign n2326 = n2325 ^ n2256 ;
  assign n2327 = n2325 ^ x75 ;
  assign n2328 = n2326 & n2327 ;
  assign n2329 = n2328 ^ x75 ;
  assign n2253 = n2174 & n2229 ;
  assign n2254 = n2253 ^ n2102 ;
  assign n2330 = n2329 ^ n2254 ;
  assign n2331 = n2329 ^ x76 ;
  assign n2332 = n2330 & n2331 ;
  assign n2333 = n2332 ^ x76 ;
  assign n2251 = n2178 & n2229 ;
  assign n2252 = n2251 ^ n2100 ;
  assign n2334 = n2333 ^ n2252 ;
  assign n2335 = n2333 ^ x77 ;
  assign n2336 = n2334 & n2335 ;
  assign n2337 = n2336 ^ x77 ;
  assign n2249 = n2182 & n2229 ;
  assign n2250 = n2249 ^ n2098 ;
  assign n2338 = n2337 ^ n2250 ;
  assign n2339 = n2337 ^ x78 ;
  assign n2340 = n2338 & n2339 ;
  assign n2341 = n2340 ^ x78 ;
  assign n2247 = n2186 & n2229 ;
  assign n2248 = n2247 ^ n2096 ;
  assign n2342 = n2341 ^ n2248 ;
  assign n2343 = n2341 ^ x79 ;
  assign n2344 = n2342 & n2343 ;
  assign n2345 = n2344 ^ x79 ;
  assign n2245 = n2190 & n2229 ;
  assign n2246 = n2245 ^ n2094 ;
  assign n2346 = n2345 ^ n2246 ;
  assign n2347 = n2345 ^ x80 ;
  assign n2348 = n2346 & n2347 ;
  assign n2349 = n2348 ^ x80 ;
  assign n2243 = n2194 & n2229 ;
  assign n2244 = n2243 ^ n2092 ;
  assign n2350 = n2349 ^ n2244 ;
  assign n2351 = n2349 ^ x81 ;
  assign n2352 = n2350 & n2351 ;
  assign n2353 = n2352 ^ x81 ;
  assign n2241 = n2198 & n2229 ;
  assign n2242 = n2241 ^ n2090 ;
  assign n2354 = n2353 ^ n2242 ;
  assign n2355 = n2353 ^ x82 ;
  assign n2356 = n2354 & n2355 ;
  assign n2357 = n2356 ^ x82 ;
  assign n2239 = n2202 & n2229 ;
  assign n2240 = n2239 ^ n2087 ;
  assign n2358 = n2357 ^ n2240 ;
  assign n2359 = n2357 ^ x83 ;
  assign n2360 = n2358 & n2359 ;
  assign n2361 = n2360 ^ x83 ;
  assign n2237 = n2206 & n2229 ;
  assign n2238 = n2237 ^ n2084 ;
  assign n2362 = n2361 ^ n2238 ;
  assign n2363 = n2361 ^ x84 ;
  assign n2364 = n2362 & n2363 ;
  assign n2365 = n2364 ^ x84 ;
  assign n2235 = n2210 & n2229 ;
  assign n2236 = n2235 ^ n2082 ;
  assign n2366 = n2365 ^ n2236 ;
  assign n2367 = n2365 ^ x85 ;
  assign n2368 = n2366 & n2367 ;
  assign n2369 = n2368 ^ x85 ;
  assign n2233 = n2214 & n2229 ;
  assign n2234 = n2233 ^ n2080 ;
  assign n2370 = n2369 ^ n2234 ;
  assign n2373 = n2234 ^ x86 ;
  assign n2374 = n2370 & ~n2373 ;
  assign n2371 = x87 ^ x86 ;
  assign n2375 = n2374 ^ n2371 ;
  assign n2378 = ~n2232 & n2375 ;
  assign n2379 = n2378 ^ x87 ;
  assign n2380 = ~n2224 & n2379 ;
  assign n2381 = n168 & ~n2380 ;
  assign n2382 = x88 & ~n2067 ;
  assign n2383 = n2381 & n2382 ;
  assign n2384 = n2383 ^ n2381 ;
  assign n2385 = n2223 & ~n2384 ;
  assign n2386 = n2385 ^ n270 ;
  assign n2387 = n270 ^ n166 ;
  assign n2388 = n2386 & n2387 ;
  assign n2728 = n2388 ^ n2386 ;
  assign n2445 = x39 & x65 ;
  assign n2440 = x65 ^ x38 ;
  assign n2441 = x64 ^ x39 ;
  assign n2442 = n2441 ^ x65 ;
  assign n2443 = n2442 ^ n2384 ;
  assign n2444 = ~n2440 & n2443 ;
  assign n2446 = n2445 ^ n2444 ;
  assign n2449 = x64 & n2446 ;
  assign n2450 = n2449 ^ n2445 ;
  assign n2451 = n2450 ^ x65 ;
  assign n2452 = n2451 ^ x66 ;
  assign n2454 = n2229 ^ x39 ;
  assign n2455 = n2454 ^ n2229 ;
  assign n2458 = n2384 & ~n2455 ;
  assign n2459 = n2458 ^ n2229 ;
  assign n2460 = x64 & n2459 ;
  assign n2461 = n2460 ^ x40 ;
  assign n2453 = x65 & n2384 ;
  assign n2462 = n2461 ^ n2453 ;
  assign n2463 = n2462 ^ n2451 ;
  assign n2464 = n2452 & n2463 ;
  assign n2465 = n2464 ^ x66 ;
  assign n2437 = n2292 ^ x66 ;
  assign n2438 = n2384 & n2437 ;
  assign n2439 = n2438 ^ n2279 ;
  assign n2466 = n2465 ^ n2439 ;
  assign n2467 = n2465 ^ x67 ;
  assign n2468 = n2466 & n2467 ;
  assign n2469 = n2468 ^ x67 ;
  assign n2435 = n2297 & n2384 ;
  assign n2436 = n2435 ^ n2276 ;
  assign n2470 = n2469 ^ n2436 ;
  assign n2471 = n2469 ^ x68 ;
  assign n2472 = n2470 & n2471 ;
  assign n2473 = n2472 ^ x68 ;
  assign n2433 = n2301 & n2384 ;
  assign n2434 = n2433 ^ n2274 ;
  assign n2474 = n2473 ^ n2434 ;
  assign n2475 = n2473 ^ x69 ;
  assign n2476 = n2474 & n2475 ;
  assign n2477 = n2476 ^ x69 ;
  assign n2431 = n2305 & n2384 ;
  assign n2432 = n2431 ^ n2272 ;
  assign n2478 = n2477 ^ n2432 ;
  assign n2479 = n2477 ^ x70 ;
  assign n2480 = n2478 & n2479 ;
  assign n2481 = n2480 ^ x70 ;
  assign n2482 = n2481 ^ x71 ;
  assign n2483 = n2309 & n2384 ;
  assign n2484 = n2483 ^ n2269 ;
  assign n2485 = n2484 ^ n2481 ;
  assign n2486 = n2482 & n2485 ;
  assign n2487 = n2486 ^ x71 ;
  assign n2489 = n2487 ^ x72 ;
  assign n2389 = n2386 ^ x89 ;
  assign n2393 = n2386 ^ x88 ;
  assign n2390 = n2375 & n2384 ;
  assign n2391 = n2390 ^ n2231 ;
  assign n2392 = n2391 ^ n2386 ;
  assign n2394 = n2393 ^ n2392 ;
  assign n2395 = n2369 ^ x86 ;
  assign n2396 = n2384 & n2395 ;
  assign n2397 = n2396 ^ n2234 ;
  assign n2398 = n2397 ^ x87 ;
  assign n2429 = n2313 & n2384 ;
  assign n2430 = n2429 ^ n2266 ;
  assign n2488 = n2487 ^ n2430 ;
  assign n2490 = n2488 & n2489 ;
  assign n2491 = n2490 ^ x72 ;
  assign n2427 = n2317 & n2384 ;
  assign n2428 = n2427 ^ n2264 ;
  assign n2492 = n2491 ^ n2428 ;
  assign n2493 = n2491 ^ x73 ;
  assign n2494 = n2492 & n2493 ;
  assign n2495 = n2494 ^ x73 ;
  assign n2424 = n2319 ^ x73 ;
  assign n2425 = n2384 & n2424 ;
  assign n2426 = n2425 ^ n2261 ;
  assign n2496 = n2495 ^ n2426 ;
  assign n2497 = n2495 ^ x74 ;
  assign n2498 = n2496 & n2497 ;
  assign n2499 = n2498 ^ x74 ;
  assign n2421 = n2322 ^ x74 ;
  assign n2422 = n2384 & n2421 ;
  assign n2423 = n2422 ^ n2258 ;
  assign n2500 = n2499 ^ n2423 ;
  assign n2501 = n2499 ^ x75 ;
  assign n2502 = n2500 & n2501 ;
  assign n2503 = n2502 ^ x75 ;
  assign n2419 = n2327 & n2384 ;
  assign n2420 = n2419 ^ n2256 ;
  assign n2504 = n2503 ^ n2420 ;
  assign n2505 = n2503 ^ x76 ;
  assign n2506 = n2504 & n2505 ;
  assign n2507 = n2506 ^ x76 ;
  assign n2417 = n2331 & n2384 ;
  assign n2418 = n2417 ^ n2254 ;
  assign n2508 = n2507 ^ n2418 ;
  assign n2509 = n2507 ^ x77 ;
  assign n2510 = n2508 & n2509 ;
  assign n2511 = n2510 ^ x77 ;
  assign n2415 = n2335 & n2384 ;
  assign n2416 = n2415 ^ n2252 ;
  assign n2512 = n2511 ^ n2416 ;
  assign n2513 = n2511 ^ x78 ;
  assign n2514 = n2512 & n2513 ;
  assign n2515 = n2514 ^ x78 ;
  assign n2413 = n2339 & n2384 ;
  assign n2414 = n2413 ^ n2250 ;
  assign n2516 = n2515 ^ n2414 ;
  assign n2517 = n2515 ^ x79 ;
  assign n2518 = n2516 & n2517 ;
  assign n2519 = n2518 ^ x79 ;
  assign n2411 = n2343 & n2384 ;
  assign n2412 = n2411 ^ n2248 ;
  assign n2520 = n2519 ^ n2412 ;
  assign n2521 = n2519 ^ x80 ;
  assign n2522 = n2520 & n2521 ;
  assign n2523 = n2522 ^ x80 ;
  assign n2409 = n2347 & n2384 ;
  assign n2410 = n2409 ^ n2246 ;
  assign n2524 = n2523 ^ n2410 ;
  assign n2525 = n2523 ^ x81 ;
  assign n2526 = n2524 & n2525 ;
  assign n2527 = n2526 ^ x81 ;
  assign n2407 = n2351 & n2384 ;
  assign n2408 = n2407 ^ n2244 ;
  assign n2528 = n2527 ^ n2408 ;
  assign n2529 = n2527 ^ x82 ;
  assign n2530 = n2528 & n2529 ;
  assign n2531 = n2530 ^ x82 ;
  assign n2405 = n2355 & n2384 ;
  assign n2406 = n2405 ^ n2242 ;
  assign n2532 = n2531 ^ n2406 ;
  assign n2533 = n2531 ^ x83 ;
  assign n2534 = n2532 & n2533 ;
  assign n2535 = n2534 ^ x83 ;
  assign n2403 = n2359 & n2384 ;
  assign n2404 = n2403 ^ n2240 ;
  assign n2536 = n2535 ^ n2404 ;
  assign n2537 = n2535 ^ x84 ;
  assign n2538 = n2536 & n2537 ;
  assign n2539 = n2538 ^ x84 ;
  assign n2401 = n2363 & n2384 ;
  assign n2402 = n2401 ^ n2238 ;
  assign n2540 = n2539 ^ n2402 ;
  assign n2541 = n2539 ^ x85 ;
  assign n2542 = n2540 & n2541 ;
  assign n2543 = n2542 ^ x85 ;
  assign n2399 = n2367 & n2384 ;
  assign n2400 = n2399 ^ n2236 ;
  assign n2544 = n2543 ^ n2400 ;
  assign n2545 = n2543 ^ x86 ;
  assign n2546 = n2544 & n2545 ;
  assign n2547 = n2546 ^ x86 ;
  assign n2548 = n2547 ^ n2397 ;
  assign n2549 = ~n2398 & n2548 ;
  assign n2550 = n2549 ^ x87 ;
  assign n2551 = n2550 ^ n2386 ;
  assign n2552 = n2551 ^ n2393 ;
  assign n2553 = ~n2394 & n2552 ;
  assign n2554 = n2553 ^ n2393 ;
  assign n2555 = ~n2389 & n2554 ;
  assign n2556 = n2555 ^ x89 ;
  assign n2557 = n167 & ~n2556 ;
  assign n2656 = n2489 & n2557 ;
  assign n2657 = n2656 ^ n2430 ;
  assign n2592 = n2482 & n2557 ;
  assign n2593 = n2592 ^ n2484 ;
  assign n2594 = n2593 ^ x72 ;
  assign n2598 = n2593 ^ x71 ;
  assign n2595 = n2479 & n2557 ;
  assign n2596 = n2595 ^ n2432 ;
  assign n2597 = n2596 ^ n2593 ;
  assign n2599 = n2598 ^ n2597 ;
  assign n2611 = n2384 ^ x38 ;
  assign n2612 = n2611 ^ n2384 ;
  assign n2613 = n2557 & ~n2612 ;
  assign n2614 = n2613 ^ n2384 ;
  assign n2615 = x64 & n2614 ;
  assign n2616 = n2615 ^ x39 ;
  assign n2608 = x65 & n2557 ;
  assign n2617 = n2616 ^ n2608 ;
  assign n2618 = n2617 ^ x66 ;
  assign n2626 = x38 & x65 ;
  assign n2623 = x65 ^ x37 ;
  assign n2619 = x64 ^ x38 ;
  assign n2620 = n2619 ^ x65 ;
  assign n2624 = n2620 ^ n2557 ;
  assign n2625 = ~n2623 & n2624 ;
  assign n2627 = n2626 ^ n2625 ;
  assign n2628 = x64 & n2627 ;
  assign n2629 = n2628 ^ n2626 ;
  assign n2630 = n2629 ^ x65 ;
  assign n2631 = n2630 ^ n2617 ;
  assign n2632 = ~n2618 & n2631 ;
  assign n2633 = n2632 ^ x66 ;
  assign n2606 = n2452 & n2557 ;
  assign n2607 = n2606 ^ n2462 ;
  assign n2634 = n2633 ^ n2607 ;
  assign n2635 = n2633 ^ x67 ;
  assign n2636 = n2634 & n2635 ;
  assign n2637 = n2636 ^ x67 ;
  assign n2604 = n2467 & n2557 ;
  assign n2605 = n2604 ^ n2439 ;
  assign n2638 = n2637 ^ n2605 ;
  assign n2639 = n2637 ^ x68 ;
  assign n2640 = n2638 & n2639 ;
  assign n2641 = n2640 ^ x68 ;
  assign n2602 = n2471 & n2557 ;
  assign n2603 = n2602 ^ n2436 ;
  assign n2642 = n2641 ^ n2603 ;
  assign n2643 = n2641 ^ x69 ;
  assign n2644 = n2642 & n2643 ;
  assign n2645 = n2644 ^ x69 ;
  assign n2600 = n2475 & n2557 ;
  assign n2601 = n2600 ^ n2434 ;
  assign n2646 = n2645 ^ n2601 ;
  assign n2647 = n2645 ^ x70 ;
  assign n2648 = n2646 & n2647 ;
  assign n2649 = n2648 ^ x70 ;
  assign n2650 = n2649 ^ n2593 ;
  assign n2651 = n2650 ^ n2598 ;
  assign n2652 = ~n2599 & n2651 ;
  assign n2653 = n2652 ^ n2598 ;
  assign n2654 = ~n2594 & n2653 ;
  assign n2655 = n2654 ^ x72 ;
  assign n2658 = n2657 ^ n2655 ;
  assign n2659 = n2657 ^ x73 ;
  assign n2660 = n2658 & ~n2659 ;
  assign n2661 = n2660 ^ x73 ;
  assign n2590 = n2493 & n2557 ;
  assign n2591 = n2590 ^ n2428 ;
  assign n2662 = n2661 ^ n2591 ;
  assign n2663 = n2661 ^ x74 ;
  assign n2664 = n2662 & n2663 ;
  assign n2665 = n2664 ^ x74 ;
  assign n2588 = n2497 & n2557 ;
  assign n2589 = n2588 ^ n2426 ;
  assign n2666 = n2665 ^ n2589 ;
  assign n2667 = n2665 ^ x75 ;
  assign n2668 = n2666 & n2667 ;
  assign n2669 = n2668 ^ x75 ;
  assign n2586 = n2501 & n2557 ;
  assign n2587 = n2586 ^ n2423 ;
  assign n2670 = n2669 ^ n2587 ;
  assign n2671 = n2669 ^ x76 ;
  assign n2672 = n2670 & n2671 ;
  assign n2673 = n2672 ^ x76 ;
  assign n2584 = n2505 & n2557 ;
  assign n2585 = n2584 ^ n2420 ;
  assign n2674 = n2673 ^ n2585 ;
  assign n2675 = n2673 ^ x77 ;
  assign n2676 = n2674 & n2675 ;
  assign n2677 = n2676 ^ x77 ;
  assign n2582 = n2509 & n2557 ;
  assign n2583 = n2582 ^ n2418 ;
  assign n2678 = n2677 ^ n2583 ;
  assign n2679 = n2677 ^ x78 ;
  assign n2680 = n2678 & n2679 ;
  assign n2681 = n2680 ^ x78 ;
  assign n2580 = n2513 & n2557 ;
  assign n2581 = n2580 ^ n2416 ;
  assign n2682 = n2681 ^ n2581 ;
  assign n2683 = n2681 ^ x79 ;
  assign n2684 = n2682 & n2683 ;
  assign n2685 = n2684 ^ x79 ;
  assign n2578 = n2517 & n2557 ;
  assign n2579 = n2578 ^ n2414 ;
  assign n2686 = n2685 ^ n2579 ;
  assign n2687 = n2685 ^ x80 ;
  assign n2688 = n2686 & n2687 ;
  assign n2689 = n2688 ^ x80 ;
  assign n2576 = n2521 & n2557 ;
  assign n2577 = n2576 ^ n2412 ;
  assign n2690 = n2689 ^ n2577 ;
  assign n2691 = n2689 ^ x81 ;
  assign n2692 = n2690 & n2691 ;
  assign n2693 = n2692 ^ x81 ;
  assign n2574 = n2525 & n2557 ;
  assign n2575 = n2574 ^ n2410 ;
  assign n2694 = n2693 ^ n2575 ;
  assign n2695 = n2693 ^ x82 ;
  assign n2696 = n2694 & n2695 ;
  assign n2697 = n2696 ^ x82 ;
  assign n2572 = n2529 & n2557 ;
  assign n2573 = n2572 ^ n2408 ;
  assign n2698 = n2697 ^ n2573 ;
  assign n2699 = n2697 ^ x83 ;
  assign n2700 = n2698 & n2699 ;
  assign n2701 = n2700 ^ x83 ;
  assign n2570 = n2533 & n2557 ;
  assign n2571 = n2570 ^ n2406 ;
  assign n2702 = n2701 ^ n2571 ;
  assign n2703 = n2701 ^ x84 ;
  assign n2704 = n2702 & n2703 ;
  assign n2705 = n2704 ^ x84 ;
  assign n2568 = n2537 & n2557 ;
  assign n2569 = n2568 ^ n2404 ;
  assign n2706 = n2705 ^ n2569 ;
  assign n2707 = n2705 ^ x85 ;
  assign n2708 = n2706 & n2707 ;
  assign n2709 = n2708 ^ x85 ;
  assign n2566 = n2541 & n2557 ;
  assign n2567 = n2566 ^ n2402 ;
  assign n2710 = n2709 ^ n2567 ;
  assign n2711 = n2709 ^ x86 ;
  assign n2712 = n2710 & n2711 ;
  assign n2713 = n2712 ^ x86 ;
  assign n2564 = n2545 & n2557 ;
  assign n2565 = n2564 ^ n2400 ;
  assign n2714 = n2713 ^ n2565 ;
  assign n2715 = n2713 ^ x87 ;
  assign n2716 = n2714 & n2715 ;
  assign n2717 = n2716 ^ x87 ;
  assign n2561 = n2547 ^ x87 ;
  assign n2562 = n2557 & n2561 ;
  assign n2563 = n2562 ^ n2397 ;
  assign n2718 = n2717 ^ n2563 ;
  assign n2719 = n2717 ^ x88 ;
  assign n2720 = n2718 & n2719 ;
  assign n2721 = n2720 ^ x88 ;
  assign n2558 = n2550 ^ x88 ;
  assign n2559 = n2557 & n2558 ;
  assign n2560 = n2559 ^ n2391 ;
  assign n2722 = n2721 ^ n2560 ;
  assign n2723 = n2721 ^ x89 ;
  assign n2724 = n2722 & n2723 ;
  assign n2725 = n2724 ^ x89 ;
  assign n2726 = x90 & n2725 ;
  assign n2727 = n2388 & n2726 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2730 = n2729 ^ x91 ;
  assign n2917 = n2729 ^ x90 ;
  assign n2731 = n2725 ^ x90 ;
  assign n2732 = n2725 ^ n270 ;
  assign n2733 = n2732 ^ n2386 ;
  assign n2734 = n2733 ^ n2732 ;
  assign n2735 = n2732 ^ n2556 ;
  assign n2736 = n2735 ^ n2725 ;
  assign n2737 = n2736 ^ n2732 ;
  assign n2738 = n2734 & ~n2737 ;
  assign n2739 = n2738 ^ n2732 ;
  assign n2740 = n2731 & n2739 ;
  assign n2741 = n2740 ^ x90 ;
  assign n2742 = n166 & ~n2741 ;
  assign n2743 = n2719 & n2742 ;
  assign n2744 = n2743 ^ n2563 ;
  assign n2745 = n2744 ^ x89 ;
  assign n2760 = n2687 & n2742 ;
  assign n2761 = n2760 ^ n2579 ;
  assign n2762 = n2761 ^ x81 ;
  assign n2763 = n2683 & n2742 ;
  assign n2764 = n2763 ^ n2581 ;
  assign n2765 = n2764 ^ x80 ;
  assign n2807 = x64 & n2557 ;
  assign n2803 = ~x37 & x64 ;
  assign n2804 = n2803 ^ x65 ;
  assign n2805 = n2742 & n2804 ;
  assign n2806 = n2805 ^ x38 ;
  assign n2808 = n2807 ^ n2806 ;
  assign n2809 = n2808 ^ x66 ;
  assign n2817 = x37 & x65 ;
  assign n2814 = x65 ^ x36 ;
  assign n2810 = x64 ^ x37 ;
  assign n2811 = n2810 ^ x65 ;
  assign n2815 = n2811 ^ n2742 ;
  assign n2816 = ~n2814 & n2815 ;
  assign n2818 = n2817 ^ n2816 ;
  assign n2819 = x64 & n2818 ;
  assign n2820 = n2819 ^ n2817 ;
  assign n2821 = n2820 ^ x65 ;
  assign n2822 = n2821 ^ n2808 ;
  assign n2823 = ~n2809 & n2822 ;
  assign n2824 = n2823 ^ x66 ;
  assign n2799 = n2630 ^ x66 ;
  assign n2800 = n2742 & n2799 ;
  assign n2801 = n2800 ^ n2617 ;
  assign n2825 = n2824 ^ n2801 ;
  assign n2826 = n2824 ^ x67 ;
  assign n2827 = n2825 & n2826 ;
  assign n2828 = n2827 ^ x67 ;
  assign n2829 = n2828 ^ x68 ;
  assign n2830 = n2635 & n2742 ;
  assign n2831 = n2830 ^ n2607 ;
  assign n2832 = n2831 ^ n2828 ;
  assign n2833 = n2829 & n2832 ;
  assign n2834 = n2833 ^ x68 ;
  assign n2797 = n2639 & n2742 ;
  assign n2798 = n2797 ^ n2605 ;
  assign n2835 = n2834 ^ n2798 ;
  assign n2836 = n2834 ^ x69 ;
  assign n2837 = n2835 & n2836 ;
  assign n2838 = n2837 ^ x69 ;
  assign n2795 = n2643 & n2742 ;
  assign n2796 = n2795 ^ n2603 ;
  assign n2839 = n2838 ^ n2796 ;
  assign n2840 = n2838 ^ x70 ;
  assign n2841 = n2839 & n2840 ;
  assign n2842 = n2841 ^ x70 ;
  assign n2793 = n2647 & n2742 ;
  assign n2794 = n2793 ^ n2601 ;
  assign n2843 = n2842 ^ n2794 ;
  assign n2844 = n2842 ^ x71 ;
  assign n2845 = n2843 & n2844 ;
  assign n2846 = n2845 ^ x71 ;
  assign n2790 = n2649 ^ x71 ;
  assign n2791 = n2742 & n2790 ;
  assign n2792 = n2791 ^ n2596 ;
  assign n2847 = n2846 ^ n2792 ;
  assign n2848 = n2846 ^ x72 ;
  assign n2849 = n2847 & n2848 ;
  assign n2850 = n2849 ^ x72 ;
  assign n2779 = n2596 ^ x72 ;
  assign n2780 = n2779 ^ n2649 ;
  assign n2781 = n2780 ^ x71 ;
  assign n2782 = n2781 ^ n2779 ;
  assign n2784 = n2649 ^ x72 ;
  assign n2785 = n2784 ^ n2779 ;
  assign n2786 = ~n2782 & ~n2785 ;
  assign n2787 = n2786 ^ n2779 ;
  assign n2788 = n2742 & ~n2787 ;
  assign n2789 = n2788 ^ n2593 ;
  assign n2851 = n2850 ^ n2789 ;
  assign n2852 = n2850 ^ x73 ;
  assign n2853 = n2851 & n2852 ;
  assign n2854 = n2853 ^ x73 ;
  assign n2776 = n2655 ^ x73 ;
  assign n2777 = n2742 & n2776 ;
  assign n2778 = n2777 ^ n2657 ;
  assign n2855 = n2854 ^ n2778 ;
  assign n2856 = n2854 ^ x74 ;
  assign n2857 = n2855 & n2856 ;
  assign n2858 = n2857 ^ x74 ;
  assign n2774 = n2663 & n2742 ;
  assign n2775 = n2774 ^ n2591 ;
  assign n2859 = n2858 ^ n2775 ;
  assign n2860 = n2858 ^ x75 ;
  assign n2861 = n2859 & n2860 ;
  assign n2862 = n2861 ^ x75 ;
  assign n2772 = n2667 & n2742 ;
  assign n2773 = n2772 ^ n2589 ;
  assign n2863 = n2862 ^ n2773 ;
  assign n2864 = n2862 ^ x76 ;
  assign n2865 = n2863 & n2864 ;
  assign n2866 = n2865 ^ x76 ;
  assign n2770 = n2671 & n2742 ;
  assign n2771 = n2770 ^ n2587 ;
  assign n2867 = n2866 ^ n2771 ;
  assign n2868 = n2866 ^ x77 ;
  assign n2869 = n2867 & n2868 ;
  assign n2870 = n2869 ^ x77 ;
  assign n2768 = n2675 & n2742 ;
  assign n2769 = n2768 ^ n2585 ;
  assign n2871 = n2870 ^ n2769 ;
  assign n2872 = n2870 ^ x78 ;
  assign n2873 = n2871 & n2872 ;
  assign n2874 = n2873 ^ x78 ;
  assign n2766 = n2679 & n2742 ;
  assign n2767 = n2766 ^ n2583 ;
  assign n2875 = n2874 ^ n2767 ;
  assign n2876 = n2874 ^ x79 ;
  assign n2877 = n2875 & n2876 ;
  assign n2878 = n2877 ^ x79 ;
  assign n2879 = n2878 ^ n2764 ;
  assign n2880 = ~n2765 & n2879 ;
  assign n2881 = n2880 ^ x80 ;
  assign n2882 = n2881 ^ n2761 ;
  assign n2883 = ~n2762 & n2882 ;
  assign n2884 = n2883 ^ x81 ;
  assign n2758 = n2691 & n2742 ;
  assign n2759 = n2758 ^ n2577 ;
  assign n2885 = n2884 ^ n2759 ;
  assign n2886 = n2884 ^ x82 ;
  assign n2887 = n2885 & n2886 ;
  assign n2888 = n2887 ^ x82 ;
  assign n2756 = n2695 & n2742 ;
  assign n2757 = n2756 ^ n2575 ;
  assign n2889 = n2888 ^ n2757 ;
  assign n2890 = n2888 ^ x83 ;
  assign n2891 = n2889 & n2890 ;
  assign n2892 = n2891 ^ x83 ;
  assign n2754 = n2699 & n2742 ;
  assign n2755 = n2754 ^ n2573 ;
  assign n2893 = n2892 ^ n2755 ;
  assign n2894 = n2892 ^ x84 ;
  assign n2895 = n2893 & n2894 ;
  assign n2896 = n2895 ^ x84 ;
  assign n2752 = n2703 & n2742 ;
  assign n2753 = n2752 ^ n2571 ;
  assign n2897 = n2896 ^ n2753 ;
  assign n2898 = n2896 ^ x85 ;
  assign n2899 = n2897 & n2898 ;
  assign n2900 = n2899 ^ x85 ;
  assign n2750 = n2707 & n2742 ;
  assign n2751 = n2750 ^ n2569 ;
  assign n2901 = n2900 ^ n2751 ;
  assign n2902 = n2900 ^ x86 ;
  assign n2903 = n2901 & n2902 ;
  assign n2904 = n2903 ^ x86 ;
  assign n2748 = n2711 & n2742 ;
  assign n2749 = n2748 ^ n2567 ;
  assign n2905 = n2904 ^ n2749 ;
  assign n2906 = n2904 ^ x87 ;
  assign n2907 = n2905 & n2906 ;
  assign n2908 = n2907 ^ x87 ;
  assign n2746 = n2715 & n2742 ;
  assign n2747 = n2746 ^ n2565 ;
  assign n2909 = n2908 ^ n2747 ;
  assign n2910 = n2908 ^ x88 ;
  assign n2911 = n2909 & n2910 ;
  assign n2912 = n2911 ^ x88 ;
  assign n2913 = n2912 ^ n2744 ;
  assign n2914 = ~n2745 & n2913 ;
  assign n2915 = n2914 ^ x89 ;
  assign n2916 = n2915 ^ n2729 ;
  assign n2918 = n2917 ^ n2916 ;
  assign n2919 = n2723 & n2742 ;
  assign n2920 = n2919 ^ n2560 ;
  assign n2921 = n2920 ^ n2729 ;
  assign n2922 = n2921 ^ n2917 ;
  assign n2923 = n2918 & ~n2922 ;
  assign n2924 = n2923 ^ n2917 ;
  assign n2925 = ~n2730 & n2924 ;
  assign n2926 = n2925 ^ x91 ;
  assign n2927 = n165 & ~n2926 ;
  assign n3094 = n2915 ^ x90 ;
  assign n3095 = n2927 & n3094 ;
  assign n3096 = n3095 ^ n2920 ;
  assign n3098 = x91 & ~n3096 ;
  assign n3097 = n3096 ^ x91 ;
  assign n3099 = n3098 ^ n3097 ;
  assign n3091 = n2729 & ~n2927 ;
  assign n3092 = n3091 ^ n270 ;
  assign n3093 = n3092 ^ x92 ;
  assign n3100 = n3099 ^ n3093 ;
  assign n2928 = n2910 & n2927 ;
  assign n2929 = n2928 ^ n2747 ;
  assign n2930 = n2929 ^ x89 ;
  assign n2931 = n2906 & n2927 ;
  assign n2932 = n2931 ^ n2749 ;
  assign n2933 = n2932 ^ x88 ;
  assign n2937 = n2932 ^ x87 ;
  assign n2934 = n2902 & n2927 ;
  assign n2935 = n2934 ^ n2751 ;
  assign n2936 = n2935 ^ n2932 ;
  assign n2938 = n2937 ^ n2936 ;
  assign n3009 = n2836 & n2927 ;
  assign n3010 = n3009 ^ n2798 ;
  assign n2971 = n2829 & n2927 ;
  assign n2972 = n2971 ^ n2831 ;
  assign n2973 = n2972 ^ x69 ;
  assign n2977 = n2972 ^ x68 ;
  assign n2974 = n2826 & n2927 ;
  assign n2975 = n2974 ^ n2801 ;
  assign n2976 = n2975 ^ n2972 ;
  assign n2978 = n2977 ^ n2976 ;
  assign n2989 = ~x35 & x64 ;
  assign n2990 = n2989 ^ x65 ;
  assign n2991 = x64 & n2927 ;
  assign n2992 = n2991 ^ n2814 ;
  assign n2993 = n2990 & ~n2992 ;
  assign n2994 = n2993 ^ x65 ;
  assign n2987 = x64 & n2742 ;
  assign n2983 = ~x36 & x64 ;
  assign n2984 = n2983 ^ x65 ;
  assign n2985 = n2927 & n2984 ;
  assign n2986 = n2985 ^ x37 ;
  assign n2988 = n2987 ^ n2986 ;
  assign n2995 = n2994 ^ n2988 ;
  assign n2996 = n2994 ^ x66 ;
  assign n2997 = n2995 & n2996 ;
  assign n2998 = n2997 ^ x66 ;
  assign n2979 = n2821 ^ x66 ;
  assign n2980 = n2927 & n2979 ;
  assign n2981 = n2980 ^ n2808 ;
  assign n2999 = n2998 ^ n2981 ;
  assign n3000 = n2998 ^ x67 ;
  assign n3001 = n2999 & n3000 ;
  assign n3002 = n3001 ^ x67 ;
  assign n3003 = n3002 ^ n2972 ;
  assign n3004 = n3003 ^ n2977 ;
  assign n3005 = ~n2978 & n3004 ;
  assign n3006 = n3005 ^ n2977 ;
  assign n3007 = ~n2973 & n3006 ;
  assign n3008 = n3007 ^ x69 ;
  assign n3011 = n3010 ^ n3008 ;
  assign n3012 = n3010 ^ x70 ;
  assign n3013 = n3011 & ~n3012 ;
  assign n3014 = n3013 ^ x70 ;
  assign n2969 = n2840 & n2927 ;
  assign n2970 = n2969 ^ n2796 ;
  assign n3015 = n3014 ^ n2970 ;
  assign n3016 = n3014 ^ x71 ;
  assign n3017 = n3015 & n3016 ;
  assign n3018 = n3017 ^ x71 ;
  assign n2967 = n2844 & n2927 ;
  assign n2968 = n2967 ^ n2794 ;
  assign n3019 = n3018 ^ n2968 ;
  assign n3020 = n3018 ^ x72 ;
  assign n3021 = n3019 & n3020 ;
  assign n3022 = n3021 ^ x72 ;
  assign n2965 = n2848 & n2927 ;
  assign n2966 = n2965 ^ n2792 ;
  assign n3023 = n3022 ^ n2966 ;
  assign n3024 = n3022 ^ x73 ;
  assign n3025 = n3023 & n3024 ;
  assign n3026 = n3025 ^ x73 ;
  assign n2963 = n2852 & n2927 ;
  assign n2964 = n2963 ^ n2789 ;
  assign n3027 = n3026 ^ n2964 ;
  assign n3028 = n3026 ^ x74 ;
  assign n3029 = n3027 & n3028 ;
  assign n3030 = n3029 ^ x74 ;
  assign n2961 = n2856 & n2927 ;
  assign n2962 = n2961 ^ n2778 ;
  assign n3031 = n3030 ^ n2962 ;
  assign n3032 = n3030 ^ x75 ;
  assign n3033 = n3031 & n3032 ;
  assign n3034 = n3033 ^ x75 ;
  assign n3035 = n3034 ^ x76 ;
  assign n3036 = n2860 & n2927 ;
  assign n3037 = n3036 ^ n2775 ;
  assign n3038 = n3037 ^ n3034 ;
  assign n3039 = n3035 & n3038 ;
  assign n3040 = n3039 ^ x76 ;
  assign n2959 = n2864 & n2927 ;
  assign n2960 = n2959 ^ n2773 ;
  assign n3041 = n3040 ^ n2960 ;
  assign n3042 = n3040 ^ x77 ;
  assign n3043 = n3041 & n3042 ;
  assign n3044 = n3043 ^ x77 ;
  assign n2957 = n2868 & n2927 ;
  assign n2958 = n2957 ^ n2771 ;
  assign n3045 = n3044 ^ n2958 ;
  assign n3046 = n3044 ^ x78 ;
  assign n3047 = n3045 & n3046 ;
  assign n3048 = n3047 ^ x78 ;
  assign n2955 = n2872 & n2927 ;
  assign n2956 = n2955 ^ n2769 ;
  assign n3049 = n3048 ^ n2956 ;
  assign n3050 = n3048 ^ x79 ;
  assign n3051 = n3049 & n3050 ;
  assign n3052 = n3051 ^ x79 ;
  assign n2953 = n2876 & n2927 ;
  assign n2954 = n2953 ^ n2767 ;
  assign n3053 = n3052 ^ n2954 ;
  assign n3054 = n3052 ^ x80 ;
  assign n3055 = n3053 & n3054 ;
  assign n3056 = n3055 ^ x80 ;
  assign n2950 = n2878 ^ x80 ;
  assign n2951 = n2927 & n2950 ;
  assign n2952 = n2951 ^ n2764 ;
  assign n3057 = n3056 ^ n2952 ;
  assign n3058 = n3056 ^ x81 ;
  assign n3059 = n3057 & n3058 ;
  assign n3060 = n3059 ^ x81 ;
  assign n2947 = n2881 ^ x81 ;
  assign n2948 = n2927 & n2947 ;
  assign n2949 = n2948 ^ n2761 ;
  assign n3061 = n3060 ^ n2949 ;
  assign n3062 = n3060 ^ x82 ;
  assign n3063 = n3061 & n3062 ;
  assign n3064 = n3063 ^ x82 ;
  assign n2945 = n2886 & n2927 ;
  assign n2946 = n2945 ^ n2759 ;
  assign n3065 = n3064 ^ n2946 ;
  assign n3066 = n3064 ^ x83 ;
  assign n3067 = n3065 & n3066 ;
  assign n3068 = n3067 ^ x83 ;
  assign n2943 = n2890 & n2927 ;
  assign n2944 = n2943 ^ n2757 ;
  assign n3069 = n3068 ^ n2944 ;
  assign n3070 = n3068 ^ x84 ;
  assign n3071 = n3069 & n3070 ;
  assign n3072 = n3071 ^ x84 ;
  assign n2941 = n2894 & n2927 ;
  assign n2942 = n2941 ^ n2755 ;
  assign n3073 = n3072 ^ n2942 ;
  assign n3074 = n3072 ^ x85 ;
  assign n3075 = n3073 & n3074 ;
  assign n3076 = n3075 ^ x85 ;
  assign n2939 = n2898 & n2927 ;
  assign n2940 = n2939 ^ n2753 ;
  assign n3077 = n3076 ^ n2940 ;
  assign n3078 = n3076 ^ x86 ;
  assign n3079 = n3077 & n3078 ;
  assign n3080 = n3079 ^ x86 ;
  assign n3081 = n3080 ^ n2932 ;
  assign n3082 = n3081 ^ n2937 ;
  assign n3083 = ~n2938 & n3082 ;
  assign n3084 = n3083 ^ n2937 ;
  assign n3085 = ~n2933 & n3084 ;
  assign n3086 = n3085 ^ x88 ;
  assign n3087 = n3086 ^ n2929 ;
  assign n3088 = ~n2930 & n3087 ;
  assign n3089 = n3088 ^ x89 ;
  assign n3090 = n3089 ^ x90 ;
  assign n3101 = n2912 ^ x89 ;
  assign n3102 = n2927 & n3101 ;
  assign n3103 = n3102 ^ n2744 ;
  assign n3104 = n3103 ^ n3089 ;
  assign n3105 = n3090 & n3104 ;
  assign n3106 = n3105 ^ x90 ;
  assign n3107 = ~n3100 & n3106 ;
  assign n3108 = n164 & ~n3107 ;
  assign n3109 = n3098 ^ n3092 ;
  assign n3110 = n3098 ^ x92 ;
  assign n3111 = ~n3109 & n3110 ;
  assign n3112 = n3111 ^ n3098 ;
  assign n3113 = n3108 & ~n3112 ;
  assign n3309 = n3106 ^ x91 ;
  assign n3310 = n3113 & n3309 ;
  assign n3311 = n3310 ^ n3096 ;
  assign n3114 = n3090 & n3113 ;
  assign n3115 = n3114 ^ n3103 ;
  assign n3116 = n3115 ^ x91 ;
  assign n3121 = n3115 ^ x90 ;
  assign n3117 = n3086 ^ x89 ;
  assign n3118 = n3113 & n3117 ;
  assign n3119 = n3118 ^ n2929 ;
  assign n3120 = n3119 ^ n3115 ;
  assign n3122 = n3121 ^ n3120 ;
  assign n3251 = n3042 & n3113 ;
  assign n3252 = n3251 ^ n2960 ;
  assign n3153 = n3035 & n3113 ;
  assign n3154 = n3153 ^ n3037 ;
  assign n3155 = n3154 ^ x77 ;
  assign n3159 = n3154 ^ x76 ;
  assign n3156 = n3032 & n3113 ;
  assign n3157 = n3156 ^ n2962 ;
  assign n3158 = n3157 ^ n3154 ;
  assign n3160 = n3159 ^ n3158 ;
  assign n3200 = x35 & x65 ;
  assign n3197 = x65 ^ x34 ;
  assign n3193 = x64 ^ x35 ;
  assign n3194 = n3193 ^ x65 ;
  assign n3198 = n3194 ^ n3113 ;
  assign n3199 = ~n3197 & n3198 ;
  assign n3201 = n3200 ^ n3199 ;
  assign n3202 = x64 & n3201 ;
  assign n3203 = n3202 ^ n3200 ;
  assign n3204 = n3203 ^ x65 ;
  assign n3191 = n2990 & n3113 ;
  assign n3190 = n2991 ^ x36 ;
  assign n3192 = n3191 ^ n3190 ;
  assign n3205 = n3204 ^ n3192 ;
  assign n3206 = n3204 ^ x66 ;
  assign n3207 = n3205 & n3206 ;
  assign n3208 = n3207 ^ x66 ;
  assign n3188 = n2996 & n3113 ;
  assign n3189 = n3188 ^ n2988 ;
  assign n3209 = n3208 ^ n3189 ;
  assign n3210 = n3208 ^ x67 ;
  assign n3211 = n3209 & n3210 ;
  assign n3212 = n3211 ^ x67 ;
  assign n3186 = n3000 & n3113 ;
  assign n3187 = n3186 ^ n2981 ;
  assign n3213 = n3212 ^ n3187 ;
  assign n3214 = n3212 ^ x68 ;
  assign n3215 = n3213 & n3214 ;
  assign n3216 = n3215 ^ x68 ;
  assign n3183 = n3002 ^ x68 ;
  assign n3184 = n3113 & n3183 ;
  assign n3185 = n3184 ^ n2975 ;
  assign n3217 = n3216 ^ n3185 ;
  assign n3218 = n3216 ^ x69 ;
  assign n3219 = n3217 & n3218 ;
  assign n3220 = n3219 ^ x69 ;
  assign n3172 = n2975 ^ x69 ;
  assign n3173 = n3172 ^ n3002 ;
  assign n3174 = n3173 ^ x68 ;
  assign n3175 = n3174 ^ n3172 ;
  assign n3177 = n3002 ^ x69 ;
  assign n3178 = n3177 ^ n3172 ;
  assign n3179 = ~n3175 & ~n3178 ;
  assign n3180 = n3179 ^ n3172 ;
  assign n3181 = n3113 & ~n3180 ;
  assign n3182 = n3181 ^ n2972 ;
  assign n3221 = n3220 ^ n3182 ;
  assign n3222 = n3220 ^ x70 ;
  assign n3223 = n3221 & n3222 ;
  assign n3224 = n3223 ^ x70 ;
  assign n3169 = n3008 ^ x70 ;
  assign n3170 = n3113 & n3169 ;
  assign n3171 = n3170 ^ n3010 ;
  assign n3225 = n3224 ^ n3171 ;
  assign n3226 = n3224 ^ x71 ;
  assign n3227 = n3225 & n3226 ;
  assign n3228 = n3227 ^ x71 ;
  assign n3167 = n3016 & n3113 ;
  assign n3168 = n3167 ^ n2970 ;
  assign n3229 = n3228 ^ n3168 ;
  assign n3230 = n3228 ^ x72 ;
  assign n3231 = n3229 & n3230 ;
  assign n3232 = n3231 ^ x72 ;
  assign n3165 = n3020 & n3113 ;
  assign n3166 = n3165 ^ n2968 ;
  assign n3233 = n3232 ^ n3166 ;
  assign n3234 = n3232 ^ x73 ;
  assign n3235 = n3233 & n3234 ;
  assign n3236 = n3235 ^ x73 ;
  assign n3163 = n3024 & n3113 ;
  assign n3164 = n3163 ^ n2966 ;
  assign n3237 = n3236 ^ n3164 ;
  assign n3238 = n3236 ^ x74 ;
  assign n3239 = n3237 & n3238 ;
  assign n3240 = n3239 ^ x74 ;
  assign n3161 = n3028 & n3113 ;
  assign n3162 = n3161 ^ n2964 ;
  assign n3241 = n3240 ^ n3162 ;
  assign n3242 = n3240 ^ x75 ;
  assign n3243 = n3241 & n3242 ;
  assign n3244 = n3243 ^ x75 ;
  assign n3245 = n3244 ^ n3154 ;
  assign n3246 = n3245 ^ n3159 ;
  assign n3247 = ~n3160 & n3246 ;
  assign n3248 = n3247 ^ n3159 ;
  assign n3249 = ~n3155 & n3248 ;
  assign n3250 = n3249 ^ x77 ;
  assign n3253 = n3252 ^ n3250 ;
  assign n3254 = n3252 ^ x78 ;
  assign n3255 = n3253 & ~n3254 ;
  assign n3256 = n3255 ^ x78 ;
  assign n3151 = n3046 & n3113 ;
  assign n3152 = n3151 ^ n2958 ;
  assign n3257 = n3256 ^ n3152 ;
  assign n3258 = n3256 ^ x79 ;
  assign n3259 = n3257 & n3258 ;
  assign n3260 = n3259 ^ x79 ;
  assign n3149 = n3050 & n3113 ;
  assign n3150 = n3149 ^ n2956 ;
  assign n3261 = n3260 ^ n3150 ;
  assign n3262 = n3260 ^ x80 ;
  assign n3263 = n3261 & n3262 ;
  assign n3264 = n3263 ^ x80 ;
  assign n3147 = n3054 & n3113 ;
  assign n3148 = n3147 ^ n2954 ;
  assign n3265 = n3264 ^ n3148 ;
  assign n3266 = n3264 ^ x81 ;
  assign n3267 = n3265 & n3266 ;
  assign n3268 = n3267 ^ x81 ;
  assign n3145 = n3058 & n3113 ;
  assign n3146 = n3145 ^ n2952 ;
  assign n3269 = n3268 ^ n3146 ;
  assign n3270 = n3268 ^ x82 ;
  assign n3271 = n3269 & n3270 ;
  assign n3272 = n3271 ^ x82 ;
  assign n3273 = n3272 ^ x83 ;
  assign n3274 = n3062 & n3113 ;
  assign n3275 = n3274 ^ n2949 ;
  assign n3276 = n3275 ^ n3272 ;
  assign n3277 = n3273 & n3276 ;
  assign n3278 = n3277 ^ x83 ;
  assign n3143 = n3066 & n3113 ;
  assign n3144 = n3143 ^ n2946 ;
  assign n3279 = n3278 ^ n3144 ;
  assign n3280 = n3278 ^ x84 ;
  assign n3281 = n3279 & n3280 ;
  assign n3282 = n3281 ^ x84 ;
  assign n3141 = n3070 & n3113 ;
  assign n3142 = n3141 ^ n2944 ;
  assign n3283 = n3282 ^ n3142 ;
  assign n3284 = n3282 ^ x85 ;
  assign n3285 = n3283 & n3284 ;
  assign n3286 = n3285 ^ x85 ;
  assign n3139 = n3074 & n3113 ;
  assign n3140 = n3139 ^ n2942 ;
  assign n3287 = n3286 ^ n3140 ;
  assign n3288 = n3286 ^ x86 ;
  assign n3289 = n3287 & n3288 ;
  assign n3290 = n3289 ^ x86 ;
  assign n3137 = n3078 & n3113 ;
  assign n3138 = n3137 ^ n2940 ;
  assign n3291 = n3290 ^ n3138 ;
  assign n3292 = n3290 ^ x87 ;
  assign n3293 = n3291 & n3292 ;
  assign n3294 = n3293 ^ x87 ;
  assign n3134 = n3080 ^ x87 ;
  assign n3135 = n3113 & n3134 ;
  assign n3136 = n3135 ^ n2935 ;
  assign n3295 = n3294 ^ n3136 ;
  assign n3296 = n3294 ^ x88 ;
  assign n3297 = n3295 & n3296 ;
  assign n3298 = n3297 ^ x88 ;
  assign n3123 = n2935 ^ x88 ;
  assign n3124 = n3123 ^ n3080 ;
  assign n3125 = n3124 ^ x87 ;
  assign n3126 = n3125 ^ n3123 ;
  assign n3128 = n3080 ^ x88 ;
  assign n3129 = n3128 ^ n3123 ;
  assign n3130 = ~n3126 & ~n3129 ;
  assign n3131 = n3130 ^ n3123 ;
  assign n3132 = n3113 & ~n3131 ;
  assign n3133 = n3132 ^ n2932 ;
  assign n3299 = n3298 ^ n3133 ;
  assign n3300 = n3298 ^ x89 ;
  assign n3301 = n3299 & n3300 ;
  assign n3302 = n3301 ^ x89 ;
  assign n3303 = n3302 ^ n3115 ;
  assign n3304 = n3303 ^ n3121 ;
  assign n3305 = ~n3122 & n3304 ;
  assign n3306 = n3305 ^ n3121 ;
  assign n3307 = ~n3116 & n3306 ;
  assign n3308 = n3307 ^ x91 ;
  assign n3312 = n3311 ^ n3308 ;
  assign n3313 = n3311 ^ x92 ;
  assign n3314 = n3312 & ~n3313 ;
  assign n3315 = n3314 ^ x92 ;
  assign n3318 = n3091 & ~n3113 ;
  assign n3319 = n3318 ^ n270 ;
  assign n3538 = n163 & n3319 ;
  assign n3539 = n3315 & n3538 ;
  assign n3540 = x93 & n3539 ;
  assign n3541 = n3540 ^ n3538 ;
  assign n3542 = n3541 ^ n3319 ;
  assign n3547 = ~x94 & ~n3542 ;
  assign n3316 = n3315 ^ x93 ;
  assign n3320 = n3319 ^ x93 ;
  assign n3321 = n3316 & ~n3320 ;
  assign n3322 = n3321 ^ x93 ;
  assign n3323 = n163 & ~n3322 ;
  assign n3529 = n3308 ^ x92 ;
  assign n3530 = n3323 & n3529 ;
  assign n3531 = n3530 ^ n3311 ;
  assign n3492 = n3280 & n3323 ;
  assign n3493 = n3492 ^ n3144 ;
  assign n3348 = n3273 & n3323 ;
  assign n3349 = n3348 ^ n3275 ;
  assign n3350 = n3349 ^ x84 ;
  assign n3354 = n3349 ^ x83 ;
  assign n3351 = n3270 & n3323 ;
  assign n3352 = n3351 ^ n3146 ;
  assign n3353 = n3352 ^ n3349 ;
  assign n3355 = n3354 ^ n3353 ;
  assign n3413 = x34 & x65 ;
  assign n3410 = x65 ^ x33 ;
  assign n3406 = x64 ^ x34 ;
  assign n3407 = n3406 ^ x65 ;
  assign n3411 = n3407 ^ n3323 ;
  assign n3412 = ~n3410 & n3411 ;
  assign n3414 = n3413 ^ n3412 ;
  assign n3415 = x64 & n3414 ;
  assign n3416 = n3415 ^ n3413 ;
  assign n3417 = n3416 ^ x65 ;
  assign n3404 = x64 & n3113 ;
  assign n3400 = ~x34 & x64 ;
  assign n3401 = n3400 ^ x65 ;
  assign n3402 = n3323 & n3401 ;
  assign n3403 = n3402 ^ x35 ;
  assign n3405 = n3404 ^ n3403 ;
  assign n3418 = n3417 ^ n3405 ;
  assign n3419 = n3417 ^ x66 ;
  assign n3420 = n3418 & n3419 ;
  assign n3421 = n3420 ^ x66 ;
  assign n3397 = n3206 & n3323 ;
  assign n3398 = n3397 ^ n3192 ;
  assign n3422 = n3421 ^ n3398 ;
  assign n3423 = n3421 ^ x67 ;
  assign n3424 = n3422 & n3423 ;
  assign n3425 = n3424 ^ x67 ;
  assign n3395 = n3210 & n3323 ;
  assign n3396 = n3395 ^ n3189 ;
  assign n3426 = n3425 ^ n3396 ;
  assign n3427 = n3425 ^ x68 ;
  assign n3428 = n3426 & n3427 ;
  assign n3429 = n3428 ^ x68 ;
  assign n3393 = n3214 & n3323 ;
  assign n3394 = n3393 ^ n3187 ;
  assign n3430 = n3429 ^ n3394 ;
  assign n3431 = n3429 ^ x69 ;
  assign n3432 = n3430 & n3431 ;
  assign n3433 = n3432 ^ x69 ;
  assign n3391 = n3218 & n3323 ;
  assign n3392 = n3391 ^ n3185 ;
  assign n3434 = n3433 ^ n3392 ;
  assign n3435 = n3433 ^ x70 ;
  assign n3436 = n3434 & n3435 ;
  assign n3437 = n3436 ^ x70 ;
  assign n3389 = n3222 & n3323 ;
  assign n3390 = n3389 ^ n3182 ;
  assign n3438 = n3437 ^ n3390 ;
  assign n3439 = n3437 ^ x71 ;
  assign n3440 = n3438 & n3439 ;
  assign n3441 = n3440 ^ x71 ;
  assign n3387 = n3226 & n3323 ;
  assign n3388 = n3387 ^ n3171 ;
  assign n3442 = n3441 ^ n3388 ;
  assign n3443 = n3441 ^ x72 ;
  assign n3444 = n3442 & n3443 ;
  assign n3445 = n3444 ^ x72 ;
  assign n3385 = n3230 & n3323 ;
  assign n3386 = n3385 ^ n3168 ;
  assign n3446 = n3445 ^ n3386 ;
  assign n3447 = n3445 ^ x73 ;
  assign n3448 = n3446 & n3447 ;
  assign n3449 = n3448 ^ x73 ;
  assign n3383 = n3234 & n3323 ;
  assign n3384 = n3383 ^ n3166 ;
  assign n3450 = n3449 ^ n3384 ;
  assign n3451 = n3449 ^ x74 ;
  assign n3452 = n3450 & n3451 ;
  assign n3453 = n3452 ^ x74 ;
  assign n3381 = n3238 & n3323 ;
  assign n3382 = n3381 ^ n3164 ;
  assign n3454 = n3453 ^ n3382 ;
  assign n3455 = n3453 ^ x75 ;
  assign n3456 = n3454 & n3455 ;
  assign n3457 = n3456 ^ x75 ;
  assign n3379 = n3242 & n3323 ;
  assign n3380 = n3379 ^ n3162 ;
  assign n3458 = n3457 ^ n3380 ;
  assign n3459 = n3457 ^ x76 ;
  assign n3460 = n3458 & n3459 ;
  assign n3461 = n3460 ^ x76 ;
  assign n3376 = n3244 ^ x76 ;
  assign n3377 = n3323 & n3376 ;
  assign n3378 = n3377 ^ n3157 ;
  assign n3462 = n3461 ^ n3378 ;
  assign n3463 = n3461 ^ x77 ;
  assign n3464 = n3462 & n3463 ;
  assign n3465 = n3464 ^ x77 ;
  assign n3365 = n3157 ^ x77 ;
  assign n3366 = n3365 ^ n3244 ;
  assign n3367 = n3366 ^ x76 ;
  assign n3368 = n3367 ^ n3365 ;
  assign n3370 = n3244 ^ x77 ;
  assign n3371 = n3370 ^ n3365 ;
  assign n3372 = ~n3368 & ~n3371 ;
  assign n3373 = n3372 ^ n3365 ;
  assign n3374 = n3323 & ~n3373 ;
  assign n3375 = n3374 ^ n3154 ;
  assign n3466 = n3465 ^ n3375 ;
  assign n3467 = n3465 ^ x78 ;
  assign n3468 = n3466 & n3467 ;
  assign n3469 = n3468 ^ x78 ;
  assign n3362 = n3250 ^ x78 ;
  assign n3363 = n3323 & n3362 ;
  assign n3364 = n3363 ^ n3252 ;
  assign n3470 = n3469 ^ n3364 ;
  assign n3471 = n3469 ^ x79 ;
  assign n3472 = n3470 & n3471 ;
  assign n3473 = n3472 ^ x79 ;
  assign n3360 = n3258 & n3323 ;
  assign n3361 = n3360 ^ n3152 ;
  assign n3474 = n3473 ^ n3361 ;
  assign n3475 = n3473 ^ x80 ;
  assign n3476 = n3474 & n3475 ;
  assign n3477 = n3476 ^ x80 ;
  assign n3358 = n3262 & n3323 ;
  assign n3359 = n3358 ^ n3150 ;
  assign n3478 = n3477 ^ n3359 ;
  assign n3479 = n3477 ^ x81 ;
  assign n3480 = n3478 & n3479 ;
  assign n3481 = n3480 ^ x81 ;
  assign n3356 = n3266 & n3323 ;
  assign n3357 = n3356 ^ n3148 ;
  assign n3482 = n3481 ^ n3357 ;
  assign n3483 = n3481 ^ x82 ;
  assign n3484 = n3482 & n3483 ;
  assign n3485 = n3484 ^ x82 ;
  assign n3486 = n3485 ^ n3349 ;
  assign n3487 = n3486 ^ n3354 ;
  assign n3488 = ~n3355 & n3487 ;
  assign n3489 = n3488 ^ n3354 ;
  assign n3490 = ~n3350 & n3489 ;
  assign n3491 = n3490 ^ x84 ;
  assign n3494 = n3493 ^ n3491 ;
  assign n3495 = n3493 ^ x85 ;
  assign n3496 = n3494 & ~n3495 ;
  assign n3497 = n3496 ^ x85 ;
  assign n3346 = n3284 & n3323 ;
  assign n3347 = n3346 ^ n3142 ;
  assign n3498 = n3497 ^ n3347 ;
  assign n3499 = n3497 ^ x86 ;
  assign n3500 = n3498 & n3499 ;
  assign n3501 = n3500 ^ x86 ;
  assign n3344 = n3288 & n3323 ;
  assign n3345 = n3344 ^ n3140 ;
  assign n3502 = n3501 ^ n3345 ;
  assign n3503 = n3501 ^ x87 ;
  assign n3504 = n3502 & n3503 ;
  assign n3505 = n3504 ^ x87 ;
  assign n3342 = n3292 & n3323 ;
  assign n3343 = n3342 ^ n3138 ;
  assign n3506 = n3505 ^ n3343 ;
  assign n3507 = n3505 ^ x88 ;
  assign n3508 = n3506 & n3507 ;
  assign n3509 = n3508 ^ x88 ;
  assign n3340 = n3296 & n3323 ;
  assign n3341 = n3340 ^ n3136 ;
  assign n3510 = n3509 ^ n3341 ;
  assign n3511 = n3509 ^ x89 ;
  assign n3512 = n3510 & n3511 ;
  assign n3513 = n3512 ^ x89 ;
  assign n3338 = n3300 & n3323 ;
  assign n3339 = n3338 ^ n3133 ;
  assign n3514 = n3513 ^ n3339 ;
  assign n3515 = n3513 ^ x90 ;
  assign n3516 = n3514 & n3515 ;
  assign n3517 = n3516 ^ x90 ;
  assign n3335 = n3302 ^ x90 ;
  assign n3336 = n3323 & n3335 ;
  assign n3337 = n3336 ^ n3119 ;
  assign n3518 = n3517 ^ n3337 ;
  assign n3519 = n3517 ^ x91 ;
  assign n3520 = n3518 & n3519 ;
  assign n3521 = n3520 ^ x91 ;
  assign n3324 = n3119 ^ x91 ;
  assign n3325 = n3324 ^ n3302 ;
  assign n3326 = n3325 ^ x90 ;
  assign n3327 = n3326 ^ n3324 ;
  assign n3329 = n3302 ^ x91 ;
  assign n3330 = n3329 ^ n3324 ;
  assign n3331 = ~n3327 & ~n3330 ;
  assign n3332 = n3331 ^ n3324 ;
  assign n3333 = n3323 & ~n3332 ;
  assign n3334 = n3333 ^ n3115 ;
  assign n3522 = n3521 ^ n3334 ;
  assign n3525 = n3334 ^ x92 ;
  assign n3526 = n3522 & ~n3525 ;
  assign n3523 = x93 ^ x92 ;
  assign n3527 = n3526 ^ n3523 ;
  assign n3532 = n3531 ^ n3527 ;
  assign n3533 = n3532 ^ x93 ;
  assign n3528 = n3527 ^ x94 ;
  assign n3534 = n3533 ^ n3528 ;
  assign n3548 = n3547 ^ n3534 ;
  assign n3550 = n3533 ^ n3531 ;
  assign n3552 = n3532 & n3550 ;
  assign n3553 = n3552 ^ n3531 ;
  assign n3554 = n3548 & ~n3553 ;
  assign n3555 = n3554 ^ n3531 ;
  assign n3556 = n162 & n3555 ;
  assign n3557 = x94 & ~n3319 ;
  assign n3558 = n3556 & n3557 ;
  assign n3559 = n3558 ^ n3556 ;
  assign n3560 = n3542 & ~n3559 ;
  assign n3561 = n3560 ^ n270 ;
  assign n3562 = n3561 ^ x95 ;
  assign n3566 = n3561 ^ x94 ;
  assign n3563 = n3527 & n3559 ;
  assign n3564 = n3563 ^ n3531 ;
  assign n3565 = n3564 ^ n3561 ;
  assign n3567 = n3566 ^ n3565 ;
  assign n3735 = n3499 & n3559 ;
  assign n3736 = n3735 ^ n3347 ;
  assign n3581 = n3491 ^ x85 ;
  assign n3582 = n3559 & n3581 ;
  assign n3583 = n3582 ^ n3493 ;
  assign n3584 = n3583 ^ x86 ;
  assign n3597 = n3583 ^ x85 ;
  assign n3585 = n3352 ^ x84 ;
  assign n3586 = n3585 ^ n3485 ;
  assign n3587 = n3586 ^ x83 ;
  assign n3588 = n3587 ^ n3585 ;
  assign n3590 = n3485 ^ x84 ;
  assign n3591 = n3590 ^ n3585 ;
  assign n3592 = ~n3588 & ~n3591 ;
  assign n3593 = n3592 ^ n3585 ;
  assign n3594 = n3559 & ~n3593 ;
  assign n3595 = n3594 ^ n3349 ;
  assign n3596 = n3595 ^ n3583 ;
  assign n3598 = n3597 ^ n3596 ;
  assign n3647 = x64 & n3559 ;
  assign n3646 = x64 & ~x65 ;
  assign n3648 = n3647 ^ n3646 ;
  assign n3649 = n3647 ^ x32 ;
  assign n3650 = n3648 & ~n3649 ;
  assign n3651 = n3650 ^ x65 ;
  assign n3643 = ~x32 & x64 ;
  assign n3644 = n3643 ^ x65 ;
  assign n3645 = x33 & n3644 ;
  assign n3652 = n3651 ^ n3645 ;
  assign n3641 = x64 & n3323 ;
  assign n3637 = ~x33 & x64 ;
  assign n3638 = n3637 ^ x65 ;
  assign n3639 = n3559 & n3638 ;
  assign n3640 = n3639 ^ x34 ;
  assign n3642 = n3641 ^ n3640 ;
  assign n3653 = n3652 ^ n3642 ;
  assign n3654 = n3652 ^ x66 ;
  assign n3655 = n3653 & n3654 ;
  assign n3656 = n3655 ^ x66 ;
  assign n3634 = n3419 & n3559 ;
  assign n3635 = n3634 ^ n3405 ;
  assign n3657 = n3656 ^ n3635 ;
  assign n3658 = n3656 ^ x67 ;
  assign n3659 = n3657 & n3658 ;
  assign n3660 = n3659 ^ x67 ;
  assign n3632 = n3423 & n3559 ;
  assign n3633 = n3632 ^ n3398 ;
  assign n3661 = n3660 ^ n3633 ;
  assign n3662 = n3660 ^ x68 ;
  assign n3663 = n3661 & n3662 ;
  assign n3664 = n3663 ^ x68 ;
  assign n3630 = n3427 & n3559 ;
  assign n3631 = n3630 ^ n3396 ;
  assign n3665 = n3664 ^ n3631 ;
  assign n3666 = n3664 ^ x69 ;
  assign n3667 = n3665 & n3666 ;
  assign n3668 = n3667 ^ x69 ;
  assign n3628 = n3431 & n3559 ;
  assign n3629 = n3628 ^ n3394 ;
  assign n3669 = n3668 ^ n3629 ;
  assign n3670 = n3668 ^ x70 ;
  assign n3671 = n3669 & n3670 ;
  assign n3672 = n3671 ^ x70 ;
  assign n3626 = n3435 & n3559 ;
  assign n3627 = n3626 ^ n3392 ;
  assign n3673 = n3672 ^ n3627 ;
  assign n3674 = n3672 ^ x71 ;
  assign n3675 = n3673 & n3674 ;
  assign n3676 = n3675 ^ x71 ;
  assign n3624 = n3439 & n3559 ;
  assign n3625 = n3624 ^ n3390 ;
  assign n3677 = n3676 ^ n3625 ;
  assign n3678 = n3676 ^ x72 ;
  assign n3679 = n3677 & n3678 ;
  assign n3680 = n3679 ^ x72 ;
  assign n3622 = n3443 & n3559 ;
  assign n3623 = n3622 ^ n3388 ;
  assign n3681 = n3680 ^ n3623 ;
  assign n3682 = n3680 ^ x73 ;
  assign n3683 = n3681 & n3682 ;
  assign n3684 = n3683 ^ x73 ;
  assign n3620 = n3447 & n3559 ;
  assign n3621 = n3620 ^ n3386 ;
  assign n3685 = n3684 ^ n3621 ;
  assign n3686 = n3684 ^ x74 ;
  assign n3687 = n3685 & n3686 ;
  assign n3688 = n3687 ^ x74 ;
  assign n3618 = n3451 & n3559 ;
  assign n3619 = n3618 ^ n3384 ;
  assign n3689 = n3688 ^ n3619 ;
  assign n3690 = n3688 ^ x75 ;
  assign n3691 = n3689 & n3690 ;
  assign n3692 = n3691 ^ x75 ;
  assign n3616 = n3455 & n3559 ;
  assign n3617 = n3616 ^ n3382 ;
  assign n3693 = n3692 ^ n3617 ;
  assign n3694 = n3692 ^ x76 ;
  assign n3695 = n3693 & n3694 ;
  assign n3696 = n3695 ^ x76 ;
  assign n3614 = n3459 & n3559 ;
  assign n3615 = n3614 ^ n3380 ;
  assign n3697 = n3696 ^ n3615 ;
  assign n3698 = n3696 ^ x77 ;
  assign n3699 = n3697 & n3698 ;
  assign n3700 = n3699 ^ x77 ;
  assign n3612 = n3463 & n3559 ;
  assign n3613 = n3612 ^ n3378 ;
  assign n3701 = n3700 ^ n3613 ;
  assign n3702 = n3700 ^ x78 ;
  assign n3703 = n3701 & n3702 ;
  assign n3704 = n3703 ^ x78 ;
  assign n3610 = n3467 & n3559 ;
  assign n3611 = n3610 ^ n3375 ;
  assign n3705 = n3704 ^ n3611 ;
  assign n3706 = n3704 ^ x79 ;
  assign n3707 = n3705 & n3706 ;
  assign n3708 = n3707 ^ x79 ;
  assign n3608 = n3471 & n3559 ;
  assign n3609 = n3608 ^ n3364 ;
  assign n3709 = n3708 ^ n3609 ;
  assign n3710 = n3708 ^ x80 ;
  assign n3711 = n3709 & n3710 ;
  assign n3712 = n3711 ^ x80 ;
  assign n3606 = n3475 & n3559 ;
  assign n3607 = n3606 ^ n3361 ;
  assign n3713 = n3712 ^ n3607 ;
  assign n3714 = n3712 ^ x81 ;
  assign n3715 = n3713 & n3714 ;
  assign n3716 = n3715 ^ x81 ;
  assign n3604 = n3479 & n3559 ;
  assign n3605 = n3604 ^ n3359 ;
  assign n3717 = n3716 ^ n3605 ;
  assign n3718 = n3716 ^ x82 ;
  assign n3719 = n3717 & n3718 ;
  assign n3720 = n3719 ^ x82 ;
  assign n3602 = n3483 & n3559 ;
  assign n3603 = n3602 ^ n3357 ;
  assign n3721 = n3720 ^ n3603 ;
  assign n3722 = n3720 ^ x83 ;
  assign n3723 = n3721 & n3722 ;
  assign n3724 = n3723 ^ x83 ;
  assign n3599 = n3485 ^ x83 ;
  assign n3600 = n3559 & n3599 ;
  assign n3601 = n3600 ^ n3352 ;
  assign n3725 = n3724 ^ n3601 ;
  assign n3726 = n3724 ^ x84 ;
  assign n3727 = n3725 & n3726 ;
  assign n3728 = n3727 ^ x84 ;
  assign n3729 = n3728 ^ n3583 ;
  assign n3730 = n3729 ^ n3597 ;
  assign n3731 = ~n3598 & n3730 ;
  assign n3732 = n3731 ^ n3597 ;
  assign n3733 = ~n3584 & n3732 ;
  assign n3734 = n3733 ^ x86 ;
  assign n3737 = n3736 ^ n3734 ;
  assign n3738 = n3736 ^ x87 ;
  assign n3739 = n3737 & ~n3738 ;
  assign n3740 = n3739 ^ x87 ;
  assign n3579 = n3503 & n3559 ;
  assign n3580 = n3579 ^ n3345 ;
  assign n3741 = n3740 ^ n3580 ;
  assign n3742 = n3740 ^ x88 ;
  assign n3743 = n3741 & n3742 ;
  assign n3744 = n3743 ^ x88 ;
  assign n3577 = n3507 & n3559 ;
  assign n3578 = n3577 ^ n3343 ;
  assign n3745 = n3744 ^ n3578 ;
  assign n3746 = n3744 ^ x89 ;
  assign n3747 = n3745 & n3746 ;
  assign n3748 = n3747 ^ x89 ;
  assign n3575 = n3511 & n3559 ;
  assign n3576 = n3575 ^ n3341 ;
  assign n3749 = n3748 ^ n3576 ;
  assign n3750 = n3748 ^ x90 ;
  assign n3751 = n3749 & n3750 ;
  assign n3752 = n3751 ^ x90 ;
  assign n3573 = n3515 & n3559 ;
  assign n3574 = n3573 ^ n3339 ;
  assign n3753 = n3752 ^ n3574 ;
  assign n3754 = n3752 ^ x91 ;
  assign n3755 = n3753 & n3754 ;
  assign n3756 = n3755 ^ x91 ;
  assign n3571 = n3519 & n3559 ;
  assign n3572 = n3571 ^ n3337 ;
  assign n3757 = n3756 ^ n3572 ;
  assign n3758 = n3756 ^ x92 ;
  assign n3759 = n3757 & n3758 ;
  assign n3760 = n3759 ^ x92 ;
  assign n3568 = n3521 ^ x92 ;
  assign n3569 = n3559 & n3568 ;
  assign n3570 = n3569 ^ n3334 ;
  assign n3761 = n3760 ^ n3570 ;
  assign n3762 = n3760 ^ x93 ;
  assign n3763 = n3761 & n3762 ;
  assign n3764 = n3763 ^ x93 ;
  assign n3765 = n3764 ^ n3561 ;
  assign n3766 = n3765 ^ n3566 ;
  assign n3767 = ~n3567 & n3766 ;
  assign n3768 = n3767 ^ n3566 ;
  assign n3769 = ~n3562 & n3768 ;
  assign n3770 = n3769 ^ x95 ;
  assign n3771 = n161 & ~n3770 ;
  assign n3772 = n3561 & ~n3771 ;
  assign n3773 = n3772 ^ n270 ;
  assign n3776 = x96 & n160 ;
  assign n3919 = n3710 & n3771 ;
  assign n3920 = n3919 ^ n3609 ;
  assign n3814 = n3706 & n3771 ;
  assign n3815 = n3814 ^ n3611 ;
  assign n3816 = n3815 ^ x80 ;
  assign n3820 = n3815 ^ x79 ;
  assign n3817 = n3702 & n3771 ;
  assign n3818 = n3817 ^ n3613 ;
  assign n3819 = n3818 ^ n3815 ;
  assign n3821 = n3820 ^ n3819 ;
  assign n3871 = n3662 & n3771 ;
  assign n3872 = n3871 ^ n3633 ;
  assign n3865 = n3658 & n3771 ;
  assign n3866 = n3865 ^ n3635 ;
  assign n3859 = n3654 & n3771 ;
  assign n3860 = n3859 ^ n3642 ;
  assign n3853 = n3647 ^ x33 ;
  assign n3852 = n3644 & n3771 ;
  assign n3854 = n3853 ^ n3852 ;
  assign n3845 = x32 & x65 ;
  assign n3840 = x65 ^ x31 ;
  assign n3841 = x64 ^ x32 ;
  assign n3842 = n3841 ^ x65 ;
  assign n3843 = n3842 ^ n3771 ;
  assign n3844 = ~n3840 & n3843 ;
  assign n3846 = n3845 ^ n3844 ;
  assign n3849 = x64 & n3846 ;
  assign n3850 = n3849 ^ n3845 ;
  assign n3851 = n3850 ^ x65 ;
  assign n3855 = n3854 ^ n3851 ;
  assign n3856 = n3854 ^ x66 ;
  assign n3857 = n3855 & ~n3856 ;
  assign n3858 = n3857 ^ x66 ;
  assign n3861 = n3860 ^ n3858 ;
  assign n3862 = n3860 ^ x67 ;
  assign n3863 = n3861 & ~n3862 ;
  assign n3864 = n3863 ^ x67 ;
  assign n3867 = n3866 ^ n3864 ;
  assign n3868 = n3866 ^ x68 ;
  assign n3869 = n3867 & ~n3868 ;
  assign n3870 = n3869 ^ x68 ;
  assign n3873 = n3872 ^ n3870 ;
  assign n3874 = n3872 ^ x69 ;
  assign n3875 = n3873 & ~n3874 ;
  assign n3876 = n3875 ^ x69 ;
  assign n3838 = n3666 & n3771 ;
  assign n3839 = n3838 ^ n3631 ;
  assign n3877 = n3876 ^ n3839 ;
  assign n3878 = n3876 ^ x70 ;
  assign n3879 = n3877 & n3878 ;
  assign n3880 = n3879 ^ x70 ;
  assign n3836 = n3670 & n3771 ;
  assign n3837 = n3836 ^ n3629 ;
  assign n3881 = n3880 ^ n3837 ;
  assign n3882 = n3880 ^ x71 ;
  assign n3883 = n3881 & n3882 ;
  assign n3884 = n3883 ^ x71 ;
  assign n3834 = n3674 & n3771 ;
  assign n3835 = n3834 ^ n3627 ;
  assign n3885 = n3884 ^ n3835 ;
  assign n3886 = n3884 ^ x72 ;
  assign n3887 = n3885 & n3886 ;
  assign n3888 = n3887 ^ x72 ;
  assign n3832 = n3678 & n3771 ;
  assign n3833 = n3832 ^ n3625 ;
  assign n3889 = n3888 ^ n3833 ;
  assign n3890 = n3888 ^ x73 ;
  assign n3891 = n3889 & n3890 ;
  assign n3892 = n3891 ^ x73 ;
  assign n3830 = n3682 & n3771 ;
  assign n3831 = n3830 ^ n3623 ;
  assign n3893 = n3892 ^ n3831 ;
  assign n3894 = n3892 ^ x74 ;
  assign n3895 = n3893 & n3894 ;
  assign n3896 = n3895 ^ x74 ;
  assign n3828 = n3686 & n3771 ;
  assign n3829 = n3828 ^ n3621 ;
  assign n3897 = n3896 ^ n3829 ;
  assign n3898 = n3896 ^ x75 ;
  assign n3899 = n3897 & n3898 ;
  assign n3900 = n3899 ^ x75 ;
  assign n3826 = n3690 & n3771 ;
  assign n3827 = n3826 ^ n3619 ;
  assign n3901 = n3900 ^ n3827 ;
  assign n3902 = n3900 ^ x76 ;
  assign n3903 = n3901 & n3902 ;
  assign n3904 = n3903 ^ x76 ;
  assign n3824 = n3694 & n3771 ;
  assign n3825 = n3824 ^ n3617 ;
  assign n3905 = n3904 ^ n3825 ;
  assign n3906 = n3904 ^ x77 ;
  assign n3907 = n3905 & n3906 ;
  assign n3908 = n3907 ^ x77 ;
  assign n3822 = n3698 & n3771 ;
  assign n3823 = n3822 ^ n3615 ;
  assign n3909 = n3908 ^ n3823 ;
  assign n3910 = n3908 ^ x78 ;
  assign n3911 = n3909 & n3910 ;
  assign n3912 = n3911 ^ x78 ;
  assign n3913 = n3912 ^ n3815 ;
  assign n3914 = n3913 ^ n3820 ;
  assign n3915 = ~n3821 & n3914 ;
  assign n3916 = n3915 ^ n3820 ;
  assign n3917 = ~n3816 & n3916 ;
  assign n3918 = n3917 ^ x80 ;
  assign n3921 = n3920 ^ n3918 ;
  assign n3922 = n3920 ^ x81 ;
  assign n3923 = n3921 & ~n3922 ;
  assign n3924 = n3923 ^ x81 ;
  assign n3812 = n3714 & n3771 ;
  assign n3813 = n3812 ^ n3607 ;
  assign n3925 = n3924 ^ n3813 ;
  assign n3926 = n3924 ^ x82 ;
  assign n3927 = n3925 & n3926 ;
  assign n3928 = n3927 ^ x82 ;
  assign n3810 = n3718 & n3771 ;
  assign n3811 = n3810 ^ n3605 ;
  assign n3929 = n3928 ^ n3811 ;
  assign n3930 = n3928 ^ x83 ;
  assign n3931 = n3929 & n3930 ;
  assign n3932 = n3931 ^ x83 ;
  assign n3808 = n3722 & n3771 ;
  assign n3809 = n3808 ^ n3603 ;
  assign n3933 = n3932 ^ n3809 ;
  assign n3934 = n3932 ^ x84 ;
  assign n3935 = n3933 & n3934 ;
  assign n3936 = n3935 ^ x84 ;
  assign n3806 = n3726 & n3771 ;
  assign n3807 = n3806 ^ n3601 ;
  assign n3937 = n3936 ^ n3807 ;
  assign n3938 = n3936 ^ x85 ;
  assign n3939 = n3937 & n3938 ;
  assign n3940 = n3939 ^ x85 ;
  assign n3803 = n3728 ^ x85 ;
  assign n3804 = n3771 & n3803 ;
  assign n3805 = n3804 ^ n3595 ;
  assign n3941 = n3940 ^ n3805 ;
  assign n3942 = n3940 ^ x86 ;
  assign n3943 = n3941 & n3942 ;
  assign n3944 = n3943 ^ x86 ;
  assign n3792 = n3595 ^ x86 ;
  assign n3793 = n3792 ^ n3728 ;
  assign n3794 = n3793 ^ x85 ;
  assign n3795 = n3794 ^ n3792 ;
  assign n3797 = n3728 ^ x86 ;
  assign n3798 = n3797 ^ n3792 ;
  assign n3799 = ~n3795 & ~n3798 ;
  assign n3800 = n3799 ^ n3792 ;
  assign n3801 = n3771 & ~n3800 ;
  assign n3802 = n3801 ^ n3583 ;
  assign n3945 = n3944 ^ n3802 ;
  assign n3946 = n3944 ^ x87 ;
  assign n3947 = n3945 & n3946 ;
  assign n3948 = n3947 ^ x87 ;
  assign n3789 = n3734 ^ x87 ;
  assign n3790 = n3771 & n3789 ;
  assign n3791 = n3790 ^ n3736 ;
  assign n3949 = n3948 ^ n3791 ;
  assign n3950 = n3948 ^ x88 ;
  assign n3951 = n3949 & n3950 ;
  assign n3952 = n3951 ^ x88 ;
  assign n3787 = n3742 & n3771 ;
  assign n3788 = n3787 ^ n3580 ;
  assign n3953 = n3952 ^ n3788 ;
  assign n3954 = n3952 ^ x89 ;
  assign n3955 = n3953 & n3954 ;
  assign n3956 = n3955 ^ x89 ;
  assign n3785 = n3746 & n3771 ;
  assign n3786 = n3785 ^ n3578 ;
  assign n3957 = n3956 ^ n3786 ;
  assign n3958 = n3956 ^ x90 ;
  assign n3959 = n3957 & n3958 ;
  assign n3960 = n3959 ^ x90 ;
  assign n3783 = n3750 & n3771 ;
  assign n3784 = n3783 ^ n3576 ;
  assign n3961 = n3960 ^ n3784 ;
  assign n3962 = n3960 ^ x91 ;
  assign n3963 = n3961 & n3962 ;
  assign n3964 = n3963 ^ x91 ;
  assign n3781 = n3754 & n3771 ;
  assign n3782 = n3781 ^ n3574 ;
  assign n3965 = n3964 ^ n3782 ;
  assign n3966 = n3964 ^ x92 ;
  assign n3967 = n3965 & n3966 ;
  assign n3968 = n3967 ^ x92 ;
  assign n3779 = n3758 & n3771 ;
  assign n3780 = n3779 ^ n3572 ;
  assign n3969 = n3968 ^ n3780 ;
  assign n3970 = n3968 ^ x93 ;
  assign n3971 = n3969 & n3970 ;
  assign n3972 = n3971 ^ x93 ;
  assign n3777 = n3762 & n3771 ;
  assign n3778 = n3777 ^ n3570 ;
  assign n3973 = n3972 ^ n3778 ;
  assign n3974 = n3972 ^ x94 ;
  assign n3975 = n3973 & n3974 ;
  assign n3976 = n3975 ^ x94 ;
  assign n3977 = n3976 ^ x95 ;
  assign n3978 = n3764 ^ x94 ;
  assign n3979 = n3771 & n3978 ;
  assign n3980 = n3979 ^ n3564 ;
  assign n3981 = n3980 ^ x95 ;
  assign n3982 = n3977 & ~n3981 ;
  assign n3983 = n3982 ^ x95 ;
  assign n3984 = n3776 & n3983 ;
  assign n3985 = n3984 ^ n160 ;
  assign n3986 = n3773 & ~n3985 ;
  assign n3987 = n3986 ^ n270 ;
  assign n3774 = x97 & ~n3773 ;
  assign n3775 = n3774 ^ x97 ;
  assign n3988 = n3987 ^ n3775 ;
  assign n3989 = n3773 ^ x96 ;
  assign n3991 = n3773 ^ x95 ;
  assign n3990 = n3976 ^ n3773 ;
  assign n3992 = n3991 ^ n3990 ;
  assign n3993 = n3980 ^ n3773 ;
  assign n3994 = n3993 ^ n3991 ;
  assign n3995 = n3992 & ~n3994 ;
  assign n3996 = n3995 ^ n3991 ;
  assign n3997 = ~n3989 & n3996 ;
  assign n3998 = n3997 ^ x96 ;
  assign n3999 = n160 & ~n3998 ;
  assign n4000 = n3977 & n3999 ;
  assign n4001 = n4000 ^ n3980 ;
  assign n4002 = n4001 ^ x96 ;
  assign n4081 = x65 & n3999 ;
  assign n4075 = n3771 ^ x31 ;
  assign n4076 = n4075 ^ n3771 ;
  assign n4077 = n3999 & ~n4076 ;
  assign n4078 = n4077 ^ n3771 ;
  assign n4079 = x64 & n4078 ;
  assign n4080 = n4079 ^ x32 ;
  assign n4082 = n4081 ^ n4080 ;
  assign n4083 = n4082 ^ x66 ;
  assign n4091 = x31 & x65 ;
  assign n4088 = x65 ^ x30 ;
  assign n4084 = x64 ^ x31 ;
  assign n4085 = n4084 ^ x65 ;
  assign n4089 = n4085 ^ n3999 ;
  assign n4090 = ~n4088 & n4089 ;
  assign n4092 = n4091 ^ n4090 ;
  assign n4093 = x64 & n4092 ;
  assign n4094 = n4093 ^ n4091 ;
  assign n4095 = n4094 ^ x65 ;
  assign n4096 = n4095 ^ n4082 ;
  assign n4097 = ~n4083 & n4096 ;
  assign n4098 = n4097 ^ x66 ;
  assign n4099 = n4098 ^ x67 ;
  assign n4100 = n3851 ^ x66 ;
  assign n4101 = n3999 & n4100 ;
  assign n4102 = n4101 ^ n3854 ;
  assign n4103 = n4102 ^ n4098 ;
  assign n4104 = n4099 & n4103 ;
  assign n4105 = n4104 ^ x67 ;
  assign n4070 = n3858 ^ x67 ;
  assign n4071 = n3999 & n4070 ;
  assign n4072 = n4071 ^ n3860 ;
  assign n4106 = n4105 ^ n4072 ;
  assign n4107 = n4105 ^ x68 ;
  assign n4108 = n4106 & n4107 ;
  assign n4109 = n4108 ^ x68 ;
  assign n4067 = n3864 ^ x68 ;
  assign n4068 = n3999 & n4067 ;
  assign n4069 = n4068 ^ n3866 ;
  assign n4110 = n4109 ^ n4069 ;
  assign n4111 = n4109 ^ x69 ;
  assign n4112 = n4110 & n4111 ;
  assign n4113 = n4112 ^ x69 ;
  assign n4064 = n3870 ^ x69 ;
  assign n4065 = n3999 & n4064 ;
  assign n4066 = n4065 ^ n3872 ;
  assign n4114 = n4113 ^ n4066 ;
  assign n4115 = n4113 ^ x70 ;
  assign n4116 = n4114 & n4115 ;
  assign n4117 = n4116 ^ x70 ;
  assign n4062 = n3878 & n3999 ;
  assign n4063 = n4062 ^ n3839 ;
  assign n4118 = n4117 ^ n4063 ;
  assign n4119 = n4117 ^ x71 ;
  assign n4120 = n4118 & n4119 ;
  assign n4121 = n4120 ^ x71 ;
  assign n4060 = n3882 & n3999 ;
  assign n4061 = n4060 ^ n3837 ;
  assign n4122 = n4121 ^ n4061 ;
  assign n4123 = n4121 ^ x72 ;
  assign n4124 = n4122 & n4123 ;
  assign n4125 = n4124 ^ x72 ;
  assign n4058 = n3886 & n3999 ;
  assign n4059 = n4058 ^ n3835 ;
  assign n4126 = n4125 ^ n4059 ;
  assign n4127 = n4125 ^ x73 ;
  assign n4128 = n4126 & n4127 ;
  assign n4129 = n4128 ^ x73 ;
  assign n4056 = n3890 & n3999 ;
  assign n4057 = n4056 ^ n3833 ;
  assign n4130 = n4129 ^ n4057 ;
  assign n4131 = n4129 ^ x74 ;
  assign n4132 = n4130 & n4131 ;
  assign n4133 = n4132 ^ x74 ;
  assign n4054 = n3894 & n3999 ;
  assign n4055 = n4054 ^ n3831 ;
  assign n4134 = n4133 ^ n4055 ;
  assign n4135 = n4133 ^ x75 ;
  assign n4136 = n4134 & n4135 ;
  assign n4137 = n4136 ^ x75 ;
  assign n4052 = n3898 & n3999 ;
  assign n4053 = n4052 ^ n3829 ;
  assign n4138 = n4137 ^ n4053 ;
  assign n4139 = n4137 ^ x76 ;
  assign n4140 = n4138 & n4139 ;
  assign n4141 = n4140 ^ x76 ;
  assign n4050 = n3902 & n3999 ;
  assign n4051 = n4050 ^ n3827 ;
  assign n4142 = n4141 ^ n4051 ;
  assign n4143 = n4141 ^ x77 ;
  assign n4144 = n4142 & n4143 ;
  assign n4145 = n4144 ^ x77 ;
  assign n4048 = n3906 & n3999 ;
  assign n4049 = n4048 ^ n3825 ;
  assign n4146 = n4145 ^ n4049 ;
  assign n4147 = n4145 ^ x78 ;
  assign n4148 = n4146 & n4147 ;
  assign n4149 = n4148 ^ x78 ;
  assign n4046 = n3910 & n3999 ;
  assign n4047 = n4046 ^ n3823 ;
  assign n4150 = n4149 ^ n4047 ;
  assign n4151 = n4149 ^ x79 ;
  assign n4152 = n4150 & n4151 ;
  assign n4153 = n4152 ^ x79 ;
  assign n4043 = n3912 ^ x79 ;
  assign n4044 = n3999 & n4043 ;
  assign n4045 = n4044 ^ n3818 ;
  assign n4154 = n4153 ^ n4045 ;
  assign n4155 = n4153 ^ x80 ;
  assign n4156 = n4154 & n4155 ;
  assign n4157 = n4156 ^ x80 ;
  assign n4032 = n3818 ^ x80 ;
  assign n4033 = n4032 ^ n3912 ;
  assign n4034 = n4033 ^ x79 ;
  assign n4035 = n4034 ^ n4032 ;
  assign n4037 = n3912 ^ x80 ;
  assign n4038 = n4037 ^ n4032 ;
  assign n4039 = ~n4035 & ~n4038 ;
  assign n4040 = n4039 ^ n4032 ;
  assign n4041 = n3999 & ~n4040 ;
  assign n4042 = n4041 ^ n3815 ;
  assign n4158 = n4157 ^ n4042 ;
  assign n4159 = n4157 ^ x81 ;
  assign n4160 = n4158 & n4159 ;
  assign n4161 = n4160 ^ x81 ;
  assign n4029 = n3918 ^ x81 ;
  assign n4030 = n3999 & n4029 ;
  assign n4031 = n4030 ^ n3920 ;
  assign n4162 = n4161 ^ n4031 ;
  assign n4163 = n4161 ^ x82 ;
  assign n4164 = n4162 & n4163 ;
  assign n4165 = n4164 ^ x82 ;
  assign n4027 = n3926 & n3999 ;
  assign n4028 = n4027 ^ n3813 ;
  assign n4166 = n4165 ^ n4028 ;
  assign n4167 = n4165 ^ x83 ;
  assign n4168 = n4166 & n4167 ;
  assign n4169 = n4168 ^ x83 ;
  assign n4025 = n3930 & n3999 ;
  assign n4026 = n4025 ^ n3811 ;
  assign n4170 = n4169 ^ n4026 ;
  assign n4171 = n4169 ^ x84 ;
  assign n4172 = n4170 & n4171 ;
  assign n4173 = n4172 ^ x84 ;
  assign n4023 = n3934 & n3999 ;
  assign n4024 = n4023 ^ n3809 ;
  assign n4174 = n4173 ^ n4024 ;
  assign n4175 = n4173 ^ x85 ;
  assign n4176 = n4174 & n4175 ;
  assign n4177 = n4176 ^ x85 ;
  assign n4021 = n3938 & n3999 ;
  assign n4022 = n4021 ^ n3807 ;
  assign n4178 = n4177 ^ n4022 ;
  assign n4179 = n4177 ^ x86 ;
  assign n4180 = n4178 & n4179 ;
  assign n4181 = n4180 ^ x86 ;
  assign n4019 = n3942 & n3999 ;
  assign n4020 = n4019 ^ n3805 ;
  assign n4182 = n4181 ^ n4020 ;
  assign n4183 = n4181 ^ x87 ;
  assign n4184 = n4182 & n4183 ;
  assign n4185 = n4184 ^ x87 ;
  assign n4017 = n3946 & n3999 ;
  assign n4018 = n4017 ^ n3802 ;
  assign n4186 = n4185 ^ n4018 ;
  assign n4187 = n4185 ^ x88 ;
  assign n4188 = n4186 & n4187 ;
  assign n4189 = n4188 ^ x88 ;
  assign n4015 = n3950 & n3999 ;
  assign n4016 = n4015 ^ n3791 ;
  assign n4190 = n4189 ^ n4016 ;
  assign n4191 = n4189 ^ x89 ;
  assign n4192 = n4190 & n4191 ;
  assign n4193 = n4192 ^ x89 ;
  assign n4013 = n3954 & n3999 ;
  assign n4014 = n4013 ^ n3788 ;
  assign n4194 = n4193 ^ n4014 ;
  assign n4195 = n4193 ^ x90 ;
  assign n4196 = n4194 & n4195 ;
  assign n4197 = n4196 ^ x90 ;
  assign n4011 = n3958 & n3999 ;
  assign n4012 = n4011 ^ n3786 ;
  assign n4198 = n4197 ^ n4012 ;
  assign n4199 = n4197 ^ x91 ;
  assign n4200 = n4198 & n4199 ;
  assign n4201 = n4200 ^ x91 ;
  assign n4009 = n3962 & n3999 ;
  assign n4010 = n4009 ^ n3784 ;
  assign n4202 = n4201 ^ n4010 ;
  assign n4203 = n4201 ^ x92 ;
  assign n4204 = n4202 & n4203 ;
  assign n4205 = n4204 ^ x92 ;
  assign n4007 = n3966 & n3999 ;
  assign n4008 = n4007 ^ n3782 ;
  assign n4206 = n4205 ^ n4008 ;
  assign n4207 = n4205 ^ x93 ;
  assign n4208 = n4206 & n4207 ;
  assign n4209 = n4208 ^ x93 ;
  assign n4005 = n3970 & n3999 ;
  assign n4006 = n4005 ^ n3780 ;
  assign n4210 = n4209 ^ n4006 ;
  assign n4211 = n4209 ^ x94 ;
  assign n4212 = n4210 & n4211 ;
  assign n4213 = n4212 ^ x94 ;
  assign n4003 = n3974 & n3999 ;
  assign n4004 = n4003 ^ n3778 ;
  assign n4214 = n4213 ^ n4004 ;
  assign n4217 = n4004 ^ x95 ;
  assign n4218 = n4214 & ~n4217 ;
  assign n4215 = x96 ^ x95 ;
  assign n4219 = n4218 ^ n4215 ;
  assign n4222 = ~n4002 & n4219 ;
  assign n4223 = n4222 ^ x96 ;
  assign n4224 = ~n3988 & n4223 ;
  assign n4225 = n4224 ^ n270 ;
  assign n4226 = n159 & ~n3774 ;
  assign n4227 = ~n4224 & n4226 ;
  assign n4228 = n4219 & n4227 ;
  assign n4229 = n4228 ^ n4001 ;
  assign n4230 = n4229 ^ x97 ;
  assign n4286 = n4099 & n4227 ;
  assign n4287 = n4286 ^ n4102 ;
  assign n4288 = n4287 ^ x68 ;
  assign n4306 = x30 & x65 ;
  assign n4303 = x65 ^ x29 ;
  assign n4299 = x64 ^ x30 ;
  assign n4300 = n4299 ^ x65 ;
  assign n4304 = n4300 ^ n4227 ;
  assign n4305 = ~n4303 & n4304 ;
  assign n4307 = n4306 ^ n4305 ;
  assign n4308 = x64 & n4307 ;
  assign n4309 = n4308 ^ n4306 ;
  assign n4310 = n4309 ^ x65 ;
  assign n4297 = x64 & n3999 ;
  assign n4293 = ~x30 & x64 ;
  assign n4294 = n4293 ^ x65 ;
  assign n4295 = n4227 & n4294 ;
  assign n4296 = n4295 ^ x31 ;
  assign n4298 = n4297 ^ n4296 ;
  assign n4311 = n4310 ^ n4298 ;
  assign n4312 = n4310 ^ x66 ;
  assign n4313 = n4311 & n4312 ;
  assign n4314 = n4313 ^ x66 ;
  assign n4289 = n4095 ^ x66 ;
  assign n4290 = n4227 & n4289 ;
  assign n4291 = n4290 ^ n4082 ;
  assign n4315 = n4314 ^ n4291 ;
  assign n4316 = n4314 ^ x67 ;
  assign n4317 = n4315 & n4316 ;
  assign n4318 = n4317 ^ x67 ;
  assign n4319 = n4318 ^ n4287 ;
  assign n4320 = ~n4288 & n4319 ;
  assign n4321 = n4320 ^ x68 ;
  assign n4322 = n4321 ^ x69 ;
  assign n4323 = n4107 & n4227 ;
  assign n4324 = n4323 ^ n4072 ;
  assign n4325 = n4324 ^ n4321 ;
  assign n4326 = n4322 & n4325 ;
  assign n4327 = n4326 ^ x69 ;
  assign n4284 = n4111 & n4227 ;
  assign n4285 = n4284 ^ n4069 ;
  assign n4328 = n4327 ^ n4285 ;
  assign n4329 = n4327 ^ x70 ;
  assign n4330 = n4328 & n4329 ;
  assign n4331 = n4330 ^ x70 ;
  assign n4282 = n4115 & n4227 ;
  assign n4283 = n4282 ^ n4066 ;
  assign n4332 = n4331 ^ n4283 ;
  assign n4333 = n4331 ^ x71 ;
  assign n4334 = n4332 & n4333 ;
  assign n4335 = n4334 ^ x71 ;
  assign n4280 = n4119 & n4227 ;
  assign n4281 = n4280 ^ n4063 ;
  assign n4336 = n4335 ^ n4281 ;
  assign n4337 = n4335 ^ x72 ;
  assign n4338 = n4336 & n4337 ;
  assign n4339 = n4338 ^ x72 ;
  assign n4278 = n4123 & n4227 ;
  assign n4279 = n4278 ^ n4061 ;
  assign n4340 = n4339 ^ n4279 ;
  assign n4341 = n4339 ^ x73 ;
  assign n4342 = n4340 & n4341 ;
  assign n4343 = n4342 ^ x73 ;
  assign n4276 = n4127 & n4227 ;
  assign n4277 = n4276 ^ n4059 ;
  assign n4344 = n4343 ^ n4277 ;
  assign n4345 = n4343 ^ x74 ;
  assign n4346 = n4344 & n4345 ;
  assign n4347 = n4346 ^ x74 ;
  assign n4274 = n4131 & n4227 ;
  assign n4275 = n4274 ^ n4057 ;
  assign n4348 = n4347 ^ n4275 ;
  assign n4349 = n4347 ^ x75 ;
  assign n4350 = n4348 & n4349 ;
  assign n4351 = n4350 ^ x75 ;
  assign n4272 = n4135 & n4227 ;
  assign n4273 = n4272 ^ n4055 ;
  assign n4352 = n4351 ^ n4273 ;
  assign n4353 = n4351 ^ x76 ;
  assign n4354 = n4352 & n4353 ;
  assign n4355 = n4354 ^ x76 ;
  assign n4270 = n4139 & n4227 ;
  assign n4271 = n4270 ^ n4053 ;
  assign n4356 = n4355 ^ n4271 ;
  assign n4357 = n4355 ^ x77 ;
  assign n4358 = n4356 & n4357 ;
  assign n4359 = n4358 ^ x77 ;
  assign n4268 = n4143 & n4227 ;
  assign n4269 = n4268 ^ n4051 ;
  assign n4360 = n4359 ^ n4269 ;
  assign n4361 = n4359 ^ x78 ;
  assign n4362 = n4360 & n4361 ;
  assign n4363 = n4362 ^ x78 ;
  assign n4266 = n4147 & n4227 ;
  assign n4267 = n4266 ^ n4049 ;
  assign n4364 = n4363 ^ n4267 ;
  assign n4365 = n4363 ^ x79 ;
  assign n4366 = n4364 & n4365 ;
  assign n4367 = n4366 ^ x79 ;
  assign n4264 = n4151 & n4227 ;
  assign n4265 = n4264 ^ n4047 ;
  assign n4368 = n4367 ^ n4265 ;
  assign n4369 = n4367 ^ x80 ;
  assign n4370 = n4368 & n4369 ;
  assign n4371 = n4370 ^ x80 ;
  assign n4262 = n4155 & n4227 ;
  assign n4263 = n4262 ^ n4045 ;
  assign n4372 = n4371 ^ n4263 ;
  assign n4373 = n4371 ^ x81 ;
  assign n4374 = n4372 & n4373 ;
  assign n4375 = n4374 ^ x81 ;
  assign n4260 = n4159 & n4227 ;
  assign n4261 = n4260 ^ n4042 ;
  assign n4376 = n4375 ^ n4261 ;
  assign n4377 = n4375 ^ x82 ;
  assign n4378 = n4376 & n4377 ;
  assign n4379 = n4378 ^ x82 ;
  assign n4258 = n4163 & n4227 ;
  assign n4259 = n4258 ^ n4031 ;
  assign n4380 = n4379 ^ n4259 ;
  assign n4381 = n4379 ^ x83 ;
  assign n4382 = n4380 & n4381 ;
  assign n4383 = n4382 ^ x83 ;
  assign n4256 = n4167 & n4227 ;
  assign n4257 = n4256 ^ n4028 ;
  assign n4384 = n4383 ^ n4257 ;
  assign n4385 = n4383 ^ x84 ;
  assign n4386 = n4384 & n4385 ;
  assign n4387 = n4386 ^ x84 ;
  assign n4254 = n4171 & n4227 ;
  assign n4255 = n4254 ^ n4026 ;
  assign n4388 = n4387 ^ n4255 ;
  assign n4389 = n4387 ^ x85 ;
  assign n4390 = n4388 & n4389 ;
  assign n4391 = n4390 ^ x85 ;
  assign n4252 = n4175 & n4227 ;
  assign n4253 = n4252 ^ n4024 ;
  assign n4392 = n4391 ^ n4253 ;
  assign n4393 = n4391 ^ x86 ;
  assign n4394 = n4392 & n4393 ;
  assign n4395 = n4394 ^ x86 ;
  assign n4250 = n4179 & n4227 ;
  assign n4251 = n4250 ^ n4022 ;
  assign n4396 = n4395 ^ n4251 ;
  assign n4397 = n4395 ^ x87 ;
  assign n4398 = n4396 & n4397 ;
  assign n4399 = n4398 ^ x87 ;
  assign n4248 = n4183 & n4227 ;
  assign n4249 = n4248 ^ n4020 ;
  assign n4400 = n4399 ^ n4249 ;
  assign n4401 = n4399 ^ x88 ;
  assign n4402 = n4400 & n4401 ;
  assign n4403 = n4402 ^ x88 ;
  assign n4246 = n4187 & n4227 ;
  assign n4247 = n4246 ^ n4018 ;
  assign n4404 = n4403 ^ n4247 ;
  assign n4405 = n4403 ^ x89 ;
  assign n4406 = n4404 & n4405 ;
  assign n4407 = n4406 ^ x89 ;
  assign n4244 = n4191 & n4227 ;
  assign n4245 = n4244 ^ n4016 ;
  assign n4408 = n4407 ^ n4245 ;
  assign n4409 = n4407 ^ x90 ;
  assign n4410 = n4408 & n4409 ;
  assign n4411 = n4410 ^ x90 ;
  assign n4242 = n4195 & n4227 ;
  assign n4243 = n4242 ^ n4014 ;
  assign n4412 = n4411 ^ n4243 ;
  assign n4413 = n4411 ^ x91 ;
  assign n4414 = n4412 & n4413 ;
  assign n4415 = n4414 ^ x91 ;
  assign n4240 = n4199 & n4227 ;
  assign n4241 = n4240 ^ n4012 ;
  assign n4416 = n4415 ^ n4241 ;
  assign n4417 = n4415 ^ x92 ;
  assign n4418 = n4416 & n4417 ;
  assign n4419 = n4418 ^ x92 ;
  assign n4238 = n4203 & n4227 ;
  assign n4239 = n4238 ^ n4010 ;
  assign n4420 = n4419 ^ n4239 ;
  assign n4421 = n4419 ^ x93 ;
  assign n4422 = n4420 & n4421 ;
  assign n4423 = n4422 ^ x93 ;
  assign n4236 = n4207 & n4227 ;
  assign n4237 = n4236 ^ n4008 ;
  assign n4424 = n4423 ^ n4237 ;
  assign n4425 = n4423 ^ x94 ;
  assign n4426 = n4424 & n4425 ;
  assign n4427 = n4426 ^ x94 ;
  assign n4234 = n4211 & n4227 ;
  assign n4235 = n4234 ^ n4006 ;
  assign n4428 = n4427 ^ n4235 ;
  assign n4429 = n4427 ^ x95 ;
  assign n4430 = n4428 & n4429 ;
  assign n4431 = n4430 ^ x95 ;
  assign n4231 = n4213 ^ x95 ;
  assign n4232 = n4227 & n4231 ;
  assign n4233 = n4232 ^ n4004 ;
  assign n4432 = n4431 ^ n4233 ;
  assign n4435 = n4233 ^ x96 ;
  assign n4436 = n4432 & ~n4435 ;
  assign n4433 = x97 ^ x96 ;
  assign n4437 = n4436 ^ n4433 ;
  assign n4438 = ~n4230 & n4437 ;
  assign n4439 = n4438 ^ x97 ;
  assign n4440 = n4439 ^ n3987 ;
  assign n4441 = n3987 ^ x98 ;
  assign n4442 = ~n4440 & n4441 ;
  assign n4443 = n4442 ^ n4439 ;
  assign n4444 = n158 & ~n4443 ;
  assign n4445 = n4442 & n4444 ;
  assign n4446 = ~n4225 & n4445 ;
  assign n4447 = n4446 ^ n4444 ;
  assign n4448 = n3986 & ~n4227 ;
  assign n4449 = ~n4447 & n4448 ;
  assign n4450 = n4449 ^ n270 ;
  assign n4451 = n4450 ^ x99 ;
  assign n4455 = n4437 & n4447 ;
  assign n4456 = n4455 ^ n4229 ;
  assign n4458 = n4456 ^ x97 ;
  assign n4452 = n4431 ^ x96 ;
  assign n4453 = n4447 & n4452 ;
  assign n4454 = n4453 ^ n4233 ;
  assign n4457 = n4456 ^ n4454 ;
  assign n4459 = n4458 ^ n4457 ;
  assign n4658 = n4425 & n4447 ;
  assign n4659 = n4658 ^ n4237 ;
  assign n4462 = n4421 & n4447 ;
  assign n4463 = n4462 ^ n4239 ;
  assign n4464 = n4463 ^ x94 ;
  assign n4468 = n4463 ^ x93 ;
  assign n4465 = n4417 & n4447 ;
  assign n4466 = n4465 ^ n4241 ;
  assign n4467 = n4466 ^ n4463 ;
  assign n4469 = n4468 ^ n4467 ;
  assign n4562 = n4329 & n4447 ;
  assign n4563 = n4562 ^ n4285 ;
  assign n4512 = n4322 & n4447 ;
  assign n4513 = n4512 ^ n4324 ;
  assign n4514 = n4513 ^ x70 ;
  assign n4519 = n4513 ^ x69 ;
  assign n4515 = n4318 ^ x68 ;
  assign n4516 = n4447 & n4515 ;
  assign n4517 = n4516 ^ n4287 ;
  assign n4518 = n4517 ^ n4513 ;
  assign n4520 = n4519 ^ n4518 ;
  assign n4539 = x29 & x65 ;
  assign n4536 = x65 ^ x28 ;
  assign n4532 = x64 ^ x29 ;
  assign n4533 = n4532 ^ x65 ;
  assign n4537 = n4533 ^ n4447 ;
  assign n4538 = ~n4536 & n4537 ;
  assign n4540 = n4539 ^ n4538 ;
  assign n4541 = x64 & n4540 ;
  assign n4542 = n4541 ^ n4539 ;
  assign n4543 = n4542 ^ x65 ;
  assign n4530 = x64 & n4227 ;
  assign n4525 = n4303 ^ x65 ;
  assign n4526 = x64 & ~n4525 ;
  assign n4527 = n4526 ^ x65 ;
  assign n4528 = n4447 & n4527 ;
  assign n4529 = n4528 ^ x30 ;
  assign n4531 = n4530 ^ n4529 ;
  assign n4544 = n4543 ^ n4531 ;
  assign n4545 = n4543 ^ x66 ;
  assign n4546 = n4544 & n4545 ;
  assign n4547 = n4546 ^ x66 ;
  assign n4523 = n4312 & n4447 ;
  assign n4524 = n4523 ^ n4298 ;
  assign n4548 = n4547 ^ n4524 ;
  assign n4549 = n4547 ^ x67 ;
  assign n4550 = n4548 & n4549 ;
  assign n4551 = n4550 ^ x67 ;
  assign n4521 = n4316 & n4447 ;
  assign n4522 = n4521 ^ n4291 ;
  assign n4552 = n4551 ^ n4522 ;
  assign n4553 = n4551 ^ x68 ;
  assign n4554 = n4552 & n4553 ;
  assign n4555 = n4554 ^ x68 ;
  assign n4556 = n4555 ^ n4513 ;
  assign n4557 = n4556 ^ n4519 ;
  assign n4558 = ~n4520 & n4557 ;
  assign n4559 = n4558 ^ n4519 ;
  assign n4560 = ~n4514 & n4559 ;
  assign n4561 = n4560 ^ x70 ;
  assign n4564 = n4563 ^ n4561 ;
  assign n4565 = n4563 ^ x71 ;
  assign n4566 = n4564 & ~n4565 ;
  assign n4567 = n4566 ^ x71 ;
  assign n4510 = n4333 & n4447 ;
  assign n4511 = n4510 ^ n4283 ;
  assign n4568 = n4567 ^ n4511 ;
  assign n4569 = n4567 ^ x72 ;
  assign n4570 = n4568 & n4569 ;
  assign n4571 = n4570 ^ x72 ;
  assign n4508 = n4337 & n4447 ;
  assign n4509 = n4508 ^ n4281 ;
  assign n4572 = n4571 ^ n4509 ;
  assign n4573 = n4571 ^ x73 ;
  assign n4574 = n4572 & n4573 ;
  assign n4575 = n4574 ^ x73 ;
  assign n4506 = n4341 & n4447 ;
  assign n4507 = n4506 ^ n4279 ;
  assign n4576 = n4575 ^ n4507 ;
  assign n4577 = n4575 ^ x74 ;
  assign n4578 = n4576 & n4577 ;
  assign n4579 = n4578 ^ x74 ;
  assign n4504 = n4345 & n4447 ;
  assign n4505 = n4504 ^ n4277 ;
  assign n4580 = n4579 ^ n4505 ;
  assign n4581 = n4579 ^ x75 ;
  assign n4582 = n4580 & n4581 ;
  assign n4583 = n4582 ^ x75 ;
  assign n4502 = n4349 & n4447 ;
  assign n4503 = n4502 ^ n4275 ;
  assign n4584 = n4583 ^ n4503 ;
  assign n4585 = n4583 ^ x76 ;
  assign n4586 = n4584 & n4585 ;
  assign n4587 = n4586 ^ x76 ;
  assign n4500 = n4353 & n4447 ;
  assign n4501 = n4500 ^ n4273 ;
  assign n4588 = n4587 ^ n4501 ;
  assign n4589 = n4587 ^ x77 ;
  assign n4590 = n4588 & n4589 ;
  assign n4591 = n4590 ^ x77 ;
  assign n4498 = n4357 & n4447 ;
  assign n4499 = n4498 ^ n4271 ;
  assign n4592 = n4591 ^ n4499 ;
  assign n4593 = n4591 ^ x78 ;
  assign n4594 = n4592 & n4593 ;
  assign n4595 = n4594 ^ x78 ;
  assign n4496 = n4361 & n4447 ;
  assign n4497 = n4496 ^ n4269 ;
  assign n4596 = n4595 ^ n4497 ;
  assign n4597 = n4595 ^ x79 ;
  assign n4598 = n4596 & n4597 ;
  assign n4599 = n4598 ^ x79 ;
  assign n4494 = n4365 & n4447 ;
  assign n4495 = n4494 ^ n4267 ;
  assign n4600 = n4599 ^ n4495 ;
  assign n4601 = n4599 ^ x80 ;
  assign n4602 = n4600 & n4601 ;
  assign n4603 = n4602 ^ x80 ;
  assign n4492 = n4369 & n4447 ;
  assign n4493 = n4492 ^ n4265 ;
  assign n4604 = n4603 ^ n4493 ;
  assign n4605 = n4603 ^ x81 ;
  assign n4606 = n4604 & n4605 ;
  assign n4607 = n4606 ^ x81 ;
  assign n4490 = n4373 & n4447 ;
  assign n4491 = n4490 ^ n4263 ;
  assign n4608 = n4607 ^ n4491 ;
  assign n4609 = n4607 ^ x82 ;
  assign n4610 = n4608 & n4609 ;
  assign n4611 = n4610 ^ x82 ;
  assign n4488 = n4377 & n4447 ;
  assign n4489 = n4488 ^ n4261 ;
  assign n4612 = n4611 ^ n4489 ;
  assign n4613 = n4611 ^ x83 ;
  assign n4614 = n4612 & n4613 ;
  assign n4615 = n4614 ^ x83 ;
  assign n4486 = n4381 & n4447 ;
  assign n4487 = n4486 ^ n4259 ;
  assign n4616 = n4615 ^ n4487 ;
  assign n4617 = n4615 ^ x84 ;
  assign n4618 = n4616 & n4617 ;
  assign n4619 = n4618 ^ x84 ;
  assign n4484 = n4385 & n4447 ;
  assign n4485 = n4484 ^ n4257 ;
  assign n4620 = n4619 ^ n4485 ;
  assign n4621 = n4619 ^ x85 ;
  assign n4622 = n4620 & n4621 ;
  assign n4623 = n4622 ^ x85 ;
  assign n4482 = n4389 & n4447 ;
  assign n4483 = n4482 ^ n4255 ;
  assign n4624 = n4623 ^ n4483 ;
  assign n4625 = n4623 ^ x86 ;
  assign n4626 = n4624 & n4625 ;
  assign n4627 = n4626 ^ x86 ;
  assign n4480 = n4393 & n4447 ;
  assign n4481 = n4480 ^ n4253 ;
  assign n4628 = n4627 ^ n4481 ;
  assign n4629 = n4627 ^ x87 ;
  assign n4630 = n4628 & n4629 ;
  assign n4631 = n4630 ^ x87 ;
  assign n4478 = n4397 & n4447 ;
  assign n4479 = n4478 ^ n4251 ;
  assign n4632 = n4631 ^ n4479 ;
  assign n4633 = n4631 ^ x88 ;
  assign n4634 = n4632 & n4633 ;
  assign n4635 = n4634 ^ x88 ;
  assign n4476 = n4401 & n4447 ;
  assign n4477 = n4476 ^ n4249 ;
  assign n4636 = n4635 ^ n4477 ;
  assign n4637 = n4635 ^ x89 ;
  assign n4638 = n4636 & n4637 ;
  assign n4639 = n4638 ^ x89 ;
  assign n4474 = n4405 & n4447 ;
  assign n4475 = n4474 ^ n4247 ;
  assign n4640 = n4639 ^ n4475 ;
  assign n4641 = n4639 ^ x90 ;
  assign n4642 = n4640 & n4641 ;
  assign n4643 = n4642 ^ x90 ;
  assign n4472 = n4409 & n4447 ;
  assign n4473 = n4472 ^ n4245 ;
  assign n4644 = n4643 ^ n4473 ;
  assign n4645 = n4643 ^ x91 ;
  assign n4646 = n4644 & n4645 ;
  assign n4647 = n4646 ^ x91 ;
  assign n4470 = n4413 & n4447 ;
  assign n4471 = n4470 ^ n4243 ;
  assign n4648 = n4647 ^ n4471 ;
  assign n4649 = n4647 ^ x92 ;
  assign n4650 = n4648 & n4649 ;
  assign n4651 = n4650 ^ x92 ;
  assign n4652 = n4651 ^ n4463 ;
  assign n4653 = n4652 ^ n4468 ;
  assign n4654 = ~n4469 & n4653 ;
  assign n4655 = n4654 ^ n4468 ;
  assign n4656 = ~n4464 & n4655 ;
  assign n4657 = n4656 ^ x94 ;
  assign n4660 = n4659 ^ n4657 ;
  assign n4661 = n4659 ^ x95 ;
  assign n4662 = n4660 & ~n4661 ;
  assign n4663 = n4662 ^ x95 ;
  assign n4460 = n4429 & n4447 ;
  assign n4461 = n4460 ^ n4235 ;
  assign n4664 = n4663 ^ n4461 ;
  assign n4665 = n4663 ^ x96 ;
  assign n4666 = n4664 & n4665 ;
  assign n4667 = n4666 ^ x96 ;
  assign n4668 = n4667 ^ n4456 ;
  assign n4669 = n4668 ^ n4458 ;
  assign n4670 = ~n4459 & n4669 ;
  assign n4671 = n4670 ^ n4458 ;
  assign n4673 = n4450 ^ x98 ;
  assign n4672 = n4456 ^ n4450 ;
  assign n4674 = n4673 ^ n4672 ;
  assign n4675 = n4671 & ~n4674 ;
  assign n4676 = n4675 ^ n4673 ;
  assign n4677 = ~n4451 & n4676 ;
  assign n4678 = n4677 ^ x99 ;
  assign n4679 = n157 & ~n4678 ;
  assign n4913 = n4651 ^ x93 ;
  assign n4914 = n4679 & n4913 ;
  assign n4915 = n4914 ^ n4466 ;
  assign n4713 = n4649 & n4679 ;
  assign n4714 = n4713 ^ n4471 ;
  assign n4715 = n4714 ^ x93 ;
  assign n4719 = n4714 ^ x92 ;
  assign n4716 = n4645 & n4679 ;
  assign n4717 = n4716 ^ n4473 ;
  assign n4718 = n4717 ^ n4714 ;
  assign n4720 = n4719 ^ n4718 ;
  assign n4893 = n4633 & n4679 ;
  assign n4894 = n4893 ^ n4479 ;
  assign n4725 = n4629 & n4679 ;
  assign n4726 = n4725 ^ n4481 ;
  assign n4727 = n4726 ^ x88 ;
  assign n4731 = n4726 ^ x87 ;
  assign n4728 = n4625 & n4679 ;
  assign n4729 = n4728 ^ n4483 ;
  assign n4730 = n4729 ^ n4726 ;
  assign n4732 = n4731 ^ n4730 ;
  assign n4877 = n4617 & n4679 ;
  assign n4878 = n4877 ^ n4487 ;
  assign n4735 = n4613 & n4679 ;
  assign n4736 = n4735 ^ n4489 ;
  assign n4737 = n4736 ^ x84 ;
  assign n4741 = n4736 ^ x83 ;
  assign n4738 = n4609 & n4679 ;
  assign n4739 = n4738 ^ n4491 ;
  assign n4740 = n4739 ^ n4736 ;
  assign n4742 = n4741 ^ n4740 ;
  assign n4743 = n4605 & n4679 ;
  assign n4744 = n4743 ^ n4493 ;
  assign n4745 = n4744 ^ x82 ;
  assign n4749 = n4744 ^ x81 ;
  assign n4746 = n4601 & n4679 ;
  assign n4747 = n4746 ^ n4495 ;
  assign n4748 = n4747 ^ n4744 ;
  assign n4750 = n4749 ^ n4748 ;
  assign n4755 = n4589 & n4679 ;
  assign n4756 = n4755 ^ n4501 ;
  assign n4757 = n4756 ^ x78 ;
  assign n4758 = n4585 & n4679 ;
  assign n4759 = n4758 ^ n4503 ;
  assign n4760 = n4759 ^ x77 ;
  assign n4799 = ~x27 & x64 ;
  assign n4804 = n4679 ^ x28 ;
  assign n4805 = n4799 & ~n4804 ;
  assign n4801 = x64 & n4679 ;
  assign n4800 = n4799 ^ x28 ;
  assign n4802 = n4801 ^ n4800 ;
  assign n4803 = x65 & ~n4802 ;
  assign n4806 = n4805 ^ n4803 ;
  assign n4797 = x64 & n4447 ;
  assign n4793 = ~x28 & x64 ;
  assign n4794 = n4793 ^ x65 ;
  assign n4795 = n4679 & n4794 ;
  assign n4796 = n4795 ^ x29 ;
  assign n4798 = n4797 ^ n4796 ;
  assign n4807 = n4806 ^ n4798 ;
  assign n4808 = n4806 ^ x66 ;
  assign n4809 = n4807 & n4808 ;
  assign n4810 = n4809 ^ x66 ;
  assign n4790 = n4545 & n4679 ;
  assign n4791 = n4790 ^ n4531 ;
  assign n4811 = n4810 ^ n4791 ;
  assign n4812 = n4810 ^ x67 ;
  assign n4813 = n4811 & n4812 ;
  assign n4814 = n4813 ^ x67 ;
  assign n4788 = n4549 & n4679 ;
  assign n4789 = n4788 ^ n4524 ;
  assign n4815 = n4814 ^ n4789 ;
  assign n4816 = n4814 ^ x68 ;
  assign n4817 = n4815 & n4816 ;
  assign n4818 = n4817 ^ x68 ;
  assign n4786 = n4553 & n4679 ;
  assign n4787 = n4786 ^ n4522 ;
  assign n4819 = n4818 ^ n4787 ;
  assign n4820 = n4818 ^ x69 ;
  assign n4821 = n4819 & n4820 ;
  assign n4822 = n4821 ^ x69 ;
  assign n4783 = n4555 ^ x69 ;
  assign n4784 = n4679 & n4783 ;
  assign n4785 = n4784 ^ n4517 ;
  assign n4823 = n4822 ^ n4785 ;
  assign n4824 = n4822 ^ x70 ;
  assign n4825 = n4823 & n4824 ;
  assign n4826 = n4825 ^ x70 ;
  assign n4772 = n4517 ^ x70 ;
  assign n4773 = n4772 ^ n4555 ;
  assign n4774 = n4773 ^ x69 ;
  assign n4775 = n4774 ^ n4772 ;
  assign n4777 = n4555 ^ x70 ;
  assign n4778 = n4777 ^ n4772 ;
  assign n4779 = ~n4775 & ~n4778 ;
  assign n4780 = n4779 ^ n4772 ;
  assign n4781 = n4679 & ~n4780 ;
  assign n4782 = n4781 ^ n4513 ;
  assign n4827 = n4826 ^ n4782 ;
  assign n4828 = n4826 ^ x71 ;
  assign n4829 = n4827 & n4828 ;
  assign n4830 = n4829 ^ x71 ;
  assign n4769 = n4561 ^ x71 ;
  assign n4770 = n4679 & n4769 ;
  assign n4771 = n4770 ^ n4563 ;
  assign n4831 = n4830 ^ n4771 ;
  assign n4832 = n4830 ^ x72 ;
  assign n4833 = n4831 & n4832 ;
  assign n4834 = n4833 ^ x72 ;
  assign n4767 = n4569 & n4679 ;
  assign n4768 = n4767 ^ n4511 ;
  assign n4835 = n4834 ^ n4768 ;
  assign n4836 = n4834 ^ x73 ;
  assign n4837 = n4835 & n4836 ;
  assign n4838 = n4837 ^ x73 ;
  assign n4765 = n4573 & n4679 ;
  assign n4766 = n4765 ^ n4509 ;
  assign n4839 = n4838 ^ n4766 ;
  assign n4840 = n4838 ^ x74 ;
  assign n4841 = n4839 & n4840 ;
  assign n4842 = n4841 ^ x74 ;
  assign n4763 = n4577 & n4679 ;
  assign n4764 = n4763 ^ n4507 ;
  assign n4843 = n4842 ^ n4764 ;
  assign n4844 = n4842 ^ x75 ;
  assign n4845 = n4843 & n4844 ;
  assign n4846 = n4845 ^ x75 ;
  assign n4761 = n4581 & n4679 ;
  assign n4762 = n4761 ^ n4505 ;
  assign n4847 = n4846 ^ n4762 ;
  assign n4848 = n4846 ^ x76 ;
  assign n4849 = n4847 & n4848 ;
  assign n4850 = n4849 ^ x76 ;
  assign n4851 = n4850 ^ n4759 ;
  assign n4852 = ~n4760 & n4851 ;
  assign n4853 = n4852 ^ x77 ;
  assign n4854 = n4853 ^ n4756 ;
  assign n4855 = ~n4757 & n4854 ;
  assign n4856 = n4855 ^ x78 ;
  assign n4753 = n4593 & n4679 ;
  assign n4754 = n4753 ^ n4499 ;
  assign n4857 = n4856 ^ n4754 ;
  assign n4858 = n4856 ^ x79 ;
  assign n4859 = n4857 & n4858 ;
  assign n4860 = n4859 ^ x79 ;
  assign n4751 = n4597 & n4679 ;
  assign n4752 = n4751 ^ n4497 ;
  assign n4861 = n4860 ^ n4752 ;
  assign n4862 = n4860 ^ x80 ;
  assign n4863 = n4861 & n4862 ;
  assign n4864 = n4863 ^ x80 ;
  assign n4865 = n4864 ^ n4744 ;
  assign n4866 = n4865 ^ n4749 ;
  assign n4867 = ~n4750 & n4866 ;
  assign n4868 = n4867 ^ n4749 ;
  assign n4869 = ~n4745 & n4868 ;
  assign n4870 = n4869 ^ x82 ;
  assign n4871 = n4870 ^ n4736 ;
  assign n4872 = n4871 ^ n4741 ;
  assign n4873 = ~n4742 & n4872 ;
  assign n4874 = n4873 ^ n4741 ;
  assign n4875 = ~n4737 & n4874 ;
  assign n4876 = n4875 ^ x84 ;
  assign n4879 = n4878 ^ n4876 ;
  assign n4880 = n4878 ^ x85 ;
  assign n4881 = n4879 & ~n4880 ;
  assign n4882 = n4881 ^ x85 ;
  assign n4733 = n4621 & n4679 ;
  assign n4734 = n4733 ^ n4485 ;
  assign n4883 = n4882 ^ n4734 ;
  assign n4884 = n4882 ^ x86 ;
  assign n4885 = n4883 & n4884 ;
  assign n4886 = n4885 ^ x86 ;
  assign n4887 = n4886 ^ n4726 ;
  assign n4888 = n4887 ^ n4731 ;
  assign n4889 = ~n4732 & n4888 ;
  assign n4890 = n4889 ^ n4731 ;
  assign n4891 = ~n4727 & n4890 ;
  assign n4892 = n4891 ^ x88 ;
  assign n4895 = n4894 ^ n4892 ;
  assign n4896 = n4894 ^ x89 ;
  assign n4897 = n4895 & ~n4896 ;
  assign n4898 = n4897 ^ x89 ;
  assign n4723 = n4637 & n4679 ;
  assign n4724 = n4723 ^ n4477 ;
  assign n4899 = n4898 ^ n4724 ;
  assign n4900 = n4898 ^ x90 ;
  assign n4901 = n4899 & n4900 ;
  assign n4902 = n4901 ^ x90 ;
  assign n4721 = n4641 & n4679 ;
  assign n4722 = n4721 ^ n4475 ;
  assign n4903 = n4902 ^ n4722 ;
  assign n4904 = n4902 ^ x91 ;
  assign n4905 = n4903 & n4904 ;
  assign n4906 = n4905 ^ x91 ;
  assign n4907 = n4906 ^ n4714 ;
  assign n4908 = n4907 ^ n4719 ;
  assign n4909 = ~n4720 & n4908 ;
  assign n4910 = n4909 ^ n4719 ;
  assign n4911 = ~n4715 & n4910 ;
  assign n4912 = n4911 ^ x93 ;
  assign n4916 = n4915 ^ n4912 ;
  assign n4917 = n4915 ^ x94 ;
  assign n4918 = n4916 & ~n4917 ;
  assign n4919 = n4918 ^ x94 ;
  assign n4702 = n4466 ^ x94 ;
  assign n4703 = n4702 ^ n4651 ;
  assign n4704 = n4703 ^ x93 ;
  assign n4705 = n4704 ^ n4702 ;
  assign n4707 = n4651 ^ x94 ;
  assign n4708 = n4707 ^ n4702 ;
  assign n4709 = ~n4705 & ~n4708 ;
  assign n4710 = n4709 ^ n4702 ;
  assign n4711 = n4679 & ~n4710 ;
  assign n4712 = n4711 ^ n4463 ;
  assign n4920 = n4919 ^ n4712 ;
  assign n4921 = n4919 ^ x95 ;
  assign n4922 = n4920 & n4921 ;
  assign n4923 = n4922 ^ x95 ;
  assign n4699 = n4657 ^ x95 ;
  assign n4700 = n4679 & n4699 ;
  assign n4701 = n4700 ^ n4659 ;
  assign n4924 = n4923 ^ n4701 ;
  assign n4925 = n4923 ^ x96 ;
  assign n4926 = n4924 & n4925 ;
  assign n4927 = n4926 ^ x96 ;
  assign n4697 = n4665 & n4679 ;
  assign n4698 = n4697 ^ n4461 ;
  assign n4928 = n4927 ^ n4698 ;
  assign n4929 = n4927 ^ x97 ;
  assign n4930 = n4928 & n4929 ;
  assign n4931 = n4930 ^ x97 ;
  assign n4694 = n4667 ^ x97 ;
  assign n4695 = n4679 & n4694 ;
  assign n4696 = n4695 ^ n4454 ;
  assign n4932 = n4931 ^ n4696 ;
  assign n4933 = n4931 ^ x98 ;
  assign n4934 = n4932 & n4933 ;
  assign n4935 = n4934 ^ x98 ;
  assign n4683 = n4667 ^ x98 ;
  assign n4684 = n4683 ^ n4454 ;
  assign n4685 = n4684 ^ x97 ;
  assign n4686 = n4685 ^ n4683 ;
  assign n4688 = n4454 ^ x98 ;
  assign n4689 = n4688 ^ n4683 ;
  assign n4690 = n4686 & ~n4689 ;
  assign n4691 = n4690 ^ n4683 ;
  assign n4692 = n4679 & n4691 ;
  assign n4693 = n4692 ^ n4456 ;
  assign n4936 = n4935 ^ n4693 ;
  assign n4939 = n4693 ^ x99 ;
  assign n4940 = n4936 & ~n4939 ;
  assign n4937 = x100 ^ x99 ;
  assign n4941 = n4940 ^ n4937 ;
  assign n4680 = n4450 & ~n4679 ;
  assign n4946 = ~n270 & ~n4680 ;
  assign n4947 = n4946 ^ x100 ;
  assign n4948 = n4941 & n4947 ;
  assign n4949 = n4948 ^ x100 ;
  assign n4950 = n156 & ~n4949 ;
  assign n5072 = x64 & n4950 ;
  assign n5359 = n5072 ^ x27 ;
  assign n5218 = n4680 & ~n4950 ;
  assign n5219 = n5218 ^ n270 ;
  assign n5243 = x100 & ~n5219 ;
  assign n5207 = n4929 & n4950 ;
  assign n5208 = n5207 ^ n4698 ;
  assign n4953 = n4925 & n4950 ;
  assign n4954 = n4953 ^ n4701 ;
  assign n4955 = n4954 ^ x97 ;
  assign n4959 = n4954 ^ x96 ;
  assign n4956 = n4921 & n4950 ;
  assign n4957 = n4956 ^ n4712 ;
  assign n4958 = n4957 ^ n4954 ;
  assign n4960 = n4959 ^ n4958 ;
  assign n4964 = n4717 ^ x93 ;
  assign n4965 = n4964 ^ n4906 ;
  assign n4966 = n4965 ^ x92 ;
  assign n4967 = n4966 ^ n4964 ;
  assign n4969 = n4906 ^ x93 ;
  assign n4970 = n4969 ^ n4964 ;
  assign n4971 = ~n4967 & ~n4970 ;
  assign n4972 = n4971 ^ n4964 ;
  assign n4973 = n4950 & ~n4972 ;
  assign n4974 = n4973 ^ n4714 ;
  assign n4975 = n4974 ^ x94 ;
  assign n4976 = n4906 ^ x92 ;
  assign n4977 = n4950 & n4976 ;
  assign n4978 = n4977 ^ n4717 ;
  assign n4979 = n4978 ^ x93 ;
  assign n5179 = n4900 & n4950 ;
  assign n5180 = n5179 ^ n4724 ;
  assign n4980 = n4892 ^ x89 ;
  assign n4981 = n4950 & n4980 ;
  assign n4982 = n4981 ^ n4894 ;
  assign n4983 = n4982 ^ x90 ;
  assign n4996 = n4982 ^ x89 ;
  assign n4984 = n4729 ^ x88 ;
  assign n4985 = n4984 ^ n4886 ;
  assign n4986 = n4985 ^ x87 ;
  assign n4987 = n4986 ^ n4984 ;
  assign n4989 = n4886 ^ x88 ;
  assign n4990 = n4989 ^ n4984 ;
  assign n4991 = ~n4987 & ~n4990 ;
  assign n4992 = n4991 ^ n4984 ;
  assign n4993 = n4950 & ~n4992 ;
  assign n4994 = n4993 ^ n4726 ;
  assign n4995 = n4994 ^ n4982 ;
  assign n4997 = n4996 ^ n4995 ;
  assign n5130 = n4853 ^ x78 ;
  assign n5131 = n4950 & n5130 ;
  assign n5132 = n5131 ^ n4756 ;
  assign n5038 = n4850 ^ x77 ;
  assign n5039 = n4950 & n5038 ;
  assign n5040 = n5039 ^ n4759 ;
  assign n5041 = n5040 ^ x78 ;
  assign n5045 = n5040 ^ x77 ;
  assign n5042 = n4848 & n4950 ;
  assign n5043 = n5042 ^ n4762 ;
  assign n5044 = n5043 ^ n5040 ;
  assign n5046 = n5045 ^ n5044 ;
  assign n5068 = n4799 ^ x65 ;
  assign n5069 = n4950 & n5068 ;
  assign n5067 = n4801 ^ x28 ;
  assign n5070 = n5069 ^ n5067 ;
  assign n5071 = n5070 ^ x66 ;
  assign n5073 = x65 ^ x27 ;
  assign n5074 = n5073 ^ n5072 ;
  assign n5077 = ~x26 & x64 ;
  assign n5078 = n5077 ^ x65 ;
  assign n5079 = ~n5074 & n5078 ;
  assign n5080 = n5079 ^ x65 ;
  assign n5081 = n5080 ^ n5070 ;
  assign n5082 = ~n5071 & n5081 ;
  assign n5083 = n5082 ^ x66 ;
  assign n5065 = n4808 & n4950 ;
  assign n5066 = n5065 ^ n4798 ;
  assign n5084 = n5083 ^ n5066 ;
  assign n5085 = n5083 ^ x67 ;
  assign n5086 = n5084 & n5085 ;
  assign n5087 = n5086 ^ x67 ;
  assign n5063 = n4812 & n4950 ;
  assign n5064 = n5063 ^ n4791 ;
  assign n5088 = n5087 ^ n5064 ;
  assign n5089 = n5087 ^ x68 ;
  assign n5090 = n5088 & n5089 ;
  assign n5091 = n5090 ^ x68 ;
  assign n5061 = n4816 & n4950 ;
  assign n5062 = n5061 ^ n4789 ;
  assign n5092 = n5091 ^ n5062 ;
  assign n5093 = n5091 ^ x69 ;
  assign n5094 = n5092 & n5093 ;
  assign n5095 = n5094 ^ x69 ;
  assign n5059 = n4820 & n4950 ;
  assign n5060 = n5059 ^ n4787 ;
  assign n5096 = n5095 ^ n5060 ;
  assign n5097 = n5095 ^ x70 ;
  assign n5098 = n5096 & n5097 ;
  assign n5099 = n5098 ^ x70 ;
  assign n5057 = n4824 & n4950 ;
  assign n5058 = n5057 ^ n4785 ;
  assign n5100 = n5099 ^ n5058 ;
  assign n5101 = n5099 ^ x71 ;
  assign n5102 = n5100 & n5101 ;
  assign n5103 = n5102 ^ x71 ;
  assign n5055 = n4828 & n4950 ;
  assign n5056 = n5055 ^ n4782 ;
  assign n5104 = n5103 ^ n5056 ;
  assign n5105 = n5103 ^ x72 ;
  assign n5106 = n5104 & n5105 ;
  assign n5107 = n5106 ^ x72 ;
  assign n5053 = n4832 & n4950 ;
  assign n5054 = n5053 ^ n4771 ;
  assign n5108 = n5107 ^ n5054 ;
  assign n5109 = n5107 ^ x73 ;
  assign n5110 = n5108 & n5109 ;
  assign n5111 = n5110 ^ x73 ;
  assign n5051 = n4836 & n4950 ;
  assign n5052 = n5051 ^ n4768 ;
  assign n5112 = n5111 ^ n5052 ;
  assign n5113 = n5111 ^ x74 ;
  assign n5114 = n5112 & n5113 ;
  assign n5115 = n5114 ^ x74 ;
  assign n5049 = n4840 & n4950 ;
  assign n5050 = n5049 ^ n4766 ;
  assign n5116 = n5115 ^ n5050 ;
  assign n5117 = n5115 ^ x75 ;
  assign n5118 = n5116 & n5117 ;
  assign n5119 = n5118 ^ x75 ;
  assign n5047 = n4844 & n4950 ;
  assign n5048 = n5047 ^ n4764 ;
  assign n5120 = n5119 ^ n5048 ;
  assign n5121 = n5119 ^ x76 ;
  assign n5122 = n5120 & n5121 ;
  assign n5123 = n5122 ^ x76 ;
  assign n5124 = n5123 ^ n5040 ;
  assign n5125 = n5124 ^ n5045 ;
  assign n5126 = ~n5046 & n5125 ;
  assign n5127 = n5126 ^ n5045 ;
  assign n5128 = ~n5041 & n5127 ;
  assign n5129 = n5128 ^ x78 ;
  assign n5133 = n5132 ^ n5129 ;
  assign n5134 = n5132 ^ x79 ;
  assign n5135 = n5133 & ~n5134 ;
  assign n5136 = n5135 ^ x79 ;
  assign n5036 = n4858 & n4950 ;
  assign n5037 = n5036 ^ n4754 ;
  assign n5137 = n5136 ^ n5037 ;
  assign n5138 = n5136 ^ x80 ;
  assign n5139 = n5137 & n5138 ;
  assign n5140 = n5139 ^ x80 ;
  assign n5034 = n4862 & n4950 ;
  assign n5035 = n5034 ^ n4752 ;
  assign n5141 = n5140 ^ n5035 ;
  assign n5142 = n5140 ^ x81 ;
  assign n5143 = n5141 & n5142 ;
  assign n5144 = n5143 ^ x81 ;
  assign n5031 = n4864 ^ x81 ;
  assign n5032 = n4950 & n5031 ;
  assign n5033 = n5032 ^ n4747 ;
  assign n5145 = n5144 ^ n5033 ;
  assign n5146 = n5144 ^ x82 ;
  assign n5147 = n5145 & n5146 ;
  assign n5148 = n5147 ^ x82 ;
  assign n5020 = n4747 ^ x82 ;
  assign n5021 = n5020 ^ n4864 ;
  assign n5022 = n5021 ^ x81 ;
  assign n5023 = n5022 ^ n5020 ;
  assign n5025 = n4864 ^ x82 ;
  assign n5026 = n5025 ^ n5020 ;
  assign n5027 = ~n5023 & ~n5026 ;
  assign n5028 = n5027 ^ n5020 ;
  assign n5029 = n4950 & ~n5028 ;
  assign n5030 = n5029 ^ n4744 ;
  assign n5149 = n5148 ^ n5030 ;
  assign n5150 = n5148 ^ x83 ;
  assign n5151 = n5149 & n5150 ;
  assign n5152 = n5151 ^ x83 ;
  assign n5017 = n4870 ^ x83 ;
  assign n5018 = n4950 & n5017 ;
  assign n5019 = n5018 ^ n4739 ;
  assign n5153 = n5152 ^ n5019 ;
  assign n5154 = n5152 ^ x84 ;
  assign n5155 = n5153 & n5154 ;
  assign n5156 = n5155 ^ x84 ;
  assign n5006 = n4739 ^ x84 ;
  assign n5007 = n5006 ^ x83 ;
  assign n5008 = n5007 ^ n4870 ;
  assign n5009 = n5008 ^ n5006 ;
  assign n5011 = x84 ^ x83 ;
  assign n5012 = n5011 ^ n5006 ;
  assign n5013 = ~n5009 & ~n5012 ;
  assign n5014 = n5013 ^ n5006 ;
  assign n5015 = n4950 & ~n5014 ;
  assign n5016 = n5015 ^ n4736 ;
  assign n5157 = n5156 ^ n5016 ;
  assign n5158 = n5156 ^ x85 ;
  assign n5159 = n5157 & n5158 ;
  assign n5160 = n5159 ^ x85 ;
  assign n5003 = n4876 ^ x85 ;
  assign n5004 = n4950 & n5003 ;
  assign n5005 = n5004 ^ n4878 ;
  assign n5161 = n5160 ^ n5005 ;
  assign n5162 = n5160 ^ x86 ;
  assign n5163 = n5161 & n5162 ;
  assign n5164 = n5163 ^ x86 ;
  assign n5001 = n4884 & n4950 ;
  assign n5002 = n5001 ^ n4734 ;
  assign n5165 = n5164 ^ n5002 ;
  assign n5166 = n5164 ^ x87 ;
  assign n5167 = n5165 & n5166 ;
  assign n5168 = n5167 ^ x87 ;
  assign n4998 = n4886 ^ x87 ;
  assign n4999 = n4950 & n4998 ;
  assign n5000 = n4999 ^ n4729 ;
  assign n5169 = n5168 ^ n5000 ;
  assign n5170 = n5168 ^ x88 ;
  assign n5171 = n5169 & n5170 ;
  assign n5172 = n5171 ^ x88 ;
  assign n5173 = n5172 ^ n4982 ;
  assign n5174 = n5173 ^ n4996 ;
  assign n5175 = ~n4997 & n5174 ;
  assign n5176 = n5175 ^ n4996 ;
  assign n5177 = ~n4983 & n5176 ;
  assign n5178 = n5177 ^ x90 ;
  assign n5181 = n5180 ^ n5178 ;
  assign n5182 = n5180 ^ x91 ;
  assign n5183 = n5181 & ~n5182 ;
  assign n5184 = n5183 ^ x91 ;
  assign n5185 = n5184 ^ x92 ;
  assign n5186 = n4904 & n4950 ;
  assign n5187 = n5186 ^ n4722 ;
  assign n5188 = n5187 ^ n5184 ;
  assign n5189 = n5185 & n5188 ;
  assign n5190 = n5189 ^ x92 ;
  assign n5191 = n5190 ^ n4978 ;
  assign n5192 = ~n4979 & n5191 ;
  assign n5193 = n5192 ^ x93 ;
  assign n5194 = n5193 ^ n4974 ;
  assign n5195 = ~n4975 & n5194 ;
  assign n5196 = n5195 ^ x94 ;
  assign n4961 = n4912 ^ x94 ;
  assign n4962 = n4950 & n4961 ;
  assign n4963 = n4962 ^ n4915 ;
  assign n5197 = n5196 ^ n4963 ;
  assign n5198 = n5196 ^ x95 ;
  assign n5199 = n5197 & n5198 ;
  assign n5200 = n5199 ^ x95 ;
  assign n5201 = n5200 ^ n4954 ;
  assign n5202 = n5201 ^ n4959 ;
  assign n5203 = ~n4960 & n5202 ;
  assign n5204 = n5203 ^ n4959 ;
  assign n5205 = ~n4955 & n5204 ;
  assign n5206 = n5205 ^ x97 ;
  assign n5209 = n5208 ^ n5206 ;
  assign n5210 = n5208 ^ x98 ;
  assign n5211 = n5209 & ~n5210 ;
  assign n5212 = n5211 ^ x98 ;
  assign n4951 = n4933 & n4950 ;
  assign n4952 = n4951 ^ n4696 ;
  assign n5213 = n5212 ^ n4952 ;
  assign n5214 = n5212 ^ x99 ;
  assign n5215 = n5213 & n5214 ;
  assign n5216 = n5215 ^ x99 ;
  assign n5220 = n5219 ^ x101 ;
  assign n5221 = n4935 ^ x99 ;
  assign n5222 = n4950 & n5221 ;
  assign n5223 = n5222 ^ n4693 ;
  assign n5226 = n5223 ^ n5219 ;
  assign n5217 = n5216 ^ x100 ;
  assign n5224 = n5223 ^ n5216 ;
  assign n5225 = ~n5217 & ~n5224 ;
  assign n5227 = n5226 ^ n5225 ;
  assign n5228 = ~n5220 & ~n5227 ;
  assign n5229 = n5228 ^ x101 ;
  assign n5230 = n5229 ^ n5216 ;
  assign n5231 = n5230 ^ n5229 ;
  assign n5234 = n5229 ^ n5225 ;
  assign n5235 = n5234 ^ n5229 ;
  assign n5236 = n5228 & n5235 ;
  assign n5237 = n5231 & n5236 ;
  assign n5238 = n5237 ^ n5231 ;
  assign n5239 = n5238 ^ n5230 ;
  assign n5240 = n155 & ~n5239 ;
  assign n5244 = n5216 & n5240 ;
  assign n5245 = n5243 & n5244 ;
  assign n5246 = n5245 ^ n5240 ;
  assign n5358 = x65 & n5246 ;
  assign n5360 = n5359 ^ n5358 ;
  assign n5356 = x64 & n5246 ;
  assign n5357 = ~x26 & n5356 ;
  assign n5361 = n5360 ^ n5357 ;
  assign n5362 = n5361 ^ x66 ;
  assign n5363 = x64 ^ x26 ;
  assign n5364 = n5363 ^ x65 ;
  assign n5365 = n5364 ^ x65 ;
  assign n5366 = n5365 ^ x26 ;
  assign n5370 = x26 & x65 ;
  assign n5367 = x65 ^ x25 ;
  assign n5368 = n5364 ^ n5246 ;
  assign n5369 = ~n5367 & n5368 ;
  assign n5371 = n5370 ^ n5369 ;
  assign n5372 = n5366 & n5371 ;
  assign n5373 = n5372 ^ n5370 ;
  assign n5374 = n5373 ^ x65 ;
  assign n5375 = n5374 ^ n5361 ;
  assign n5376 = ~n5362 & n5375 ;
  assign n5377 = n5376 ^ x66 ;
  assign n5353 = n5080 ^ x66 ;
  assign n5354 = n5246 & n5353 ;
  assign n5355 = n5354 ^ n5070 ;
  assign n5378 = n5377 ^ n5355 ;
  assign n5379 = n5377 ^ x67 ;
  assign n5380 = n5378 & n5379 ;
  assign n5381 = n5380 ^ x67 ;
  assign n5351 = n5085 & n5246 ;
  assign n5352 = n5351 ^ n5066 ;
  assign n5382 = n5381 ^ n5352 ;
  assign n5383 = n5381 ^ x68 ;
  assign n5384 = n5382 & n5383 ;
  assign n5385 = n5384 ^ x68 ;
  assign n5349 = n5089 & n5246 ;
  assign n5350 = n5349 ^ n5064 ;
  assign n5386 = n5385 ^ n5350 ;
  assign n5387 = n5385 ^ x69 ;
  assign n5388 = n5386 & n5387 ;
  assign n5389 = n5388 ^ x69 ;
  assign n5347 = n5093 & n5246 ;
  assign n5348 = n5347 ^ n5062 ;
  assign n5390 = n5389 ^ n5348 ;
  assign n5391 = n5389 ^ x70 ;
  assign n5392 = n5390 & n5391 ;
  assign n5393 = n5392 ^ x70 ;
  assign n5345 = n5097 & n5246 ;
  assign n5346 = n5345 ^ n5060 ;
  assign n5394 = n5393 ^ n5346 ;
  assign n5395 = n5393 ^ x71 ;
  assign n5396 = n5394 & n5395 ;
  assign n5397 = n5396 ^ x71 ;
  assign n5343 = n5101 & n5246 ;
  assign n5344 = n5343 ^ n5058 ;
  assign n5398 = n5397 ^ n5344 ;
  assign n5399 = n5397 ^ x72 ;
  assign n5400 = n5398 & n5399 ;
  assign n5401 = n5400 ^ x72 ;
  assign n5341 = n5105 & n5246 ;
  assign n5342 = n5341 ^ n5056 ;
  assign n5402 = n5401 ^ n5342 ;
  assign n5403 = n5401 ^ x73 ;
  assign n5404 = n5402 & n5403 ;
  assign n5405 = n5404 ^ x73 ;
  assign n5407 = n5405 ^ x74 ;
  assign n5482 = n5190 ^ x93 ;
  assign n5483 = n5246 & n5482 ;
  assign n5484 = n5483 ^ n4978 ;
  assign n5271 = n5185 & n5246 ;
  assign n5272 = n5271 ^ n5187 ;
  assign n5273 = n5272 ^ x93 ;
  assign n5278 = n5272 ^ x92 ;
  assign n5274 = n5178 ^ x91 ;
  assign n5275 = n5246 & n5274 ;
  assign n5276 = n5275 ^ n5180 ;
  assign n5277 = n5276 ^ n5272 ;
  assign n5279 = n5278 ^ n5277 ;
  assign n5280 = n4994 ^ x90 ;
  assign n5281 = n5280 ^ n5172 ;
  assign n5282 = n5281 ^ x89 ;
  assign n5283 = n5282 ^ n5280 ;
  assign n5285 = n5172 ^ x90 ;
  assign n5286 = n5285 ^ n5280 ;
  assign n5287 = ~n5283 & ~n5286 ;
  assign n5288 = n5287 ^ n5280 ;
  assign n5289 = n5246 & ~n5288 ;
  assign n5290 = n5289 ^ n4982 ;
  assign n5291 = n5290 ^ x91 ;
  assign n5296 = n5290 ^ x90 ;
  assign n5292 = n5172 ^ x89 ;
  assign n5293 = n5246 & n5292 ;
  assign n5294 = n5293 ^ n4994 ;
  assign n5295 = n5294 ^ n5290 ;
  assign n5297 = n5296 ^ n5295 ;
  assign n5339 = n5109 & n5246 ;
  assign n5340 = n5339 ^ n5054 ;
  assign n5406 = n5405 ^ n5340 ;
  assign n5408 = n5406 & n5407 ;
  assign n5409 = n5408 ^ x74 ;
  assign n5337 = n5113 & n5246 ;
  assign n5338 = n5337 ^ n5052 ;
  assign n5410 = n5409 ^ n5338 ;
  assign n5411 = n5409 ^ x75 ;
  assign n5412 = n5410 & n5411 ;
  assign n5413 = n5412 ^ x75 ;
  assign n5335 = n5117 & n5246 ;
  assign n5336 = n5335 ^ n5050 ;
  assign n5414 = n5413 ^ n5336 ;
  assign n5415 = n5413 ^ x76 ;
  assign n5416 = n5414 & n5415 ;
  assign n5417 = n5416 ^ x76 ;
  assign n5333 = n5121 & n5246 ;
  assign n5334 = n5333 ^ n5048 ;
  assign n5418 = n5417 ^ n5334 ;
  assign n5419 = n5417 ^ x77 ;
  assign n5420 = n5418 & n5419 ;
  assign n5421 = n5420 ^ x77 ;
  assign n5330 = n5123 ^ x77 ;
  assign n5331 = n5246 & n5330 ;
  assign n5332 = n5331 ^ n5043 ;
  assign n5422 = n5421 ^ n5332 ;
  assign n5423 = n5421 ^ x78 ;
  assign n5424 = n5422 & n5423 ;
  assign n5425 = n5424 ^ x78 ;
  assign n5319 = n5043 ^ x78 ;
  assign n5320 = n5319 ^ n5123 ;
  assign n5321 = n5320 ^ x77 ;
  assign n5322 = n5321 ^ n5319 ;
  assign n5324 = n5123 ^ x78 ;
  assign n5325 = n5324 ^ n5319 ;
  assign n5326 = ~n5322 & ~n5325 ;
  assign n5327 = n5326 ^ n5319 ;
  assign n5328 = n5246 & ~n5327 ;
  assign n5329 = n5328 ^ n5040 ;
  assign n5426 = n5425 ^ n5329 ;
  assign n5427 = n5425 ^ x79 ;
  assign n5428 = n5426 & n5427 ;
  assign n5429 = n5428 ^ x79 ;
  assign n5316 = n5129 ^ x79 ;
  assign n5317 = n5246 & n5316 ;
  assign n5318 = n5317 ^ n5132 ;
  assign n5430 = n5429 ^ n5318 ;
  assign n5431 = n5429 ^ x80 ;
  assign n5432 = n5430 & n5431 ;
  assign n5433 = n5432 ^ x80 ;
  assign n5314 = n5138 & n5246 ;
  assign n5315 = n5314 ^ n5037 ;
  assign n5434 = n5433 ^ n5315 ;
  assign n5435 = n5433 ^ x81 ;
  assign n5436 = n5434 & n5435 ;
  assign n5437 = n5436 ^ x81 ;
  assign n5312 = n5142 & n5246 ;
  assign n5313 = n5312 ^ n5035 ;
  assign n5438 = n5437 ^ n5313 ;
  assign n5439 = n5437 ^ x82 ;
  assign n5440 = n5438 & n5439 ;
  assign n5441 = n5440 ^ x82 ;
  assign n5310 = n5146 & n5246 ;
  assign n5311 = n5310 ^ n5033 ;
  assign n5442 = n5441 ^ n5311 ;
  assign n5443 = n5441 ^ x83 ;
  assign n5444 = n5442 & n5443 ;
  assign n5445 = n5444 ^ x83 ;
  assign n5308 = n5150 & n5246 ;
  assign n5309 = n5308 ^ n5030 ;
  assign n5446 = n5445 ^ n5309 ;
  assign n5447 = n5445 ^ x84 ;
  assign n5448 = n5446 & n5447 ;
  assign n5449 = n5448 ^ x84 ;
  assign n5306 = n5154 & n5246 ;
  assign n5307 = n5306 ^ n5019 ;
  assign n5450 = n5449 ^ n5307 ;
  assign n5451 = n5449 ^ x85 ;
  assign n5452 = n5450 & n5451 ;
  assign n5453 = n5452 ^ x85 ;
  assign n5304 = n5158 & n5246 ;
  assign n5305 = n5304 ^ n5016 ;
  assign n5454 = n5453 ^ n5305 ;
  assign n5455 = n5453 ^ x86 ;
  assign n5456 = n5454 & n5455 ;
  assign n5457 = n5456 ^ x86 ;
  assign n5302 = n5162 & n5246 ;
  assign n5303 = n5302 ^ n5005 ;
  assign n5458 = n5457 ^ n5303 ;
  assign n5459 = n5457 ^ x87 ;
  assign n5460 = n5458 & n5459 ;
  assign n5461 = n5460 ^ x87 ;
  assign n5300 = n5166 & n5246 ;
  assign n5301 = n5300 ^ n5002 ;
  assign n5462 = n5461 ^ n5301 ;
  assign n5463 = n5461 ^ x88 ;
  assign n5464 = n5462 & n5463 ;
  assign n5465 = n5464 ^ x88 ;
  assign n5298 = n5170 & n5246 ;
  assign n5299 = n5298 ^ n5000 ;
  assign n5466 = n5465 ^ n5299 ;
  assign n5467 = n5465 ^ x89 ;
  assign n5468 = n5466 & n5467 ;
  assign n5469 = n5468 ^ x89 ;
  assign n5470 = n5469 ^ n5290 ;
  assign n5471 = n5470 ^ n5296 ;
  assign n5472 = ~n5297 & n5471 ;
  assign n5473 = n5472 ^ n5296 ;
  assign n5474 = ~n5291 & n5473 ;
  assign n5475 = n5474 ^ x91 ;
  assign n5476 = n5475 ^ n5272 ;
  assign n5477 = n5476 ^ n5278 ;
  assign n5478 = ~n5279 & n5477 ;
  assign n5479 = n5478 ^ n5278 ;
  assign n5480 = ~n5273 & n5479 ;
  assign n5481 = n5480 ^ x93 ;
  assign n5485 = n5484 ^ n5481 ;
  assign n5486 = n5484 ^ x94 ;
  assign n5487 = n5485 & ~n5486 ;
  assign n5488 = n5487 ^ x94 ;
  assign n5268 = n5193 ^ x94 ;
  assign n5269 = n5246 & n5268 ;
  assign n5270 = n5269 ^ n4974 ;
  assign n5489 = n5488 ^ n5270 ;
  assign n5490 = n5488 ^ x95 ;
  assign n5491 = n5489 & n5490 ;
  assign n5492 = n5491 ^ x95 ;
  assign n5266 = n5198 & n5246 ;
  assign n5267 = n5266 ^ n4963 ;
  assign n5493 = n5492 ^ n5267 ;
  assign n5494 = n5492 ^ x96 ;
  assign n5495 = n5493 & n5494 ;
  assign n5496 = n5495 ^ x96 ;
  assign n5263 = n5200 ^ x96 ;
  assign n5264 = n5246 & n5263 ;
  assign n5265 = n5264 ^ n4957 ;
  assign n5497 = n5496 ^ n5265 ;
  assign n5498 = n5496 ^ x97 ;
  assign n5499 = n5497 & n5498 ;
  assign n5500 = n5499 ^ x97 ;
  assign n5252 = n4957 ^ x97 ;
  assign n5253 = n5252 ^ n5200 ;
  assign n5254 = n5253 ^ x96 ;
  assign n5255 = n5254 ^ n5252 ;
  assign n5257 = n5200 ^ x97 ;
  assign n5258 = n5257 ^ n5252 ;
  assign n5259 = ~n5255 & ~n5258 ;
  assign n5260 = n5259 ^ n5252 ;
  assign n5261 = n5246 & ~n5260 ;
  assign n5262 = n5261 ^ n4954 ;
  assign n5501 = n5500 ^ n5262 ;
  assign n5502 = n5500 ^ x98 ;
  assign n5503 = n5501 & n5502 ;
  assign n5504 = n5503 ^ x98 ;
  assign n5249 = n5206 ^ x98 ;
  assign n5250 = n5246 & n5249 ;
  assign n5251 = n5250 ^ n5208 ;
  assign n5505 = n5504 ^ n5251 ;
  assign n5506 = n5504 ^ x99 ;
  assign n5507 = n5505 & n5506 ;
  assign n5508 = n5507 ^ x99 ;
  assign n5247 = n5214 & n5246 ;
  assign n5248 = n5247 ^ n4952 ;
  assign n5509 = n5508 ^ n5248 ;
  assign n5510 = n5508 ^ x100 ;
  assign n5511 = n5509 & n5510 ;
  assign n5512 = n5511 ^ x100 ;
  assign n5241 = n5217 & n5240 ;
  assign n5242 = n5241 ^ n5223 ;
  assign n5513 = n5512 ^ n5242 ;
  assign n5514 = n5512 ^ x101 ;
  assign n5515 = n5513 & n5514 ;
  assign n5516 = n5515 ^ x101 ;
  assign n5523 = n5516 ^ x102 ;
  assign n5524 = n5516 ^ n5219 ;
  assign n5526 = n5524 ^ n5240 ;
  assign n5527 = n5526 ^ n5524 ;
  assign n5530 = ~n270 & n5527 ;
  assign n5531 = n5219 & n5530 ;
  assign n5532 = n5531 ^ n5219 ;
  assign n5533 = n5532 ^ n5516 ;
  assign n5534 = n5523 & n5533 ;
  assign n5535 = n5534 ^ x102 ;
  assign n5536 = n154 & ~n5535 ;
  assign n5689 = n5407 & n5536 ;
  assign n5690 = n5689 ^ n5340 ;
  assign n5683 = n5403 & n5536 ;
  assign n5684 = n5683 ^ n5342 ;
  assign n5677 = n5399 & n5536 ;
  assign n5678 = n5677 ^ n5344 ;
  assign n5616 = n5395 & n5536 ;
  assign n5617 = n5616 ^ n5346 ;
  assign n5618 = n5617 ^ x72 ;
  assign n5622 = n5617 ^ x71 ;
  assign n5619 = n5391 & n5536 ;
  assign n5620 = n5619 ^ n5348 ;
  assign n5621 = n5620 ^ n5617 ;
  assign n5623 = n5622 ^ n5621 ;
  assign n5637 = n5356 ^ x26 ;
  assign n5634 = ~x25 & x64 ;
  assign n5635 = n5634 ^ x65 ;
  assign n5636 = n5536 & n5635 ;
  assign n5638 = n5637 ^ n5636 ;
  assign n5639 = n5638 ^ x66 ;
  assign n5647 = x25 & x65 ;
  assign n5644 = x65 ^ x24 ;
  assign n5640 = x64 ^ x25 ;
  assign n5641 = n5640 ^ x65 ;
  assign n5645 = n5641 ^ n5536 ;
  assign n5646 = ~n5644 & n5645 ;
  assign n5648 = n5647 ^ n5646 ;
  assign n5649 = x64 & n5648 ;
  assign n5650 = n5649 ^ n5647 ;
  assign n5651 = n5650 ^ x65 ;
  assign n5652 = n5651 ^ n5638 ;
  assign n5653 = ~n5639 & n5652 ;
  assign n5654 = n5653 ^ x66 ;
  assign n5630 = n5374 ^ x66 ;
  assign n5631 = n5536 & n5630 ;
  assign n5632 = n5631 ^ n5361 ;
  assign n5655 = n5654 ^ n5632 ;
  assign n5656 = n5654 ^ x67 ;
  assign n5657 = n5655 & n5656 ;
  assign n5658 = n5657 ^ x67 ;
  assign n5628 = n5379 & n5536 ;
  assign n5629 = n5628 ^ n5355 ;
  assign n5659 = n5658 ^ n5629 ;
  assign n5660 = n5658 ^ x68 ;
  assign n5661 = n5659 & n5660 ;
  assign n5662 = n5661 ^ x68 ;
  assign n5626 = n5383 & n5536 ;
  assign n5627 = n5626 ^ n5352 ;
  assign n5663 = n5662 ^ n5627 ;
  assign n5664 = n5662 ^ x69 ;
  assign n5665 = n5663 & n5664 ;
  assign n5666 = n5665 ^ x69 ;
  assign n5624 = n5387 & n5536 ;
  assign n5625 = n5624 ^ n5350 ;
  assign n5667 = n5666 ^ n5625 ;
  assign n5668 = n5666 ^ x70 ;
  assign n5669 = n5667 & n5668 ;
  assign n5670 = n5669 ^ x70 ;
  assign n5671 = n5670 ^ n5617 ;
  assign n5672 = n5671 ^ n5622 ;
  assign n5673 = ~n5623 & n5672 ;
  assign n5674 = n5673 ^ n5622 ;
  assign n5675 = ~n5618 & n5674 ;
  assign n5676 = n5675 ^ x72 ;
  assign n5679 = n5678 ^ n5676 ;
  assign n5680 = n5678 ^ x73 ;
  assign n5681 = n5679 & ~n5680 ;
  assign n5682 = n5681 ^ x73 ;
  assign n5685 = n5684 ^ n5682 ;
  assign n5686 = n5684 ^ x74 ;
  assign n5687 = n5685 & ~n5686 ;
  assign n5688 = n5687 ^ x74 ;
  assign n5691 = n5690 ^ n5688 ;
  assign n5692 = n5690 ^ x75 ;
  assign n5693 = n5691 & ~n5692 ;
  assign n5694 = n5693 ^ x75 ;
  assign n5614 = n5411 & n5536 ;
  assign n5615 = n5614 ^ n5338 ;
  assign n5695 = n5694 ^ n5615 ;
  assign n5696 = n5694 ^ x76 ;
  assign n5697 = n5695 & n5696 ;
  assign n5698 = n5697 ^ x76 ;
  assign n5612 = n5415 & n5536 ;
  assign n5613 = n5612 ^ n5336 ;
  assign n5699 = n5698 ^ n5613 ;
  assign n5700 = n5698 ^ x77 ;
  assign n5701 = n5699 & n5700 ;
  assign n5702 = n5701 ^ x77 ;
  assign n5610 = n5419 & n5536 ;
  assign n5611 = n5610 ^ n5334 ;
  assign n5703 = n5702 ^ n5611 ;
  assign n5704 = n5702 ^ x78 ;
  assign n5705 = n5703 & n5704 ;
  assign n5706 = n5705 ^ x78 ;
  assign n5608 = n5423 & n5536 ;
  assign n5609 = n5608 ^ n5332 ;
  assign n5707 = n5706 ^ n5609 ;
  assign n5708 = n5706 ^ x79 ;
  assign n5709 = n5707 & n5708 ;
  assign n5710 = n5709 ^ x79 ;
  assign n5606 = n5427 & n5536 ;
  assign n5607 = n5606 ^ n5329 ;
  assign n5711 = n5710 ^ n5607 ;
  assign n5712 = n5710 ^ x80 ;
  assign n5713 = n5711 & n5712 ;
  assign n5714 = n5713 ^ x80 ;
  assign n5604 = n5431 & n5536 ;
  assign n5605 = n5604 ^ n5318 ;
  assign n5715 = n5714 ^ n5605 ;
  assign n5716 = n5714 ^ x81 ;
  assign n5717 = n5715 & n5716 ;
  assign n5718 = n5717 ^ x81 ;
  assign n5602 = n5435 & n5536 ;
  assign n5603 = n5602 ^ n5315 ;
  assign n5719 = n5718 ^ n5603 ;
  assign n5720 = n5718 ^ x82 ;
  assign n5721 = n5719 & n5720 ;
  assign n5722 = n5721 ^ x82 ;
  assign n5600 = n5439 & n5536 ;
  assign n5601 = n5600 ^ n5313 ;
  assign n5723 = n5722 ^ n5601 ;
  assign n5724 = n5722 ^ x83 ;
  assign n5725 = n5723 & n5724 ;
  assign n5726 = n5725 ^ x83 ;
  assign n5598 = n5443 & n5536 ;
  assign n5599 = n5598 ^ n5311 ;
  assign n5727 = n5726 ^ n5599 ;
  assign n5728 = n5726 ^ x84 ;
  assign n5729 = n5727 & n5728 ;
  assign n5730 = n5729 ^ x84 ;
  assign n5596 = n5447 & n5536 ;
  assign n5597 = n5596 ^ n5309 ;
  assign n5731 = n5730 ^ n5597 ;
  assign n5732 = n5730 ^ x85 ;
  assign n5733 = n5731 & n5732 ;
  assign n5734 = n5733 ^ x85 ;
  assign n5594 = n5451 & n5536 ;
  assign n5595 = n5594 ^ n5307 ;
  assign n5735 = n5734 ^ n5595 ;
  assign n5736 = n5734 ^ x86 ;
  assign n5737 = n5735 & n5736 ;
  assign n5738 = n5737 ^ x86 ;
  assign n5592 = n5455 & n5536 ;
  assign n5593 = n5592 ^ n5305 ;
  assign n5739 = n5738 ^ n5593 ;
  assign n5740 = n5738 ^ x87 ;
  assign n5741 = n5739 & n5740 ;
  assign n5742 = n5741 ^ x87 ;
  assign n5590 = n5459 & n5536 ;
  assign n5591 = n5590 ^ n5303 ;
  assign n5743 = n5742 ^ n5591 ;
  assign n5744 = n5742 ^ x88 ;
  assign n5745 = n5743 & n5744 ;
  assign n5746 = n5745 ^ x88 ;
  assign n5588 = n5463 & n5536 ;
  assign n5589 = n5588 ^ n5301 ;
  assign n5747 = n5746 ^ n5589 ;
  assign n5748 = n5746 ^ x89 ;
  assign n5749 = n5747 & n5748 ;
  assign n5750 = n5749 ^ x89 ;
  assign n5586 = n5467 & n5536 ;
  assign n5587 = n5586 ^ n5299 ;
  assign n5751 = n5750 ^ n5587 ;
  assign n5752 = n5750 ^ x90 ;
  assign n5753 = n5751 & n5752 ;
  assign n5754 = n5753 ^ x90 ;
  assign n5583 = n5469 ^ x90 ;
  assign n5584 = n5536 & n5583 ;
  assign n5585 = n5584 ^ n5294 ;
  assign n5755 = n5754 ^ n5585 ;
  assign n5756 = n5754 ^ x91 ;
  assign n5757 = n5755 & n5756 ;
  assign n5758 = n5757 ^ x91 ;
  assign n5572 = n5294 ^ x91 ;
  assign n5573 = n5572 ^ n5469 ;
  assign n5574 = n5573 ^ x90 ;
  assign n5575 = n5574 ^ n5572 ;
  assign n5577 = n5469 ^ x91 ;
  assign n5578 = n5577 ^ n5572 ;
  assign n5579 = ~n5575 & ~n5578 ;
  assign n5580 = n5579 ^ n5572 ;
  assign n5581 = n5536 & ~n5580 ;
  assign n5582 = n5581 ^ n5290 ;
  assign n5759 = n5758 ^ n5582 ;
  assign n5760 = n5758 ^ x92 ;
  assign n5761 = n5759 & n5760 ;
  assign n5762 = n5761 ^ x92 ;
  assign n5569 = n5475 ^ x92 ;
  assign n5570 = n5536 & n5569 ;
  assign n5571 = n5570 ^ n5276 ;
  assign n5763 = n5762 ^ n5571 ;
  assign n5764 = n5762 ^ x93 ;
  assign n5765 = n5763 & n5764 ;
  assign n5766 = n5765 ^ x93 ;
  assign n5558 = n5276 ^ x93 ;
  assign n5559 = n5558 ^ x92 ;
  assign n5560 = n5559 ^ n5475 ;
  assign n5561 = n5560 ^ n5558 ;
  assign n5564 = n5558 ^ n3523 ;
  assign n5565 = ~n5561 & ~n5564 ;
  assign n5566 = n5565 ^ n5558 ;
  assign n5567 = n5536 & ~n5566 ;
  assign n5568 = n5567 ^ n5272 ;
  assign n5767 = n5766 ^ n5568 ;
  assign n5768 = n5766 ^ x94 ;
  assign n5769 = n5767 & n5768 ;
  assign n5770 = n5769 ^ x94 ;
  assign n5555 = n5481 ^ x94 ;
  assign n5556 = n5536 & n5555 ;
  assign n5557 = n5556 ^ n5484 ;
  assign n5771 = n5770 ^ n5557 ;
  assign n5772 = n5770 ^ x95 ;
  assign n5773 = n5771 & n5772 ;
  assign n5774 = n5773 ^ x95 ;
  assign n5776 = n5774 ^ x96 ;
  assign n5537 = n5514 & n5536 ;
  assign n5538 = n5537 ^ n5242 ;
  assign n5520 = x103 ^ x102 ;
  assign n5521 = n5520 ^ n153 ;
  assign n5522 = n5521 ^ x102 ;
  assign n5539 = n5538 ^ n5522 ;
  assign n5540 = n5539 ^ n5521 ;
  assign n5547 = n5498 & n5536 ;
  assign n5548 = n5547 ^ n5265 ;
  assign n5549 = n5548 ^ x98 ;
  assign n5550 = n5494 & n5536 ;
  assign n5551 = n5550 ^ n5267 ;
  assign n5552 = n5551 ^ x97 ;
  assign n5553 = n5490 & n5536 ;
  assign n5554 = n5553 ^ n5270 ;
  assign n5775 = n5774 ^ n5554 ;
  assign n5777 = n5775 & n5776 ;
  assign n5778 = n5777 ^ x96 ;
  assign n5779 = n5778 ^ n5551 ;
  assign n5780 = ~n5552 & n5779 ;
  assign n5781 = n5780 ^ x97 ;
  assign n5782 = n5781 ^ n5548 ;
  assign n5783 = ~n5549 & n5782 ;
  assign n5784 = n5783 ^ x98 ;
  assign n5545 = n5502 & n5536 ;
  assign n5546 = n5545 ^ n5262 ;
  assign n5785 = n5784 ^ n5546 ;
  assign n5786 = n5784 ^ x99 ;
  assign n5787 = n5785 & n5786 ;
  assign n5788 = n5787 ^ x99 ;
  assign n5543 = n5506 & n5536 ;
  assign n5544 = n5543 ^ n5251 ;
  assign n5789 = n5788 ^ n5544 ;
  assign n5790 = n5788 ^ x100 ;
  assign n5791 = n5789 & n5790 ;
  assign n5792 = n5791 ^ x100 ;
  assign n5541 = n5510 & n5536 ;
  assign n5542 = n5541 ^ n5248 ;
  assign n5793 = n5792 ^ n5542 ;
  assign n5796 = n5542 ^ x101 ;
  assign n5797 = n5793 & ~n5796 ;
  assign n5794 = x102 ^ x101 ;
  assign n5798 = n5797 ^ n5794 ;
  assign n5801 = ~n5540 & n5798 ;
  assign n5802 = n5801 ^ n5521 ;
  assign n4681 = n154 & n4680 ;
  assign n4682 = x102 & n4681 ;
  assign n5517 = n4682 & n5516 ;
  assign n5518 = n5517 ^ n4681 ;
  assign n5519 = n5518 ^ n4680 ;
  assign n5805 = n5519 ^ n270 ;
  assign n5806 = n5805 ^ n5219 ;
  assign n5807 = ~x103 & ~n5806 ;
  assign n5808 = n5807 ^ n5219 ;
  assign n5809 = ~n5802 & n5808 ;
  assign n5810 = n5809 ^ x103 ;
  assign n5811 = n153 & ~n5810 ;
  assign n5836 = n5776 & n5811 ;
  assign n5837 = n5836 ^ n5554 ;
  assign n5838 = n5837 ^ x97 ;
  assign n5839 = n5772 & n5811 ;
  assign n5840 = n5839 ^ n5557 ;
  assign n5841 = n5840 ^ x96 ;
  assign n6045 = n5764 & n5811 ;
  assign n6046 = n6045 ^ n5571 ;
  assign n5844 = n5760 & n5811 ;
  assign n5845 = n5844 ^ n5582 ;
  assign n5846 = n5845 ^ x93 ;
  assign n5850 = n5845 ^ x92 ;
  assign n5847 = n5756 & n5811 ;
  assign n5848 = n5847 ^ n5585 ;
  assign n5849 = n5848 ^ n5845 ;
  assign n5851 = n5850 ^ n5849 ;
  assign n6029 = n5748 & n5811 ;
  assign n6030 = n6029 ^ n5589 ;
  assign n5854 = n5744 & n5811 ;
  assign n5855 = n5854 ^ n5591 ;
  assign n5856 = n5855 ^ x89 ;
  assign n5860 = n5855 ^ x88 ;
  assign n5857 = n5740 & n5811 ;
  assign n5858 = n5857 ^ n5593 ;
  assign n5859 = n5858 ^ n5855 ;
  assign n5861 = n5860 ^ n5859 ;
  assign n5862 = n5736 & n5811 ;
  assign n5863 = n5862 ^ n5595 ;
  assign n5864 = n5863 ^ x87 ;
  assign n5868 = n5863 ^ x86 ;
  assign n5865 = n5732 & n5811 ;
  assign n5866 = n5865 ^ n5597 ;
  assign n5867 = n5866 ^ n5863 ;
  assign n5869 = n5868 ^ n5867 ;
  assign n5927 = x64 & n5536 ;
  assign n5923 = ~x24 & x64 ;
  assign n5924 = n5923 ^ x65 ;
  assign n5925 = n5811 & n5924 ;
  assign n5926 = n5925 ^ x25 ;
  assign n5928 = n5927 ^ n5926 ;
  assign n5929 = n5928 ^ x66 ;
  assign n5933 = x64 & n5811 ;
  assign n5934 = n5933 ^ x24 ;
  assign n5930 = ~x23 & x64 ;
  assign n5935 = n5934 ^ n5930 ;
  assign n5936 = x65 & ~n5935 ;
  assign n5931 = n5811 ^ x24 ;
  assign n5932 = n5930 & ~n5931 ;
  assign n5937 = n5936 ^ n5932 ;
  assign n5938 = n5937 ^ n5928 ;
  assign n5939 = ~n5929 & n5938 ;
  assign n5940 = n5939 ^ x66 ;
  assign n5919 = n5651 ^ x66 ;
  assign n5920 = n5811 & n5919 ;
  assign n5921 = n5920 ^ n5638 ;
  assign n5941 = n5940 ^ n5921 ;
  assign n5942 = n5940 ^ x67 ;
  assign n5943 = n5941 & n5942 ;
  assign n5944 = n5943 ^ x67 ;
  assign n5917 = n5656 & n5811 ;
  assign n5918 = n5917 ^ n5632 ;
  assign n5945 = n5944 ^ n5918 ;
  assign n5946 = n5944 ^ x68 ;
  assign n5947 = n5945 & n5946 ;
  assign n5948 = n5947 ^ x68 ;
  assign n5915 = n5660 & n5811 ;
  assign n5916 = n5915 ^ n5629 ;
  assign n5949 = n5948 ^ n5916 ;
  assign n5950 = n5948 ^ x69 ;
  assign n5951 = n5949 & n5950 ;
  assign n5952 = n5951 ^ x69 ;
  assign n5913 = n5664 & n5811 ;
  assign n5914 = n5913 ^ n5627 ;
  assign n5953 = n5952 ^ n5914 ;
  assign n5954 = n5952 ^ x70 ;
  assign n5955 = n5953 & n5954 ;
  assign n5956 = n5955 ^ x70 ;
  assign n5911 = n5668 & n5811 ;
  assign n5912 = n5911 ^ n5625 ;
  assign n5957 = n5956 ^ n5912 ;
  assign n5958 = n5956 ^ x71 ;
  assign n5959 = n5957 & n5958 ;
  assign n5960 = n5959 ^ x71 ;
  assign n5908 = n5670 ^ x71 ;
  assign n5909 = n5811 & n5908 ;
  assign n5910 = n5909 ^ n5620 ;
  assign n5961 = n5960 ^ n5910 ;
  assign n5962 = n5960 ^ x72 ;
  assign n5963 = n5961 & n5962 ;
  assign n5964 = n5963 ^ x72 ;
  assign n5897 = n5620 ^ x72 ;
  assign n5898 = n5897 ^ n5670 ;
  assign n5899 = n5898 ^ x71 ;
  assign n5900 = n5899 ^ n5897 ;
  assign n5902 = n5670 ^ x72 ;
  assign n5903 = n5902 ^ n5897 ;
  assign n5904 = ~n5900 & ~n5903 ;
  assign n5905 = n5904 ^ n5897 ;
  assign n5906 = n5811 & ~n5905 ;
  assign n5907 = n5906 ^ n5617 ;
  assign n5965 = n5964 ^ n5907 ;
  assign n5966 = n5964 ^ x73 ;
  assign n5967 = n5965 & n5966 ;
  assign n5968 = n5967 ^ x73 ;
  assign n5894 = n5676 ^ x73 ;
  assign n5895 = n5811 & n5894 ;
  assign n5896 = n5895 ^ n5678 ;
  assign n5969 = n5968 ^ n5896 ;
  assign n5970 = n5968 ^ x74 ;
  assign n5971 = n5969 & n5970 ;
  assign n5972 = n5971 ^ x74 ;
  assign n5891 = n5682 ^ x74 ;
  assign n5892 = n5811 & n5891 ;
  assign n5893 = n5892 ^ n5684 ;
  assign n5973 = n5972 ^ n5893 ;
  assign n5974 = n5972 ^ x75 ;
  assign n5975 = n5973 & n5974 ;
  assign n5976 = n5975 ^ x75 ;
  assign n5888 = n5688 ^ x75 ;
  assign n5889 = n5811 & n5888 ;
  assign n5890 = n5889 ^ n5690 ;
  assign n5977 = n5976 ^ n5890 ;
  assign n5978 = n5976 ^ x76 ;
  assign n5979 = n5977 & n5978 ;
  assign n5980 = n5979 ^ x76 ;
  assign n5886 = n5696 & n5811 ;
  assign n5887 = n5886 ^ n5615 ;
  assign n5981 = n5980 ^ n5887 ;
  assign n5982 = n5980 ^ x77 ;
  assign n5983 = n5981 & n5982 ;
  assign n5984 = n5983 ^ x77 ;
  assign n5884 = n5700 & n5811 ;
  assign n5885 = n5884 ^ n5613 ;
  assign n5985 = n5984 ^ n5885 ;
  assign n5986 = n5984 ^ x78 ;
  assign n5987 = n5985 & n5986 ;
  assign n5988 = n5987 ^ x78 ;
  assign n5882 = n5704 & n5811 ;
  assign n5883 = n5882 ^ n5611 ;
  assign n5989 = n5988 ^ n5883 ;
  assign n5990 = n5988 ^ x79 ;
  assign n5991 = n5989 & n5990 ;
  assign n5992 = n5991 ^ x79 ;
  assign n5880 = n5708 & n5811 ;
  assign n5881 = n5880 ^ n5609 ;
  assign n5993 = n5992 ^ n5881 ;
  assign n5994 = n5992 ^ x80 ;
  assign n5995 = n5993 & n5994 ;
  assign n5996 = n5995 ^ x80 ;
  assign n5878 = n5712 & n5811 ;
  assign n5879 = n5878 ^ n5607 ;
  assign n5997 = n5996 ^ n5879 ;
  assign n5998 = n5996 ^ x81 ;
  assign n5999 = n5997 & n5998 ;
  assign n6000 = n5999 ^ x81 ;
  assign n5876 = n5716 & n5811 ;
  assign n5877 = n5876 ^ n5605 ;
  assign n6001 = n6000 ^ n5877 ;
  assign n6002 = n6000 ^ x82 ;
  assign n6003 = n6001 & n6002 ;
  assign n6004 = n6003 ^ x82 ;
  assign n5874 = n5720 & n5811 ;
  assign n5875 = n5874 ^ n5603 ;
  assign n6005 = n6004 ^ n5875 ;
  assign n6006 = n6004 ^ x83 ;
  assign n6007 = n6005 & n6006 ;
  assign n6008 = n6007 ^ x83 ;
  assign n5872 = n5724 & n5811 ;
  assign n5873 = n5872 ^ n5601 ;
  assign n6009 = n6008 ^ n5873 ;
  assign n6010 = n6008 ^ x84 ;
  assign n6011 = n6009 & n6010 ;
  assign n6012 = n6011 ^ x84 ;
  assign n5870 = n5728 & n5811 ;
  assign n5871 = n5870 ^ n5599 ;
  assign n6013 = n6012 ^ n5871 ;
  assign n6014 = n6012 ^ x85 ;
  assign n6015 = n6013 & n6014 ;
  assign n6016 = n6015 ^ x85 ;
  assign n6017 = n6016 ^ n5863 ;
  assign n6018 = n6017 ^ n5868 ;
  assign n6019 = ~n5869 & n6018 ;
  assign n6020 = n6019 ^ n5868 ;
  assign n6021 = ~n5864 & n6020 ;
  assign n6022 = n6021 ^ x87 ;
  assign n6023 = n6022 ^ n5855 ;
  assign n6024 = n6023 ^ n5860 ;
  assign n6025 = ~n5861 & n6024 ;
  assign n6026 = n6025 ^ n5860 ;
  assign n6027 = ~n5856 & n6026 ;
  assign n6028 = n6027 ^ x89 ;
  assign n6031 = n6030 ^ n6028 ;
  assign n6032 = n6030 ^ x90 ;
  assign n6033 = n6031 & ~n6032 ;
  assign n6034 = n6033 ^ x90 ;
  assign n5852 = n5752 & n5811 ;
  assign n5853 = n5852 ^ n5587 ;
  assign n6035 = n6034 ^ n5853 ;
  assign n6036 = n6034 ^ x91 ;
  assign n6037 = n6035 & n6036 ;
  assign n6038 = n6037 ^ x91 ;
  assign n6039 = n6038 ^ n5845 ;
  assign n6040 = n6039 ^ n5850 ;
  assign n6041 = ~n5851 & n6040 ;
  assign n6042 = n6041 ^ n5850 ;
  assign n6043 = ~n5846 & n6042 ;
  assign n6044 = n6043 ^ x93 ;
  assign n6047 = n6046 ^ n6044 ;
  assign n6048 = n6046 ^ x94 ;
  assign n6049 = n6047 & ~n6048 ;
  assign n6050 = n6049 ^ x94 ;
  assign n5842 = n5768 & n5811 ;
  assign n5843 = n5842 ^ n5568 ;
  assign n6051 = n6050 ^ n5843 ;
  assign n6052 = n6050 ^ x95 ;
  assign n6053 = n6051 & n6052 ;
  assign n6054 = n6053 ^ x95 ;
  assign n6055 = n6054 ^ n5840 ;
  assign n6056 = ~n5841 & n6055 ;
  assign n6057 = n6056 ^ x96 ;
  assign n6058 = n6057 ^ n5837 ;
  assign n6059 = ~n5838 & n6058 ;
  assign n6060 = n6059 ^ x97 ;
  assign n6062 = n6060 ^ x98 ;
  assign n5814 = n150 & n5813 ;
  assign n5815 = ~x105 & n5814 ;
  assign n5812 = n5519 & ~n5811 ;
  assign n5816 = n5812 ^ n270 ;
  assign n5817 = n5816 ^ x104 ;
  assign n5821 = n5816 ^ x103 ;
  assign n5818 = n5798 & n5811 ;
  assign n5819 = n5818 ^ n5538 ;
  assign n5820 = n5819 ^ n5816 ;
  assign n5822 = n5821 ^ n5820 ;
  assign n5833 = n5778 ^ x97 ;
  assign n5834 = n5811 & n5833 ;
  assign n5835 = n5834 ^ n5551 ;
  assign n6061 = n6060 ^ n5835 ;
  assign n6063 = n6061 & n6062 ;
  assign n6064 = n6063 ^ x98 ;
  assign n5830 = n5781 ^ x98 ;
  assign n5831 = n5811 & n5830 ;
  assign n5832 = n5831 ^ n5548 ;
  assign n6065 = n6064 ^ n5832 ;
  assign n6066 = n6064 ^ x99 ;
  assign n6067 = n6065 & n6066 ;
  assign n6068 = n6067 ^ x99 ;
  assign n5828 = n5786 & n5811 ;
  assign n5829 = n5828 ^ n5546 ;
  assign n6069 = n6068 ^ n5829 ;
  assign n6070 = n6068 ^ x100 ;
  assign n6071 = n6069 & n6070 ;
  assign n6072 = n6071 ^ x100 ;
  assign n5826 = n5790 & n5811 ;
  assign n5827 = n5826 ^ n5544 ;
  assign n6073 = n6072 ^ n5827 ;
  assign n6074 = n6072 ^ x101 ;
  assign n6075 = n6073 & n6074 ;
  assign n6076 = n6075 ^ x101 ;
  assign n5823 = n5792 ^ x101 ;
  assign n5824 = n5811 & n5823 ;
  assign n5825 = n5824 ^ n5542 ;
  assign n6077 = n6076 ^ n5825 ;
  assign n6078 = n6076 ^ x102 ;
  assign n6079 = n6077 & n6078 ;
  assign n6080 = n6079 ^ x102 ;
  assign n6081 = n6080 ^ n5816 ;
  assign n6082 = n6081 ^ n5821 ;
  assign n6083 = ~n5822 & n6082 ;
  assign n6084 = n6083 ^ n5821 ;
  assign n6085 = ~n5817 & n6084 ;
  assign n6086 = n6085 ^ x104 ;
  assign n6087 = n5815 & ~n6086 ;
  assign n6097 = n6062 & n6087 ;
  assign n6098 = n6097 ^ n5835 ;
  assign n6099 = n6098 ^ x99 ;
  assign n6235 = n5962 & n6087 ;
  assign n6236 = n6235 ^ n5910 ;
  assign n6182 = n5958 & n6087 ;
  assign n6183 = n6182 ^ n5912 ;
  assign n6184 = n6183 ^ x72 ;
  assign n6188 = n6183 ^ x71 ;
  assign n6185 = n5954 & n6087 ;
  assign n6186 = n6185 ^ n5914 ;
  assign n6187 = n6186 ^ n6183 ;
  assign n6189 = n6188 ^ n6187 ;
  assign n6199 = n5930 ^ x65 ;
  assign n6200 = n6087 & n6199 ;
  assign n6201 = n6200 ^ n5934 ;
  assign n6202 = n6201 ^ x66 ;
  assign n6203 = ~x22 & x64 ;
  assign n6204 = n6203 ^ x65 ;
  assign n6205 = x64 & n6087 ;
  assign n6206 = n6205 ^ x23 ;
  assign n6207 = n6206 ^ n6203 ;
  assign n6208 = n6204 & n6207 ;
  assign n6209 = n6208 ^ x65 ;
  assign n6210 = n6209 ^ n6201 ;
  assign n6211 = ~n6202 & n6210 ;
  assign n6212 = n6211 ^ x66 ;
  assign n6196 = n5937 ^ x66 ;
  assign n6197 = n6087 & n6196 ;
  assign n6198 = n6197 ^ n5928 ;
  assign n6213 = n6212 ^ n6198 ;
  assign n6214 = n6212 ^ x67 ;
  assign n6215 = n6213 & n6214 ;
  assign n6216 = n6215 ^ x67 ;
  assign n6194 = n5942 & n6087 ;
  assign n6195 = n6194 ^ n5921 ;
  assign n6217 = n6216 ^ n6195 ;
  assign n6218 = n6216 ^ x68 ;
  assign n6219 = n6217 & n6218 ;
  assign n6220 = n6219 ^ x68 ;
  assign n6192 = n5946 & n6087 ;
  assign n6193 = n6192 ^ n5918 ;
  assign n6221 = n6220 ^ n6193 ;
  assign n6222 = n6220 ^ x69 ;
  assign n6223 = n6221 & n6222 ;
  assign n6224 = n6223 ^ x69 ;
  assign n6190 = n5950 & n6087 ;
  assign n6191 = n6190 ^ n5916 ;
  assign n6225 = n6224 ^ n6191 ;
  assign n6226 = n6224 ^ x70 ;
  assign n6227 = n6225 & n6226 ;
  assign n6228 = n6227 ^ x70 ;
  assign n6229 = n6228 ^ n6183 ;
  assign n6230 = n6229 ^ n6188 ;
  assign n6231 = ~n6189 & n6230 ;
  assign n6232 = n6231 ^ n6188 ;
  assign n6233 = ~n6184 & n6232 ;
  assign n6234 = n6233 ^ x72 ;
  assign n6237 = n6236 ^ n6234 ;
  assign n6238 = n6236 ^ x73 ;
  assign n6239 = n6237 & ~n6238 ;
  assign n6240 = n6239 ^ x73 ;
  assign n6180 = n5966 & n6087 ;
  assign n6181 = n6180 ^ n5907 ;
  assign n6241 = n6240 ^ n6181 ;
  assign n6242 = n6240 ^ x74 ;
  assign n6243 = n6241 & n6242 ;
  assign n6244 = n6243 ^ x74 ;
  assign n6178 = n5970 & n6087 ;
  assign n6179 = n6178 ^ n5896 ;
  assign n6245 = n6244 ^ n6179 ;
  assign n6246 = n6244 ^ x75 ;
  assign n6247 = n6245 & n6246 ;
  assign n6248 = n6247 ^ x75 ;
  assign n6176 = n5974 & n6087 ;
  assign n6177 = n6176 ^ n5893 ;
  assign n6249 = n6248 ^ n6177 ;
  assign n6250 = n6248 ^ x76 ;
  assign n6251 = n6249 & n6250 ;
  assign n6252 = n6251 ^ x76 ;
  assign n6174 = n5978 & n6087 ;
  assign n6175 = n6174 ^ n5890 ;
  assign n6253 = n6252 ^ n6175 ;
  assign n6254 = n6252 ^ x77 ;
  assign n6255 = n6253 & n6254 ;
  assign n6256 = n6255 ^ x77 ;
  assign n6172 = n5982 & n6087 ;
  assign n6173 = n6172 ^ n5887 ;
  assign n6257 = n6256 ^ n6173 ;
  assign n6258 = n6256 ^ x78 ;
  assign n6259 = n6257 & n6258 ;
  assign n6260 = n6259 ^ x78 ;
  assign n6170 = n5986 & n6087 ;
  assign n6171 = n6170 ^ n5885 ;
  assign n6261 = n6260 ^ n6171 ;
  assign n6262 = n6260 ^ x79 ;
  assign n6263 = n6261 & n6262 ;
  assign n6264 = n6263 ^ x79 ;
  assign n6168 = n5990 & n6087 ;
  assign n6169 = n6168 ^ n5883 ;
  assign n6265 = n6264 ^ n6169 ;
  assign n6266 = n6264 ^ x80 ;
  assign n6267 = n6265 & n6266 ;
  assign n6268 = n6267 ^ x80 ;
  assign n6166 = n5994 & n6087 ;
  assign n6167 = n6166 ^ n5881 ;
  assign n6269 = n6268 ^ n6167 ;
  assign n6270 = n6268 ^ x81 ;
  assign n6271 = n6269 & n6270 ;
  assign n6272 = n6271 ^ x81 ;
  assign n6164 = n5998 & n6087 ;
  assign n6165 = n6164 ^ n5879 ;
  assign n6273 = n6272 ^ n6165 ;
  assign n6274 = n6272 ^ x82 ;
  assign n6275 = n6273 & n6274 ;
  assign n6276 = n6275 ^ x82 ;
  assign n6162 = n6002 & n6087 ;
  assign n6163 = n6162 ^ n5877 ;
  assign n6277 = n6276 ^ n6163 ;
  assign n6278 = n6276 ^ x83 ;
  assign n6279 = n6277 & n6278 ;
  assign n6280 = n6279 ^ x83 ;
  assign n6160 = n6006 & n6087 ;
  assign n6161 = n6160 ^ n5875 ;
  assign n6281 = n6280 ^ n6161 ;
  assign n6282 = n6280 ^ x84 ;
  assign n6283 = n6281 & n6282 ;
  assign n6284 = n6283 ^ x84 ;
  assign n6158 = n6010 & n6087 ;
  assign n6159 = n6158 ^ n5873 ;
  assign n6285 = n6284 ^ n6159 ;
  assign n6286 = n6284 ^ x85 ;
  assign n6287 = n6285 & n6286 ;
  assign n6288 = n6287 ^ x85 ;
  assign n6156 = n6014 & n6087 ;
  assign n6157 = n6156 ^ n5871 ;
  assign n6289 = n6288 ^ n6157 ;
  assign n6290 = n6288 ^ x86 ;
  assign n6291 = n6289 & n6290 ;
  assign n6292 = n6291 ^ x86 ;
  assign n6153 = n6016 ^ x86 ;
  assign n6154 = n6087 & n6153 ;
  assign n6155 = n6154 ^ n5866 ;
  assign n6293 = n6292 ^ n6155 ;
  assign n6294 = n6292 ^ x87 ;
  assign n6295 = n6293 & n6294 ;
  assign n6296 = n6295 ^ x87 ;
  assign n6142 = n5866 ^ x87 ;
  assign n6143 = n6142 ^ n6016 ;
  assign n6144 = n6143 ^ x86 ;
  assign n6145 = n6144 ^ n6142 ;
  assign n6147 = n6016 ^ x87 ;
  assign n6148 = n6147 ^ n6142 ;
  assign n6149 = ~n6145 & ~n6148 ;
  assign n6150 = n6149 ^ n6142 ;
  assign n6151 = n6087 & ~n6150 ;
  assign n6152 = n6151 ^ n5863 ;
  assign n6297 = n6296 ^ n6152 ;
  assign n6298 = n6296 ^ x88 ;
  assign n6299 = n6297 & n6298 ;
  assign n6300 = n6299 ^ x88 ;
  assign n6139 = n6022 ^ x88 ;
  assign n6140 = n6087 & n6139 ;
  assign n6141 = n6140 ^ n5858 ;
  assign n6301 = n6300 ^ n6141 ;
  assign n6302 = n6300 ^ x89 ;
  assign n6303 = n6301 & n6302 ;
  assign n6304 = n6303 ^ x89 ;
  assign n6128 = n5858 ^ x89 ;
  assign n6129 = n6128 ^ x88 ;
  assign n6130 = n6129 ^ n6022 ;
  assign n6131 = n6130 ^ n6128 ;
  assign n6133 = x89 ^ x88 ;
  assign n6134 = n6133 ^ n6128 ;
  assign n6135 = ~n6131 & ~n6134 ;
  assign n6136 = n6135 ^ n6128 ;
  assign n6137 = n6087 & ~n6136 ;
  assign n6138 = n6137 ^ n5855 ;
  assign n6305 = n6304 ^ n6138 ;
  assign n6306 = n6304 ^ x90 ;
  assign n6307 = n6305 & n6306 ;
  assign n6308 = n6307 ^ x90 ;
  assign n6125 = n6028 ^ x90 ;
  assign n6126 = n6087 & n6125 ;
  assign n6127 = n6126 ^ n6030 ;
  assign n6309 = n6308 ^ n6127 ;
  assign n6310 = n6308 ^ x91 ;
  assign n6311 = n6309 & n6310 ;
  assign n6312 = n6311 ^ x91 ;
  assign n6123 = n6036 & n6087 ;
  assign n6124 = n6123 ^ n5853 ;
  assign n6313 = n6312 ^ n6124 ;
  assign n6314 = n6312 ^ x92 ;
  assign n6315 = n6313 & n6314 ;
  assign n6316 = n6315 ^ x92 ;
  assign n6120 = n6038 ^ x92 ;
  assign n6121 = n6087 & n6120 ;
  assign n6122 = n6121 ^ n5848 ;
  assign n6317 = n6316 ^ n6122 ;
  assign n6318 = n6316 ^ x93 ;
  assign n6319 = n6317 & n6318 ;
  assign n6320 = n6319 ^ x93 ;
  assign n6109 = n5848 ^ x93 ;
  assign n6110 = n6109 ^ n6038 ;
  assign n6111 = n6110 ^ x92 ;
  assign n6112 = n6111 ^ n6109 ;
  assign n6114 = n6038 ^ x93 ;
  assign n6115 = n6114 ^ n6109 ;
  assign n6116 = ~n6112 & ~n6115 ;
  assign n6117 = n6116 ^ n6109 ;
  assign n6118 = n6087 & ~n6117 ;
  assign n6119 = n6118 ^ n5845 ;
  assign n6321 = n6320 ^ n6119 ;
  assign n6322 = n6320 ^ x94 ;
  assign n6323 = n6321 & n6322 ;
  assign n6324 = n6323 ^ x94 ;
  assign n6106 = n6044 ^ x94 ;
  assign n6107 = n6087 & n6106 ;
  assign n6108 = n6107 ^ n6046 ;
  assign n6325 = n6324 ^ n6108 ;
  assign n6326 = n6324 ^ x95 ;
  assign n6327 = n6325 & n6326 ;
  assign n6328 = n6327 ^ x95 ;
  assign n6104 = n6052 & n6087 ;
  assign n6105 = n6104 ^ n5843 ;
  assign n6329 = n6328 ^ n6105 ;
  assign n6330 = n6328 ^ x96 ;
  assign n6331 = n6329 & n6330 ;
  assign n6332 = n6331 ^ x96 ;
  assign n6101 = n6054 ^ x96 ;
  assign n6102 = n6087 & n6101 ;
  assign n6103 = n6102 ^ n5840 ;
  assign n6333 = n6332 ^ n6103 ;
  assign n6334 = n6332 ^ x97 ;
  assign n6335 = n6333 & n6334 ;
  assign n6336 = n6335 ^ x97 ;
  assign n6337 = n6336 ^ x98 ;
  assign n6338 = n6057 ^ x97 ;
  assign n6339 = n6087 & n6338 ;
  assign n6340 = n6339 ^ n5837 ;
  assign n6341 = n6340 ^ n6336 ;
  assign n6342 = n6337 & n6341 ;
  assign n6100 = n6098 ^ x98 ;
  assign n6343 = n6342 ^ n6100 ;
  assign n6344 = ~n6099 & n6343 ;
  assign n6345 = n6344 ^ x99 ;
  assign n6095 = n6066 & n6087 ;
  assign n6096 = n6095 ^ n5832 ;
  assign n6346 = n6345 ^ n6096 ;
  assign n6347 = n6345 ^ x100 ;
  assign n6348 = n6346 & n6347 ;
  assign n6349 = n6348 ^ x100 ;
  assign n6350 = n6349 ^ x101 ;
  assign n6351 = n6070 & n6087 ;
  assign n6352 = n6351 ^ n5829 ;
  assign n6353 = n6352 ^ n6349 ;
  assign n6354 = n6350 & n6353 ;
  assign n6355 = n6354 ^ x101 ;
  assign n6357 = n6355 ^ x102 ;
  assign n6088 = n5812 & ~n6087 ;
  assign n6089 = n6088 ^ n270 ;
  assign n6365 = n6089 ^ x105 ;
  assign n6366 = n6080 ^ x103 ;
  assign n6367 = n6087 & n6366 ;
  assign n6368 = n6367 ^ n5819 ;
  assign n6093 = n6074 & n6087 ;
  assign n6094 = n6093 ^ n5827 ;
  assign n6356 = n6355 ^ n6094 ;
  assign n6358 = n6356 & n6357 ;
  assign n6359 = n6358 ^ x102 ;
  assign n6091 = n6078 & n6087 ;
  assign n6092 = n6091 ^ n5825 ;
  assign n6360 = n6359 ^ n6092 ;
  assign n6361 = n6359 ^ x103 ;
  assign n6362 = n6360 & n6361 ;
  assign n6363 = n6362 ^ x103 ;
  assign n6369 = n6368 ^ n6363 ;
  assign n6372 = n6368 ^ x104 ;
  assign n6373 = n6369 & ~n6372 ;
  assign n6370 = x105 ^ x104 ;
  assign n6374 = n6373 ^ n6370 ;
  assign n6377 = ~n6365 & n6374 ;
  assign n6378 = n6377 ^ x105 ;
  assign n6379 = n5814 & ~n6378 ;
  assign n6676 = n6357 & n6379 ;
  assign n6677 = n6676 ^ n6094 ;
  assign n6384 = n6350 & n6379 ;
  assign n6385 = n6384 ^ n6352 ;
  assign n6386 = n6385 ^ x102 ;
  assign n6390 = n6385 ^ x101 ;
  assign n6387 = n6347 & n6379 ;
  assign n6388 = n6387 ^ n6096 ;
  assign n6389 = n6388 ^ n6385 ;
  assign n6391 = n6390 ^ n6389 ;
  assign n6392 = n6342 ^ x99 ;
  assign n6393 = n6392 ^ x98 ;
  assign n6394 = n6379 & n6393 ;
  assign n6395 = n6394 ^ n6098 ;
  assign n6396 = n6395 ^ x100 ;
  assign n6400 = n6395 ^ x99 ;
  assign n6397 = n6337 & n6379 ;
  assign n6398 = n6397 ^ n6340 ;
  assign n6399 = n6398 ^ n6395 ;
  assign n6401 = n6400 ^ n6399 ;
  assign n6650 = n6326 & n6379 ;
  assign n6651 = n6650 ^ n6108 ;
  assign n6406 = n6322 & n6379 ;
  assign n6407 = n6406 ^ n6119 ;
  assign n6408 = n6407 ^ x95 ;
  assign n6412 = n6407 ^ x94 ;
  assign n6409 = n6318 & n6379 ;
  assign n6410 = n6409 ^ n6122 ;
  assign n6411 = n6410 ^ n6407 ;
  assign n6413 = n6412 ^ n6411 ;
  assign n6414 = n6314 & n6379 ;
  assign n6415 = n6414 ^ n6124 ;
  assign n6416 = n6415 ^ x93 ;
  assign n6420 = n6415 ^ x92 ;
  assign n6417 = n6310 & n6379 ;
  assign n6418 = n6417 ^ n6127 ;
  assign n6419 = n6418 ^ n6415 ;
  assign n6421 = n6420 ^ n6419 ;
  assign n6507 = x64 ^ x22 ;
  assign n6508 = n6206 ^ n191 ;
  assign n6509 = n6507 & n6508 ;
  assign n6510 = n6206 ^ x65 ;
  assign n6485 = ~x21 & x65 ;
  assign n6511 = n6485 ^ x65 ;
  assign n6512 = ~n6510 & ~n6511 ;
  assign n6513 = n6512 ^ x65 ;
  assign n6514 = n6509 & n6513 ;
  assign n6515 = n6379 & n6514 ;
  assign n6491 = x64 & n6379 ;
  assign n6492 = ~x21 & n6491 ;
  assign n6484 = ~x22 & x65 ;
  assign n6486 = n6485 ^ x21 ;
  assign n6487 = x22 & ~n6486 ;
  assign n6488 = n6487 ^ x21 ;
  assign n6489 = x64 & ~n6488 ;
  assign n6490 = ~n6484 & ~n6489 ;
  assign n6493 = n6492 ^ n6490 ;
  assign n6494 = n6206 & n6379 ;
  assign n6495 = n6494 ^ n6206 ;
  assign n6496 = n6495 ^ n6203 ;
  assign n6497 = n6496 ^ n6495 ;
  assign n6502 = ~x65 & n6494 ;
  assign n6503 = ~n6497 & n6502 ;
  assign n6504 = n6503 ^ n6497 ;
  assign n6505 = n6504 ^ n6496 ;
  assign n6506 = n6493 & n6505 ;
  assign n6516 = n6515 ^ n6506 ;
  assign n6532 = n6484 & ~n6491 ;
  assign n6517 = ~n6206 & n6489 ;
  assign n6518 = ~x66 & n6491 ;
  assign n6520 = n6488 ^ n6484 ;
  assign n6519 = x65 ^ x21 ;
  assign n6521 = n6520 ^ n6519 ;
  assign n6522 = ~n6510 & n6521 ;
  assign n6523 = n6518 & n6522 ;
  assign n6524 = n6523 ^ x66 ;
  assign n6525 = n6517 & ~n6524 ;
  assign n6530 = n6525 ^ n6524 ;
  assign n6526 = n6379 & n6525 ;
  assign n6527 = ~x22 & n6526 ;
  assign n6528 = n6485 & n6527 ;
  assign n6529 = n6528 ^ n6526 ;
  assign n6531 = n6530 ^ n6529 ;
  assign n6533 = n6379 ^ n6206 ;
  assign n6534 = ~n6531 & ~n6533 ;
  assign n6535 = n6532 & n6534 ;
  assign n6536 = n6535 ^ n6531 ;
  assign n6537 = ~n6516 & n6536 ;
  assign n6481 = n6209 ^ x66 ;
  assign n6482 = n6379 & n6481 ;
  assign n6483 = n6482 ^ n6201 ;
  assign n6538 = n6537 ^ n6483 ;
  assign n6539 = n6537 ^ x67 ;
  assign n6540 = n6538 & n6539 ;
  assign n6541 = n6540 ^ x67 ;
  assign n6479 = n6214 & n6379 ;
  assign n6480 = n6479 ^ n6198 ;
  assign n6542 = n6541 ^ n6480 ;
  assign n6543 = n6541 ^ x68 ;
  assign n6544 = n6542 & n6543 ;
  assign n6545 = n6544 ^ x68 ;
  assign n6477 = n6218 & n6379 ;
  assign n6478 = n6477 ^ n6195 ;
  assign n6546 = n6545 ^ n6478 ;
  assign n6547 = n6545 ^ x69 ;
  assign n6548 = n6546 & n6547 ;
  assign n6549 = n6548 ^ x69 ;
  assign n6475 = n6222 & n6379 ;
  assign n6476 = n6475 ^ n6193 ;
  assign n6550 = n6549 ^ n6476 ;
  assign n6551 = n6549 ^ x70 ;
  assign n6552 = n6550 & n6551 ;
  assign n6553 = n6552 ^ x70 ;
  assign n6473 = n6226 & n6379 ;
  assign n6474 = n6473 ^ n6191 ;
  assign n6554 = n6553 ^ n6474 ;
  assign n6555 = n6553 ^ x71 ;
  assign n6556 = n6554 & n6555 ;
  assign n6557 = n6556 ^ x71 ;
  assign n6470 = n6228 ^ x71 ;
  assign n6471 = n6379 & n6470 ;
  assign n6472 = n6471 ^ n6186 ;
  assign n6558 = n6557 ^ n6472 ;
  assign n6559 = n6557 ^ x72 ;
  assign n6560 = n6558 & n6559 ;
  assign n6561 = n6560 ^ x72 ;
  assign n6459 = n6186 ^ x72 ;
  assign n6460 = n6459 ^ n6228 ;
  assign n6461 = n6460 ^ x71 ;
  assign n6462 = n6461 ^ n6459 ;
  assign n6464 = n6228 ^ x72 ;
  assign n6465 = n6464 ^ n6459 ;
  assign n6466 = ~n6462 & ~n6465 ;
  assign n6467 = n6466 ^ n6459 ;
  assign n6468 = n6379 & ~n6467 ;
  assign n6469 = n6468 ^ n6183 ;
  assign n6562 = n6561 ^ n6469 ;
  assign n6563 = n6561 ^ x73 ;
  assign n6564 = n6562 & n6563 ;
  assign n6565 = n6564 ^ x73 ;
  assign n6456 = n6234 ^ x73 ;
  assign n6457 = n6379 & n6456 ;
  assign n6458 = n6457 ^ n6236 ;
  assign n6566 = n6565 ^ n6458 ;
  assign n6567 = n6565 ^ x74 ;
  assign n6568 = n6566 & n6567 ;
  assign n6569 = n6568 ^ x74 ;
  assign n6454 = n6242 & n6379 ;
  assign n6455 = n6454 ^ n6181 ;
  assign n6570 = n6569 ^ n6455 ;
  assign n6571 = n6569 ^ x75 ;
  assign n6572 = n6570 & n6571 ;
  assign n6573 = n6572 ^ x75 ;
  assign n6452 = n6246 & n6379 ;
  assign n6453 = n6452 ^ n6179 ;
  assign n6574 = n6573 ^ n6453 ;
  assign n6575 = n6573 ^ x76 ;
  assign n6576 = n6574 & n6575 ;
  assign n6577 = n6576 ^ x76 ;
  assign n6450 = n6250 & n6379 ;
  assign n6451 = n6450 ^ n6177 ;
  assign n6578 = n6577 ^ n6451 ;
  assign n6579 = n6577 ^ x77 ;
  assign n6580 = n6578 & n6579 ;
  assign n6581 = n6580 ^ x77 ;
  assign n6448 = n6254 & n6379 ;
  assign n6449 = n6448 ^ n6175 ;
  assign n6582 = n6581 ^ n6449 ;
  assign n6583 = n6581 ^ x78 ;
  assign n6584 = n6582 & n6583 ;
  assign n6585 = n6584 ^ x78 ;
  assign n6446 = n6258 & n6379 ;
  assign n6447 = n6446 ^ n6173 ;
  assign n6586 = n6585 ^ n6447 ;
  assign n6587 = n6585 ^ x79 ;
  assign n6588 = n6586 & n6587 ;
  assign n6589 = n6588 ^ x79 ;
  assign n6444 = n6262 & n6379 ;
  assign n6445 = n6444 ^ n6171 ;
  assign n6590 = n6589 ^ n6445 ;
  assign n6591 = n6589 ^ x80 ;
  assign n6592 = n6590 & n6591 ;
  assign n6593 = n6592 ^ x80 ;
  assign n6442 = n6266 & n6379 ;
  assign n6443 = n6442 ^ n6169 ;
  assign n6594 = n6593 ^ n6443 ;
  assign n6595 = n6593 ^ x81 ;
  assign n6596 = n6594 & n6595 ;
  assign n6597 = n6596 ^ x81 ;
  assign n6440 = n6270 & n6379 ;
  assign n6441 = n6440 ^ n6167 ;
  assign n6598 = n6597 ^ n6441 ;
  assign n6599 = n6597 ^ x82 ;
  assign n6600 = n6598 & n6599 ;
  assign n6601 = n6600 ^ x82 ;
  assign n6438 = n6274 & n6379 ;
  assign n6439 = n6438 ^ n6165 ;
  assign n6602 = n6601 ^ n6439 ;
  assign n6603 = n6601 ^ x83 ;
  assign n6604 = n6602 & n6603 ;
  assign n6605 = n6604 ^ x83 ;
  assign n6436 = n6278 & n6379 ;
  assign n6437 = n6436 ^ n6163 ;
  assign n6606 = n6605 ^ n6437 ;
  assign n6607 = n6605 ^ x84 ;
  assign n6608 = n6606 & n6607 ;
  assign n6609 = n6608 ^ x84 ;
  assign n6434 = n6282 & n6379 ;
  assign n6435 = n6434 ^ n6161 ;
  assign n6610 = n6609 ^ n6435 ;
  assign n6611 = n6609 ^ x85 ;
  assign n6612 = n6610 & n6611 ;
  assign n6613 = n6612 ^ x85 ;
  assign n6432 = n6286 & n6379 ;
  assign n6433 = n6432 ^ n6159 ;
  assign n6614 = n6613 ^ n6433 ;
  assign n6615 = n6613 ^ x86 ;
  assign n6616 = n6614 & n6615 ;
  assign n6617 = n6616 ^ x86 ;
  assign n6430 = n6290 & n6379 ;
  assign n6431 = n6430 ^ n6157 ;
  assign n6618 = n6617 ^ n6431 ;
  assign n6619 = n6617 ^ x87 ;
  assign n6620 = n6618 & n6619 ;
  assign n6621 = n6620 ^ x87 ;
  assign n6428 = n6294 & n6379 ;
  assign n6429 = n6428 ^ n6155 ;
  assign n6622 = n6621 ^ n6429 ;
  assign n6623 = n6621 ^ x88 ;
  assign n6624 = n6622 & n6623 ;
  assign n6625 = n6624 ^ x88 ;
  assign n6426 = n6298 & n6379 ;
  assign n6427 = n6426 ^ n6152 ;
  assign n6626 = n6625 ^ n6427 ;
  assign n6627 = n6625 ^ x89 ;
  assign n6628 = n6626 & n6627 ;
  assign n6629 = n6628 ^ x89 ;
  assign n6424 = n6302 & n6379 ;
  assign n6425 = n6424 ^ n6141 ;
  assign n6630 = n6629 ^ n6425 ;
  assign n6631 = n6629 ^ x90 ;
  assign n6632 = n6630 & n6631 ;
  assign n6633 = n6632 ^ x90 ;
  assign n6422 = n6306 & n6379 ;
  assign n6423 = n6422 ^ n6138 ;
  assign n6634 = n6633 ^ n6423 ;
  assign n6635 = n6633 ^ x91 ;
  assign n6636 = n6634 & n6635 ;
  assign n6637 = n6636 ^ x91 ;
  assign n6638 = n6637 ^ n6415 ;
  assign n6639 = n6638 ^ n6420 ;
  assign n6640 = ~n6421 & n6639 ;
  assign n6641 = n6640 ^ n6420 ;
  assign n6642 = ~n6416 & n6641 ;
  assign n6643 = n6642 ^ x93 ;
  assign n6644 = n6643 ^ n6407 ;
  assign n6645 = n6644 ^ n6412 ;
  assign n6646 = ~n6413 & n6645 ;
  assign n6647 = n6646 ^ n6412 ;
  assign n6648 = ~n6408 & n6647 ;
  assign n6649 = n6648 ^ x95 ;
  assign n6652 = n6651 ^ n6649 ;
  assign n6653 = n6651 ^ x96 ;
  assign n6654 = n6652 & ~n6653 ;
  assign n6655 = n6654 ^ x96 ;
  assign n6404 = n6330 & n6379 ;
  assign n6405 = n6404 ^ n6105 ;
  assign n6656 = n6655 ^ n6405 ;
  assign n6657 = n6655 ^ x97 ;
  assign n6658 = n6656 & n6657 ;
  assign n6659 = n6658 ^ x97 ;
  assign n6402 = n6334 & n6379 ;
  assign n6403 = n6402 ^ n6103 ;
  assign n6660 = n6659 ^ n6403 ;
  assign n6661 = n6659 ^ x98 ;
  assign n6662 = n6660 & n6661 ;
  assign n6663 = n6662 ^ x98 ;
  assign n6664 = n6663 ^ n6395 ;
  assign n6665 = n6664 ^ n6400 ;
  assign n6666 = ~n6401 & n6665 ;
  assign n6667 = n6666 ^ n6400 ;
  assign n6668 = ~n6396 & n6667 ;
  assign n6669 = n6668 ^ x100 ;
  assign n6670 = n6669 ^ n6385 ;
  assign n6671 = n6670 ^ n6390 ;
  assign n6672 = ~n6391 & n6671 ;
  assign n6673 = n6672 ^ n6390 ;
  assign n6674 = ~n6386 & n6673 ;
  assign n6675 = n6674 ^ x102 ;
  assign n6678 = n6677 ^ n6675 ;
  assign n6679 = n6677 ^ x103 ;
  assign n6680 = n6678 & ~n6679 ;
  assign n6681 = n6680 ^ x103 ;
  assign n6683 = n6681 ^ x104 ;
  assign n6090 = n6089 ^ x106 ;
  assign n6382 = n6361 & n6379 ;
  assign n6383 = n6382 ^ n6092 ;
  assign n6682 = n6681 ^ n6383 ;
  assign n6684 = n6682 & n6683 ;
  assign n6685 = n6684 ^ x104 ;
  assign n6364 = n6363 ^ x104 ;
  assign n6380 = n6364 & n6379 ;
  assign n6381 = n6380 ^ n6368 ;
  assign n6686 = n6685 ^ n6381 ;
  assign n6687 = n6685 ^ x105 ;
  assign n6688 = n6686 & n6687 ;
  assign n6689 = n6688 ^ x105 ;
  assign n6690 = n6689 ^ n6089 ;
  assign n6691 = n6090 & ~n6690 ;
  assign n6692 = ~x107 & n5813 ;
  assign n6693 = n6691 ^ n6689 ;
  assign n6694 = n6692 & ~n6693 ;
  assign n6695 = n6691 & n6694 ;
  assign n6696 = n6374 & n6695 ;
  assign n6697 = n6696 ^ n6694 ;
  assign n6997 = n6683 & n6697 ;
  assign n6998 = n6997 ^ n6383 ;
  assign n6999 = n6998 ^ x105 ;
  assign n6698 = n6388 ^ x102 ;
  assign n6699 = n6698 ^ x101 ;
  assign n6700 = n6699 ^ n6669 ;
  assign n6701 = n6700 ^ n6698 ;
  assign n6704 = n6698 ^ n5794 ;
  assign n6705 = ~n6701 & ~n6704 ;
  assign n6706 = n6705 ^ n6698 ;
  assign n6707 = n6697 & ~n6706 ;
  assign n6708 = n6707 ^ n6385 ;
  assign n6709 = n6708 ^ x103 ;
  assign n6710 = n6669 ^ x101 ;
  assign n6711 = n6697 & n6710 ;
  assign n6712 = n6711 ^ n6388 ;
  assign n6713 = n6712 ^ x102 ;
  assign n6979 = n6663 ^ x99 ;
  assign n6980 = n6697 & n6979 ;
  assign n6981 = n6980 ^ n6398 ;
  assign n6725 = n6661 & n6697 ;
  assign n6726 = n6725 ^ n6403 ;
  assign n6727 = n6726 ^ x99 ;
  assign n6731 = n6726 ^ x98 ;
  assign n6728 = n6657 & n6697 ;
  assign n6729 = n6728 ^ n6405 ;
  assign n6730 = n6729 ^ n6726 ;
  assign n6732 = n6731 ^ n6730 ;
  assign n6911 = n6599 & n6697 ;
  assign n6912 = n6911 ^ n6441 ;
  assign n6782 = n6595 & n6697 ;
  assign n6783 = n6782 ^ n6443 ;
  assign n6784 = n6783 ^ x82 ;
  assign n6788 = n6783 ^ x81 ;
  assign n6785 = n6591 & n6697 ;
  assign n6786 = n6785 ^ n6445 ;
  assign n6787 = n6786 ^ n6783 ;
  assign n6789 = n6788 ^ n6787 ;
  assign n6808 = n6551 & n6697 ;
  assign n6809 = n6808 ^ n6476 ;
  assign n6810 = n6809 ^ x71 ;
  assign n6811 = n6547 & n6697 ;
  assign n6812 = n6811 ^ n6478 ;
  assign n6813 = n6812 ^ x70 ;
  assign n6857 = n6543 & n6697 ;
  assign n6858 = n6857 ^ n6480 ;
  assign n6851 = n6539 & n6697 ;
  assign n6852 = n6851 ^ n6483 ;
  assign n6840 = x22 & x65 ;
  assign n6831 = n6507 ^ x65 ;
  assign n6832 = n6831 ^ n6379 ;
  assign n6833 = ~n6519 & n6832 ;
  assign n6841 = n6840 ^ n6833 ;
  assign n6842 = ~x64 & n6841 ;
  assign n6836 = x66 ^ x65 ;
  assign n6837 = n6836 ^ n6833 ;
  assign n6843 = n6842 ^ n6837 ;
  assign n6844 = n6697 & n6843 ;
  assign n6845 = n6844 ^ n6206 ;
  assign n6830 = n6204 & n6379 ;
  assign n6846 = n6845 ^ n6830 ;
  assign n6823 = n6491 ^ x22 ;
  assign n6815 = x64 & n6697 ;
  assign n6822 = ~x21 & n6815 ;
  assign n6824 = n6823 ^ n6822 ;
  assign n6821 = x65 & n6697 ;
  assign n6825 = n6824 ^ n6821 ;
  assign n6816 = n6815 ^ x21 ;
  assign n6814 = ~x20 & x64 ;
  assign n6817 = n6816 ^ n6814 ;
  assign n6818 = n6816 ^ x65 ;
  assign n6819 = n6817 & ~n6818 ;
  assign n6820 = n6819 ^ x65 ;
  assign n6826 = n6825 ^ n6820 ;
  assign n6827 = n6825 ^ x66 ;
  assign n6828 = n6826 & ~n6827 ;
  assign n6829 = n6828 ^ x66 ;
  assign n6847 = n6846 ^ n6829 ;
  assign n6848 = n6846 ^ x67 ;
  assign n6849 = n6847 & ~n6848 ;
  assign n6850 = n6849 ^ x67 ;
  assign n6853 = n6852 ^ n6850 ;
  assign n6854 = n6852 ^ x68 ;
  assign n6855 = n6853 & ~n6854 ;
  assign n6856 = n6855 ^ x68 ;
  assign n6859 = n6858 ^ n6856 ;
  assign n6860 = n6858 ^ x69 ;
  assign n6861 = n6859 & ~n6860 ;
  assign n6862 = n6861 ^ x69 ;
  assign n6863 = n6862 ^ n6812 ;
  assign n6864 = ~n6813 & n6863 ;
  assign n6865 = n6864 ^ x70 ;
  assign n6866 = n6865 ^ n6809 ;
  assign n6867 = ~n6810 & n6866 ;
  assign n6868 = n6867 ^ x71 ;
  assign n6806 = n6555 & n6697 ;
  assign n6807 = n6806 ^ n6474 ;
  assign n6869 = n6868 ^ n6807 ;
  assign n6870 = n6868 ^ x72 ;
  assign n6871 = n6869 & n6870 ;
  assign n6872 = n6871 ^ x72 ;
  assign n6804 = n6559 & n6697 ;
  assign n6805 = n6804 ^ n6472 ;
  assign n6873 = n6872 ^ n6805 ;
  assign n6874 = n6872 ^ x73 ;
  assign n6875 = n6873 & n6874 ;
  assign n6876 = n6875 ^ x73 ;
  assign n6802 = n6563 & n6697 ;
  assign n6803 = n6802 ^ n6469 ;
  assign n6877 = n6876 ^ n6803 ;
  assign n6878 = n6876 ^ x74 ;
  assign n6879 = n6877 & n6878 ;
  assign n6880 = n6879 ^ x74 ;
  assign n6800 = n6567 & n6697 ;
  assign n6801 = n6800 ^ n6458 ;
  assign n6881 = n6880 ^ n6801 ;
  assign n6882 = n6880 ^ x75 ;
  assign n6883 = n6881 & n6882 ;
  assign n6884 = n6883 ^ x75 ;
  assign n6798 = n6571 & n6697 ;
  assign n6799 = n6798 ^ n6455 ;
  assign n6885 = n6884 ^ n6799 ;
  assign n6886 = n6884 ^ x76 ;
  assign n6887 = n6885 & n6886 ;
  assign n6888 = n6887 ^ x76 ;
  assign n6796 = n6575 & n6697 ;
  assign n6797 = n6796 ^ n6453 ;
  assign n6889 = n6888 ^ n6797 ;
  assign n6890 = n6888 ^ x77 ;
  assign n6891 = n6889 & n6890 ;
  assign n6892 = n6891 ^ x77 ;
  assign n6794 = n6579 & n6697 ;
  assign n6795 = n6794 ^ n6451 ;
  assign n6893 = n6892 ^ n6795 ;
  assign n6894 = n6892 ^ x78 ;
  assign n6895 = n6893 & n6894 ;
  assign n6896 = n6895 ^ x78 ;
  assign n6792 = n6583 & n6697 ;
  assign n6793 = n6792 ^ n6449 ;
  assign n6897 = n6896 ^ n6793 ;
  assign n6898 = n6896 ^ x79 ;
  assign n6899 = n6897 & n6898 ;
  assign n6900 = n6899 ^ x79 ;
  assign n6790 = n6587 & n6697 ;
  assign n6791 = n6790 ^ n6447 ;
  assign n6901 = n6900 ^ n6791 ;
  assign n6902 = n6900 ^ x80 ;
  assign n6903 = n6901 & n6902 ;
  assign n6904 = n6903 ^ x80 ;
  assign n6905 = n6904 ^ n6783 ;
  assign n6906 = n6905 ^ n6788 ;
  assign n6907 = ~n6789 & n6906 ;
  assign n6908 = n6907 ^ n6788 ;
  assign n6909 = ~n6784 & n6908 ;
  assign n6910 = n6909 ^ x82 ;
  assign n6913 = n6912 ^ n6910 ;
  assign n6914 = n6912 ^ x83 ;
  assign n6915 = n6913 & ~n6914 ;
  assign n6916 = n6915 ^ x83 ;
  assign n6780 = n6603 & n6697 ;
  assign n6781 = n6780 ^ n6439 ;
  assign n6917 = n6916 ^ n6781 ;
  assign n6918 = n6916 ^ x84 ;
  assign n6919 = n6917 & n6918 ;
  assign n6920 = n6919 ^ x84 ;
  assign n6778 = n6607 & n6697 ;
  assign n6779 = n6778 ^ n6437 ;
  assign n6921 = n6920 ^ n6779 ;
  assign n6922 = n6920 ^ x85 ;
  assign n6923 = n6921 & n6922 ;
  assign n6924 = n6923 ^ x85 ;
  assign n6776 = n6611 & n6697 ;
  assign n6777 = n6776 ^ n6435 ;
  assign n6925 = n6924 ^ n6777 ;
  assign n6926 = n6924 ^ x86 ;
  assign n6927 = n6925 & n6926 ;
  assign n6928 = n6927 ^ x86 ;
  assign n6774 = n6615 & n6697 ;
  assign n6775 = n6774 ^ n6433 ;
  assign n6929 = n6928 ^ n6775 ;
  assign n6930 = n6928 ^ x87 ;
  assign n6931 = n6929 & n6930 ;
  assign n6932 = n6931 ^ x87 ;
  assign n6772 = n6619 & n6697 ;
  assign n6773 = n6772 ^ n6431 ;
  assign n6933 = n6932 ^ n6773 ;
  assign n6934 = n6932 ^ x88 ;
  assign n6935 = n6933 & n6934 ;
  assign n6936 = n6935 ^ x88 ;
  assign n6770 = n6623 & n6697 ;
  assign n6771 = n6770 ^ n6429 ;
  assign n6937 = n6936 ^ n6771 ;
  assign n6938 = n6936 ^ x89 ;
  assign n6939 = n6937 & n6938 ;
  assign n6940 = n6939 ^ x89 ;
  assign n6768 = n6627 & n6697 ;
  assign n6769 = n6768 ^ n6427 ;
  assign n6941 = n6940 ^ n6769 ;
  assign n6942 = n6940 ^ x90 ;
  assign n6943 = n6941 & n6942 ;
  assign n6944 = n6943 ^ x90 ;
  assign n6766 = n6631 & n6697 ;
  assign n6767 = n6766 ^ n6425 ;
  assign n6945 = n6944 ^ n6767 ;
  assign n6946 = n6944 ^ x91 ;
  assign n6947 = n6945 & n6946 ;
  assign n6948 = n6947 ^ x91 ;
  assign n6764 = n6635 & n6697 ;
  assign n6765 = n6764 ^ n6423 ;
  assign n6949 = n6948 ^ n6765 ;
  assign n6950 = n6948 ^ x92 ;
  assign n6951 = n6949 & n6950 ;
  assign n6952 = n6951 ^ x92 ;
  assign n6761 = n6637 ^ x92 ;
  assign n6762 = n6697 & n6761 ;
  assign n6763 = n6762 ^ n6418 ;
  assign n6953 = n6952 ^ n6763 ;
  assign n6954 = n6952 ^ x93 ;
  assign n6955 = n6953 & n6954 ;
  assign n6956 = n6955 ^ x93 ;
  assign n6750 = n6418 ^ x93 ;
  assign n6751 = n6750 ^ n6637 ;
  assign n6752 = n6751 ^ x92 ;
  assign n6753 = n6752 ^ n6750 ;
  assign n6755 = n6637 ^ x93 ;
  assign n6756 = n6755 ^ n6750 ;
  assign n6757 = ~n6753 & ~n6756 ;
  assign n6758 = n6757 ^ n6750 ;
  assign n6759 = n6697 & ~n6758 ;
  assign n6760 = n6759 ^ n6415 ;
  assign n6957 = n6956 ^ n6760 ;
  assign n6958 = n6956 ^ x94 ;
  assign n6959 = n6957 & n6958 ;
  assign n6960 = n6959 ^ x94 ;
  assign n6747 = n6643 ^ x94 ;
  assign n6748 = n6697 & n6747 ;
  assign n6749 = n6748 ^ n6410 ;
  assign n6961 = n6960 ^ n6749 ;
  assign n6962 = n6960 ^ x95 ;
  assign n6963 = n6961 & n6962 ;
  assign n6964 = n6963 ^ x95 ;
  assign n6736 = n6410 ^ x95 ;
  assign n6737 = n6736 ^ x94 ;
  assign n6738 = n6737 ^ n6643 ;
  assign n6739 = n6738 ^ n6736 ;
  assign n6741 = x95 ^ x94 ;
  assign n6742 = n6741 ^ n6736 ;
  assign n6743 = ~n6739 & ~n6742 ;
  assign n6744 = n6743 ^ n6736 ;
  assign n6745 = n6697 & ~n6744 ;
  assign n6746 = n6745 ^ n6407 ;
  assign n6965 = n6964 ^ n6746 ;
  assign n6966 = n6964 ^ x96 ;
  assign n6967 = n6965 & n6966 ;
  assign n6968 = n6967 ^ x96 ;
  assign n6733 = n6649 ^ x96 ;
  assign n6734 = n6697 & n6733 ;
  assign n6735 = n6734 ^ n6651 ;
  assign n6969 = n6968 ^ n6735 ;
  assign n6970 = n6968 ^ x97 ;
  assign n6971 = n6969 & n6970 ;
  assign n6972 = n6971 ^ x97 ;
  assign n6973 = n6972 ^ n6726 ;
  assign n6974 = n6973 ^ n6731 ;
  assign n6975 = ~n6732 & n6974 ;
  assign n6976 = n6975 ^ n6731 ;
  assign n6977 = ~n6727 & n6976 ;
  assign n6978 = n6977 ^ x99 ;
  assign n6982 = n6981 ^ n6978 ;
  assign n6983 = n6981 ^ x100 ;
  assign n6984 = n6982 & ~n6983 ;
  assign n6985 = n6984 ^ x100 ;
  assign n6714 = n6398 ^ x100 ;
  assign n6715 = n6714 ^ n6663 ;
  assign n6716 = n6715 ^ x99 ;
  assign n6717 = n6716 ^ n6714 ;
  assign n6719 = n6663 ^ x100 ;
  assign n6720 = n6719 ^ n6714 ;
  assign n6721 = ~n6717 & ~n6720 ;
  assign n6722 = n6721 ^ n6714 ;
  assign n6723 = n6697 & ~n6722 ;
  assign n6724 = n6723 ^ n6395 ;
  assign n6986 = n6985 ^ n6724 ;
  assign n6987 = n6985 ^ x101 ;
  assign n6988 = n6986 & n6987 ;
  assign n6989 = n6988 ^ x101 ;
  assign n6990 = n6989 ^ n6712 ;
  assign n6991 = ~n6713 & n6990 ;
  assign n6992 = n6991 ^ x102 ;
  assign n6993 = n6992 ^ n6708 ;
  assign n6994 = ~n6709 & n6993 ;
  assign n6995 = n6994 ^ x103 ;
  assign n6996 = n6995 ^ x104 ;
  assign n7000 = n6675 ^ x103 ;
  assign n7001 = n6697 & n7000 ;
  assign n7002 = n7001 ^ n6677 ;
  assign n7003 = n7002 ^ n6995 ;
  assign n7004 = n6996 & n7003 ;
  assign n7005 = n7004 ^ x104 ;
  assign n7006 = n7005 ^ n6998 ;
  assign n7007 = ~n6999 & n7006 ;
  assign n7008 = n7007 ^ x105 ;
  assign n7009 = n7008 ^ x106 ;
  assign n7010 = n6687 & n6697 ;
  assign n7011 = n7010 ^ n6381 ;
  assign n7012 = n7011 ^ n7008 ;
  assign n7013 = n7009 & n7012 ;
  assign n7014 = n7013 ^ x106 ;
  assign n7015 = n7014 ^ n6089 ;
  assign n7017 = n6689 ^ x106 ;
  assign n7018 = n6692 & ~n7017 ;
  assign n7019 = ~x106 & n7018 ;
  assign n7020 = n6374 & n7019 ;
  assign n7021 = n7020 ^ n7018 ;
  assign n7022 = n7021 ^ n6692 ;
  assign n7023 = n6089 & ~n7022 ;
  assign n7016 = n6089 ^ x107 ;
  assign n7024 = n7023 ^ n7016 ;
  assign n7025 = n7024 ^ n6089 ;
  assign n7026 = ~n7015 & ~n7025 ;
  assign n7027 = n7026 ^ n6089 ;
  assign n7028 = n5813 & n7027 ;
  assign n7334 = n7009 & n7028 ;
  assign n7335 = n7334 ^ n7011 ;
  assign n7336 = ~x107 & n7335 ;
  assign n7337 = n7335 ^ x107 ;
  assign n7338 = n7337 ^ n7336 ;
  assign n7149 = ~x19 & x65 ;
  assign n7150 = n6814 & ~n7149 ;
  assign n7151 = x64 & n7028 ;
  assign n7152 = ~n6818 & n7151 ;
  assign n7153 = n7150 & n7152 ;
  assign n7146 = x20 & ~x21 ;
  assign n7147 = n911 & n7028 ;
  assign n7148 = n7146 & n7147 ;
  assign n7154 = n7153 ^ n7148 ;
  assign n7137 = ~x20 & x65 ;
  assign n7138 = n6816 & ~n7137 ;
  assign n7140 = n6814 ^ x65 ;
  assign n7139 = ~x19 & x64 ;
  assign n7141 = n7140 ^ n7139 ;
  assign n7142 = n7140 ^ n7028 ;
  assign n7143 = n7141 & n7142 ;
  assign n7144 = n7143 ^ n7140 ;
  assign n7145 = n7138 & ~n7144 ;
  assign n7155 = n7154 ^ n7145 ;
  assign n7156 = n6816 ^ x19 ;
  assign n7157 = n7156 ^ x65 ;
  assign n7158 = n7157 ^ x20 ;
  assign n7159 = n7158 ^ n7028 ;
  assign n7160 = ~x19 & ~n7159 ;
  assign n7161 = n7160 ^ n7156 ;
  assign n7162 = n7028 ^ x20 ;
  assign n7163 = n7156 ^ n7028 ;
  assign n7164 = n7163 ^ x19 ;
  assign n7165 = ~n7162 & ~n7164 ;
  assign n7166 = n7165 ^ n7156 ;
  assign n7167 = ~n7161 & ~n7166 ;
  assign n7168 = n7167 ^ n7156 ;
  assign n7169 = x64 & ~n7168 ;
  assign n7170 = ~x66 & n7137 ;
  assign n7171 = n7028 ^ n6816 ;
  assign n7172 = ~n7151 & ~n7171 ;
  assign n7173 = n7170 & n7172 ;
  assign n7174 = n7173 ^ x66 ;
  assign n7175 = ~n7169 & ~n7174 ;
  assign n7176 = ~n7155 & ~n7175 ;
  assign n7134 = n6820 ^ x66 ;
  assign n7135 = n7028 & n7134 ;
  assign n7136 = n7135 ^ n6825 ;
  assign n7177 = n7176 ^ n7136 ;
  assign n7178 = n7176 ^ x67 ;
  assign n7179 = n7177 & n7178 ;
  assign n7180 = n7179 ^ x67 ;
  assign n7131 = n6829 ^ x67 ;
  assign n7132 = n7028 & n7131 ;
  assign n7133 = n7132 ^ n6846 ;
  assign n7181 = n7180 ^ n7133 ;
  assign n7182 = n7180 ^ x68 ;
  assign n7183 = n7181 & n7182 ;
  assign n7184 = n7183 ^ x68 ;
  assign n7128 = n6850 ^ x68 ;
  assign n7129 = n7028 & n7128 ;
  assign n7130 = n7129 ^ n6852 ;
  assign n7185 = n7184 ^ n7130 ;
  assign n7186 = n7184 ^ x69 ;
  assign n7187 = n7185 & n7186 ;
  assign n7188 = n7187 ^ x69 ;
  assign n7125 = n6856 ^ x69 ;
  assign n7126 = n7028 & n7125 ;
  assign n7127 = n7126 ^ n6858 ;
  assign n7189 = n7188 ^ n7127 ;
  assign n7190 = n7188 ^ x70 ;
  assign n7191 = n7189 & n7190 ;
  assign n7192 = n7191 ^ x70 ;
  assign n7122 = n6862 ^ x70 ;
  assign n7123 = n7028 & n7122 ;
  assign n7124 = n7123 ^ n6812 ;
  assign n7193 = n7192 ^ n7124 ;
  assign n7194 = n7192 ^ x71 ;
  assign n7195 = n7193 & n7194 ;
  assign n7196 = n7195 ^ x71 ;
  assign n7119 = n6865 ^ x71 ;
  assign n7120 = n7028 & n7119 ;
  assign n7121 = n7120 ^ n6809 ;
  assign n7197 = n7196 ^ n7121 ;
  assign n7198 = n7196 ^ x72 ;
  assign n7199 = n7197 & n7198 ;
  assign n7200 = n7199 ^ x72 ;
  assign n7117 = n6870 & n7028 ;
  assign n7118 = n7117 ^ n6807 ;
  assign n7201 = n7200 ^ n7118 ;
  assign n7202 = n7200 ^ x73 ;
  assign n7203 = n7201 & n7202 ;
  assign n7204 = n7203 ^ x73 ;
  assign n7115 = n6874 & n7028 ;
  assign n7116 = n7115 ^ n6805 ;
  assign n7205 = n7204 ^ n7116 ;
  assign n7206 = n7204 ^ x74 ;
  assign n7207 = n7205 & n7206 ;
  assign n7208 = n7207 ^ x74 ;
  assign n7113 = n6878 & n7028 ;
  assign n7114 = n7113 ^ n6803 ;
  assign n7209 = n7208 ^ n7114 ;
  assign n7210 = n7208 ^ x75 ;
  assign n7211 = n7209 & n7210 ;
  assign n7212 = n7211 ^ x75 ;
  assign n7111 = n6882 & n7028 ;
  assign n7112 = n7111 ^ n6801 ;
  assign n7213 = n7212 ^ n7112 ;
  assign n7214 = n7212 ^ x76 ;
  assign n7215 = n7213 & n7214 ;
  assign n7216 = n7215 ^ x76 ;
  assign n7109 = n6886 & n7028 ;
  assign n7110 = n7109 ^ n6799 ;
  assign n7217 = n7216 ^ n7110 ;
  assign n7218 = n7216 ^ x77 ;
  assign n7219 = n7217 & n7218 ;
  assign n7220 = n7219 ^ x77 ;
  assign n7107 = n6890 & n7028 ;
  assign n7108 = n7107 ^ n6797 ;
  assign n7221 = n7220 ^ n7108 ;
  assign n7222 = n7220 ^ x78 ;
  assign n7223 = n7221 & n7222 ;
  assign n7224 = n7223 ^ x78 ;
  assign n7105 = n6894 & n7028 ;
  assign n7106 = n7105 ^ n6795 ;
  assign n7225 = n7224 ^ n7106 ;
  assign n7226 = n7224 ^ x79 ;
  assign n7227 = n7225 & n7226 ;
  assign n7228 = n7227 ^ x79 ;
  assign n7103 = n6898 & n7028 ;
  assign n7104 = n7103 ^ n6793 ;
  assign n7229 = n7228 ^ n7104 ;
  assign n7230 = n7228 ^ x80 ;
  assign n7231 = n7229 & n7230 ;
  assign n7232 = n7231 ^ x80 ;
  assign n7101 = n6902 & n7028 ;
  assign n7102 = n7101 ^ n6791 ;
  assign n7233 = n7232 ^ n7102 ;
  assign n7234 = n7232 ^ x81 ;
  assign n7235 = n7233 & n7234 ;
  assign n7236 = n7235 ^ x81 ;
  assign n7098 = n6904 ^ x81 ;
  assign n7099 = n7028 & n7098 ;
  assign n7100 = n7099 ^ n6786 ;
  assign n7237 = n7236 ^ n7100 ;
  assign n7238 = n7236 ^ x82 ;
  assign n7239 = n7237 & n7238 ;
  assign n7240 = n7239 ^ x82 ;
  assign n7087 = n6786 ^ x82 ;
  assign n7088 = n7087 ^ n6904 ;
  assign n7089 = n7088 ^ x81 ;
  assign n7090 = n7089 ^ n7087 ;
  assign n7092 = n6904 ^ x82 ;
  assign n7093 = n7092 ^ n7087 ;
  assign n7094 = ~n7090 & ~n7093 ;
  assign n7095 = n7094 ^ n7087 ;
  assign n7096 = n7028 & ~n7095 ;
  assign n7097 = n7096 ^ n6783 ;
  assign n7241 = n7240 ^ n7097 ;
  assign n7242 = n7240 ^ x83 ;
  assign n7243 = n7241 & n7242 ;
  assign n7244 = n7243 ^ x83 ;
  assign n7084 = n6910 ^ x83 ;
  assign n7085 = n7028 & n7084 ;
  assign n7086 = n7085 ^ n6912 ;
  assign n7245 = n7244 ^ n7086 ;
  assign n7246 = n7244 ^ x84 ;
  assign n7247 = n7245 & n7246 ;
  assign n7248 = n7247 ^ x84 ;
  assign n7082 = n6918 & n7028 ;
  assign n7083 = n7082 ^ n6781 ;
  assign n7249 = n7248 ^ n7083 ;
  assign n7250 = n7248 ^ x85 ;
  assign n7251 = n7249 & n7250 ;
  assign n7252 = n7251 ^ x85 ;
  assign n7080 = n6922 & n7028 ;
  assign n7081 = n7080 ^ n6779 ;
  assign n7253 = n7252 ^ n7081 ;
  assign n7254 = n7252 ^ x86 ;
  assign n7255 = n7253 & n7254 ;
  assign n7256 = n7255 ^ x86 ;
  assign n7078 = n6926 & n7028 ;
  assign n7079 = n7078 ^ n6777 ;
  assign n7257 = n7256 ^ n7079 ;
  assign n7258 = n7256 ^ x87 ;
  assign n7259 = n7257 & n7258 ;
  assign n7260 = n7259 ^ x87 ;
  assign n7076 = n6930 & n7028 ;
  assign n7077 = n7076 ^ n6775 ;
  assign n7261 = n7260 ^ n7077 ;
  assign n7262 = n7260 ^ x88 ;
  assign n7263 = n7261 & n7262 ;
  assign n7264 = n7263 ^ x88 ;
  assign n7074 = n6934 & n7028 ;
  assign n7075 = n7074 ^ n6773 ;
  assign n7265 = n7264 ^ n7075 ;
  assign n7266 = n7264 ^ x89 ;
  assign n7267 = n7265 & n7266 ;
  assign n7268 = n7267 ^ x89 ;
  assign n7072 = n6938 & n7028 ;
  assign n7073 = n7072 ^ n6771 ;
  assign n7269 = n7268 ^ n7073 ;
  assign n7270 = n7268 ^ x90 ;
  assign n7271 = n7269 & n7270 ;
  assign n7272 = n7271 ^ x90 ;
  assign n7070 = n6942 & n7028 ;
  assign n7071 = n7070 ^ n6769 ;
  assign n7273 = n7272 ^ n7071 ;
  assign n7274 = n7272 ^ x91 ;
  assign n7275 = n7273 & n7274 ;
  assign n7276 = n7275 ^ x91 ;
  assign n7068 = n6946 & n7028 ;
  assign n7069 = n7068 ^ n6767 ;
  assign n7277 = n7276 ^ n7069 ;
  assign n7278 = n7276 ^ x92 ;
  assign n7279 = n7277 & n7278 ;
  assign n7280 = n7279 ^ x92 ;
  assign n7066 = n6950 & n7028 ;
  assign n7067 = n7066 ^ n6765 ;
  assign n7281 = n7280 ^ n7067 ;
  assign n7282 = n7280 ^ x93 ;
  assign n7283 = n7281 & n7282 ;
  assign n7284 = n7283 ^ x93 ;
  assign n7064 = n6954 & n7028 ;
  assign n7065 = n7064 ^ n6763 ;
  assign n7285 = n7284 ^ n7065 ;
  assign n7286 = n7284 ^ x94 ;
  assign n7287 = n7285 & n7286 ;
  assign n7288 = n7287 ^ x94 ;
  assign n7062 = n6958 & n7028 ;
  assign n7063 = n7062 ^ n6760 ;
  assign n7289 = n7288 ^ n7063 ;
  assign n7290 = n7288 ^ x95 ;
  assign n7291 = n7289 & n7290 ;
  assign n7292 = n7291 ^ x95 ;
  assign n7060 = n6962 & n7028 ;
  assign n7061 = n7060 ^ n6749 ;
  assign n7293 = n7292 ^ n7061 ;
  assign n7294 = n7292 ^ x96 ;
  assign n7295 = n7293 & n7294 ;
  assign n7296 = n7295 ^ x96 ;
  assign n7058 = n6966 & n7028 ;
  assign n7059 = n7058 ^ n6746 ;
  assign n7297 = n7296 ^ n7059 ;
  assign n7298 = n7296 ^ x97 ;
  assign n7299 = n7297 & n7298 ;
  assign n7300 = n7299 ^ x97 ;
  assign n7056 = n6970 & n7028 ;
  assign n7057 = n7056 ^ n6735 ;
  assign n7301 = n7300 ^ n7057 ;
  assign n7302 = n7300 ^ x98 ;
  assign n7303 = n7301 & n7302 ;
  assign n7304 = n7303 ^ x98 ;
  assign n7053 = n6972 ^ x98 ;
  assign n7054 = n7028 & n7053 ;
  assign n7055 = n7054 ^ n6729 ;
  assign n7305 = n7304 ^ n7055 ;
  assign n7306 = n7304 ^ x99 ;
  assign n7307 = n7305 & n7306 ;
  assign n7308 = n7307 ^ x99 ;
  assign n7042 = n6729 ^ x99 ;
  assign n7043 = n7042 ^ n6972 ;
  assign n7044 = n7043 ^ x98 ;
  assign n7045 = n7044 ^ n7042 ;
  assign n7047 = n6972 ^ x99 ;
  assign n7048 = n7047 ^ n7042 ;
  assign n7049 = ~n7045 & ~n7048 ;
  assign n7050 = n7049 ^ n7042 ;
  assign n7051 = n7028 & ~n7050 ;
  assign n7052 = n7051 ^ n6726 ;
  assign n7309 = n7308 ^ n7052 ;
  assign n7310 = n7308 ^ x100 ;
  assign n7311 = n7309 & n7310 ;
  assign n7312 = n7311 ^ x100 ;
  assign n7039 = n6978 ^ x100 ;
  assign n7040 = n7028 & n7039 ;
  assign n7041 = n7040 ^ n6981 ;
  assign n7313 = n7312 ^ n7041 ;
  assign n7314 = n7312 ^ x101 ;
  assign n7315 = n7313 & n7314 ;
  assign n7316 = n7315 ^ x101 ;
  assign n7037 = n6987 & n7028 ;
  assign n7038 = n7037 ^ n6724 ;
  assign n7317 = n7316 ^ n7038 ;
  assign n7318 = n7316 ^ x102 ;
  assign n7319 = n7317 & n7318 ;
  assign n7320 = n7319 ^ x102 ;
  assign n7034 = n6989 ^ x102 ;
  assign n7035 = n7028 & n7034 ;
  assign n7036 = n7035 ^ n6712 ;
  assign n7321 = n7320 ^ n7036 ;
  assign n7322 = n7320 ^ x103 ;
  assign n7323 = n7321 & n7322 ;
  assign n7324 = n7323 ^ x103 ;
  assign n7031 = n6992 ^ x103 ;
  assign n7032 = n7028 & n7031 ;
  assign n7033 = n7032 ^ n6708 ;
  assign n7325 = n7324 ^ n7033 ;
  assign n7326 = n7324 ^ x104 ;
  assign n7327 = n7325 & n7326 ;
  assign n7328 = n7327 ^ x104 ;
  assign n7029 = n6996 & n7028 ;
  assign n7030 = n7029 ^ n7002 ;
  assign n7329 = n7328 ^ n7030 ;
  assign n7330 = n7328 ^ x105 ;
  assign n7331 = n7329 & n7330 ;
  assign n7332 = n7331 ^ x105 ;
  assign n7333 = n7332 ^ x106 ;
  assign n7339 = n7005 ^ x105 ;
  assign n7340 = n7028 & n7339 ;
  assign n7341 = n7340 ^ n6998 ;
  assign n7342 = n7341 ^ n7332 ;
  assign n7343 = n7333 & n7342 ;
  assign n7344 = n7343 ^ x106 ;
  assign n7345 = ~n7338 & ~n7344 ;
  assign n7346 = ~n7336 & ~n7345 ;
  assign n7347 = n5813 & ~n7346 ;
  assign n7348 = n148 & n6089 ;
  assign n7349 = n7336 ^ n7022 ;
  assign n7350 = n7349 ^ n7336 ;
  assign n7351 = n7014 ^ x107 ;
  assign n7352 = ~x108 & ~n7351 ;
  assign n7355 = ~n7350 & n7352 ;
  assign n7356 = n7355 ^ n7336 ;
  assign n7357 = ~n7345 & ~n7356 ;
  assign n7358 = n7348 & ~n7357 ;
  assign n7359 = n7347 & ~n7358 ;
  assign n7360 = n7359 ^ n7358 ;
  assign n7666 = n7344 ^ x107 ;
  assign n7667 = n7360 & n7666 ;
  assign n7668 = n7667 ^ n7335 ;
  assign n7361 = n7333 & n7360 ;
  assign n7362 = n7361 ^ n7341 ;
  assign n7363 = n7362 ^ x107 ;
  assign n7367 = n7362 ^ x106 ;
  assign n7364 = n7330 & n7360 ;
  assign n7365 = n7364 ^ n7030 ;
  assign n7366 = n7365 ^ n7362 ;
  assign n7368 = n7367 ^ n7366 ;
  assign n7638 = n7310 & n7360 ;
  assign n7639 = n7638 ^ n7052 ;
  assign n7377 = n7306 & n7360 ;
  assign n7378 = n7377 ^ n7055 ;
  assign n7379 = n7378 ^ x100 ;
  assign n7383 = n7378 ^ x99 ;
  assign n7380 = n7302 & n7360 ;
  assign n7381 = n7380 ^ n7057 ;
  assign n7382 = n7381 ^ n7378 ;
  assign n7384 = n7383 ^ n7382 ;
  assign n7385 = n7298 & n7360 ;
  assign n7386 = n7385 ^ n7059 ;
  assign n7387 = n7386 ^ x98 ;
  assign n7391 = n7386 ^ x97 ;
  assign n7388 = n7294 & n7360 ;
  assign n7389 = n7388 ^ n7061 ;
  assign n7390 = n7389 ^ n7386 ;
  assign n7392 = n7391 ^ n7390 ;
  assign n7564 = n7234 & n7360 ;
  assign n7565 = n7564 ^ n7102 ;
  assign n7421 = n7230 & n7360 ;
  assign n7422 = n7421 ^ n7104 ;
  assign n7423 = n7422 ^ x81 ;
  assign n7427 = n7422 ^ x80 ;
  assign n7424 = n7226 & n7360 ;
  assign n7425 = n7424 ^ n7106 ;
  assign n7426 = n7425 ^ n7422 ;
  assign n7428 = n7427 ^ n7426 ;
  assign n7455 = n7151 ^ x20 ;
  assign n7453 = n7139 ^ x65 ;
  assign n7454 = n7360 & n7453 ;
  assign n7456 = n7455 ^ n7454 ;
  assign n7457 = n7456 ^ x66 ;
  assign n7458 = x64 & n7360 ;
  assign n7460 = x65 ^ x19 ;
  assign n7459 = n7149 ^ x19 ;
  assign n7461 = n7460 ^ n7459 ;
  assign n7462 = n7461 ^ x19 ;
  assign n7465 = x18 & n7462 ;
  assign n7466 = n7465 ^ x19 ;
  assign n7467 = n7458 & n7466 ;
  assign n7468 = x65 ^ x18 ;
  assign n7469 = n7468 ^ n7460 ;
  assign n7470 = n7469 ^ x65 ;
  assign n7477 = x64 & n7470 ;
  assign n7472 = n7460 ^ n191 ;
  assign n7478 = n7477 ^ n7472 ;
  assign n7481 = n7477 ^ x64 ;
  assign n7482 = ~n7360 & n7481 ;
  assign n7483 = n7482 ^ x65 ;
  assign n7484 = n7478 & n7483 ;
  assign n7485 = n7484 ^ x65 ;
  assign n7486 = ~n7467 & ~n7485 ;
  assign n7487 = n7486 ^ n7456 ;
  assign n7488 = ~n7457 & ~n7487 ;
  assign n7489 = n7488 ^ x66 ;
  assign n7490 = n7489 ^ x67 ;
  assign n7500 = x20 & x65 ;
  assign n7492 = n191 ^ x20 ;
  assign n7493 = n7492 ^ n7028 ;
  assign n7494 = ~n7460 & n7493 ;
  assign n7501 = n7500 ^ n7494 ;
  assign n7502 = ~x64 & n7501 ;
  assign n7497 = n7494 ^ n6836 ;
  assign n7503 = n7502 ^ n7497 ;
  assign n7504 = n7360 & n7503 ;
  assign n7505 = n7504 ^ n6816 ;
  assign n7491 = n7028 & n7140 ;
  assign n7506 = n7505 ^ n7491 ;
  assign n7507 = n7506 ^ n7489 ;
  assign n7508 = n7490 & n7507 ;
  assign n7509 = n7508 ^ x67 ;
  assign n7451 = n7178 & n7360 ;
  assign n7452 = n7451 ^ n7136 ;
  assign n7510 = n7509 ^ n7452 ;
  assign n7511 = n7509 ^ x68 ;
  assign n7512 = n7510 & n7511 ;
  assign n7513 = n7512 ^ x68 ;
  assign n7449 = n7182 & n7360 ;
  assign n7450 = n7449 ^ n7133 ;
  assign n7514 = n7513 ^ n7450 ;
  assign n7515 = n7513 ^ x69 ;
  assign n7516 = n7514 & n7515 ;
  assign n7517 = n7516 ^ x69 ;
  assign n7447 = n7186 & n7360 ;
  assign n7448 = n7447 ^ n7130 ;
  assign n7518 = n7517 ^ n7448 ;
  assign n7519 = n7517 ^ x70 ;
  assign n7520 = n7518 & n7519 ;
  assign n7521 = n7520 ^ x70 ;
  assign n7445 = n7190 & n7360 ;
  assign n7446 = n7445 ^ n7127 ;
  assign n7522 = n7521 ^ n7446 ;
  assign n7523 = n7521 ^ x71 ;
  assign n7524 = n7522 & n7523 ;
  assign n7525 = n7524 ^ x71 ;
  assign n7443 = n7194 & n7360 ;
  assign n7444 = n7443 ^ n7124 ;
  assign n7526 = n7525 ^ n7444 ;
  assign n7527 = n7525 ^ x72 ;
  assign n7528 = n7526 & n7527 ;
  assign n7529 = n7528 ^ x72 ;
  assign n7441 = n7198 & n7360 ;
  assign n7442 = n7441 ^ n7121 ;
  assign n7530 = n7529 ^ n7442 ;
  assign n7531 = n7529 ^ x73 ;
  assign n7532 = n7530 & n7531 ;
  assign n7533 = n7532 ^ x73 ;
  assign n7439 = n7202 & n7360 ;
  assign n7440 = n7439 ^ n7118 ;
  assign n7534 = n7533 ^ n7440 ;
  assign n7535 = n7533 ^ x74 ;
  assign n7536 = n7534 & n7535 ;
  assign n7537 = n7536 ^ x74 ;
  assign n7437 = n7206 & n7360 ;
  assign n7438 = n7437 ^ n7116 ;
  assign n7538 = n7537 ^ n7438 ;
  assign n7539 = n7537 ^ x75 ;
  assign n7540 = n7538 & n7539 ;
  assign n7541 = n7540 ^ x75 ;
  assign n7435 = n7210 & n7360 ;
  assign n7436 = n7435 ^ n7114 ;
  assign n7542 = n7541 ^ n7436 ;
  assign n7543 = n7541 ^ x76 ;
  assign n7544 = n7542 & n7543 ;
  assign n7545 = n7544 ^ x76 ;
  assign n7433 = n7214 & n7360 ;
  assign n7434 = n7433 ^ n7112 ;
  assign n7546 = n7545 ^ n7434 ;
  assign n7547 = n7545 ^ x77 ;
  assign n7548 = n7546 & n7547 ;
  assign n7549 = n7548 ^ x77 ;
  assign n7431 = n7218 & n7360 ;
  assign n7432 = n7431 ^ n7110 ;
  assign n7550 = n7549 ^ n7432 ;
  assign n7551 = n7549 ^ x78 ;
  assign n7552 = n7550 & n7551 ;
  assign n7553 = n7552 ^ x78 ;
  assign n7429 = n7222 & n7360 ;
  assign n7430 = n7429 ^ n7108 ;
  assign n7554 = n7553 ^ n7430 ;
  assign n7555 = n7553 ^ x79 ;
  assign n7556 = n7554 & n7555 ;
  assign n7557 = n7556 ^ x79 ;
  assign n7558 = n7557 ^ n7422 ;
  assign n7559 = n7558 ^ n7427 ;
  assign n7560 = ~n7428 & n7559 ;
  assign n7561 = n7560 ^ n7427 ;
  assign n7562 = ~n7423 & n7561 ;
  assign n7563 = n7562 ^ x81 ;
  assign n7566 = n7565 ^ n7563 ;
  assign n7567 = n7565 ^ x82 ;
  assign n7568 = n7566 & ~n7567 ;
  assign n7569 = n7568 ^ x82 ;
  assign n7419 = n7238 & n7360 ;
  assign n7420 = n7419 ^ n7100 ;
  assign n7570 = n7569 ^ n7420 ;
  assign n7571 = n7569 ^ x83 ;
  assign n7572 = n7570 & n7571 ;
  assign n7573 = n7572 ^ x83 ;
  assign n7417 = n7242 & n7360 ;
  assign n7418 = n7417 ^ n7097 ;
  assign n7574 = n7573 ^ n7418 ;
  assign n7575 = n7573 ^ x84 ;
  assign n7576 = n7574 & n7575 ;
  assign n7577 = n7576 ^ x84 ;
  assign n7415 = n7246 & n7360 ;
  assign n7416 = n7415 ^ n7086 ;
  assign n7578 = n7577 ^ n7416 ;
  assign n7579 = n7577 ^ x85 ;
  assign n7580 = n7578 & n7579 ;
  assign n7581 = n7580 ^ x85 ;
  assign n7413 = n7250 & n7360 ;
  assign n7414 = n7413 ^ n7083 ;
  assign n7582 = n7581 ^ n7414 ;
  assign n7583 = n7581 ^ x86 ;
  assign n7584 = n7582 & n7583 ;
  assign n7585 = n7584 ^ x86 ;
  assign n7411 = n7254 & n7360 ;
  assign n7412 = n7411 ^ n7081 ;
  assign n7586 = n7585 ^ n7412 ;
  assign n7587 = n7585 ^ x87 ;
  assign n7588 = n7586 & n7587 ;
  assign n7589 = n7588 ^ x87 ;
  assign n7409 = n7258 & n7360 ;
  assign n7410 = n7409 ^ n7079 ;
  assign n7590 = n7589 ^ n7410 ;
  assign n7591 = n7589 ^ x88 ;
  assign n7592 = n7590 & n7591 ;
  assign n7593 = n7592 ^ x88 ;
  assign n7407 = n7262 & n7360 ;
  assign n7408 = n7407 ^ n7077 ;
  assign n7594 = n7593 ^ n7408 ;
  assign n7595 = n7593 ^ x89 ;
  assign n7596 = n7594 & n7595 ;
  assign n7597 = n7596 ^ x89 ;
  assign n7405 = n7266 & n7360 ;
  assign n7406 = n7405 ^ n7075 ;
  assign n7598 = n7597 ^ n7406 ;
  assign n7599 = n7597 ^ x90 ;
  assign n7600 = n7598 & n7599 ;
  assign n7601 = n7600 ^ x90 ;
  assign n7403 = n7270 & n7360 ;
  assign n7404 = n7403 ^ n7073 ;
  assign n7602 = n7601 ^ n7404 ;
  assign n7603 = n7601 ^ x91 ;
  assign n7604 = n7602 & n7603 ;
  assign n7605 = n7604 ^ x91 ;
  assign n7401 = n7274 & n7360 ;
  assign n7402 = n7401 ^ n7071 ;
  assign n7606 = n7605 ^ n7402 ;
  assign n7607 = n7605 ^ x92 ;
  assign n7608 = n7606 & n7607 ;
  assign n7609 = n7608 ^ x92 ;
  assign n7399 = n7278 & n7360 ;
  assign n7400 = n7399 ^ n7069 ;
  assign n7610 = n7609 ^ n7400 ;
  assign n7611 = n7609 ^ x93 ;
  assign n7612 = n7610 & n7611 ;
  assign n7613 = n7612 ^ x93 ;
  assign n7397 = n7282 & n7360 ;
  assign n7398 = n7397 ^ n7067 ;
  assign n7614 = n7613 ^ n7398 ;
  assign n7615 = n7613 ^ x94 ;
  assign n7616 = n7614 & n7615 ;
  assign n7617 = n7616 ^ x94 ;
  assign n7395 = n7286 & n7360 ;
  assign n7396 = n7395 ^ n7065 ;
  assign n7618 = n7617 ^ n7396 ;
  assign n7619 = n7617 ^ x95 ;
  assign n7620 = n7618 & n7619 ;
  assign n7621 = n7620 ^ x95 ;
  assign n7393 = n7290 & n7360 ;
  assign n7394 = n7393 ^ n7063 ;
  assign n7622 = n7621 ^ n7394 ;
  assign n7623 = n7621 ^ x96 ;
  assign n7624 = n7622 & n7623 ;
  assign n7625 = n7624 ^ x96 ;
  assign n7626 = n7625 ^ n7386 ;
  assign n7627 = n7626 ^ n7391 ;
  assign n7628 = ~n7392 & n7627 ;
  assign n7629 = n7628 ^ n7391 ;
  assign n7630 = ~n7387 & n7629 ;
  assign n7631 = n7630 ^ x98 ;
  assign n7632 = n7631 ^ n7378 ;
  assign n7633 = n7632 ^ n7383 ;
  assign n7634 = ~n7384 & n7633 ;
  assign n7635 = n7634 ^ n7383 ;
  assign n7636 = ~n7379 & n7635 ;
  assign n7637 = n7636 ^ x100 ;
  assign n7640 = n7639 ^ n7637 ;
  assign n7641 = n7639 ^ x101 ;
  assign n7642 = n7640 & ~n7641 ;
  assign n7643 = n7642 ^ x101 ;
  assign n7375 = n7314 & n7360 ;
  assign n7376 = n7375 ^ n7041 ;
  assign n7644 = n7643 ^ n7376 ;
  assign n7645 = n7643 ^ x102 ;
  assign n7646 = n7644 & n7645 ;
  assign n7647 = n7646 ^ x102 ;
  assign n7373 = n7318 & n7360 ;
  assign n7374 = n7373 ^ n7038 ;
  assign n7648 = n7647 ^ n7374 ;
  assign n7649 = n7647 ^ x103 ;
  assign n7650 = n7648 & n7649 ;
  assign n7651 = n7650 ^ x103 ;
  assign n7371 = n7322 & n7360 ;
  assign n7372 = n7371 ^ n7036 ;
  assign n7652 = n7651 ^ n7372 ;
  assign n7653 = n7651 ^ x104 ;
  assign n7654 = n7652 & n7653 ;
  assign n7655 = n7654 ^ x104 ;
  assign n7369 = n7326 & n7360 ;
  assign n7370 = n7369 ^ n7033 ;
  assign n7656 = n7655 ^ n7370 ;
  assign n7657 = n7655 ^ x105 ;
  assign n7658 = n7656 & n7657 ;
  assign n7659 = n7658 ^ x105 ;
  assign n7660 = n7659 ^ n7362 ;
  assign n7661 = n7660 ^ n7367 ;
  assign n7662 = ~n7368 & n7661 ;
  assign n7663 = n7662 ^ n7367 ;
  assign n7664 = ~n7363 & n7663 ;
  assign n7665 = n7664 ^ x107 ;
  assign n7669 = n7668 ^ n7665 ;
  assign n7670 = n7668 ^ x108 ;
  assign n7671 = n7669 & ~n7670 ;
  assign n7672 = n7671 ^ x108 ;
  assign n7687 = x109 & n147 ;
  assign n7688 = ~n6089 & n7687 ;
  assign n7689 = n7688 ^ n147 ;
  assign n7674 = n148 & n7023 ;
  assign n7675 = n7352 ^ x108 ;
  assign n7678 = ~n7346 & n7675 ;
  assign n7679 = n7678 ^ x108 ;
  assign n7680 = n7674 & ~n7679 ;
  assign n7681 = n7680 ^ n7023 ;
  assign n7690 = n7681 ^ x109 ;
  assign n7691 = n7690 ^ n7672 ;
  assign n7692 = n7691 ^ n147 ;
  assign n7693 = n7689 & ~n7692 ;
  assign n7694 = n7672 & n7693 ;
  assign n7695 = n7694 ^ n7688 ;
  assign n7696 = n7695 ^ n147 ;
  assign n7830 = x64 & n7696 ;
  assign n7831 = n7830 ^ x18 ;
  assign n7832 = n7831 ^ n7828 ;
  assign n7833 = n7829 & n7832 ;
  assign n7834 = n7833 ^ x65 ;
  assign n7835 = n7834 ^ x66 ;
  assign n7840 = n7458 ^ x19 ;
  assign n7837 = ~x18 & x64 ;
  assign n7838 = n7837 ^ x65 ;
  assign n7839 = n7696 & n7838 ;
  assign n7841 = n7840 ^ n7839 ;
  assign n7842 = n7841 ^ n7834 ;
  assign n7843 = n7835 & n7842 ;
  assign n7844 = n7843 ^ x66 ;
  assign n7825 = n7486 ^ x66 ;
  assign n7826 = n7696 & ~n7825 ;
  assign n7827 = n7826 ^ n7456 ;
  assign n7845 = n7844 ^ n7827 ;
  assign n7846 = n7844 ^ x67 ;
  assign n7847 = n7845 & n7846 ;
  assign n7848 = n7847 ^ x67 ;
  assign n7823 = n7490 & n7696 ;
  assign n7824 = n7823 ^ n7506 ;
  assign n7849 = n7848 ^ n7824 ;
  assign n7850 = n7848 ^ x68 ;
  assign n7851 = n7849 & n7850 ;
  assign n7852 = n7851 ^ x68 ;
  assign n7854 = n7852 ^ x69 ;
  assign n7923 = n7583 & n7696 ;
  assign n7924 = n7923 ^ n7414 ;
  assign n7772 = n7579 & n7696 ;
  assign n7773 = n7772 ^ n7416 ;
  assign n7774 = n7773 ^ x86 ;
  assign n7778 = n7773 ^ x85 ;
  assign n7775 = n7575 & n7696 ;
  assign n7776 = n7775 ^ n7418 ;
  assign n7777 = n7776 ^ n7773 ;
  assign n7779 = n7778 ^ n7777 ;
  assign n7821 = n7511 & n7696 ;
  assign n7822 = n7821 ^ n7452 ;
  assign n7853 = n7852 ^ n7822 ;
  assign n7855 = n7853 & n7854 ;
  assign n7856 = n7855 ^ x69 ;
  assign n7819 = n7515 & n7696 ;
  assign n7820 = n7819 ^ n7450 ;
  assign n7857 = n7856 ^ n7820 ;
  assign n7858 = n7856 ^ x70 ;
  assign n7859 = n7857 & n7858 ;
  assign n7860 = n7859 ^ x70 ;
  assign n7817 = n7519 & n7696 ;
  assign n7818 = n7817 ^ n7448 ;
  assign n7861 = n7860 ^ n7818 ;
  assign n7862 = n7860 ^ x71 ;
  assign n7863 = n7861 & n7862 ;
  assign n7864 = n7863 ^ x71 ;
  assign n7815 = n7523 & n7696 ;
  assign n7816 = n7815 ^ n7446 ;
  assign n7865 = n7864 ^ n7816 ;
  assign n7866 = n7864 ^ x72 ;
  assign n7867 = n7865 & n7866 ;
  assign n7868 = n7867 ^ x72 ;
  assign n7813 = n7527 & n7696 ;
  assign n7814 = n7813 ^ n7444 ;
  assign n7869 = n7868 ^ n7814 ;
  assign n7870 = n7868 ^ x73 ;
  assign n7871 = n7869 & n7870 ;
  assign n7872 = n7871 ^ x73 ;
  assign n7811 = n7531 & n7696 ;
  assign n7812 = n7811 ^ n7442 ;
  assign n7873 = n7872 ^ n7812 ;
  assign n7874 = n7872 ^ x74 ;
  assign n7875 = n7873 & n7874 ;
  assign n7876 = n7875 ^ x74 ;
  assign n7809 = n7535 & n7696 ;
  assign n7810 = n7809 ^ n7440 ;
  assign n7877 = n7876 ^ n7810 ;
  assign n7878 = n7876 ^ x75 ;
  assign n7879 = n7877 & n7878 ;
  assign n7880 = n7879 ^ x75 ;
  assign n7807 = n7539 & n7696 ;
  assign n7808 = n7807 ^ n7438 ;
  assign n7881 = n7880 ^ n7808 ;
  assign n7882 = n7880 ^ x76 ;
  assign n7883 = n7881 & n7882 ;
  assign n7884 = n7883 ^ x76 ;
  assign n7805 = n7543 & n7696 ;
  assign n7806 = n7805 ^ n7436 ;
  assign n7885 = n7884 ^ n7806 ;
  assign n7886 = n7884 ^ x77 ;
  assign n7887 = n7885 & n7886 ;
  assign n7888 = n7887 ^ x77 ;
  assign n7803 = n7547 & n7696 ;
  assign n7804 = n7803 ^ n7434 ;
  assign n7889 = n7888 ^ n7804 ;
  assign n7890 = n7888 ^ x78 ;
  assign n7891 = n7889 & n7890 ;
  assign n7892 = n7891 ^ x78 ;
  assign n7801 = n7551 & n7696 ;
  assign n7802 = n7801 ^ n7432 ;
  assign n7893 = n7892 ^ n7802 ;
  assign n7894 = n7892 ^ x79 ;
  assign n7895 = n7893 & n7894 ;
  assign n7896 = n7895 ^ x79 ;
  assign n7799 = n7555 & n7696 ;
  assign n7800 = n7799 ^ n7430 ;
  assign n7897 = n7896 ^ n7800 ;
  assign n7898 = n7896 ^ x80 ;
  assign n7899 = n7897 & n7898 ;
  assign n7900 = n7899 ^ x80 ;
  assign n7796 = n7557 ^ x80 ;
  assign n7797 = n7696 & n7796 ;
  assign n7798 = n7797 ^ n7425 ;
  assign n7901 = n7900 ^ n7798 ;
  assign n7902 = n7900 ^ x81 ;
  assign n7903 = n7901 & n7902 ;
  assign n7904 = n7903 ^ x81 ;
  assign n7785 = n7425 ^ x81 ;
  assign n7786 = n7785 ^ n7557 ;
  assign n7787 = n7786 ^ x80 ;
  assign n7788 = n7787 ^ n7785 ;
  assign n7790 = n7557 ^ x81 ;
  assign n7791 = n7790 ^ n7785 ;
  assign n7792 = ~n7788 & ~n7791 ;
  assign n7793 = n7792 ^ n7785 ;
  assign n7794 = n7696 & ~n7793 ;
  assign n7795 = n7794 ^ n7422 ;
  assign n7905 = n7904 ^ n7795 ;
  assign n7906 = n7904 ^ x82 ;
  assign n7907 = n7905 & n7906 ;
  assign n7908 = n7907 ^ x82 ;
  assign n7782 = n7563 ^ x82 ;
  assign n7783 = n7696 & n7782 ;
  assign n7784 = n7783 ^ n7565 ;
  assign n7909 = n7908 ^ n7784 ;
  assign n7910 = n7908 ^ x83 ;
  assign n7911 = n7909 & n7910 ;
  assign n7912 = n7911 ^ x83 ;
  assign n7780 = n7571 & n7696 ;
  assign n7781 = n7780 ^ n7420 ;
  assign n7913 = n7912 ^ n7781 ;
  assign n7914 = n7912 ^ x84 ;
  assign n7915 = n7913 & n7914 ;
  assign n7916 = n7915 ^ x84 ;
  assign n7917 = n7916 ^ n7773 ;
  assign n7918 = n7917 ^ n7778 ;
  assign n7919 = ~n7779 & n7918 ;
  assign n7920 = n7919 ^ n7778 ;
  assign n7921 = ~n7774 & n7920 ;
  assign n7922 = n7921 ^ x86 ;
  assign n7925 = n7924 ^ n7922 ;
  assign n7926 = n7924 ^ x87 ;
  assign n7927 = n7925 & ~n7926 ;
  assign n7928 = n7927 ^ x87 ;
  assign n7770 = n7587 & n7696 ;
  assign n7771 = n7770 ^ n7412 ;
  assign n7929 = n7928 ^ n7771 ;
  assign n7930 = n7928 ^ x88 ;
  assign n7931 = n7929 & n7930 ;
  assign n7932 = n7931 ^ x88 ;
  assign n7768 = n7591 & n7696 ;
  assign n7769 = n7768 ^ n7410 ;
  assign n7933 = n7932 ^ n7769 ;
  assign n7934 = n7932 ^ x89 ;
  assign n7935 = n7933 & n7934 ;
  assign n7936 = n7935 ^ x89 ;
  assign n7766 = n7595 & n7696 ;
  assign n7767 = n7766 ^ n7408 ;
  assign n7937 = n7936 ^ n7767 ;
  assign n7938 = n7936 ^ x90 ;
  assign n7939 = n7937 & n7938 ;
  assign n7940 = n7939 ^ x90 ;
  assign n7764 = n7599 & n7696 ;
  assign n7765 = n7764 ^ n7406 ;
  assign n7941 = n7940 ^ n7765 ;
  assign n7942 = n7940 ^ x91 ;
  assign n7943 = n7941 & n7942 ;
  assign n7944 = n7943 ^ x91 ;
  assign n7762 = n7603 & n7696 ;
  assign n7763 = n7762 ^ n7404 ;
  assign n7945 = n7944 ^ n7763 ;
  assign n7946 = n7944 ^ x92 ;
  assign n7947 = n7945 & n7946 ;
  assign n7948 = n7947 ^ x92 ;
  assign n7760 = n7607 & n7696 ;
  assign n7761 = n7760 ^ n7402 ;
  assign n7949 = n7948 ^ n7761 ;
  assign n7950 = n7948 ^ x93 ;
  assign n7951 = n7949 & n7950 ;
  assign n7952 = n7951 ^ x93 ;
  assign n7758 = n7611 & n7696 ;
  assign n7759 = n7758 ^ n7400 ;
  assign n7953 = n7952 ^ n7759 ;
  assign n7954 = n7952 ^ x94 ;
  assign n7955 = n7953 & n7954 ;
  assign n7956 = n7955 ^ x94 ;
  assign n7756 = n7615 & n7696 ;
  assign n7757 = n7756 ^ n7398 ;
  assign n7957 = n7956 ^ n7757 ;
  assign n7958 = n7956 ^ x95 ;
  assign n7959 = n7957 & n7958 ;
  assign n7960 = n7959 ^ x95 ;
  assign n7754 = n7619 & n7696 ;
  assign n7755 = n7754 ^ n7396 ;
  assign n7961 = n7960 ^ n7755 ;
  assign n7962 = n7960 ^ x96 ;
  assign n7963 = n7961 & n7962 ;
  assign n7964 = n7963 ^ x96 ;
  assign n7752 = n7623 & n7696 ;
  assign n7753 = n7752 ^ n7394 ;
  assign n7965 = n7964 ^ n7753 ;
  assign n7966 = n7964 ^ x97 ;
  assign n7967 = n7965 & n7966 ;
  assign n7968 = n7967 ^ x97 ;
  assign n7749 = n7625 ^ x97 ;
  assign n7750 = n7696 & n7749 ;
  assign n7751 = n7750 ^ n7389 ;
  assign n7969 = n7968 ^ n7751 ;
  assign n7970 = n7968 ^ x98 ;
  assign n7971 = n7969 & n7970 ;
  assign n7972 = n7971 ^ x98 ;
  assign n7738 = n7389 ^ x98 ;
  assign n7739 = n7738 ^ n7625 ;
  assign n7740 = n7739 ^ x97 ;
  assign n7741 = n7740 ^ n7738 ;
  assign n7743 = n7625 ^ x98 ;
  assign n7744 = n7743 ^ n7738 ;
  assign n7745 = ~n7741 & ~n7744 ;
  assign n7746 = n7745 ^ n7738 ;
  assign n7747 = n7696 & ~n7746 ;
  assign n7748 = n7747 ^ n7386 ;
  assign n7973 = n7972 ^ n7748 ;
  assign n7974 = n7972 ^ x99 ;
  assign n7975 = n7973 & n7974 ;
  assign n7976 = n7975 ^ x99 ;
  assign n7735 = n7631 ^ x99 ;
  assign n7736 = n7696 & n7735 ;
  assign n7737 = n7736 ^ n7381 ;
  assign n7977 = n7976 ^ n7737 ;
  assign n7978 = n7976 ^ x100 ;
  assign n7979 = n7977 & n7978 ;
  assign n7980 = n7979 ^ x100 ;
  assign n7724 = n7381 ^ x100 ;
  assign n7725 = n7724 ^ n7631 ;
  assign n7726 = n7725 ^ x99 ;
  assign n7727 = n7726 ^ n7724 ;
  assign n7729 = n7631 ^ x100 ;
  assign n7730 = n7729 ^ n7724 ;
  assign n7731 = ~n7727 & ~n7730 ;
  assign n7732 = n7731 ^ n7724 ;
  assign n7733 = n7696 & ~n7732 ;
  assign n7734 = n7733 ^ n7378 ;
  assign n7981 = n7980 ^ n7734 ;
  assign n7982 = n7980 ^ x101 ;
  assign n7983 = n7981 & n7982 ;
  assign n7984 = n7983 ^ x101 ;
  assign n7721 = n7637 ^ x101 ;
  assign n7722 = n7696 & n7721 ;
  assign n7723 = n7722 ^ n7639 ;
  assign n7985 = n7984 ^ n7723 ;
  assign n7986 = n7984 ^ x102 ;
  assign n7987 = n7985 & n7986 ;
  assign n7988 = n7987 ^ x102 ;
  assign n7719 = n7645 & n7696 ;
  assign n7720 = n7719 ^ n7376 ;
  assign n7989 = n7988 ^ n7720 ;
  assign n7990 = n7988 ^ x103 ;
  assign n7991 = n7989 & n7990 ;
  assign n7992 = n7991 ^ x103 ;
  assign n7717 = n7649 & n7696 ;
  assign n7718 = n7717 ^ n7374 ;
  assign n7993 = n7992 ^ n7718 ;
  assign n7994 = n7992 ^ x104 ;
  assign n7995 = n7993 & n7994 ;
  assign n7996 = n7995 ^ x104 ;
  assign n7715 = n7653 & n7696 ;
  assign n7716 = n7715 ^ n7372 ;
  assign n7997 = n7996 ^ n7716 ;
  assign n7998 = n7996 ^ x105 ;
  assign n7999 = n7997 & n7998 ;
  assign n8000 = n7999 ^ x105 ;
  assign n7713 = n7657 & n7696 ;
  assign n7714 = n7713 ^ n7370 ;
  assign n8001 = n8000 ^ n7714 ;
  assign n8002 = n8000 ^ x106 ;
  assign n8003 = n8001 & n8002 ;
  assign n8004 = n8003 ^ x106 ;
  assign n7710 = n7659 ^ x106 ;
  assign n7711 = n7696 & n7710 ;
  assign n7712 = n7711 ^ n7365 ;
  assign n8005 = n8004 ^ n7712 ;
  assign n8006 = n8004 ^ x107 ;
  assign n8007 = n8005 & n8006 ;
  assign n8008 = n8007 ^ x107 ;
  assign n7699 = n7365 ^ x107 ;
  assign n7700 = n7699 ^ n7659 ;
  assign n7701 = n7700 ^ x106 ;
  assign n7702 = n7701 ^ n7699 ;
  assign n7704 = n7659 ^ x107 ;
  assign n7705 = n7704 ^ n7699 ;
  assign n7706 = ~n7702 & ~n7705 ;
  assign n7707 = n7706 ^ n7699 ;
  assign n7708 = n7696 & ~n7707 ;
  assign n7709 = n7708 ^ n7362 ;
  assign n8009 = n8008 ^ n7709 ;
  assign n8010 = n8008 ^ x108 ;
  assign n8011 = n8009 & n8010 ;
  assign n8012 = n8011 ^ x108 ;
  assign n7686 = n7665 ^ x108 ;
  assign n7697 = n7686 & n7696 ;
  assign n7698 = n7697 ^ n7668 ;
  assign n8013 = n8012 ^ n7698 ;
  assign n8016 = n7698 ^ x109 ;
  assign n8017 = n8013 & ~n8016 ;
  assign n8014 = x110 ^ x109 ;
  assign n8018 = n8017 ^ n8014 ;
  assign n7673 = n7672 ^ x109 ;
  assign n7682 = n147 & n7681 ;
  assign n7683 = n7673 & n7682 ;
  assign n7684 = n7683 ^ n7681 ;
  assign n8021 = n7684 ^ x110 ;
  assign n8024 = n8018 & ~n8021 ;
  assign n8025 = n8024 ^ x110 ;
  assign n8026 = n145 & ~n8025 ;
  assign n8122 = n7854 & n8026 ;
  assign n8123 = n8122 ^ n7822 ;
  assign n8124 = n8123 ^ x70 ;
  assign n8125 = n7850 & n8026 ;
  assign n8126 = n8125 ^ n7824 ;
  assign n8127 = n8126 ^ x69 ;
  assign n8183 = n7846 & n8026 ;
  assign n8184 = n8183 ^ n7827 ;
  assign n8177 = n7835 & n8026 ;
  assign n8178 = n8177 ^ n7841 ;
  assign n8151 = ~x17 & x65 ;
  assign n8159 = n7829 & n8026 ;
  assign n8139 = ~x16 & x64 ;
  assign n8154 = n8026 ^ x17 ;
  assign n8155 = n8154 ^ n8026 ;
  assign n8156 = ~x65 & n8155 ;
  assign n8157 = n8156 ^ n8026 ;
  assign n8158 = n8139 & ~n8157 ;
  assign n8160 = n8159 ^ n8158 ;
  assign n8161 = n7831 & ~n8160 ;
  assign n8162 = ~n8151 & n8161 ;
  assign n8144 = x64 ^ x17 ;
  assign n8145 = n7831 ^ n191 ;
  assign n8146 = n8144 & n8145 ;
  assign n8147 = n8026 & n8146 ;
  assign n8163 = n8162 ^ n8147 ;
  assign n8148 = x16 & x65 ;
  assign n8149 = ~n191 & ~n8148 ;
  assign n8150 = n8147 & n8149 ;
  assign n8164 = n8163 ^ n8150 ;
  assign n8140 = ~n7831 & n8139 ;
  assign n8128 = n7831 ^ x65 ;
  assign n8129 = n8128 ^ n8026 ;
  assign n8131 = x17 ^ x16 ;
  assign n8130 = n8026 ^ n7831 ;
  assign n8132 = n8131 ^ n8130 ;
  assign n8133 = n7831 ^ x16 ;
  assign n8134 = n8133 ^ n8131 ;
  assign n8135 = ~n8132 & ~n8134 ;
  assign n8136 = n8135 ^ n8131 ;
  assign n8137 = n8129 & n8136 ;
  assign n8138 = x64 & n8137 ;
  assign n8141 = n8140 ^ n8138 ;
  assign n8165 = n8141 ^ n8140 ;
  assign n8142 = ~x17 & n8141 ;
  assign n8166 = n8165 ^ n8142 ;
  assign n8167 = ~x66 & ~n8166 ;
  assign n8168 = x64 & n8026 ;
  assign n8169 = n8151 & ~n8168 ;
  assign n8170 = ~n8130 & n8169 ;
  assign n8171 = n8170 ^ n8167 ;
  assign n8172 = n8167 & n8171 ;
  assign n8173 = ~n8164 & n8172 ;
  assign n8175 = n8173 ^ n8164 ;
  assign n8179 = n8178 ^ n8175 ;
  assign n8180 = n8178 ^ x67 ;
  assign n8181 = ~n8179 & ~n8180 ;
  assign n8182 = n8181 ^ x67 ;
  assign n8185 = n8184 ^ n8182 ;
  assign n8186 = n8184 ^ x68 ;
  assign n8187 = n8185 & ~n8186 ;
  assign n8188 = n8187 ^ x68 ;
  assign n8189 = n8188 ^ n8126 ;
  assign n8190 = ~n8127 & n8189 ;
  assign n8191 = n8190 ^ x69 ;
  assign n8192 = n8191 ^ n8123 ;
  assign n8193 = ~n8124 & n8192 ;
  assign n8194 = n8193 ^ x70 ;
  assign n8120 = n7858 & n8026 ;
  assign n8121 = n8120 ^ n7820 ;
  assign n8195 = n8194 ^ n8121 ;
  assign n8196 = n8194 ^ x71 ;
  assign n8197 = n8195 & n8196 ;
  assign n8198 = n8197 ^ x71 ;
  assign n8118 = n7862 & n8026 ;
  assign n8119 = n8118 ^ n7818 ;
  assign n8199 = n8198 ^ n8119 ;
  assign n8200 = n8198 ^ x72 ;
  assign n8201 = n8199 & n8200 ;
  assign n8202 = n8201 ^ x72 ;
  assign n8116 = n7866 & n8026 ;
  assign n8117 = n8116 ^ n7816 ;
  assign n8203 = n8202 ^ n8117 ;
  assign n8204 = n8202 ^ x73 ;
  assign n8205 = n8203 & n8204 ;
  assign n8206 = n8205 ^ x73 ;
  assign n8114 = n7870 & n8026 ;
  assign n8115 = n8114 ^ n7814 ;
  assign n8207 = n8206 ^ n8115 ;
  assign n8208 = n8206 ^ x74 ;
  assign n8209 = n8207 & n8208 ;
  assign n8210 = n8209 ^ x74 ;
  assign n8112 = n7874 & n8026 ;
  assign n8113 = n8112 ^ n7812 ;
  assign n8211 = n8210 ^ n8113 ;
  assign n8212 = n8210 ^ x75 ;
  assign n8213 = n8211 & n8212 ;
  assign n8214 = n8213 ^ x75 ;
  assign n8110 = n7878 & n8026 ;
  assign n8111 = n8110 ^ n7810 ;
  assign n8215 = n8214 ^ n8111 ;
  assign n8216 = n8214 ^ x76 ;
  assign n8217 = n8215 & n8216 ;
  assign n8218 = n8217 ^ x76 ;
  assign n8108 = n7882 & n8026 ;
  assign n8109 = n8108 ^ n7808 ;
  assign n8219 = n8218 ^ n8109 ;
  assign n8220 = n8218 ^ x77 ;
  assign n8221 = n8219 & n8220 ;
  assign n8222 = n8221 ^ x77 ;
  assign n8106 = n7886 & n8026 ;
  assign n8107 = n8106 ^ n7806 ;
  assign n8223 = n8222 ^ n8107 ;
  assign n8224 = n8222 ^ x78 ;
  assign n8225 = n8223 & n8224 ;
  assign n8226 = n8225 ^ x78 ;
  assign n8104 = n7890 & n8026 ;
  assign n8105 = n8104 ^ n7804 ;
  assign n8227 = n8226 ^ n8105 ;
  assign n8228 = n8226 ^ x79 ;
  assign n8229 = n8227 & n8228 ;
  assign n8230 = n8229 ^ x79 ;
  assign n8102 = n7894 & n8026 ;
  assign n8103 = n8102 ^ n7802 ;
  assign n8231 = n8230 ^ n8103 ;
  assign n8232 = n8230 ^ x80 ;
  assign n8233 = n8231 & n8232 ;
  assign n8234 = n8233 ^ x80 ;
  assign n8100 = n7898 & n8026 ;
  assign n8101 = n8100 ^ n7800 ;
  assign n8235 = n8234 ^ n8101 ;
  assign n8236 = n8234 ^ x81 ;
  assign n8237 = n8235 & n8236 ;
  assign n8238 = n8237 ^ x81 ;
  assign n8240 = n8238 ^ x82 ;
  assign n8346 = ~x112 & n144 ;
  assign n7685 = n145 & n7684 ;
  assign n8019 = n7685 & n8018 ;
  assign n8020 = n8019 ^ n7684 ;
  assign n8347 = n8020 ^ x111 ;
  assign n8031 = n8002 & n8026 ;
  assign n8032 = n8031 ^ n7714 ;
  assign n8033 = n8032 ^ x107 ;
  assign n8034 = n7998 & n8026 ;
  assign n8035 = n8034 ^ n7716 ;
  assign n8036 = n8035 ^ x106 ;
  assign n8045 = n7978 & n8026 ;
  assign n8046 = n8045 ^ n7737 ;
  assign n8047 = n8046 ^ x101 ;
  assign n8048 = n7974 & n8026 ;
  assign n8049 = n8048 ^ n7748 ;
  assign n8050 = n8049 ^ x100 ;
  assign n8059 = n7954 & n8026 ;
  assign n8060 = n8059 ^ n7759 ;
  assign n8061 = n8060 ^ x95 ;
  assign n8062 = n7950 & n8026 ;
  assign n8063 = n8062 ^ n7761 ;
  assign n8064 = n8063 ^ x94 ;
  assign n8098 = n7902 & n8026 ;
  assign n8099 = n8098 ^ n7798 ;
  assign n8239 = n8238 ^ n8099 ;
  assign n8241 = n8239 & n8240 ;
  assign n8242 = n8241 ^ x82 ;
  assign n8096 = n7906 & n8026 ;
  assign n8097 = n8096 ^ n7795 ;
  assign n8243 = n8242 ^ n8097 ;
  assign n8244 = n8242 ^ x83 ;
  assign n8245 = n8243 & n8244 ;
  assign n8246 = n8245 ^ x83 ;
  assign n8094 = n7910 & n8026 ;
  assign n8095 = n8094 ^ n7784 ;
  assign n8247 = n8246 ^ n8095 ;
  assign n8248 = n8246 ^ x84 ;
  assign n8249 = n8247 & n8248 ;
  assign n8250 = n8249 ^ x84 ;
  assign n8092 = n7914 & n8026 ;
  assign n8093 = n8092 ^ n7781 ;
  assign n8251 = n8250 ^ n8093 ;
  assign n8252 = n8250 ^ x85 ;
  assign n8253 = n8251 & n8252 ;
  assign n8254 = n8253 ^ x85 ;
  assign n8089 = n7916 ^ x85 ;
  assign n8090 = n8026 & n8089 ;
  assign n8091 = n8090 ^ n7776 ;
  assign n8255 = n8254 ^ n8091 ;
  assign n8256 = n8254 ^ x86 ;
  assign n8257 = n8255 & n8256 ;
  assign n8258 = n8257 ^ x86 ;
  assign n8078 = n7776 ^ x86 ;
  assign n8079 = n8078 ^ n7916 ;
  assign n8080 = n8079 ^ x85 ;
  assign n8081 = n8080 ^ n8078 ;
  assign n8083 = n7916 ^ x86 ;
  assign n8084 = n8083 ^ n8078 ;
  assign n8085 = ~n8081 & ~n8084 ;
  assign n8086 = n8085 ^ n8078 ;
  assign n8087 = n8026 & ~n8086 ;
  assign n8088 = n8087 ^ n7773 ;
  assign n8259 = n8258 ^ n8088 ;
  assign n8260 = n8258 ^ x87 ;
  assign n8261 = n8259 & n8260 ;
  assign n8262 = n8261 ^ x87 ;
  assign n8075 = n7922 ^ x87 ;
  assign n8076 = n8026 & n8075 ;
  assign n8077 = n8076 ^ n7924 ;
  assign n8263 = n8262 ^ n8077 ;
  assign n8264 = n8262 ^ x88 ;
  assign n8265 = n8263 & n8264 ;
  assign n8266 = n8265 ^ x88 ;
  assign n8073 = n7930 & n8026 ;
  assign n8074 = n8073 ^ n7771 ;
  assign n8267 = n8266 ^ n8074 ;
  assign n8268 = n8266 ^ x89 ;
  assign n8269 = n8267 & n8268 ;
  assign n8270 = n8269 ^ x89 ;
  assign n8071 = n7934 & n8026 ;
  assign n8072 = n8071 ^ n7769 ;
  assign n8271 = n8270 ^ n8072 ;
  assign n8272 = n8270 ^ x90 ;
  assign n8273 = n8271 & n8272 ;
  assign n8274 = n8273 ^ x90 ;
  assign n8069 = n7938 & n8026 ;
  assign n8070 = n8069 ^ n7767 ;
  assign n8275 = n8274 ^ n8070 ;
  assign n8276 = n8274 ^ x91 ;
  assign n8277 = n8275 & n8276 ;
  assign n8278 = n8277 ^ x91 ;
  assign n8067 = n7942 & n8026 ;
  assign n8068 = n8067 ^ n7765 ;
  assign n8279 = n8278 ^ n8068 ;
  assign n8280 = n8278 ^ x92 ;
  assign n8281 = n8279 & n8280 ;
  assign n8282 = n8281 ^ x92 ;
  assign n8065 = n7946 & n8026 ;
  assign n8066 = n8065 ^ n7763 ;
  assign n8283 = n8282 ^ n8066 ;
  assign n8284 = n8282 ^ x93 ;
  assign n8285 = n8283 & n8284 ;
  assign n8286 = n8285 ^ x93 ;
  assign n8287 = n8286 ^ n8063 ;
  assign n8288 = ~n8064 & n8287 ;
  assign n8289 = n8288 ^ x94 ;
  assign n8290 = n8289 ^ n8060 ;
  assign n8291 = ~n8061 & n8290 ;
  assign n8292 = n8291 ^ x95 ;
  assign n8057 = n7958 & n8026 ;
  assign n8058 = n8057 ^ n7757 ;
  assign n8293 = n8292 ^ n8058 ;
  assign n8294 = n8292 ^ x96 ;
  assign n8295 = n8293 & n8294 ;
  assign n8296 = n8295 ^ x96 ;
  assign n8055 = n7962 & n8026 ;
  assign n8056 = n8055 ^ n7755 ;
  assign n8297 = n8296 ^ n8056 ;
  assign n8298 = n8296 ^ x97 ;
  assign n8299 = n8297 & n8298 ;
  assign n8300 = n8299 ^ x97 ;
  assign n8053 = n7966 & n8026 ;
  assign n8054 = n8053 ^ n7753 ;
  assign n8301 = n8300 ^ n8054 ;
  assign n8302 = n8300 ^ x98 ;
  assign n8303 = n8301 & n8302 ;
  assign n8304 = n8303 ^ x98 ;
  assign n8051 = n7970 & n8026 ;
  assign n8052 = n8051 ^ n7751 ;
  assign n8305 = n8304 ^ n8052 ;
  assign n8306 = n8304 ^ x99 ;
  assign n8307 = n8305 & n8306 ;
  assign n8308 = n8307 ^ x99 ;
  assign n8309 = n8308 ^ n8049 ;
  assign n8310 = ~n8050 & n8309 ;
  assign n8311 = n8310 ^ x100 ;
  assign n8312 = n8311 ^ n8046 ;
  assign n8313 = ~n8047 & n8312 ;
  assign n8314 = n8313 ^ x101 ;
  assign n8043 = n7982 & n8026 ;
  assign n8044 = n8043 ^ n7734 ;
  assign n8315 = n8314 ^ n8044 ;
  assign n8316 = n8314 ^ x102 ;
  assign n8317 = n8315 & n8316 ;
  assign n8318 = n8317 ^ x102 ;
  assign n8041 = n7986 & n8026 ;
  assign n8042 = n8041 ^ n7723 ;
  assign n8319 = n8318 ^ n8042 ;
  assign n8320 = n8318 ^ x103 ;
  assign n8321 = n8319 & n8320 ;
  assign n8322 = n8321 ^ x103 ;
  assign n8039 = n7990 & n8026 ;
  assign n8040 = n8039 ^ n7720 ;
  assign n8323 = n8322 ^ n8040 ;
  assign n8324 = n8322 ^ x104 ;
  assign n8325 = n8323 & n8324 ;
  assign n8326 = n8325 ^ x104 ;
  assign n8037 = n7994 & n8026 ;
  assign n8038 = n8037 ^ n7718 ;
  assign n8327 = n8326 ^ n8038 ;
  assign n8328 = n8326 ^ x105 ;
  assign n8329 = n8327 & n8328 ;
  assign n8330 = n8329 ^ x105 ;
  assign n8331 = n8330 ^ n8035 ;
  assign n8332 = ~n8036 & n8331 ;
  assign n8333 = n8332 ^ x106 ;
  assign n8334 = n8333 ^ n8032 ;
  assign n8335 = ~n8033 & n8334 ;
  assign n8336 = n8335 ^ x107 ;
  assign n8029 = n8006 & n8026 ;
  assign n8030 = n8029 ^ n7712 ;
  assign n8337 = n8336 ^ n8030 ;
  assign n8338 = n8336 ^ x108 ;
  assign n8339 = n8337 & n8338 ;
  assign n8340 = n8339 ^ x108 ;
  assign n8027 = n8010 & n8026 ;
  assign n8028 = n8027 ^ n7709 ;
  assign n8341 = n8340 ^ n8028 ;
  assign n8342 = n8340 ^ x109 ;
  assign n8343 = n8341 & n8342 ;
  assign n8344 = n8343 ^ x109 ;
  assign n8345 = n8344 ^ x110 ;
  assign n8348 = n8012 ^ x109 ;
  assign n8349 = n8026 & n8348 ;
  assign n8350 = n8349 ^ n7698 ;
  assign n8351 = n8350 ^ n8344 ;
  assign n8352 = n8345 & n8351 ;
  assign n8353 = n8352 ^ x110 ;
  assign n8354 = n8353 ^ x111 ;
  assign n8355 = ~n8347 & n8354 ;
  assign n8356 = n8355 ^ x111 ;
  assign n8357 = n8346 & ~n8356 ;
  assign n8561 = n8240 & n8357 ;
  assign n8562 = n8561 ^ n8099 ;
  assign n8424 = n8236 & n8357 ;
  assign n8425 = n8424 ^ n8101 ;
  assign n8426 = n8425 ^ x82 ;
  assign n8430 = n8425 ^ x81 ;
  assign n8427 = n8232 & n8357 ;
  assign n8428 = n8427 ^ n8103 ;
  assign n8429 = n8428 ^ n8425 ;
  assign n8431 = n8430 ^ n8429 ;
  assign n8480 = n8168 ^ x17 ;
  assign n8478 = n8139 ^ x65 ;
  assign n8479 = n8357 & n8478 ;
  assign n8481 = n8480 ^ n8479 ;
  assign n8482 = n8481 ^ x66 ;
  assign n8484 = x64 ^ x16 ;
  assign n8485 = n8484 ^ x65 ;
  assign n8486 = n8485 ^ n8148 ;
  assign n8487 = n8486 ^ n8357 ;
  assign n8488 = n8487 ^ n8148 ;
  assign n8489 = x65 ^ x15 ;
  assign n8492 = n8488 & ~n8489 ;
  assign n8493 = n8492 ^ n8148 ;
  assign n8494 = x64 & n8493 ;
  assign n8483 = n8148 ^ x65 ;
  assign n8495 = n8494 ^ n8483 ;
  assign n8496 = n8495 ^ n8481 ;
  assign n8497 = ~n8482 & n8496 ;
  assign n8498 = n8497 ^ x66 ;
  assign n8472 = x17 & x65 ;
  assign n8463 = x65 ^ x16 ;
  assign n8464 = n8144 ^ x65 ;
  assign n8465 = n8464 ^ n8026 ;
  assign n8466 = ~n8463 & n8465 ;
  assign n8473 = n8472 ^ n8466 ;
  assign n8474 = ~x64 & n8473 ;
  assign n8469 = n8466 ^ n6836 ;
  assign n8475 = n8474 ^ n8469 ;
  assign n8476 = n8357 & n8475 ;
  assign n8462 = n8159 ^ n7831 ;
  assign n8477 = n8476 ^ n8462 ;
  assign n8499 = n8498 ^ n8477 ;
  assign n8500 = n8498 ^ x67 ;
  assign n8501 = n8499 & n8500 ;
  assign n8502 = n8501 ^ x67 ;
  assign n8459 = n8175 ^ x67 ;
  assign n8460 = n8357 & ~n8459 ;
  assign n8461 = n8460 ^ n8178 ;
  assign n8503 = n8502 ^ n8461 ;
  assign n8504 = n8502 ^ x68 ;
  assign n8505 = n8503 & n8504 ;
  assign n8506 = n8505 ^ x68 ;
  assign n8456 = n8182 ^ x68 ;
  assign n8457 = n8357 & n8456 ;
  assign n8458 = n8457 ^ n8184 ;
  assign n8507 = n8506 ^ n8458 ;
  assign n8508 = n8506 ^ x69 ;
  assign n8509 = n8507 & n8508 ;
  assign n8510 = n8509 ^ x69 ;
  assign n8453 = n8188 ^ x69 ;
  assign n8454 = n8357 & n8453 ;
  assign n8455 = n8454 ^ n8126 ;
  assign n8511 = n8510 ^ n8455 ;
  assign n8512 = n8510 ^ x70 ;
  assign n8513 = n8511 & n8512 ;
  assign n8514 = n8513 ^ x70 ;
  assign n8450 = n8191 ^ x70 ;
  assign n8451 = n8357 & n8450 ;
  assign n8452 = n8451 ^ n8123 ;
  assign n8515 = n8514 ^ n8452 ;
  assign n8516 = n8514 ^ x71 ;
  assign n8517 = n8515 & n8516 ;
  assign n8518 = n8517 ^ x71 ;
  assign n8448 = n8196 & n8357 ;
  assign n8449 = n8448 ^ n8121 ;
  assign n8519 = n8518 ^ n8449 ;
  assign n8520 = n8518 ^ x72 ;
  assign n8521 = n8519 & n8520 ;
  assign n8522 = n8521 ^ x72 ;
  assign n8446 = n8200 & n8357 ;
  assign n8447 = n8446 ^ n8119 ;
  assign n8523 = n8522 ^ n8447 ;
  assign n8524 = n8522 ^ x73 ;
  assign n8525 = n8523 & n8524 ;
  assign n8526 = n8525 ^ x73 ;
  assign n8444 = n8204 & n8357 ;
  assign n8445 = n8444 ^ n8117 ;
  assign n8527 = n8526 ^ n8445 ;
  assign n8528 = n8526 ^ x74 ;
  assign n8529 = n8527 & n8528 ;
  assign n8530 = n8529 ^ x74 ;
  assign n8442 = n8208 & n8357 ;
  assign n8443 = n8442 ^ n8115 ;
  assign n8531 = n8530 ^ n8443 ;
  assign n8532 = n8530 ^ x75 ;
  assign n8533 = n8531 & n8532 ;
  assign n8534 = n8533 ^ x75 ;
  assign n8440 = n8212 & n8357 ;
  assign n8441 = n8440 ^ n8113 ;
  assign n8535 = n8534 ^ n8441 ;
  assign n8536 = n8534 ^ x76 ;
  assign n8537 = n8535 & n8536 ;
  assign n8538 = n8537 ^ x76 ;
  assign n8438 = n8216 & n8357 ;
  assign n8439 = n8438 ^ n8111 ;
  assign n8539 = n8538 ^ n8439 ;
  assign n8540 = n8538 ^ x77 ;
  assign n8541 = n8539 & n8540 ;
  assign n8542 = n8541 ^ x77 ;
  assign n8436 = n8220 & n8357 ;
  assign n8437 = n8436 ^ n8109 ;
  assign n8543 = n8542 ^ n8437 ;
  assign n8544 = n8542 ^ x78 ;
  assign n8545 = n8543 & n8544 ;
  assign n8546 = n8545 ^ x78 ;
  assign n8434 = n8224 & n8357 ;
  assign n8435 = n8434 ^ n8107 ;
  assign n8547 = n8546 ^ n8435 ;
  assign n8548 = n8546 ^ x79 ;
  assign n8549 = n8547 & n8548 ;
  assign n8550 = n8549 ^ x79 ;
  assign n8432 = n8228 & n8357 ;
  assign n8433 = n8432 ^ n8105 ;
  assign n8551 = n8550 ^ n8433 ;
  assign n8552 = n8550 ^ x80 ;
  assign n8553 = n8551 & n8552 ;
  assign n8554 = n8553 ^ x80 ;
  assign n8555 = n8554 ^ n8425 ;
  assign n8556 = n8555 ^ n8430 ;
  assign n8557 = ~n8431 & n8556 ;
  assign n8558 = n8557 ^ n8430 ;
  assign n8559 = ~n8426 & n8558 ;
  assign n8560 = n8559 ^ x82 ;
  assign n8563 = n8562 ^ n8560 ;
  assign n8564 = n8562 ^ x83 ;
  assign n8565 = n8563 & ~n8564 ;
  assign n8566 = n8565 ^ x83 ;
  assign n8422 = n8244 & n8357 ;
  assign n8423 = n8422 ^ n8097 ;
  assign n8567 = n8566 ^ n8423 ;
  assign n8568 = n8566 ^ x84 ;
  assign n8569 = n8567 & n8568 ;
  assign n8570 = n8569 ^ x84 ;
  assign n8420 = n8248 & n8357 ;
  assign n8421 = n8420 ^ n8095 ;
  assign n8571 = n8570 ^ n8421 ;
  assign n8572 = n8570 ^ x85 ;
  assign n8573 = n8571 & n8572 ;
  assign n8574 = n8573 ^ x85 ;
  assign n8418 = n8252 & n8357 ;
  assign n8419 = n8418 ^ n8093 ;
  assign n8575 = n8574 ^ n8419 ;
  assign n8576 = n8574 ^ x86 ;
  assign n8577 = n8575 & n8576 ;
  assign n8578 = n8577 ^ x86 ;
  assign n8416 = n8256 & n8357 ;
  assign n8417 = n8416 ^ n8091 ;
  assign n8579 = n8578 ^ n8417 ;
  assign n8580 = n8578 ^ x87 ;
  assign n8581 = n8579 & n8580 ;
  assign n8582 = n8581 ^ x87 ;
  assign n8414 = n8260 & n8357 ;
  assign n8415 = n8414 ^ n8088 ;
  assign n8583 = n8582 ^ n8415 ;
  assign n8584 = n8582 ^ x88 ;
  assign n8585 = n8583 & n8584 ;
  assign n8586 = n8585 ^ x88 ;
  assign n8412 = n8264 & n8357 ;
  assign n8413 = n8412 ^ n8077 ;
  assign n8587 = n8586 ^ n8413 ;
  assign n8588 = n8586 ^ x89 ;
  assign n8589 = n8587 & n8588 ;
  assign n8590 = n8589 ^ x89 ;
  assign n8410 = n8268 & n8357 ;
  assign n8411 = n8410 ^ n8074 ;
  assign n8591 = n8590 ^ n8411 ;
  assign n8592 = n8590 ^ x90 ;
  assign n8593 = n8591 & n8592 ;
  assign n8594 = n8593 ^ x90 ;
  assign n8596 = n8594 ^ x91 ;
  assign n8360 = n8342 & n8357 ;
  assign n8361 = n8360 ^ n8028 ;
  assign n8362 = n8361 ^ x110 ;
  assign n8363 = n8338 & n8357 ;
  assign n8364 = n8363 ^ n8030 ;
  assign n8365 = n8364 ^ x109 ;
  assign n8653 = n8328 & n8357 ;
  assign n8654 = n8653 ^ n8038 ;
  assign n8372 = n8324 & n8357 ;
  assign n8373 = n8372 ^ n8040 ;
  assign n8374 = n8373 ^ x105 ;
  assign n8378 = n8373 ^ x104 ;
  assign n8375 = n8320 & n8357 ;
  assign n8376 = n8375 ^ n8042 ;
  assign n8377 = n8376 ^ n8373 ;
  assign n8379 = n8378 ^ n8377 ;
  assign n8408 = n8272 & n8357 ;
  assign n8409 = n8408 ^ n8072 ;
  assign n8595 = n8594 ^ n8409 ;
  assign n8597 = n8595 & n8596 ;
  assign n8598 = n8597 ^ x91 ;
  assign n8406 = n8276 & n8357 ;
  assign n8407 = n8406 ^ n8070 ;
  assign n8599 = n8598 ^ n8407 ;
  assign n8600 = n8598 ^ x92 ;
  assign n8601 = n8599 & n8600 ;
  assign n8602 = n8601 ^ x92 ;
  assign n8404 = n8280 & n8357 ;
  assign n8405 = n8404 ^ n8068 ;
  assign n8603 = n8602 ^ n8405 ;
  assign n8604 = n8602 ^ x93 ;
  assign n8605 = n8603 & n8604 ;
  assign n8606 = n8605 ^ x93 ;
  assign n8402 = n8284 & n8357 ;
  assign n8403 = n8402 ^ n8066 ;
  assign n8607 = n8606 ^ n8403 ;
  assign n8608 = n8606 ^ x94 ;
  assign n8609 = n8607 & n8608 ;
  assign n8610 = n8609 ^ x94 ;
  assign n8399 = n8286 ^ x94 ;
  assign n8400 = n8357 & n8399 ;
  assign n8401 = n8400 ^ n8063 ;
  assign n8611 = n8610 ^ n8401 ;
  assign n8612 = n8610 ^ x95 ;
  assign n8613 = n8611 & n8612 ;
  assign n8614 = n8613 ^ x95 ;
  assign n8396 = n8289 ^ x95 ;
  assign n8397 = n8357 & n8396 ;
  assign n8398 = n8397 ^ n8060 ;
  assign n8615 = n8614 ^ n8398 ;
  assign n8616 = n8614 ^ x96 ;
  assign n8617 = n8615 & n8616 ;
  assign n8618 = n8617 ^ x96 ;
  assign n8394 = n8294 & n8357 ;
  assign n8395 = n8394 ^ n8058 ;
  assign n8619 = n8618 ^ n8395 ;
  assign n8620 = n8618 ^ x97 ;
  assign n8621 = n8619 & n8620 ;
  assign n8622 = n8621 ^ x97 ;
  assign n8392 = n8298 & n8357 ;
  assign n8393 = n8392 ^ n8056 ;
  assign n8623 = n8622 ^ n8393 ;
  assign n8624 = n8622 ^ x98 ;
  assign n8625 = n8623 & n8624 ;
  assign n8626 = n8625 ^ x98 ;
  assign n8390 = n8302 & n8357 ;
  assign n8391 = n8390 ^ n8054 ;
  assign n8627 = n8626 ^ n8391 ;
  assign n8628 = n8626 ^ x99 ;
  assign n8629 = n8627 & n8628 ;
  assign n8630 = n8629 ^ x99 ;
  assign n8388 = n8306 & n8357 ;
  assign n8389 = n8388 ^ n8052 ;
  assign n8631 = n8630 ^ n8389 ;
  assign n8632 = n8630 ^ x100 ;
  assign n8633 = n8631 & n8632 ;
  assign n8634 = n8633 ^ x100 ;
  assign n8385 = n8308 ^ x100 ;
  assign n8386 = n8357 & n8385 ;
  assign n8387 = n8386 ^ n8049 ;
  assign n8635 = n8634 ^ n8387 ;
  assign n8636 = n8634 ^ x101 ;
  assign n8637 = n8635 & n8636 ;
  assign n8638 = n8637 ^ x101 ;
  assign n8382 = n8311 ^ x101 ;
  assign n8383 = n8357 & n8382 ;
  assign n8384 = n8383 ^ n8046 ;
  assign n8639 = n8638 ^ n8384 ;
  assign n8640 = n8638 ^ x102 ;
  assign n8641 = n8639 & n8640 ;
  assign n8642 = n8641 ^ x102 ;
  assign n8380 = n8316 & n8357 ;
  assign n8381 = n8380 ^ n8044 ;
  assign n8643 = n8642 ^ n8381 ;
  assign n8644 = n8642 ^ x103 ;
  assign n8645 = n8643 & n8644 ;
  assign n8646 = n8645 ^ x103 ;
  assign n8647 = n8646 ^ n8373 ;
  assign n8648 = n8647 ^ n8378 ;
  assign n8649 = ~n8379 & n8648 ;
  assign n8650 = n8649 ^ n8378 ;
  assign n8651 = ~n8374 & n8650 ;
  assign n8652 = n8651 ^ x105 ;
  assign n8655 = n8654 ^ n8652 ;
  assign n8656 = n8654 ^ x106 ;
  assign n8657 = n8655 & ~n8656 ;
  assign n8658 = n8657 ^ x106 ;
  assign n8369 = n8330 ^ x106 ;
  assign n8370 = n8357 & n8369 ;
  assign n8371 = n8370 ^ n8035 ;
  assign n8659 = n8658 ^ n8371 ;
  assign n8660 = n8658 ^ x107 ;
  assign n8661 = n8659 & n8660 ;
  assign n8662 = n8661 ^ x107 ;
  assign n8366 = n8333 ^ x107 ;
  assign n8367 = n8357 & n8366 ;
  assign n8368 = n8367 ^ n8032 ;
  assign n8663 = n8662 ^ n8368 ;
  assign n8664 = n8662 ^ x108 ;
  assign n8665 = n8663 & n8664 ;
  assign n8666 = n8665 ^ x108 ;
  assign n8667 = n8666 ^ n8364 ;
  assign n8668 = ~n8365 & n8667 ;
  assign n8669 = n8668 ^ x109 ;
  assign n8670 = n8669 ^ n8361 ;
  assign n8671 = ~n8362 & n8670 ;
  assign n8672 = n8671 ^ x110 ;
  assign n8358 = n8345 & n8357 ;
  assign n8359 = n8358 ^ n8350 ;
  assign n8674 = n8672 ^ n8359 ;
  assign n8673 = n8359 & ~n8672 ;
  assign n8675 = n8674 ^ n8673 ;
  assign n8676 = ~x111 & ~n8675 ;
  assign n8697 = n8676 ^ x111 ;
  assign n8689 = ~n8673 & ~n8676 ;
  assign n8698 = n8697 ^ n8689 ;
  assign n8699 = n8698 ^ n8697 ;
  assign n8700 = n8697 ^ n8353 ;
  assign n8701 = n8700 ^ n8697 ;
  assign n8702 = n8699 & ~n8701 ;
  assign n8703 = n8702 ^ n8697 ;
  assign n8704 = n8357 & ~n8703 ;
  assign n8705 = n8704 ^ n7681 ;
  assign n8696 = n8020 & n8689 ;
  assign n8706 = n8705 ^ n8696 ;
  assign n8688 = n7681 ^ n144 ;
  assign n8690 = n8689 ^ n8688 ;
  assign n8691 = n7681 ^ x112 ;
  assign n8692 = n8689 ^ x112 ;
  assign n8693 = ~n8691 & n8692 ;
  assign n8694 = n8693 ^ x112 ;
  assign n8695 = n8690 & ~n8694 ;
  assign n8707 = n8706 ^ n8695 ;
  assign n8948 = n8596 & n8707 ;
  assign n8949 = n8948 ^ n8409 ;
  assign n8762 = n8592 & n8707 ;
  assign n8763 = n8762 ^ n8411 ;
  assign n8764 = n8763 ^ x91 ;
  assign n8768 = n8763 ^ x90 ;
  assign n8765 = n8588 & n8707 ;
  assign n8766 = n8765 ^ n8413 ;
  assign n8767 = n8766 ^ n8763 ;
  assign n8769 = n8768 ^ n8767 ;
  assign n8770 = n8584 & n8707 ;
  assign n8771 = n8770 ^ n8415 ;
  assign n8772 = n8771 ^ x89 ;
  assign n8776 = n8771 ^ x88 ;
  assign n8773 = n8580 & n8707 ;
  assign n8774 = n8773 ^ n8417 ;
  assign n8775 = n8774 ^ n8771 ;
  assign n8777 = n8776 ^ n8775 ;
  assign n8780 = n8572 & n8707 ;
  assign n8781 = n8780 ^ n8421 ;
  assign n8782 = n8781 ^ x86 ;
  assign n8783 = n8568 & n8707 ;
  assign n8784 = n8783 ^ n8423 ;
  assign n8785 = n8784 ^ x85 ;
  assign n8896 = n8540 & n8707 ;
  assign n8897 = n8896 ^ n8439 ;
  assign n8809 = n8536 & n8707 ;
  assign n8810 = n8809 ^ n8441 ;
  assign n8811 = n8810 ^ x77 ;
  assign n8815 = n8810 ^ x76 ;
  assign n8812 = n8532 & n8707 ;
  assign n8813 = n8812 ^ n8443 ;
  assign n8814 = n8813 ^ n8810 ;
  assign n8816 = n8815 ^ n8814 ;
  assign n8836 = ~x14 & x64 ;
  assign n8837 = n8836 ^ x65 ;
  assign n8838 = x64 & n8707 ;
  assign n8839 = n8838 ^ x15 ;
  assign n8840 = n8839 ^ n8836 ;
  assign n8841 = n8837 & n8840 ;
  assign n8842 = n8841 ^ x65 ;
  assign n8843 = n8842 ^ x66 ;
  assign n8849 = x64 & n8357 ;
  assign n8845 = ~x15 & x64 ;
  assign n8846 = n8845 ^ x65 ;
  assign n8847 = n8707 & n8846 ;
  assign n8848 = n8847 ^ x16 ;
  assign n8850 = n8849 ^ n8848 ;
  assign n8851 = n8850 ^ n8842 ;
  assign n8852 = n8843 & n8851 ;
  assign n8853 = n8852 ^ x66 ;
  assign n8833 = n8495 ^ x66 ;
  assign n8834 = n8707 & n8833 ;
  assign n8835 = n8834 ^ n8481 ;
  assign n8854 = n8853 ^ n8835 ;
  assign n8855 = n8853 ^ x67 ;
  assign n8856 = n8854 & n8855 ;
  assign n8857 = n8856 ^ x67 ;
  assign n8831 = n8500 & n8707 ;
  assign n8832 = n8831 ^ n8477 ;
  assign n8858 = n8857 ^ n8832 ;
  assign n8859 = n8857 ^ x68 ;
  assign n8860 = n8858 & n8859 ;
  assign n8861 = n8860 ^ x68 ;
  assign n8829 = n8504 & n8707 ;
  assign n8830 = n8829 ^ n8461 ;
  assign n8862 = n8861 ^ n8830 ;
  assign n8863 = n8861 ^ x69 ;
  assign n8864 = n8862 & n8863 ;
  assign n8865 = n8864 ^ x69 ;
  assign n8827 = n8508 & n8707 ;
  assign n8828 = n8827 ^ n8458 ;
  assign n8866 = n8865 ^ n8828 ;
  assign n8867 = n8865 ^ x70 ;
  assign n8868 = n8866 & n8867 ;
  assign n8869 = n8868 ^ x70 ;
  assign n8825 = n8512 & n8707 ;
  assign n8826 = n8825 ^ n8455 ;
  assign n8870 = n8869 ^ n8826 ;
  assign n8871 = n8869 ^ x71 ;
  assign n8872 = n8870 & n8871 ;
  assign n8873 = n8872 ^ x71 ;
  assign n8823 = n8516 & n8707 ;
  assign n8824 = n8823 ^ n8452 ;
  assign n8874 = n8873 ^ n8824 ;
  assign n8875 = n8873 ^ x72 ;
  assign n8876 = n8874 & n8875 ;
  assign n8877 = n8876 ^ x72 ;
  assign n8821 = n8520 & n8707 ;
  assign n8822 = n8821 ^ n8449 ;
  assign n8878 = n8877 ^ n8822 ;
  assign n8879 = n8877 ^ x73 ;
  assign n8880 = n8878 & n8879 ;
  assign n8881 = n8880 ^ x73 ;
  assign n8819 = n8524 & n8707 ;
  assign n8820 = n8819 ^ n8447 ;
  assign n8882 = n8881 ^ n8820 ;
  assign n8883 = n8881 ^ x74 ;
  assign n8884 = n8882 & n8883 ;
  assign n8885 = n8884 ^ x74 ;
  assign n8817 = n8528 & n8707 ;
  assign n8818 = n8817 ^ n8445 ;
  assign n8886 = n8885 ^ n8818 ;
  assign n8887 = n8885 ^ x75 ;
  assign n8888 = n8886 & n8887 ;
  assign n8889 = n8888 ^ x75 ;
  assign n8890 = n8889 ^ n8810 ;
  assign n8891 = n8890 ^ n8815 ;
  assign n8892 = ~n8816 & n8891 ;
  assign n8893 = n8892 ^ n8815 ;
  assign n8894 = ~n8811 & n8893 ;
  assign n8895 = n8894 ^ x77 ;
  assign n8898 = n8897 ^ n8895 ;
  assign n8899 = n8897 ^ x78 ;
  assign n8900 = n8898 & ~n8899 ;
  assign n8901 = n8900 ^ x78 ;
  assign n8807 = n8544 & n8707 ;
  assign n8808 = n8807 ^ n8437 ;
  assign n8902 = n8901 ^ n8808 ;
  assign n8903 = n8901 ^ x79 ;
  assign n8904 = n8902 & n8903 ;
  assign n8905 = n8904 ^ x79 ;
  assign n8805 = n8548 & n8707 ;
  assign n8806 = n8805 ^ n8435 ;
  assign n8906 = n8905 ^ n8806 ;
  assign n8907 = n8905 ^ x80 ;
  assign n8908 = n8906 & n8907 ;
  assign n8909 = n8908 ^ x80 ;
  assign n8803 = n8552 & n8707 ;
  assign n8804 = n8803 ^ n8433 ;
  assign n8910 = n8909 ^ n8804 ;
  assign n8911 = n8909 ^ x81 ;
  assign n8912 = n8910 & n8911 ;
  assign n8913 = n8912 ^ x81 ;
  assign n8800 = n8554 ^ x81 ;
  assign n8801 = n8707 & n8800 ;
  assign n8802 = n8801 ^ n8428 ;
  assign n8914 = n8913 ^ n8802 ;
  assign n8915 = n8913 ^ x82 ;
  assign n8916 = n8914 & n8915 ;
  assign n8917 = n8916 ^ x82 ;
  assign n8789 = n8428 ^ x82 ;
  assign n8790 = n8789 ^ n8554 ;
  assign n8791 = n8790 ^ x81 ;
  assign n8792 = n8791 ^ n8789 ;
  assign n8794 = n8554 ^ x82 ;
  assign n8795 = n8794 ^ n8789 ;
  assign n8796 = ~n8792 & ~n8795 ;
  assign n8797 = n8796 ^ n8789 ;
  assign n8798 = n8707 & ~n8797 ;
  assign n8799 = n8798 ^ n8425 ;
  assign n8918 = n8917 ^ n8799 ;
  assign n8919 = n8917 ^ x83 ;
  assign n8920 = n8918 & n8919 ;
  assign n8921 = n8920 ^ x83 ;
  assign n8786 = n8560 ^ x83 ;
  assign n8787 = n8707 & n8786 ;
  assign n8788 = n8787 ^ n8562 ;
  assign n8922 = n8921 ^ n8788 ;
  assign n8923 = n8921 ^ x84 ;
  assign n8924 = n8922 & n8923 ;
  assign n8925 = n8924 ^ x84 ;
  assign n8926 = n8925 ^ n8784 ;
  assign n8927 = ~n8785 & n8926 ;
  assign n8928 = n8927 ^ x85 ;
  assign n8929 = n8928 ^ n8781 ;
  assign n8930 = ~n8782 & n8929 ;
  assign n8931 = n8930 ^ x86 ;
  assign n8778 = n8576 & n8707 ;
  assign n8779 = n8778 ^ n8419 ;
  assign n8932 = n8931 ^ n8779 ;
  assign n8933 = n8931 ^ x87 ;
  assign n8934 = n8932 & n8933 ;
  assign n8935 = n8934 ^ x87 ;
  assign n8936 = n8935 ^ n8771 ;
  assign n8937 = n8936 ^ n8776 ;
  assign n8938 = ~n8777 & n8937 ;
  assign n8939 = n8938 ^ n8776 ;
  assign n8940 = ~n8772 & n8939 ;
  assign n8941 = n8940 ^ x89 ;
  assign n8942 = n8941 ^ n8763 ;
  assign n8943 = n8942 ^ n8768 ;
  assign n8944 = ~n8769 & n8943 ;
  assign n8945 = n8944 ^ n8768 ;
  assign n8946 = ~n8764 & n8945 ;
  assign n8947 = n8946 ^ x91 ;
  assign n8950 = n8949 ^ n8947 ;
  assign n8951 = n8949 ^ x92 ;
  assign n8952 = n8950 & ~n8951 ;
  assign n8953 = n8952 ^ x92 ;
  assign n8760 = n8600 & n8707 ;
  assign n8761 = n8760 ^ n8407 ;
  assign n8954 = n8953 ^ n8761 ;
  assign n8955 = n8953 ^ x93 ;
  assign n8956 = n8954 & n8955 ;
  assign n8957 = n8956 ^ x93 ;
  assign n8758 = n8604 & n8707 ;
  assign n8759 = n8758 ^ n8405 ;
  assign n8958 = n8957 ^ n8759 ;
  assign n8959 = n8957 ^ x94 ;
  assign n8960 = n8958 & n8959 ;
  assign n8961 = n8960 ^ x94 ;
  assign n8756 = n8608 & n8707 ;
  assign n8757 = n8756 ^ n8403 ;
  assign n8962 = n8961 ^ n8757 ;
  assign n8963 = n8961 ^ x95 ;
  assign n8964 = n8962 & n8963 ;
  assign n8965 = n8964 ^ x95 ;
  assign n8967 = n8965 ^ x96 ;
  assign n141 = ~x114 & n140 ;
  assign n8754 = n8612 & n8707 ;
  assign n8755 = n8754 ^ n8401 ;
  assign n8966 = n8965 ^ n8755 ;
  assign n8968 = n8966 & n8967 ;
  assign n8969 = n8968 ^ x96 ;
  assign n8752 = n8616 & n8707 ;
  assign n8753 = n8752 ^ n8398 ;
  assign n8970 = n8969 ^ n8753 ;
  assign n8971 = n8969 ^ x97 ;
  assign n8972 = n8970 & n8971 ;
  assign n8973 = n8972 ^ x97 ;
  assign n8750 = n8620 & n8707 ;
  assign n8751 = n8750 ^ n8395 ;
  assign n8974 = n8973 ^ n8751 ;
  assign n8975 = n8973 ^ x98 ;
  assign n8976 = n8974 & n8975 ;
  assign n8977 = n8976 ^ x98 ;
  assign n8748 = n8624 & n8707 ;
  assign n8749 = n8748 ^ n8393 ;
  assign n8978 = n8977 ^ n8749 ;
  assign n8979 = n8977 ^ x99 ;
  assign n8980 = n8978 & n8979 ;
  assign n8981 = n8980 ^ x99 ;
  assign n8746 = n8628 & n8707 ;
  assign n8747 = n8746 ^ n8391 ;
  assign n8982 = n8981 ^ n8747 ;
  assign n8983 = n8981 ^ x100 ;
  assign n8984 = n8982 & n8983 ;
  assign n8985 = n8984 ^ x100 ;
  assign n8744 = n8632 & n8707 ;
  assign n8745 = n8744 ^ n8389 ;
  assign n8986 = n8985 ^ n8745 ;
  assign n8987 = n8985 ^ x101 ;
  assign n8988 = n8986 & n8987 ;
  assign n8989 = n8988 ^ x101 ;
  assign n8742 = n8636 & n8707 ;
  assign n8743 = n8742 ^ n8387 ;
  assign n8990 = n8989 ^ n8743 ;
  assign n8991 = n8989 ^ x102 ;
  assign n8992 = n8990 & n8991 ;
  assign n8993 = n8992 ^ x102 ;
  assign n8740 = n8640 & n8707 ;
  assign n8741 = n8740 ^ n8384 ;
  assign n8994 = n8993 ^ n8741 ;
  assign n8995 = n8993 ^ x103 ;
  assign n8996 = n8994 & n8995 ;
  assign n8997 = n8996 ^ x103 ;
  assign n8738 = n8644 & n8707 ;
  assign n8739 = n8738 ^ n8381 ;
  assign n8998 = n8997 ^ n8739 ;
  assign n8999 = n8997 ^ x104 ;
  assign n9000 = n8998 & n8999 ;
  assign n9001 = n9000 ^ x104 ;
  assign n8735 = n8646 ^ x104 ;
  assign n8736 = n8707 & n8735 ;
  assign n8737 = n8736 ^ n8376 ;
  assign n9002 = n9001 ^ n8737 ;
  assign n9003 = n9001 ^ x105 ;
  assign n9004 = n9002 & n9003 ;
  assign n9005 = n9004 ^ x105 ;
  assign n8724 = n8376 ^ x105 ;
  assign n8725 = n8724 ^ n8646 ;
  assign n8726 = n8725 ^ x104 ;
  assign n8727 = n8726 ^ n8724 ;
  assign n8729 = n8646 ^ x105 ;
  assign n8730 = n8729 ^ n8724 ;
  assign n8731 = ~n8727 & ~n8730 ;
  assign n8732 = n8731 ^ n8724 ;
  assign n8733 = n8707 & ~n8732 ;
  assign n8734 = n8733 ^ n8373 ;
  assign n9006 = n9005 ^ n8734 ;
  assign n9007 = n9005 ^ x106 ;
  assign n9008 = n9006 & n9007 ;
  assign n9009 = n9008 ^ x106 ;
  assign n8721 = n8652 ^ x106 ;
  assign n8722 = n8707 & n8721 ;
  assign n8723 = n8722 ^ n8654 ;
  assign n9010 = n9009 ^ n8723 ;
  assign n9011 = n9009 ^ x107 ;
  assign n9012 = n9010 & n9011 ;
  assign n9013 = n9012 ^ x107 ;
  assign n8719 = n8660 & n8707 ;
  assign n8720 = n8719 ^ n8371 ;
  assign n9014 = n9013 ^ n8720 ;
  assign n9015 = n9013 ^ x108 ;
  assign n9016 = n9014 & n9015 ;
  assign n9017 = n9016 ^ x108 ;
  assign n8717 = n8664 & n8707 ;
  assign n8718 = n8717 ^ n8368 ;
  assign n9018 = n9017 ^ n8718 ;
  assign n9019 = n9017 ^ x109 ;
  assign n9020 = n9018 & n9019 ;
  assign n9021 = n9020 ^ x109 ;
  assign n8714 = n8666 ^ x109 ;
  assign n8715 = n8707 & n8714 ;
  assign n8716 = n8715 ^ n8364 ;
  assign n9022 = n9021 ^ n8716 ;
  assign n9023 = n9021 ^ x110 ;
  assign n9024 = n9022 & n9023 ;
  assign n9025 = n9024 ^ x110 ;
  assign n8711 = n8669 ^ x110 ;
  assign n8712 = n8707 & n8711 ;
  assign n8713 = n8712 ^ n8361 ;
  assign n9026 = n9025 ^ n8713 ;
  assign n9027 = n9025 ^ x111 ;
  assign n9028 = n9026 & n9027 ;
  assign n9029 = n9028 ^ x111 ;
  assign n8708 = n8672 ^ x111 ;
  assign n8709 = n8707 & n8708 ;
  assign n8710 = n8709 ^ n8359 ;
  assign n9030 = n9029 ^ n8710 ;
  assign n9033 = n8710 ^ x112 ;
  assign n9034 = n9030 & ~n9033 ;
  assign n9031 = x113 ^ x112 ;
  assign n9035 = n9034 ^ n9031 ;
  assign n8677 = n8676 ^ x112 ;
  assign n8678 = n144 & n8677 ;
  assign n8679 = n8673 ^ n8353 ;
  assign n8682 = ~n8676 & n8679 ;
  assign n8683 = n8682 ^ n8353 ;
  assign n8684 = n8678 & ~n8683 ;
  assign n8685 = n8684 ^ n144 ;
  assign n8686 = n8020 & ~n8685 ;
  assign n9040 = n8686 ^ x113 ;
  assign n9043 = n9035 & ~n9040 ;
  assign n9044 = n9043 ^ x113 ;
  assign n9045 = n141 & ~n9044 ;
  assign n9080 = n8967 & n9045 ;
  assign n9081 = n9080 ^ n8755 ;
  assign n9082 = n9081 ^ x97 ;
  assign n9083 = n8963 & n9045 ;
  assign n9084 = n9083 ^ n8757 ;
  assign n9085 = n9084 ^ x96 ;
  assign n9306 = n8925 ^ x85 ;
  assign n9307 = n9045 & n9306 ;
  assign n9308 = n9307 ^ n8784 ;
  assign n9126 = n8923 & n9045 ;
  assign n9127 = n9126 ^ n8788 ;
  assign n9128 = n9127 ^ x85 ;
  assign n9132 = n9127 ^ x84 ;
  assign n9129 = n8919 & n9045 ;
  assign n9130 = n9129 ^ n8799 ;
  assign n9131 = n9130 ^ n9127 ;
  assign n9133 = n9132 ^ n9131 ;
  assign n9230 = n8843 & n9045 ;
  assign n9231 = n9230 ^ n8850 ;
  assign n9187 = x64 ^ x14 ;
  assign n9188 = n191 & n9187 ;
  assign n9184 = n191 ^ x13 ;
  assign n9185 = x64 & n8839 ;
  assign n9186 = n9184 & n9185 ;
  assign n9189 = n9188 ^ n9186 ;
  assign n9190 = n9045 & n9189 ;
  assign n9177 = x14 & ~x65 ;
  assign n9178 = ~x13 & x64 ;
  assign n9179 = ~n9177 & n9178 ;
  assign n9180 = x65 ^ x14 ;
  assign n9181 = n9180 ^ n9177 ;
  assign n9182 = n8839 & ~n9181 ;
  assign n9183 = ~n9179 & n9182 ;
  assign n9191 = n9190 ^ n9183 ;
  assign n9192 = n9045 ^ n8839 ;
  assign n9193 = n9192 ^ n9179 ;
  assign n9194 = n9193 ^ x66 ;
  assign n9195 = x64 & n9045 ;
  assign n9196 = n9181 & ~n9195 ;
  assign n9197 = n9196 ^ n9179 ;
  assign n9198 = n9197 ^ x66 ;
  assign n9199 = n9196 ^ n9045 ;
  assign n9200 = n9199 ^ n9192 ;
  assign n9201 = n9198 & ~n9200 ;
  assign n9202 = n9194 & n9201 ;
  assign n9203 = n9202 ^ n9196 ;
  assign n9204 = n9203 ^ n9192 ;
  assign n9205 = ~x66 & n9204 ;
  assign n9206 = ~n9192 & n9205 ;
  assign n9207 = n9206 ^ x66 ;
  assign n9208 = n9180 ^ n8839 ;
  assign n9209 = n8839 ^ x13 ;
  assign n9210 = n9209 ^ n9045 ;
  assign n9211 = x65 ^ x13 ;
  assign n9212 = n9211 ^ n9045 ;
  assign n9213 = ~n9210 & n9212 ;
  assign n9214 = n9213 ^ n9045 ;
  assign n9215 = n9208 & n9214 ;
  assign n9216 = x64 & n9215 ;
  assign n9217 = ~n9207 & n9216 ;
  assign n9218 = n9217 ^ n9207 ;
  assign n9219 = n9218 ^ x13 ;
  assign n9220 = n9219 ^ n9218 ;
  assign n9225 = ~x65 & n9217 ;
  assign n9226 = n9220 & n9225 ;
  assign n9227 = n9226 ^ n9220 ;
  assign n9228 = n9227 ^ n9219 ;
  assign n9229 = ~n9191 & n9228 ;
  assign n9232 = n9231 ^ n9229 ;
  assign n9233 = n9231 ^ x67 ;
  assign n9234 = n9232 & ~n9233 ;
  assign n9235 = n9234 ^ x67 ;
  assign n9175 = n8855 & n9045 ;
  assign n9176 = n9175 ^ n8835 ;
  assign n9236 = n9235 ^ n9176 ;
  assign n9237 = n9235 ^ x68 ;
  assign n9238 = n9236 & n9237 ;
  assign n9239 = n9238 ^ x68 ;
  assign n9173 = n8859 & n9045 ;
  assign n9174 = n9173 ^ n8832 ;
  assign n9240 = n9239 ^ n9174 ;
  assign n9241 = n9239 ^ x69 ;
  assign n9242 = n9240 & n9241 ;
  assign n9243 = n9242 ^ x69 ;
  assign n9171 = n8863 & n9045 ;
  assign n9172 = n9171 ^ n8830 ;
  assign n9244 = n9243 ^ n9172 ;
  assign n9245 = n9243 ^ x70 ;
  assign n9246 = n9244 & n9245 ;
  assign n9247 = n9246 ^ x70 ;
  assign n9169 = n8867 & n9045 ;
  assign n9170 = n9169 ^ n8828 ;
  assign n9248 = n9247 ^ n9170 ;
  assign n9249 = n9247 ^ x71 ;
  assign n9250 = n9248 & n9249 ;
  assign n9251 = n9250 ^ x71 ;
  assign n9167 = n8871 & n9045 ;
  assign n9168 = n9167 ^ n8826 ;
  assign n9252 = n9251 ^ n9168 ;
  assign n9253 = n9251 ^ x72 ;
  assign n9254 = n9252 & n9253 ;
  assign n9255 = n9254 ^ x72 ;
  assign n9165 = n8875 & n9045 ;
  assign n9166 = n9165 ^ n8824 ;
  assign n9256 = n9255 ^ n9166 ;
  assign n9257 = n9255 ^ x73 ;
  assign n9258 = n9256 & n9257 ;
  assign n9259 = n9258 ^ x73 ;
  assign n9163 = n8879 & n9045 ;
  assign n9164 = n9163 ^ n8822 ;
  assign n9260 = n9259 ^ n9164 ;
  assign n9261 = n9259 ^ x74 ;
  assign n9262 = n9260 & n9261 ;
  assign n9263 = n9262 ^ x74 ;
  assign n9161 = n8883 & n9045 ;
  assign n9162 = n9161 ^ n8820 ;
  assign n9264 = n9263 ^ n9162 ;
  assign n9265 = n9263 ^ x75 ;
  assign n9266 = n9264 & n9265 ;
  assign n9267 = n9266 ^ x75 ;
  assign n9159 = n8887 & n9045 ;
  assign n9160 = n9159 ^ n8818 ;
  assign n9268 = n9267 ^ n9160 ;
  assign n9269 = n9267 ^ x76 ;
  assign n9270 = n9268 & n9269 ;
  assign n9271 = n9270 ^ x76 ;
  assign n9156 = n8889 ^ x76 ;
  assign n9157 = n9045 & n9156 ;
  assign n9158 = n9157 ^ n8813 ;
  assign n9272 = n9271 ^ n9158 ;
  assign n9273 = n9271 ^ x77 ;
  assign n9274 = n9272 & n9273 ;
  assign n9275 = n9274 ^ x77 ;
  assign n9145 = n8813 ^ x77 ;
  assign n9146 = n9145 ^ n8889 ;
  assign n9147 = n9146 ^ x76 ;
  assign n9148 = n9147 ^ n9145 ;
  assign n9150 = n8889 ^ x77 ;
  assign n9151 = n9150 ^ n9145 ;
  assign n9152 = ~n9148 & ~n9151 ;
  assign n9153 = n9152 ^ n9145 ;
  assign n9154 = n9045 & ~n9153 ;
  assign n9155 = n9154 ^ n8810 ;
  assign n9276 = n9275 ^ n9155 ;
  assign n9277 = n9275 ^ x78 ;
  assign n9278 = n9276 & n9277 ;
  assign n9279 = n9278 ^ x78 ;
  assign n9142 = n8895 ^ x78 ;
  assign n9143 = n9045 & n9142 ;
  assign n9144 = n9143 ^ n8897 ;
  assign n9280 = n9279 ^ n9144 ;
  assign n9281 = n9279 ^ x79 ;
  assign n9282 = n9280 & n9281 ;
  assign n9283 = n9282 ^ x79 ;
  assign n9140 = n8903 & n9045 ;
  assign n9141 = n9140 ^ n8808 ;
  assign n9284 = n9283 ^ n9141 ;
  assign n9285 = n9283 ^ x80 ;
  assign n9286 = n9284 & n9285 ;
  assign n9287 = n9286 ^ x80 ;
  assign n9138 = n8907 & n9045 ;
  assign n9139 = n9138 ^ n8806 ;
  assign n9288 = n9287 ^ n9139 ;
  assign n9289 = n9287 ^ x81 ;
  assign n9290 = n9288 & n9289 ;
  assign n9291 = n9290 ^ x81 ;
  assign n9136 = n8911 & n9045 ;
  assign n9137 = n9136 ^ n8804 ;
  assign n9292 = n9291 ^ n9137 ;
  assign n9293 = n9291 ^ x82 ;
  assign n9294 = n9292 & n9293 ;
  assign n9295 = n9294 ^ x82 ;
  assign n9134 = n8915 & n9045 ;
  assign n9135 = n9134 ^ n8802 ;
  assign n9296 = n9295 ^ n9135 ;
  assign n9297 = n9295 ^ x83 ;
  assign n9298 = n9296 & n9297 ;
  assign n9299 = n9298 ^ x83 ;
  assign n9300 = n9299 ^ n9127 ;
  assign n9301 = n9300 ^ n9132 ;
  assign n9302 = ~n9133 & n9301 ;
  assign n9303 = n9302 ^ n9132 ;
  assign n9304 = ~n9128 & n9303 ;
  assign n9305 = n9304 ^ x85 ;
  assign n9309 = n9308 ^ n9305 ;
  assign n9310 = n9308 ^ x86 ;
  assign n9311 = n9309 & ~n9310 ;
  assign n9312 = n9311 ^ x86 ;
  assign n9123 = n8928 ^ x86 ;
  assign n9124 = n9045 & n9123 ;
  assign n9125 = n9124 ^ n8781 ;
  assign n9313 = n9312 ^ n9125 ;
  assign n9314 = n9312 ^ x87 ;
  assign n9315 = n9313 & n9314 ;
  assign n9316 = n9315 ^ x87 ;
  assign n9121 = n8933 & n9045 ;
  assign n9122 = n9121 ^ n8779 ;
  assign n9317 = n9316 ^ n9122 ;
  assign n9318 = n9316 ^ x88 ;
  assign n9319 = n9317 & n9318 ;
  assign n9320 = n9319 ^ x88 ;
  assign n9118 = n8935 ^ x88 ;
  assign n9119 = n9045 & n9118 ;
  assign n9120 = n9119 ^ n8774 ;
  assign n9321 = n9320 ^ n9120 ;
  assign n9322 = n9320 ^ x89 ;
  assign n9323 = n9321 & n9322 ;
  assign n9324 = n9323 ^ x89 ;
  assign n9107 = n8774 ^ x89 ;
  assign n9108 = n9107 ^ n8935 ;
  assign n9109 = n9108 ^ x88 ;
  assign n9110 = n9109 ^ n9107 ;
  assign n9112 = n8935 ^ x89 ;
  assign n9113 = n9112 ^ n9107 ;
  assign n9114 = ~n9110 & ~n9113 ;
  assign n9115 = n9114 ^ n9107 ;
  assign n9116 = n9045 & ~n9115 ;
  assign n9117 = n9116 ^ n8771 ;
  assign n9325 = n9324 ^ n9117 ;
  assign n9326 = n9324 ^ x90 ;
  assign n9327 = n9325 & n9326 ;
  assign n9328 = n9327 ^ x90 ;
  assign n9104 = n8941 ^ x90 ;
  assign n9105 = n9045 & n9104 ;
  assign n9106 = n9105 ^ n8766 ;
  assign n9329 = n9328 ^ n9106 ;
  assign n9330 = n9328 ^ x91 ;
  assign n9331 = n9329 & n9330 ;
  assign n9332 = n9331 ^ x91 ;
  assign n9093 = n8766 ^ x91 ;
  assign n9094 = n9093 ^ n8941 ;
  assign n9095 = n9094 ^ x90 ;
  assign n9096 = n9095 ^ n9093 ;
  assign n9098 = n8941 ^ x91 ;
  assign n9099 = n9098 ^ n9093 ;
  assign n9100 = ~n9096 & ~n9099 ;
  assign n9101 = n9100 ^ n9093 ;
  assign n9102 = n9045 & ~n9101 ;
  assign n9103 = n9102 ^ n8763 ;
  assign n9333 = n9332 ^ n9103 ;
  assign n9334 = n9332 ^ x92 ;
  assign n9335 = n9333 & n9334 ;
  assign n9336 = n9335 ^ x92 ;
  assign n9090 = n8947 ^ x92 ;
  assign n9091 = n9045 & n9090 ;
  assign n9092 = n9091 ^ n8949 ;
  assign n9337 = n9336 ^ n9092 ;
  assign n9338 = n9336 ^ x93 ;
  assign n9339 = n9337 & n9338 ;
  assign n9340 = n9339 ^ x93 ;
  assign n9088 = n8955 & n9045 ;
  assign n9089 = n9088 ^ n8761 ;
  assign n9341 = n9340 ^ n9089 ;
  assign n9342 = n9340 ^ x94 ;
  assign n9343 = n9341 & n9342 ;
  assign n9344 = n9343 ^ x94 ;
  assign n9086 = n8959 & n9045 ;
  assign n9087 = n9086 ^ n8759 ;
  assign n9345 = n9344 ^ n9087 ;
  assign n9346 = n9344 ^ x95 ;
  assign n9347 = n9345 & n9346 ;
  assign n9348 = n9347 ^ x95 ;
  assign n9349 = n9348 ^ n9084 ;
  assign n9350 = ~n9085 & n9349 ;
  assign n9351 = n9350 ^ x96 ;
  assign n9352 = n9351 ^ n9081 ;
  assign n9353 = ~n9082 & n9352 ;
  assign n9354 = n9353 ^ x97 ;
  assign n9078 = n8971 & n9045 ;
  assign n9079 = n9078 ^ n8753 ;
  assign n9355 = n9354 ^ n9079 ;
  assign n9356 = n9354 ^ x98 ;
  assign n9357 = n9355 & n9356 ;
  assign n9358 = n9357 ^ x98 ;
  assign n9076 = n8975 & n9045 ;
  assign n9077 = n9076 ^ n8751 ;
  assign n9359 = n9358 ^ n9077 ;
  assign n9360 = n9358 ^ x99 ;
  assign n9361 = n9359 & n9360 ;
  assign n9362 = n9361 ^ x99 ;
  assign n9074 = n8979 & n9045 ;
  assign n9075 = n9074 ^ n8749 ;
  assign n9363 = n9362 ^ n9075 ;
  assign n9364 = n9362 ^ x100 ;
  assign n9365 = n9363 & n9364 ;
  assign n9366 = n9365 ^ x100 ;
  assign n9368 = n9366 ^ x101 ;
  assign n9393 = n9011 & n9045 ;
  assign n9394 = n9393 ^ n8723 ;
  assign n9056 = n9007 & n9045 ;
  assign n9057 = n9056 ^ n8734 ;
  assign n9058 = n9057 ^ x107 ;
  assign n9062 = n9057 ^ x106 ;
  assign n9059 = n9003 & n9045 ;
  assign n9060 = n9059 ^ n8737 ;
  assign n9061 = n9060 ^ n9057 ;
  assign n9063 = n9062 ^ n9061 ;
  assign n9072 = n8983 & n9045 ;
  assign n9073 = n9072 ^ n8747 ;
  assign n9367 = n9366 ^ n9073 ;
  assign n9369 = n9367 & n9368 ;
  assign n9370 = n9369 ^ x101 ;
  assign n9070 = n8987 & n9045 ;
  assign n9071 = n9070 ^ n8745 ;
  assign n9371 = n9370 ^ n9071 ;
  assign n9372 = n9370 ^ x102 ;
  assign n9373 = n9371 & n9372 ;
  assign n9374 = n9373 ^ x102 ;
  assign n9068 = n8991 & n9045 ;
  assign n9069 = n9068 ^ n8743 ;
  assign n9375 = n9374 ^ n9069 ;
  assign n9376 = n9374 ^ x103 ;
  assign n9377 = n9375 & n9376 ;
  assign n9378 = n9377 ^ x103 ;
  assign n9066 = n8995 & n9045 ;
  assign n9067 = n9066 ^ n8741 ;
  assign n9379 = n9378 ^ n9067 ;
  assign n9380 = n9378 ^ x104 ;
  assign n9381 = n9379 & n9380 ;
  assign n9382 = n9381 ^ x104 ;
  assign n9064 = n8999 & n9045 ;
  assign n9065 = n9064 ^ n8739 ;
  assign n9383 = n9382 ^ n9065 ;
  assign n9384 = n9382 ^ x105 ;
  assign n9385 = n9383 & n9384 ;
  assign n9386 = n9385 ^ x105 ;
  assign n9387 = n9386 ^ n9057 ;
  assign n9388 = n9387 ^ n9062 ;
  assign n9389 = ~n9063 & n9388 ;
  assign n9390 = n9389 ^ n9062 ;
  assign n9391 = ~n9058 & n9390 ;
  assign n9392 = n9391 ^ x107 ;
  assign n9395 = n9394 ^ n9392 ;
  assign n9396 = n9394 ^ x108 ;
  assign n9397 = n9395 & ~n9396 ;
  assign n9398 = n9397 ^ x108 ;
  assign n9054 = n9015 & n9045 ;
  assign n9055 = n9054 ^ n8720 ;
  assign n9399 = n9398 ^ n9055 ;
  assign n9400 = n9398 ^ x109 ;
  assign n9401 = n9399 & n9400 ;
  assign n9402 = n9401 ^ x109 ;
  assign n9052 = n9019 & n9045 ;
  assign n9053 = n9052 ^ n8718 ;
  assign n9403 = n9402 ^ n9053 ;
  assign n9404 = n9402 ^ x110 ;
  assign n9405 = n9403 & n9404 ;
  assign n9406 = n9405 ^ x110 ;
  assign n9050 = n9023 & n9045 ;
  assign n9051 = n9050 ^ n8716 ;
  assign n9407 = n9406 ^ n9051 ;
  assign n9408 = n9406 ^ x111 ;
  assign n9409 = n9407 & n9408 ;
  assign n9410 = n9409 ^ x111 ;
  assign n9048 = n9027 & n9045 ;
  assign n9049 = n9048 ^ n8713 ;
  assign n9411 = n9410 ^ n9049 ;
  assign n9412 = n9410 ^ x112 ;
  assign n9413 = n9411 & n9412 ;
  assign n9414 = n9413 ^ x112 ;
  assign n9039 = n9029 ^ x112 ;
  assign n9046 = n9039 & n9045 ;
  assign n9047 = n9046 ^ n8710 ;
  assign n9415 = n9414 ^ n9047 ;
  assign n9418 = n9047 ^ x113 ;
  assign n9419 = n9415 & ~n9418 ;
  assign n9416 = x114 ^ x113 ;
  assign n9420 = n9419 ^ n9416 ;
  assign n8687 = n141 & n8686 ;
  assign n9036 = n8687 & n9035 ;
  assign n9037 = n9036 ^ n8686 ;
  assign n9423 = n9037 ^ x114 ;
  assign n9426 = n9420 & ~n9423 ;
  assign n9427 = n9426 ^ x114 ;
  assign n9428 = n140 & ~n9427 ;
  assign n9724 = n9368 & n9428 ;
  assign n9725 = n9724 ^ n9073 ;
  assign n9462 = n9364 & n9428 ;
  assign n9463 = n9462 ^ n9075 ;
  assign n9464 = n9463 ^ x101 ;
  assign n9468 = n9463 ^ x100 ;
  assign n9465 = n9360 & n9428 ;
  assign n9466 = n9465 ^ n9077 ;
  assign n9467 = n9466 ^ n9463 ;
  assign n9469 = n9468 ^ n9467 ;
  assign n9624 = n9269 & n9428 ;
  assign n9625 = n9624 ^ n9160 ;
  assign n9527 = n9265 & n9428 ;
  assign n9528 = n9527 ^ n9162 ;
  assign n9529 = n9528 ^ x76 ;
  assign n9533 = n9528 ^ x75 ;
  assign n9530 = n9261 & n9428 ;
  assign n9531 = n9530 ^ n9164 ;
  assign n9532 = n9531 ^ n9528 ;
  assign n9534 = n9533 ^ n9532 ;
  assign n9551 = n9178 ^ x65 ;
  assign n9552 = n9428 & n9551 ;
  assign n9550 = n9195 ^ x14 ;
  assign n9553 = n9552 ^ n9550 ;
  assign n9554 = n9553 ^ x66 ;
  assign n9562 = x13 & x65 ;
  assign n9559 = x65 ^ x12 ;
  assign n9555 = x64 ^ x13 ;
  assign n9556 = n9555 ^ x65 ;
  assign n9560 = n9556 ^ n9428 ;
  assign n9561 = ~n9559 & n9560 ;
  assign n9563 = n9562 ^ n9561 ;
  assign n9564 = x64 & n9563 ;
  assign n9565 = n9564 ^ n9562 ;
  assign n9566 = n9565 ^ x65 ;
  assign n9567 = n9566 ^ n9553 ;
  assign n9568 = ~n9554 & n9567 ;
  assign n9569 = n9568 ^ x66 ;
  assign n9570 = n9569 ^ x67 ;
  assign n9580 = x14 & x65 ;
  assign n9572 = n9187 ^ x65 ;
  assign n9573 = n9572 ^ n9045 ;
  assign n9574 = ~n9211 & n9573 ;
  assign n9581 = n9580 ^ n9574 ;
  assign n9582 = ~x64 & n9581 ;
  assign n9577 = n9574 ^ n6836 ;
  assign n9583 = n9582 ^ n9577 ;
  assign n9584 = n9428 & n9583 ;
  assign n9585 = n9584 ^ n8839 ;
  assign n9571 = n8837 & n9045 ;
  assign n9586 = n9585 ^ n9571 ;
  assign n9587 = n9586 ^ n9569 ;
  assign n9588 = n9570 & n9587 ;
  assign n9589 = n9588 ^ x67 ;
  assign n9547 = n9229 ^ x67 ;
  assign n9548 = n9428 & n9547 ;
  assign n9549 = n9548 ^ n9231 ;
  assign n9590 = n9589 ^ n9549 ;
  assign n9591 = n9589 ^ x68 ;
  assign n9592 = n9590 & n9591 ;
  assign n9593 = n9592 ^ x68 ;
  assign n9545 = n9237 & n9428 ;
  assign n9546 = n9545 ^ n9176 ;
  assign n9594 = n9593 ^ n9546 ;
  assign n9595 = n9593 ^ x69 ;
  assign n9596 = n9594 & n9595 ;
  assign n9597 = n9596 ^ x69 ;
  assign n9543 = n9241 & n9428 ;
  assign n9544 = n9543 ^ n9174 ;
  assign n9598 = n9597 ^ n9544 ;
  assign n9599 = n9597 ^ x70 ;
  assign n9600 = n9598 & n9599 ;
  assign n9601 = n9600 ^ x70 ;
  assign n9541 = n9245 & n9428 ;
  assign n9542 = n9541 ^ n9172 ;
  assign n9602 = n9601 ^ n9542 ;
  assign n9603 = n9601 ^ x71 ;
  assign n9604 = n9602 & n9603 ;
  assign n9605 = n9604 ^ x71 ;
  assign n9539 = n9249 & n9428 ;
  assign n9540 = n9539 ^ n9170 ;
  assign n9606 = n9605 ^ n9540 ;
  assign n9607 = n9605 ^ x72 ;
  assign n9608 = n9606 & n9607 ;
  assign n9609 = n9608 ^ x72 ;
  assign n9537 = n9253 & n9428 ;
  assign n9538 = n9537 ^ n9168 ;
  assign n9610 = n9609 ^ n9538 ;
  assign n9611 = n9609 ^ x73 ;
  assign n9612 = n9610 & n9611 ;
  assign n9613 = n9612 ^ x73 ;
  assign n9535 = n9257 & n9428 ;
  assign n9536 = n9535 ^ n9166 ;
  assign n9614 = n9613 ^ n9536 ;
  assign n9615 = n9613 ^ x74 ;
  assign n9616 = n9614 & n9615 ;
  assign n9617 = n9616 ^ x74 ;
  assign n9618 = n9617 ^ n9528 ;
  assign n9619 = n9618 ^ n9533 ;
  assign n9620 = ~n9534 & n9619 ;
  assign n9621 = n9620 ^ n9533 ;
  assign n9622 = ~n9529 & n9621 ;
  assign n9623 = n9622 ^ x76 ;
  assign n9626 = n9625 ^ n9623 ;
  assign n9627 = n9625 ^ x77 ;
  assign n9628 = n9626 & ~n9627 ;
  assign n9629 = n9628 ^ x77 ;
  assign n9525 = n9273 & n9428 ;
  assign n9526 = n9525 ^ n9158 ;
  assign n9630 = n9629 ^ n9526 ;
  assign n9631 = n9629 ^ x78 ;
  assign n9632 = n9630 & n9631 ;
  assign n9633 = n9632 ^ x78 ;
  assign n9523 = n9277 & n9428 ;
  assign n9524 = n9523 ^ n9155 ;
  assign n9634 = n9633 ^ n9524 ;
  assign n9635 = n9633 ^ x79 ;
  assign n9636 = n9634 & n9635 ;
  assign n9637 = n9636 ^ x79 ;
  assign n9521 = n9281 & n9428 ;
  assign n9522 = n9521 ^ n9144 ;
  assign n9638 = n9637 ^ n9522 ;
  assign n9639 = n9637 ^ x80 ;
  assign n9640 = n9638 & n9639 ;
  assign n9641 = n9640 ^ x80 ;
  assign n9519 = n9285 & n9428 ;
  assign n9520 = n9519 ^ n9141 ;
  assign n9642 = n9641 ^ n9520 ;
  assign n9643 = n9641 ^ x81 ;
  assign n9644 = n9642 & n9643 ;
  assign n9645 = n9644 ^ x81 ;
  assign n9517 = n9289 & n9428 ;
  assign n9518 = n9517 ^ n9139 ;
  assign n9646 = n9645 ^ n9518 ;
  assign n9647 = n9645 ^ x82 ;
  assign n9648 = n9646 & n9647 ;
  assign n9649 = n9648 ^ x82 ;
  assign n9515 = n9293 & n9428 ;
  assign n9516 = n9515 ^ n9137 ;
  assign n9650 = n9649 ^ n9516 ;
  assign n9651 = n9649 ^ x83 ;
  assign n9652 = n9650 & n9651 ;
  assign n9653 = n9652 ^ x83 ;
  assign n9513 = n9297 & n9428 ;
  assign n9514 = n9513 ^ n9135 ;
  assign n9654 = n9653 ^ n9514 ;
  assign n9655 = n9653 ^ x84 ;
  assign n9656 = n9654 & n9655 ;
  assign n9657 = n9656 ^ x84 ;
  assign n9510 = n9299 ^ x84 ;
  assign n9511 = n9428 & n9510 ;
  assign n9512 = n9511 ^ n9130 ;
  assign n9658 = n9657 ^ n9512 ;
  assign n9659 = n9657 ^ x85 ;
  assign n9660 = n9658 & n9659 ;
  assign n9661 = n9660 ^ x85 ;
  assign n9499 = n9130 ^ x85 ;
  assign n9500 = n9499 ^ n9299 ;
  assign n9501 = n9500 ^ x84 ;
  assign n9502 = n9501 ^ n9499 ;
  assign n9504 = n9299 ^ x85 ;
  assign n9505 = n9504 ^ n9499 ;
  assign n9506 = ~n9502 & ~n9505 ;
  assign n9507 = n9506 ^ n9499 ;
  assign n9508 = n9428 & ~n9507 ;
  assign n9509 = n9508 ^ n9127 ;
  assign n9662 = n9661 ^ n9509 ;
  assign n9663 = n9661 ^ x86 ;
  assign n9664 = n9662 & n9663 ;
  assign n9665 = n9664 ^ x86 ;
  assign n9496 = n9305 ^ x86 ;
  assign n9497 = n9428 & n9496 ;
  assign n9498 = n9497 ^ n9308 ;
  assign n9666 = n9665 ^ n9498 ;
  assign n9667 = n9665 ^ x87 ;
  assign n9668 = n9666 & n9667 ;
  assign n9669 = n9668 ^ x87 ;
  assign n9494 = n9314 & n9428 ;
  assign n9495 = n9494 ^ n9125 ;
  assign n9670 = n9669 ^ n9495 ;
  assign n9671 = n9669 ^ x88 ;
  assign n9672 = n9670 & n9671 ;
  assign n9673 = n9672 ^ x88 ;
  assign n9492 = n9318 & n9428 ;
  assign n9493 = n9492 ^ n9122 ;
  assign n9674 = n9673 ^ n9493 ;
  assign n9675 = n9673 ^ x89 ;
  assign n9676 = n9674 & n9675 ;
  assign n9677 = n9676 ^ x89 ;
  assign n9490 = n9322 & n9428 ;
  assign n9491 = n9490 ^ n9120 ;
  assign n9678 = n9677 ^ n9491 ;
  assign n9679 = n9677 ^ x90 ;
  assign n9680 = n9678 & n9679 ;
  assign n9681 = n9680 ^ x90 ;
  assign n9488 = n9326 & n9428 ;
  assign n9489 = n9488 ^ n9117 ;
  assign n9682 = n9681 ^ n9489 ;
  assign n9683 = n9681 ^ x91 ;
  assign n9684 = n9682 & n9683 ;
  assign n9685 = n9684 ^ x91 ;
  assign n9486 = n9330 & n9428 ;
  assign n9487 = n9486 ^ n9106 ;
  assign n9686 = n9685 ^ n9487 ;
  assign n9687 = n9685 ^ x92 ;
  assign n9688 = n9686 & n9687 ;
  assign n9689 = n9688 ^ x92 ;
  assign n9484 = n9334 & n9428 ;
  assign n9485 = n9484 ^ n9103 ;
  assign n9690 = n9689 ^ n9485 ;
  assign n9691 = n9689 ^ x93 ;
  assign n9692 = n9690 & n9691 ;
  assign n9693 = n9692 ^ x93 ;
  assign n9482 = n9338 & n9428 ;
  assign n9483 = n9482 ^ n9092 ;
  assign n9694 = n9693 ^ n9483 ;
  assign n9695 = n9693 ^ x94 ;
  assign n9696 = n9694 & n9695 ;
  assign n9697 = n9696 ^ x94 ;
  assign n9480 = n9342 & n9428 ;
  assign n9481 = n9480 ^ n9089 ;
  assign n9698 = n9697 ^ n9481 ;
  assign n9699 = n9697 ^ x95 ;
  assign n9700 = n9698 & n9699 ;
  assign n9701 = n9700 ^ x95 ;
  assign n9478 = n9346 & n9428 ;
  assign n9479 = n9478 ^ n9087 ;
  assign n9702 = n9701 ^ n9479 ;
  assign n9703 = n9701 ^ x96 ;
  assign n9704 = n9702 & n9703 ;
  assign n9705 = n9704 ^ x96 ;
  assign n9475 = n9348 ^ x96 ;
  assign n9476 = n9428 & n9475 ;
  assign n9477 = n9476 ^ n9084 ;
  assign n9706 = n9705 ^ n9477 ;
  assign n9707 = n9705 ^ x97 ;
  assign n9708 = n9706 & n9707 ;
  assign n9709 = n9708 ^ x97 ;
  assign n9472 = n9351 ^ x97 ;
  assign n9473 = n9428 & n9472 ;
  assign n9474 = n9473 ^ n9081 ;
  assign n9710 = n9709 ^ n9474 ;
  assign n9711 = n9709 ^ x98 ;
  assign n9712 = n9710 & n9711 ;
  assign n9713 = n9712 ^ x98 ;
  assign n9470 = n9356 & n9428 ;
  assign n9471 = n9470 ^ n9079 ;
  assign n9714 = n9713 ^ n9471 ;
  assign n9715 = n9713 ^ x99 ;
  assign n9716 = n9714 & n9715 ;
  assign n9717 = n9716 ^ x99 ;
  assign n9718 = n9717 ^ n9463 ;
  assign n9719 = n9718 ^ n9468 ;
  assign n9720 = ~n9469 & n9719 ;
  assign n9721 = n9720 ^ n9468 ;
  assign n9722 = ~n9464 & n9721 ;
  assign n9723 = n9722 ^ x101 ;
  assign n9726 = n9725 ^ n9723 ;
  assign n9727 = n9725 ^ x102 ;
  assign n9728 = n9726 & ~n9727 ;
  assign n9729 = n9728 ^ x102 ;
  assign n9460 = n9372 & n9428 ;
  assign n9461 = n9460 ^ n9071 ;
  assign n9730 = n9729 ^ n9461 ;
  assign n9731 = n9729 ^ x103 ;
  assign n9732 = n9730 & n9731 ;
  assign n9733 = n9732 ^ x103 ;
  assign n9458 = n9376 & n9428 ;
  assign n9459 = n9458 ^ n9069 ;
  assign n9734 = n9733 ^ n9459 ;
  assign n9735 = n9733 ^ x104 ;
  assign n9736 = n9734 & n9735 ;
  assign n9737 = n9736 ^ x104 ;
  assign n9456 = n9380 & n9428 ;
  assign n9457 = n9456 ^ n9067 ;
  assign n9738 = n9737 ^ n9457 ;
  assign n9739 = n9737 ^ x105 ;
  assign n9740 = n9738 & n9739 ;
  assign n9741 = n9740 ^ x105 ;
  assign n9454 = n9384 & n9428 ;
  assign n9455 = n9454 ^ n9065 ;
  assign n9742 = n9741 ^ n9455 ;
  assign n9743 = n9741 ^ x106 ;
  assign n9744 = n9742 & n9743 ;
  assign n9745 = n9744 ^ x106 ;
  assign n9451 = n9386 ^ x106 ;
  assign n9452 = n9428 & n9451 ;
  assign n9453 = n9452 ^ n9060 ;
  assign n9746 = n9745 ^ n9453 ;
  assign n9747 = n9745 ^ x107 ;
  assign n9748 = n9746 & n9747 ;
  assign n9749 = n9748 ^ x107 ;
  assign n9440 = n9060 ^ x107 ;
  assign n9441 = n9440 ^ n9386 ;
  assign n9442 = n9441 ^ x106 ;
  assign n9443 = n9442 ^ n9440 ;
  assign n9445 = n9386 ^ x107 ;
  assign n9446 = n9445 ^ n9440 ;
  assign n9447 = ~n9443 & ~n9446 ;
  assign n9448 = n9447 ^ n9440 ;
  assign n9449 = n9428 & ~n9448 ;
  assign n9450 = n9449 ^ n9057 ;
  assign n9750 = n9749 ^ n9450 ;
  assign n9751 = n9749 ^ x108 ;
  assign n9752 = n9750 & n9751 ;
  assign n9753 = n9752 ^ x108 ;
  assign n9437 = n9392 ^ x108 ;
  assign n9438 = n9428 & n9437 ;
  assign n9439 = n9438 ^ n9394 ;
  assign n9754 = n9753 ^ n9439 ;
  assign n9755 = n9753 ^ x109 ;
  assign n9756 = n9754 & n9755 ;
  assign n9757 = n9756 ^ x109 ;
  assign n9435 = n9400 & n9428 ;
  assign n9436 = n9435 ^ n9055 ;
  assign n9758 = n9757 ^ n9436 ;
  assign n9759 = n9757 ^ x110 ;
  assign n9760 = n9758 & n9759 ;
  assign n9761 = n9760 ^ x110 ;
  assign n9433 = n9404 & n9428 ;
  assign n9434 = n9433 ^ n9053 ;
  assign n9762 = n9761 ^ n9434 ;
  assign n9763 = n9761 ^ x111 ;
  assign n9764 = n9762 & n9763 ;
  assign n9765 = n9764 ^ x111 ;
  assign n9431 = n9408 & n9428 ;
  assign n9432 = n9431 ^ n9051 ;
  assign n9766 = n9765 ^ n9432 ;
  assign n9767 = n9765 ^ x112 ;
  assign n9768 = n9766 & n9767 ;
  assign n9769 = n9768 ^ x112 ;
  assign n9429 = n9412 & n9428 ;
  assign n9430 = n9429 ^ n9049 ;
  assign n9770 = n9769 ^ n9430 ;
  assign n9771 = n9769 ^ x113 ;
  assign n9772 = n9770 & n9771 ;
  assign n9773 = n9772 ^ x113 ;
  assign n9038 = n140 & n9037 ;
  assign n9421 = n9038 & n9420 ;
  assign n9422 = n9421 ^ n9037 ;
  assign n9775 = n9422 ^ x115 ;
  assign n9776 = n9414 ^ x113 ;
  assign n9777 = n9428 & n9776 ;
  assign n9778 = n9777 ^ n9047 ;
  assign n9780 = x114 & ~n9778 ;
  assign n9779 = n9778 ^ x114 ;
  assign n9781 = n9780 ^ n9779 ;
  assign n9782 = ~n9775 & ~n9781 ;
  assign n9783 = n9773 & n9782 ;
  assign n9784 = n139 & ~n9783 ;
  assign n9785 = n9780 ^ n9422 ;
  assign n9786 = ~n9775 & ~n9785 ;
  assign n9787 = n9786 ^ n9422 ;
  assign n9788 = n9784 & n9787 ;
  assign n9921 = n9917 ^ n9788 ;
  assign n9922 = ~n9920 & n9921 ;
  assign n9924 = n9923 ^ n9922 ;
  assign n9925 = x64 & n9924 ;
  assign n9926 = n9925 ^ n9923 ;
  assign n9927 = n9926 ^ x65 ;
  assign n9914 = x64 & n9428 ;
  assign n9910 = ~x12 & x64 ;
  assign n9911 = n9910 ^ x65 ;
  assign n9912 = n9788 & n9911 ;
  assign n9913 = n9912 ^ x13 ;
  assign n9915 = n9914 ^ n9913 ;
  assign n9928 = n9927 ^ n9915 ;
  assign n9929 = n9927 ^ x66 ;
  assign n9930 = n9928 & n9929 ;
  assign n9931 = n9930 ^ x66 ;
  assign n9906 = n9566 ^ x66 ;
  assign n9907 = n9788 & n9906 ;
  assign n9908 = n9907 ^ n9553 ;
  assign n9932 = n9931 ^ n9908 ;
  assign n9933 = n9931 ^ x67 ;
  assign n9934 = n9932 & n9933 ;
  assign n9935 = n9934 ^ x67 ;
  assign n9936 = n9935 ^ x68 ;
  assign n9774 = n9773 ^ x114 ;
  assign n10139 = n9778 ^ n9773 ;
  assign n10143 = n9774 & n10139 ;
  assign n10140 = x115 ^ x114 ;
  assign n10144 = n10143 ^ n10140 ;
  assign n9789 = n9774 & n9788 ;
  assign n9790 = n9789 ^ n9778 ;
  assign n9791 = ~x115 & n9790 ;
  assign n10207 = n10144 ^ n9791 ;
  assign n9792 = n9790 ^ x115 ;
  assign n9793 = n9792 ^ n9791 ;
  assign n10069 = n9466 ^ x101 ;
  assign n10070 = n10069 ^ n9717 ;
  assign n10071 = n10070 ^ x100 ;
  assign n10072 = n10071 ^ n10069 ;
  assign n10074 = n9717 ^ x101 ;
  assign n10075 = n10074 ^ n10069 ;
  assign n10076 = ~n10072 & ~n10075 ;
  assign n10077 = n10076 ^ n10069 ;
  assign n10078 = n9788 & ~n10077 ;
  assign n10079 = n10078 ^ n9463 ;
  assign n9819 = n9717 ^ x100 ;
  assign n9820 = n9788 & n9819 ;
  assign n9821 = n9820 ^ n9466 ;
  assign n9822 = n9821 ^ x101 ;
  assign n9826 = n9821 ^ x100 ;
  assign n9823 = n9715 & n9788 ;
  assign n9824 = n9823 ^ n9471 ;
  assign n9825 = n9824 ^ n9821 ;
  assign n9827 = n9826 ^ n9825 ;
  assign n9981 = n9635 & n9788 ;
  assign n9982 = n9981 ^ n9524 ;
  assign n9866 = n9631 & n9788 ;
  assign n9867 = n9866 ^ n9526 ;
  assign n9868 = n9867 ^ x79 ;
  assign n9873 = n9867 ^ x78 ;
  assign n9869 = n9623 ^ x77 ;
  assign n9870 = n9788 & n9869 ;
  assign n9871 = n9870 ^ n9625 ;
  assign n9872 = n9871 ^ n9867 ;
  assign n9874 = n9873 ^ n9872 ;
  assign n9875 = n9531 ^ x76 ;
  assign n9876 = n9875 ^ n9617 ;
  assign n9877 = n9876 ^ x75 ;
  assign n9878 = n9877 ^ n9875 ;
  assign n9880 = n9617 ^ x76 ;
  assign n9881 = n9880 ^ n9875 ;
  assign n9882 = ~n9878 & ~n9881 ;
  assign n9883 = n9882 ^ n9875 ;
  assign n9884 = n9788 & ~n9883 ;
  assign n9885 = n9884 ^ n9528 ;
  assign n9886 = n9885 ^ x77 ;
  assign n9894 = n9607 & n9788 ;
  assign n9895 = n9894 ^ n9540 ;
  assign n9896 = n9895 ^ x73 ;
  assign n9897 = n9603 & n9788 ;
  assign n9898 = n9897 ^ n9542 ;
  assign n9899 = n9898 ^ x72 ;
  assign n9937 = n9570 & n9788 ;
  assign n9938 = n9937 ^ n9586 ;
  assign n9939 = n9938 ^ n9935 ;
  assign n9940 = n9936 & n9939 ;
  assign n9941 = n9940 ^ x68 ;
  assign n9904 = n9591 & n9788 ;
  assign n9905 = n9904 ^ n9549 ;
  assign n9942 = n9941 ^ n9905 ;
  assign n9943 = n9941 ^ x69 ;
  assign n9944 = n9942 & n9943 ;
  assign n9945 = n9944 ^ x69 ;
  assign n9902 = n9595 & n9788 ;
  assign n9903 = n9902 ^ n9546 ;
  assign n9946 = n9945 ^ n9903 ;
  assign n9947 = n9945 ^ x70 ;
  assign n9948 = n9946 & n9947 ;
  assign n9949 = n9948 ^ x70 ;
  assign n9900 = n9599 & n9788 ;
  assign n9901 = n9900 ^ n9544 ;
  assign n9950 = n9949 ^ n9901 ;
  assign n9951 = n9949 ^ x71 ;
  assign n9952 = n9950 & n9951 ;
  assign n9953 = n9952 ^ x71 ;
  assign n9954 = n9953 ^ n9898 ;
  assign n9955 = ~n9899 & n9954 ;
  assign n9956 = n9955 ^ x72 ;
  assign n9957 = n9956 ^ n9895 ;
  assign n9958 = ~n9896 & n9957 ;
  assign n9959 = n9958 ^ x73 ;
  assign n9892 = n9611 & n9788 ;
  assign n9893 = n9892 ^ n9538 ;
  assign n9960 = n9959 ^ n9893 ;
  assign n9961 = n9959 ^ x74 ;
  assign n9962 = n9960 & n9961 ;
  assign n9963 = n9962 ^ x74 ;
  assign n9890 = n9615 & n9788 ;
  assign n9891 = n9890 ^ n9536 ;
  assign n9964 = n9963 ^ n9891 ;
  assign n9965 = n9963 ^ x75 ;
  assign n9966 = n9964 & n9965 ;
  assign n9967 = n9966 ^ x75 ;
  assign n9887 = n9617 ^ x75 ;
  assign n9888 = n9788 & n9887 ;
  assign n9889 = n9888 ^ n9531 ;
  assign n9968 = n9967 ^ n9889 ;
  assign n9969 = n9967 ^ x76 ;
  assign n9970 = n9968 & n9969 ;
  assign n9971 = n9970 ^ x76 ;
  assign n9972 = n9971 ^ n9885 ;
  assign n9973 = ~n9886 & n9972 ;
  assign n9974 = n9973 ^ x77 ;
  assign n9975 = n9974 ^ n9867 ;
  assign n9976 = n9975 ^ n9873 ;
  assign n9977 = ~n9874 & n9976 ;
  assign n9978 = n9977 ^ n9873 ;
  assign n9979 = ~n9868 & n9978 ;
  assign n9980 = n9979 ^ x79 ;
  assign n9983 = n9982 ^ n9980 ;
  assign n9984 = n9982 ^ x80 ;
  assign n9985 = n9983 & ~n9984 ;
  assign n9986 = n9985 ^ x80 ;
  assign n9864 = n9639 & n9788 ;
  assign n9865 = n9864 ^ n9522 ;
  assign n9987 = n9986 ^ n9865 ;
  assign n9988 = n9986 ^ x81 ;
  assign n9989 = n9987 & n9988 ;
  assign n9990 = n9989 ^ x81 ;
  assign n9862 = n9643 & n9788 ;
  assign n9863 = n9862 ^ n9520 ;
  assign n9991 = n9990 ^ n9863 ;
  assign n9992 = n9990 ^ x82 ;
  assign n9993 = n9991 & n9992 ;
  assign n9994 = n9993 ^ x82 ;
  assign n9860 = n9647 & n9788 ;
  assign n9861 = n9860 ^ n9518 ;
  assign n9995 = n9994 ^ n9861 ;
  assign n9996 = n9994 ^ x83 ;
  assign n9997 = n9995 & n9996 ;
  assign n9998 = n9997 ^ x83 ;
  assign n9858 = n9651 & n9788 ;
  assign n9859 = n9858 ^ n9516 ;
  assign n9999 = n9998 ^ n9859 ;
  assign n10000 = n9998 ^ x84 ;
  assign n10001 = n9999 & n10000 ;
  assign n10002 = n10001 ^ x84 ;
  assign n9856 = n9655 & n9788 ;
  assign n9857 = n9856 ^ n9514 ;
  assign n10003 = n10002 ^ n9857 ;
  assign n10004 = n10002 ^ x85 ;
  assign n10005 = n10003 & n10004 ;
  assign n10006 = n10005 ^ x85 ;
  assign n9854 = n9659 & n9788 ;
  assign n9855 = n9854 ^ n9512 ;
  assign n10007 = n10006 ^ n9855 ;
  assign n10008 = n10006 ^ x86 ;
  assign n10009 = n10007 & n10008 ;
  assign n10010 = n10009 ^ x86 ;
  assign n9852 = n9663 & n9788 ;
  assign n9853 = n9852 ^ n9509 ;
  assign n10011 = n10010 ^ n9853 ;
  assign n10012 = n10010 ^ x87 ;
  assign n10013 = n10011 & n10012 ;
  assign n10014 = n10013 ^ x87 ;
  assign n9850 = n9667 & n9788 ;
  assign n9851 = n9850 ^ n9498 ;
  assign n10015 = n10014 ^ n9851 ;
  assign n10016 = n10014 ^ x88 ;
  assign n10017 = n10015 & n10016 ;
  assign n10018 = n10017 ^ x88 ;
  assign n9848 = n9671 & n9788 ;
  assign n9849 = n9848 ^ n9495 ;
  assign n10019 = n10018 ^ n9849 ;
  assign n10020 = n10018 ^ x89 ;
  assign n10021 = n10019 & n10020 ;
  assign n10022 = n10021 ^ x89 ;
  assign n9846 = n9675 & n9788 ;
  assign n9847 = n9846 ^ n9493 ;
  assign n10023 = n10022 ^ n9847 ;
  assign n10024 = n10022 ^ x90 ;
  assign n10025 = n10023 & n10024 ;
  assign n10026 = n10025 ^ x90 ;
  assign n9844 = n9679 & n9788 ;
  assign n9845 = n9844 ^ n9491 ;
  assign n10027 = n10026 ^ n9845 ;
  assign n10028 = n10026 ^ x91 ;
  assign n10029 = n10027 & n10028 ;
  assign n10030 = n10029 ^ x91 ;
  assign n9842 = n9683 & n9788 ;
  assign n9843 = n9842 ^ n9489 ;
  assign n10031 = n10030 ^ n9843 ;
  assign n10032 = n10030 ^ x92 ;
  assign n10033 = n10031 & n10032 ;
  assign n10034 = n10033 ^ x92 ;
  assign n9840 = n9687 & n9788 ;
  assign n9841 = n9840 ^ n9487 ;
  assign n10035 = n10034 ^ n9841 ;
  assign n10036 = n10034 ^ x93 ;
  assign n10037 = n10035 & n10036 ;
  assign n10038 = n10037 ^ x93 ;
  assign n9838 = n9691 & n9788 ;
  assign n9839 = n9838 ^ n9485 ;
  assign n10039 = n10038 ^ n9839 ;
  assign n10040 = n10038 ^ x94 ;
  assign n10041 = n10039 & n10040 ;
  assign n10042 = n10041 ^ x94 ;
  assign n9836 = n9695 & n9788 ;
  assign n9837 = n9836 ^ n9483 ;
  assign n10043 = n10042 ^ n9837 ;
  assign n10044 = n10042 ^ x95 ;
  assign n10045 = n10043 & n10044 ;
  assign n10046 = n10045 ^ x95 ;
  assign n9834 = n9699 & n9788 ;
  assign n9835 = n9834 ^ n9481 ;
  assign n10047 = n10046 ^ n9835 ;
  assign n10048 = n10046 ^ x96 ;
  assign n10049 = n10047 & n10048 ;
  assign n10050 = n10049 ^ x96 ;
  assign n9832 = n9703 & n9788 ;
  assign n9833 = n9832 ^ n9479 ;
  assign n10051 = n10050 ^ n9833 ;
  assign n10052 = n10050 ^ x97 ;
  assign n10053 = n10051 & n10052 ;
  assign n10054 = n10053 ^ x97 ;
  assign n9830 = n9707 & n9788 ;
  assign n9831 = n9830 ^ n9477 ;
  assign n10055 = n10054 ^ n9831 ;
  assign n10056 = n10054 ^ x98 ;
  assign n10057 = n10055 & n10056 ;
  assign n10058 = n10057 ^ x98 ;
  assign n9828 = n9711 & n9788 ;
  assign n9829 = n9828 ^ n9474 ;
  assign n10059 = n10058 ^ n9829 ;
  assign n10060 = n10058 ^ x99 ;
  assign n10061 = n10059 & n10060 ;
  assign n10062 = n10061 ^ x99 ;
  assign n10063 = n10062 ^ n9821 ;
  assign n10064 = n10063 ^ n9826 ;
  assign n10065 = ~n9827 & n10064 ;
  assign n10066 = n10065 ^ n9826 ;
  assign n10067 = ~n9822 & n10066 ;
  assign n10068 = n10067 ^ x101 ;
  assign n10080 = n10079 ^ n10068 ;
  assign n10081 = n10079 ^ x102 ;
  assign n10082 = n10080 & ~n10081 ;
  assign n10083 = n10082 ^ x102 ;
  assign n9816 = n9723 ^ x102 ;
  assign n9817 = n9788 & n9816 ;
  assign n9818 = n9817 ^ n9725 ;
  assign n10084 = n10083 ^ n9818 ;
  assign n10085 = n10083 ^ x103 ;
  assign n10086 = n10084 & n10085 ;
  assign n10087 = n10086 ^ x103 ;
  assign n9814 = n9731 & n9788 ;
  assign n9815 = n9814 ^ n9461 ;
  assign n10088 = n10087 ^ n9815 ;
  assign n10089 = n10087 ^ x104 ;
  assign n10090 = n10088 & n10089 ;
  assign n10091 = n10090 ^ x104 ;
  assign n9812 = n9735 & n9788 ;
  assign n9813 = n9812 ^ n9459 ;
  assign n10092 = n10091 ^ n9813 ;
  assign n10093 = n10091 ^ x105 ;
  assign n10094 = n10092 & n10093 ;
  assign n10095 = n10094 ^ x105 ;
  assign n9810 = n9739 & n9788 ;
  assign n9811 = n9810 ^ n9457 ;
  assign n10096 = n10095 ^ n9811 ;
  assign n10097 = n10095 ^ x106 ;
  assign n10098 = n10096 & n10097 ;
  assign n10099 = n10098 ^ x106 ;
  assign n9808 = n9743 & n9788 ;
  assign n9809 = n9808 ^ n9455 ;
  assign n10100 = n10099 ^ n9809 ;
  assign n10101 = n10099 ^ x107 ;
  assign n10102 = n10100 & n10101 ;
  assign n10103 = n10102 ^ x107 ;
  assign n9806 = n9747 & n9788 ;
  assign n9807 = n9806 ^ n9453 ;
  assign n10104 = n10103 ^ n9807 ;
  assign n10105 = n10103 ^ x108 ;
  assign n10106 = n10104 & n10105 ;
  assign n10107 = n10106 ^ x108 ;
  assign n9804 = n9751 & n9788 ;
  assign n9805 = n9804 ^ n9450 ;
  assign n10108 = n10107 ^ n9805 ;
  assign n10109 = n10107 ^ x109 ;
  assign n10110 = n10108 & n10109 ;
  assign n10111 = n10110 ^ x109 ;
  assign n9802 = n9755 & n9788 ;
  assign n9803 = n9802 ^ n9439 ;
  assign n10112 = n10111 ^ n9803 ;
  assign n10113 = n10111 ^ x110 ;
  assign n10114 = n10112 & n10113 ;
  assign n10115 = n10114 ^ x110 ;
  assign n9800 = n9759 & n9788 ;
  assign n9801 = n9800 ^ n9436 ;
  assign n10116 = n10115 ^ n9801 ;
  assign n10117 = n10115 ^ x111 ;
  assign n10118 = n10116 & n10117 ;
  assign n10119 = n10118 ^ x111 ;
  assign n9798 = n9763 & n9788 ;
  assign n9799 = n9798 ^ n9434 ;
  assign n10120 = n10119 ^ n9799 ;
  assign n10121 = n10119 ^ x112 ;
  assign n10122 = n10120 & n10121 ;
  assign n10123 = n10122 ^ x112 ;
  assign n9796 = n9767 & n9788 ;
  assign n9797 = n9796 ^ n9432 ;
  assign n10124 = n10123 ^ n9797 ;
  assign n10125 = n10123 ^ x113 ;
  assign n10126 = n10124 & n10125 ;
  assign n10127 = n10126 ^ x113 ;
  assign n9794 = n9771 & n9788 ;
  assign n9795 = n9794 ^ n9430 ;
  assign n10128 = n10127 ^ n9795 ;
  assign n10129 = n10127 ^ x114 ;
  assign n10130 = n10128 & n10129 ;
  assign n10131 = n10130 ^ x114 ;
  assign n10132 = ~n9793 & ~n10131 ;
  assign n10163 = n10132 ^ x116 ;
  assign n10164 = n10163 ^ n10144 ;
  assign n10165 = n10164 ^ n9422 ;
  assign n10166 = n10165 ^ n10132 ;
  assign n10167 = n10166 ^ n10144 ;
  assign n10169 = n10167 ^ n10132 ;
  assign n10170 = n10169 ^ x116 ;
  assign n10171 = n10170 ^ n9791 ;
  assign n10172 = n10171 ^ n10170 ;
  assign n10200 = n10172 ^ n10132 ;
  assign n10201 = n10200 ^ n10167 ;
  assign n10175 = n10171 ^ n10132 ;
  assign n10176 = n10175 ^ n10170 ;
  assign n10184 = n10176 ^ n10169 ;
  assign n10185 = n10184 ^ n10167 ;
  assign n10187 = ~n10169 & n10185 ;
  assign n10177 = n10176 ^ n10144 ;
  assign n10180 = n10176 ^ n10167 ;
  assign n10178 = n10175 ^ n10167 ;
  assign n10179 = n10178 ^ n10144 ;
  assign n10181 = n10180 ^ n10179 ;
  assign n10182 = ~n10177 & n10181 ;
  assign n10188 = n10187 ^ n10182 ;
  assign n10189 = n10188 ^ n10180 ;
  assign n10190 = n10187 ^ n10178 ;
  assign n10191 = n10190 ^ n10180 ;
  assign n10192 = ~n10189 & n10191 ;
  assign n10193 = n10167 & n10192 ;
  assign n10194 = n10193 ^ n10187 ;
  assign n10195 = n10194 ^ n10185 ;
  assign n10202 = n10201 ^ n10195 ;
  assign n10205 = n10202 ^ n10164 ;
  assign n10206 = n10205 ^ n9422 ;
  assign n10208 = n10207 ^ n10206 ;
  assign n10154 = n9422 ^ x116 ;
  assign n10155 = n10154 ^ n10132 ;
  assign n10156 = n10155 ^ n9422 ;
  assign n10159 = n10156 ^ n9791 ;
  assign n10160 = n10159 ^ n10156 ;
  assign n10157 = n10156 ^ n10154 ;
  assign n10158 = n10157 ^ n9422 ;
  assign n10161 = n10160 ^ n10158 ;
  assign n10162 = n10161 ^ n10154 ;
  assign n10209 = n10208 ^ n10162 ;
  assign n10210 = n10209 ^ x116 ;
  assign n10211 = n10210 ^ n9422 ;
  assign n10212 = n138 & n10211 ;
  assign n10334 = n9936 & n10212 ;
  assign n10335 = n10334 ^ n9938 ;
  assign n10336 = n10335 ^ x69 ;
  assign n10346 = x64 & n9788 ;
  assign n10342 = ~x11 & x64 ;
  assign n10343 = n10342 ^ x65 ;
  assign n10344 = n10212 & n10343 ;
  assign n10345 = n10344 ^ x12 ;
  assign n10347 = n10346 ^ n10345 ;
  assign n10348 = n10347 ^ x66 ;
  assign n10357 = ~x11 & n911 ;
  assign n10358 = x10 & n10357 ;
  assign n10359 = n10358 ^ n10357 ;
  assign n10353 = ~x10 & x65 ;
  assign n10354 = ~x64 & n10353 ;
  assign n10360 = n10359 ^ n10354 ;
  assign n10361 = n10360 ^ n10353 ;
  assign n10349 = x64 & n10212 ;
  assign n10350 = n10349 ^ x11 ;
  assign n10351 = ~x10 & x64 ;
  assign n10352 = n10351 ^ x65 ;
  assign n10355 = n10354 ^ n10352 ;
  assign n10356 = ~n10350 & n10355 ;
  assign n10362 = n10361 ^ n10356 ;
  assign n10363 = n10362 ^ n10347 ;
  assign n10364 = ~n10348 & n10363 ;
  assign n10365 = n10364 ^ x66 ;
  assign n10339 = n9929 & n10212 ;
  assign n10340 = n10339 ^ n9915 ;
  assign n10366 = n10365 ^ n10340 ;
  assign n10367 = n10365 ^ x67 ;
  assign n10368 = n10366 & n10367 ;
  assign n10369 = n10368 ^ x67 ;
  assign n10337 = n9933 & n10212 ;
  assign n10338 = n10337 ^ n9908 ;
  assign n10370 = n10369 ^ n10338 ;
  assign n10371 = n10369 ^ x68 ;
  assign n10372 = n10370 & n10371 ;
  assign n10373 = n10372 ^ x68 ;
  assign n10374 = n10373 ^ n10335 ;
  assign n10375 = ~n10336 & n10374 ;
  assign n10376 = n10375 ^ x69 ;
  assign n10377 = n10376 ^ x70 ;
  assign n10378 = n9943 & n10212 ;
  assign n10379 = n10378 ^ n9905 ;
  assign n10380 = n10379 ^ n10376 ;
  assign n10381 = n10377 & n10380 ;
  assign n10382 = n10381 ^ x70 ;
  assign n10384 = n10382 ^ x71 ;
  assign n10554 = n10125 & n10212 ;
  assign n10555 = n10554 ^ n9797 ;
  assign n10218 = n10121 & n10212 ;
  assign n10219 = n10218 ^ n9799 ;
  assign n10220 = n10219 ^ x113 ;
  assign n10224 = n10219 ^ x112 ;
  assign n10221 = n10117 & n10212 ;
  assign n10222 = n10221 ^ n9801 ;
  assign n10223 = n10222 ^ n10219 ;
  assign n10225 = n10224 ^ n10223 ;
  assign n10409 = n9971 ^ x77 ;
  assign n10410 = n10212 & n10409 ;
  assign n10411 = n10410 ^ n9885 ;
  assign n10314 = n9969 & n10212 ;
  assign n10315 = n10314 ^ n9889 ;
  assign n10316 = n10315 ^ x77 ;
  assign n10320 = n10315 ^ x76 ;
  assign n10317 = n9965 & n10212 ;
  assign n10318 = n10317 ^ n9891 ;
  assign n10319 = n10318 ^ n10315 ;
  assign n10321 = n10320 ^ n10319 ;
  assign n10332 = n9947 & n10212 ;
  assign n10333 = n10332 ^ n9903 ;
  assign n10383 = n10382 ^ n10333 ;
  assign n10385 = n10383 & n10384 ;
  assign n10386 = n10385 ^ x71 ;
  assign n10330 = n9951 & n10212 ;
  assign n10331 = n10330 ^ n9901 ;
  assign n10387 = n10386 ^ n10331 ;
  assign n10388 = n10386 ^ x72 ;
  assign n10389 = n10387 & n10388 ;
  assign n10390 = n10389 ^ x72 ;
  assign n10327 = n9953 ^ x72 ;
  assign n10328 = n10212 & n10327 ;
  assign n10329 = n10328 ^ n9898 ;
  assign n10391 = n10390 ^ n10329 ;
  assign n10392 = n10390 ^ x73 ;
  assign n10393 = n10391 & n10392 ;
  assign n10394 = n10393 ^ x73 ;
  assign n10324 = n9956 ^ x73 ;
  assign n10325 = n10212 & n10324 ;
  assign n10326 = n10325 ^ n9895 ;
  assign n10395 = n10394 ^ n10326 ;
  assign n10396 = n10394 ^ x74 ;
  assign n10397 = n10395 & n10396 ;
  assign n10398 = n10397 ^ x74 ;
  assign n10322 = n9961 & n10212 ;
  assign n10323 = n10322 ^ n9893 ;
  assign n10399 = n10398 ^ n10323 ;
  assign n10400 = n10398 ^ x75 ;
  assign n10401 = n10399 & n10400 ;
  assign n10402 = n10401 ^ x75 ;
  assign n10403 = n10402 ^ n10315 ;
  assign n10404 = n10403 ^ n10320 ;
  assign n10405 = ~n10321 & n10404 ;
  assign n10406 = n10405 ^ n10320 ;
  assign n10407 = ~n10316 & n10406 ;
  assign n10408 = n10407 ^ x77 ;
  assign n10412 = n10411 ^ n10408 ;
  assign n10413 = n10411 ^ x78 ;
  assign n10414 = n10412 & ~n10413 ;
  assign n10415 = n10414 ^ x78 ;
  assign n10311 = n9974 ^ x78 ;
  assign n10312 = n10212 & n10311 ;
  assign n10313 = n10312 ^ n9871 ;
  assign n10416 = n10415 ^ n10313 ;
  assign n10417 = n10415 ^ x79 ;
  assign n10418 = n10416 & n10417 ;
  assign n10419 = n10418 ^ x79 ;
  assign n10300 = n9871 ^ x79 ;
  assign n10301 = n10300 ^ n9974 ;
  assign n10302 = n10301 ^ x78 ;
  assign n10303 = n10302 ^ n10300 ;
  assign n10305 = n9974 ^ x79 ;
  assign n10306 = n10305 ^ n10300 ;
  assign n10307 = ~n10303 & ~n10306 ;
  assign n10308 = n10307 ^ n10300 ;
  assign n10309 = n10212 & ~n10308 ;
  assign n10310 = n10309 ^ n9867 ;
  assign n10420 = n10419 ^ n10310 ;
  assign n10421 = n10419 ^ x80 ;
  assign n10422 = n10420 & n10421 ;
  assign n10423 = n10422 ^ x80 ;
  assign n10297 = n9980 ^ x80 ;
  assign n10298 = n10212 & n10297 ;
  assign n10299 = n10298 ^ n9982 ;
  assign n10424 = n10423 ^ n10299 ;
  assign n10425 = n10423 ^ x81 ;
  assign n10426 = n10424 & n10425 ;
  assign n10427 = n10426 ^ x81 ;
  assign n10295 = n9988 & n10212 ;
  assign n10296 = n10295 ^ n9865 ;
  assign n10428 = n10427 ^ n10296 ;
  assign n10429 = n10427 ^ x82 ;
  assign n10430 = n10428 & n10429 ;
  assign n10431 = n10430 ^ x82 ;
  assign n10293 = n9992 & n10212 ;
  assign n10294 = n10293 ^ n9863 ;
  assign n10432 = n10431 ^ n10294 ;
  assign n10433 = n10431 ^ x83 ;
  assign n10434 = n10432 & n10433 ;
  assign n10435 = n10434 ^ x83 ;
  assign n10291 = n9996 & n10212 ;
  assign n10292 = n10291 ^ n9861 ;
  assign n10436 = n10435 ^ n10292 ;
  assign n10437 = n10435 ^ x84 ;
  assign n10438 = n10436 & n10437 ;
  assign n10439 = n10438 ^ x84 ;
  assign n10289 = n10000 & n10212 ;
  assign n10290 = n10289 ^ n9859 ;
  assign n10440 = n10439 ^ n10290 ;
  assign n10441 = n10439 ^ x85 ;
  assign n10442 = n10440 & n10441 ;
  assign n10443 = n10442 ^ x85 ;
  assign n10287 = n10004 & n10212 ;
  assign n10288 = n10287 ^ n9857 ;
  assign n10444 = n10443 ^ n10288 ;
  assign n10445 = n10443 ^ x86 ;
  assign n10446 = n10444 & n10445 ;
  assign n10447 = n10446 ^ x86 ;
  assign n10285 = n10008 & n10212 ;
  assign n10286 = n10285 ^ n9855 ;
  assign n10448 = n10447 ^ n10286 ;
  assign n10449 = n10447 ^ x87 ;
  assign n10450 = n10448 & n10449 ;
  assign n10451 = n10450 ^ x87 ;
  assign n10283 = n10012 & n10212 ;
  assign n10284 = n10283 ^ n9853 ;
  assign n10452 = n10451 ^ n10284 ;
  assign n10453 = n10451 ^ x88 ;
  assign n10454 = n10452 & n10453 ;
  assign n10455 = n10454 ^ x88 ;
  assign n10281 = n10016 & n10212 ;
  assign n10282 = n10281 ^ n9851 ;
  assign n10456 = n10455 ^ n10282 ;
  assign n10457 = n10455 ^ x89 ;
  assign n10458 = n10456 & n10457 ;
  assign n10459 = n10458 ^ x89 ;
  assign n10279 = n10020 & n10212 ;
  assign n10280 = n10279 ^ n9849 ;
  assign n10460 = n10459 ^ n10280 ;
  assign n10461 = n10459 ^ x90 ;
  assign n10462 = n10460 & n10461 ;
  assign n10463 = n10462 ^ x90 ;
  assign n10277 = n10024 & n10212 ;
  assign n10278 = n10277 ^ n9847 ;
  assign n10464 = n10463 ^ n10278 ;
  assign n10465 = n10463 ^ x91 ;
  assign n10466 = n10464 & n10465 ;
  assign n10467 = n10466 ^ x91 ;
  assign n10275 = n10028 & n10212 ;
  assign n10276 = n10275 ^ n9845 ;
  assign n10468 = n10467 ^ n10276 ;
  assign n10469 = n10467 ^ x92 ;
  assign n10470 = n10468 & n10469 ;
  assign n10471 = n10470 ^ x92 ;
  assign n10273 = n10032 & n10212 ;
  assign n10274 = n10273 ^ n9843 ;
  assign n10472 = n10471 ^ n10274 ;
  assign n10473 = n10471 ^ x93 ;
  assign n10474 = n10472 & n10473 ;
  assign n10475 = n10474 ^ x93 ;
  assign n10271 = n10036 & n10212 ;
  assign n10272 = n10271 ^ n9841 ;
  assign n10476 = n10475 ^ n10272 ;
  assign n10477 = n10475 ^ x94 ;
  assign n10478 = n10476 & n10477 ;
  assign n10479 = n10478 ^ x94 ;
  assign n10269 = n10040 & n10212 ;
  assign n10270 = n10269 ^ n9839 ;
  assign n10480 = n10479 ^ n10270 ;
  assign n10481 = n10479 ^ x95 ;
  assign n10482 = n10480 & n10481 ;
  assign n10483 = n10482 ^ x95 ;
  assign n10267 = n10044 & n10212 ;
  assign n10268 = n10267 ^ n9837 ;
  assign n10484 = n10483 ^ n10268 ;
  assign n10485 = n10483 ^ x96 ;
  assign n10486 = n10484 & n10485 ;
  assign n10487 = n10486 ^ x96 ;
  assign n10265 = n10048 & n10212 ;
  assign n10266 = n10265 ^ n9835 ;
  assign n10488 = n10487 ^ n10266 ;
  assign n10489 = n10487 ^ x97 ;
  assign n10490 = n10488 & n10489 ;
  assign n10491 = n10490 ^ x97 ;
  assign n10263 = n10052 & n10212 ;
  assign n10264 = n10263 ^ n9833 ;
  assign n10492 = n10491 ^ n10264 ;
  assign n10493 = n10491 ^ x98 ;
  assign n10494 = n10492 & n10493 ;
  assign n10495 = n10494 ^ x98 ;
  assign n10261 = n10056 & n10212 ;
  assign n10262 = n10261 ^ n9831 ;
  assign n10496 = n10495 ^ n10262 ;
  assign n10497 = n10495 ^ x99 ;
  assign n10498 = n10496 & n10497 ;
  assign n10499 = n10498 ^ x99 ;
  assign n10259 = n10060 & n10212 ;
  assign n10260 = n10259 ^ n9829 ;
  assign n10500 = n10499 ^ n10260 ;
  assign n10501 = n10499 ^ x100 ;
  assign n10502 = n10500 & n10501 ;
  assign n10503 = n10502 ^ x100 ;
  assign n10256 = n10062 ^ x100 ;
  assign n10257 = n10212 & n10256 ;
  assign n10258 = n10257 ^ n9824 ;
  assign n10504 = n10503 ^ n10258 ;
  assign n10505 = n10503 ^ x101 ;
  assign n10506 = n10504 & n10505 ;
  assign n10507 = n10506 ^ x101 ;
  assign n10245 = n9824 ^ x101 ;
  assign n10246 = n10245 ^ n10062 ;
  assign n10247 = n10246 ^ x100 ;
  assign n10248 = n10247 ^ n10245 ;
  assign n10250 = n10062 ^ x101 ;
  assign n10251 = n10250 ^ n10245 ;
  assign n10252 = ~n10248 & ~n10251 ;
  assign n10253 = n10252 ^ n10245 ;
  assign n10254 = n10212 & ~n10253 ;
  assign n10255 = n10254 ^ n9821 ;
  assign n10508 = n10507 ^ n10255 ;
  assign n10509 = n10507 ^ x102 ;
  assign n10510 = n10508 & n10509 ;
  assign n10511 = n10510 ^ x102 ;
  assign n10242 = n10068 ^ x102 ;
  assign n10243 = n10212 & n10242 ;
  assign n10244 = n10243 ^ n10079 ;
  assign n10512 = n10511 ^ n10244 ;
  assign n10513 = n10511 ^ x103 ;
  assign n10514 = n10512 & n10513 ;
  assign n10515 = n10514 ^ x103 ;
  assign n10240 = n10085 & n10212 ;
  assign n10241 = n10240 ^ n9818 ;
  assign n10516 = n10515 ^ n10241 ;
  assign n10517 = n10515 ^ x104 ;
  assign n10518 = n10516 & n10517 ;
  assign n10519 = n10518 ^ x104 ;
  assign n10238 = n10089 & n10212 ;
  assign n10239 = n10238 ^ n9815 ;
  assign n10520 = n10519 ^ n10239 ;
  assign n10521 = n10519 ^ x105 ;
  assign n10522 = n10520 & n10521 ;
  assign n10523 = n10522 ^ x105 ;
  assign n10236 = n10093 & n10212 ;
  assign n10237 = n10236 ^ n9813 ;
  assign n10524 = n10523 ^ n10237 ;
  assign n10525 = n10523 ^ x106 ;
  assign n10526 = n10524 & n10525 ;
  assign n10527 = n10526 ^ x106 ;
  assign n10234 = n10097 & n10212 ;
  assign n10235 = n10234 ^ n9811 ;
  assign n10528 = n10527 ^ n10235 ;
  assign n10529 = n10527 ^ x107 ;
  assign n10530 = n10528 & n10529 ;
  assign n10531 = n10530 ^ x107 ;
  assign n10232 = n10101 & n10212 ;
  assign n10233 = n10232 ^ n9809 ;
  assign n10532 = n10531 ^ n10233 ;
  assign n10533 = n10531 ^ x108 ;
  assign n10534 = n10532 & n10533 ;
  assign n10535 = n10534 ^ x108 ;
  assign n10230 = n10105 & n10212 ;
  assign n10231 = n10230 ^ n9807 ;
  assign n10536 = n10535 ^ n10231 ;
  assign n10537 = n10535 ^ x109 ;
  assign n10538 = n10536 & n10537 ;
  assign n10539 = n10538 ^ x109 ;
  assign n10228 = n10109 & n10212 ;
  assign n10229 = n10228 ^ n9805 ;
  assign n10540 = n10539 ^ n10229 ;
  assign n10541 = n10539 ^ x110 ;
  assign n10542 = n10540 & n10541 ;
  assign n10543 = n10542 ^ x110 ;
  assign n10226 = n10113 & n10212 ;
  assign n10227 = n10226 ^ n9803 ;
  assign n10544 = n10543 ^ n10227 ;
  assign n10545 = n10543 ^ x111 ;
  assign n10546 = n10544 & n10545 ;
  assign n10547 = n10546 ^ x111 ;
  assign n10548 = n10547 ^ n10219 ;
  assign n10549 = n10548 ^ n10224 ;
  assign n10550 = ~n10225 & n10549 ;
  assign n10551 = n10550 ^ n10224 ;
  assign n10552 = ~n10220 & n10551 ;
  assign n10553 = n10552 ^ x113 ;
  assign n10556 = n10555 ^ n10553 ;
  assign n10557 = n10555 ^ x114 ;
  assign n10558 = n10556 & ~n10557 ;
  assign n10559 = n10558 ^ x114 ;
  assign n10216 = n10129 & n10212 ;
  assign n10217 = n10216 ^ n9795 ;
  assign n10560 = n10559 ^ n10217 ;
  assign n10561 = n10559 ^ x115 ;
  assign n10562 = n10560 & n10561 ;
  assign n10563 = n10562 ^ x115 ;
  assign n10213 = n10131 ^ x115 ;
  assign n10214 = n10212 & n10213 ;
  assign n10215 = n10214 ^ n9790 ;
  assign n10564 = n10563 ^ n10215 ;
  assign n10567 = n10215 ^ x116 ;
  assign n10568 = n10564 & ~n10567 ;
  assign n10565 = x117 ^ x116 ;
  assign n10569 = n10568 ^ n10565 ;
  assign n10133 = ~n9791 & ~n10132 ;
  assign n10134 = n10133 ^ x116 ;
  assign n10135 = n138 & ~n10134 ;
  assign n10149 = n10135 & n10144 ;
  assign n10150 = ~n10133 & n10149 ;
  assign n10151 = n10150 ^ n10133 ;
  assign n10136 = n10135 ^ n138 ;
  assign n10137 = n10136 ^ n10133 ;
  assign n10152 = n10151 ^ n10137 ;
  assign n10153 = n9422 & ~n10152 ;
  assign n10570 = n10153 ^ x117 ;
  assign n10573 = n10569 & ~n10570 ;
  assign n10574 = n10573 ^ x117 ;
  assign n10575 = n137 & ~n10574 ;
  assign n10787 = n10384 & n10575 ;
  assign n10788 = n10787 ^ n10333 ;
  assign n10698 = n10377 & n10575 ;
  assign n10699 = n10698 ^ n10379 ;
  assign n10700 = n10699 ^ x71 ;
  assign n10705 = n10699 ^ x70 ;
  assign n10701 = n10373 ^ x69 ;
  assign n10702 = n10575 & n10701 ;
  assign n10703 = n10702 ^ n10335 ;
  assign n10704 = n10703 ^ n10699 ;
  assign n10706 = n10705 ^ n10704 ;
  assign n10766 = n10362 ^ x66 ;
  assign n10767 = n10575 & n10766 ;
  assign n10768 = n10767 ^ n10347 ;
  assign n10711 = n10354 ^ n10353 ;
  assign n10712 = n10711 ^ n10352 ;
  assign n10713 = ~x9 & x64 ;
  assign n10714 = ~n10712 & ~n10713 ;
  assign n10720 = n10350 ^ x65 ;
  assign n10715 = n10713 ^ n10712 ;
  assign n10716 = n10715 ^ n10714 ;
  assign n10717 = ~n10353 & n10716 ;
  assign n10722 = n10717 ^ n10351 ;
  assign n10721 = n10716 ^ n10353 ;
  assign n10723 = n10722 ^ n10721 ;
  assign n10724 = ~n10720 & n10723 ;
  assign n10718 = n10350 & n10717 ;
  assign n10719 = n10718 ^ n10358 ;
  assign n10725 = n10724 ^ n10719 ;
  assign n10726 = ~n10714 & n10725 ;
  assign n10727 = n10575 & n10726 ;
  assign n10728 = n10727 ^ n10718 ;
  assign n10740 = x65 ^ x9 ;
  assign n10731 = n10350 ^ x9 ;
  assign n10741 = n10740 ^ n10731 ;
  assign n10742 = n10741 ^ x10 ;
  assign n10743 = n10742 ^ n10575 ;
  assign n10744 = n10743 ^ x9 ;
  assign n10729 = x65 ^ x10 ;
  assign n10730 = n10729 ^ n10575 ;
  assign n10732 = n10731 ^ n10350 ;
  assign n10733 = n10732 ^ n10575 ;
  assign n10734 = n10733 ^ n10731 ;
  assign n10737 = x65 & ~n10734 ;
  assign n10738 = n10737 ^ n10731 ;
  assign n10739 = n10730 & n10738 ;
  assign n10745 = n10744 ^ n10739 ;
  assign n10746 = ~x66 & n10353 ;
  assign n10747 = x64 & n10575 ;
  assign n10748 = n10575 ^ n10350 ;
  assign n10749 = ~n10747 & ~n10748 ;
  assign n10750 = n10746 & n10749 ;
  assign n10751 = n10750 ^ x66 ;
  assign n10752 = x64 & ~n10751 ;
  assign n10753 = ~n10745 & n10752 ;
  assign n10754 = n10753 ^ n10751 ;
  assign n10757 = n10754 ^ n10739 ;
  assign n10758 = n10757 ^ n10754 ;
  assign n10761 = n10753 & ~n10758 ;
  assign n10762 = n10743 & n10761 ;
  assign n10763 = n10762 ^ n10743 ;
  assign n10755 = n10754 ^ n10743 ;
  assign n10764 = n10763 ^ n10755 ;
  assign n10765 = ~n10728 & n10764 ;
  assign n10769 = n10768 ^ n10765 ;
  assign n10770 = n10768 ^ x67 ;
  assign n10771 = n10769 & ~n10770 ;
  assign n10772 = n10771 ^ x67 ;
  assign n10709 = n10367 & n10575 ;
  assign n10710 = n10709 ^ n10340 ;
  assign n10773 = n10772 ^ n10710 ;
  assign n10774 = n10772 ^ x68 ;
  assign n10775 = n10773 & n10774 ;
  assign n10776 = n10775 ^ x68 ;
  assign n10707 = n10371 & n10575 ;
  assign n10708 = n10707 ^ n10338 ;
  assign n10777 = n10776 ^ n10708 ;
  assign n10778 = n10776 ^ x69 ;
  assign n10779 = n10777 & n10778 ;
  assign n10780 = n10779 ^ x69 ;
  assign n10781 = n10780 ^ n10699 ;
  assign n10782 = n10781 ^ n10705 ;
  assign n10783 = ~n10706 & n10782 ;
  assign n10784 = n10783 ^ n10705 ;
  assign n10785 = ~n10700 & n10784 ;
  assign n10786 = n10785 ^ x71 ;
  assign n10789 = n10788 ^ n10786 ;
  assign n10790 = n10788 ^ x72 ;
  assign n10791 = n10789 & ~n10790 ;
  assign n10792 = n10791 ^ x72 ;
  assign n10696 = n10388 & n10575 ;
  assign n10697 = n10696 ^ n10331 ;
  assign n10793 = n10792 ^ n10697 ;
  assign n10794 = n10792 ^ x73 ;
  assign n10795 = n10793 & n10794 ;
  assign n10796 = n10795 ^ x73 ;
  assign n10694 = n10392 & n10575 ;
  assign n10695 = n10694 ^ n10329 ;
  assign n10797 = n10796 ^ n10695 ;
  assign n10798 = n10796 ^ x74 ;
  assign n10799 = n10797 & n10798 ;
  assign n10800 = n10799 ^ x74 ;
  assign n10692 = n10396 & n10575 ;
  assign n10693 = n10692 ^ n10326 ;
  assign n10801 = n10800 ^ n10693 ;
  assign n10802 = n10800 ^ x75 ;
  assign n10803 = n10801 & n10802 ;
  assign n10804 = n10803 ^ x75 ;
  assign n10690 = n10400 & n10575 ;
  assign n10691 = n10690 ^ n10323 ;
  assign n10805 = n10804 ^ n10691 ;
  assign n10806 = n10804 ^ x76 ;
  assign n10807 = n10805 & n10806 ;
  assign n10808 = n10807 ^ x76 ;
  assign n10687 = n10402 ^ x76 ;
  assign n10688 = n10575 & n10687 ;
  assign n10689 = n10688 ^ n10318 ;
  assign n10809 = n10808 ^ n10689 ;
  assign n10810 = n10808 ^ x77 ;
  assign n10811 = n10809 & n10810 ;
  assign n10812 = n10811 ^ x77 ;
  assign n10676 = n10318 ^ x77 ;
  assign n10677 = n10676 ^ n10402 ;
  assign n10678 = n10677 ^ x76 ;
  assign n10679 = n10678 ^ n10676 ;
  assign n10681 = n10402 ^ x77 ;
  assign n10682 = n10681 ^ n10676 ;
  assign n10683 = ~n10679 & ~n10682 ;
  assign n10684 = n10683 ^ n10676 ;
  assign n10685 = n10575 & ~n10684 ;
  assign n10686 = n10685 ^ n10315 ;
  assign n10813 = n10812 ^ n10686 ;
  assign n10814 = n10812 ^ x78 ;
  assign n10815 = n10813 & n10814 ;
  assign n10816 = n10815 ^ x78 ;
  assign n10673 = n10408 ^ x78 ;
  assign n10674 = n10575 & n10673 ;
  assign n10675 = n10674 ^ n10411 ;
  assign n10817 = n10816 ^ n10675 ;
  assign n10818 = n10816 ^ x79 ;
  assign n10819 = n10817 & n10818 ;
  assign n10820 = n10819 ^ x79 ;
  assign n10671 = n10417 & n10575 ;
  assign n10672 = n10671 ^ n10313 ;
  assign n10821 = n10820 ^ n10672 ;
  assign n10822 = n10820 ^ x80 ;
  assign n10823 = n10821 & n10822 ;
  assign n10824 = n10823 ^ x80 ;
  assign n10669 = n10421 & n10575 ;
  assign n10670 = n10669 ^ n10310 ;
  assign n10825 = n10824 ^ n10670 ;
  assign n10826 = n10824 ^ x81 ;
  assign n10827 = n10825 & n10826 ;
  assign n10828 = n10827 ^ x81 ;
  assign n10667 = n10425 & n10575 ;
  assign n10668 = n10667 ^ n10299 ;
  assign n10829 = n10828 ^ n10668 ;
  assign n10830 = n10828 ^ x82 ;
  assign n10831 = n10829 & n10830 ;
  assign n10832 = n10831 ^ x82 ;
  assign n10665 = n10429 & n10575 ;
  assign n10666 = n10665 ^ n10296 ;
  assign n10833 = n10832 ^ n10666 ;
  assign n10834 = n10832 ^ x83 ;
  assign n10835 = n10833 & n10834 ;
  assign n10836 = n10835 ^ x83 ;
  assign n10663 = n10433 & n10575 ;
  assign n10664 = n10663 ^ n10294 ;
  assign n10837 = n10836 ^ n10664 ;
  assign n10838 = n10836 ^ x84 ;
  assign n10839 = n10837 & n10838 ;
  assign n10840 = n10839 ^ x84 ;
  assign n10661 = n10437 & n10575 ;
  assign n10662 = n10661 ^ n10292 ;
  assign n10841 = n10840 ^ n10662 ;
  assign n10842 = n10840 ^ x85 ;
  assign n10843 = n10841 & n10842 ;
  assign n10844 = n10843 ^ x85 ;
  assign n10659 = n10441 & n10575 ;
  assign n10660 = n10659 ^ n10290 ;
  assign n10845 = n10844 ^ n10660 ;
  assign n10846 = n10844 ^ x86 ;
  assign n10847 = n10845 & n10846 ;
  assign n10848 = n10847 ^ x86 ;
  assign n10657 = n10445 & n10575 ;
  assign n10658 = n10657 ^ n10288 ;
  assign n10849 = n10848 ^ n10658 ;
  assign n10850 = n10848 ^ x87 ;
  assign n10851 = n10849 & n10850 ;
  assign n10852 = n10851 ^ x87 ;
  assign n10655 = n10449 & n10575 ;
  assign n10656 = n10655 ^ n10286 ;
  assign n10853 = n10852 ^ n10656 ;
  assign n10854 = n10852 ^ x88 ;
  assign n10855 = n10853 & n10854 ;
  assign n10856 = n10855 ^ x88 ;
  assign n10653 = n10453 & n10575 ;
  assign n10654 = n10653 ^ n10284 ;
  assign n10857 = n10856 ^ n10654 ;
  assign n10858 = n10856 ^ x89 ;
  assign n10859 = n10857 & n10858 ;
  assign n10860 = n10859 ^ x89 ;
  assign n10651 = n10457 & n10575 ;
  assign n10652 = n10651 ^ n10282 ;
  assign n10861 = n10860 ^ n10652 ;
  assign n10862 = n10860 ^ x90 ;
  assign n10863 = n10861 & n10862 ;
  assign n10864 = n10863 ^ x90 ;
  assign n10649 = n10461 & n10575 ;
  assign n10650 = n10649 ^ n10280 ;
  assign n10865 = n10864 ^ n10650 ;
  assign n10866 = n10864 ^ x91 ;
  assign n10867 = n10865 & n10866 ;
  assign n10868 = n10867 ^ x91 ;
  assign n10647 = n10465 & n10575 ;
  assign n10648 = n10647 ^ n10278 ;
  assign n10869 = n10868 ^ n10648 ;
  assign n10870 = n10868 ^ x92 ;
  assign n10871 = n10869 & n10870 ;
  assign n10872 = n10871 ^ x92 ;
  assign n10873 = n10872 ^ x93 ;
  assign n10874 = n10469 & n10575 ;
  assign n10875 = n10874 ^ n10276 ;
  assign n10876 = n10875 ^ n10872 ;
  assign n10877 = n10873 & n10876 ;
  assign n10878 = n10877 ^ x93 ;
  assign n10880 = n10878 ^ x94 ;
  assign n10576 = n10569 & n10575 ;
  assign n10577 = n10576 ^ n10153 ;
  assign n10998 = x117 & ~n10577 ;
  assign n10580 = n10561 & n10575 ;
  assign n10581 = n10580 ^ n10217 ;
  assign n10582 = n10581 ^ x116 ;
  assign n10587 = n10581 ^ x115 ;
  assign n10583 = n10553 ^ x114 ;
  assign n10584 = n10575 & n10583 ;
  assign n10585 = n10584 ^ n10555 ;
  assign n10586 = n10585 ^ n10581 ;
  assign n10588 = n10587 ^ n10586 ;
  assign n10589 = n10222 ^ x113 ;
  assign n10590 = n10589 ^ n10547 ;
  assign n10591 = n10590 ^ x112 ;
  assign n10592 = n10591 ^ n10589 ;
  assign n10594 = n10547 ^ x113 ;
  assign n10595 = n10594 ^ n10589 ;
  assign n10596 = ~n10592 & ~n10595 ;
  assign n10597 = n10596 ^ n10589 ;
  assign n10598 = n10575 & ~n10597 ;
  assign n10599 = n10598 ^ n10219 ;
  assign n10600 = n10599 ^ x114 ;
  assign n10605 = n10599 ^ x113 ;
  assign n10601 = n10547 ^ x112 ;
  assign n10602 = n10575 & n10601 ;
  assign n10603 = n10602 ^ n10222 ;
  assign n10604 = n10603 ^ n10599 ;
  assign n10606 = n10605 ^ n10604 ;
  assign n10937 = n10533 & n10575 ;
  assign n10938 = n10937 ^ n10233 ;
  assign n10613 = n10529 & n10575 ;
  assign n10614 = n10613 ^ n10235 ;
  assign n10615 = n10614 ^ x108 ;
  assign n10619 = n10614 ^ x107 ;
  assign n10616 = n10525 & n10575 ;
  assign n10617 = n10616 ^ n10237 ;
  assign n10618 = n10617 ^ n10614 ;
  assign n10620 = n10619 ^ n10618 ;
  assign n10645 = n10473 & n10575 ;
  assign n10646 = n10645 ^ n10274 ;
  assign n10879 = n10878 ^ n10646 ;
  assign n10881 = n10879 & n10880 ;
  assign n10882 = n10881 ^ x94 ;
  assign n10643 = n10477 & n10575 ;
  assign n10644 = n10643 ^ n10272 ;
  assign n10883 = n10882 ^ n10644 ;
  assign n10884 = n10882 ^ x95 ;
  assign n10885 = n10883 & n10884 ;
  assign n10886 = n10885 ^ x95 ;
  assign n10641 = n10481 & n10575 ;
  assign n10642 = n10641 ^ n10270 ;
  assign n10887 = n10886 ^ n10642 ;
  assign n10888 = n10886 ^ x96 ;
  assign n10889 = n10887 & n10888 ;
  assign n10890 = n10889 ^ x96 ;
  assign n10639 = n10485 & n10575 ;
  assign n10640 = n10639 ^ n10268 ;
  assign n10891 = n10890 ^ n10640 ;
  assign n10892 = n10890 ^ x97 ;
  assign n10893 = n10891 & n10892 ;
  assign n10894 = n10893 ^ x97 ;
  assign n10637 = n10489 & n10575 ;
  assign n10638 = n10637 ^ n10266 ;
  assign n10895 = n10894 ^ n10638 ;
  assign n10896 = n10894 ^ x98 ;
  assign n10897 = n10895 & n10896 ;
  assign n10898 = n10897 ^ x98 ;
  assign n10635 = n10493 & n10575 ;
  assign n10636 = n10635 ^ n10264 ;
  assign n10899 = n10898 ^ n10636 ;
  assign n10900 = n10898 ^ x99 ;
  assign n10901 = n10899 & n10900 ;
  assign n10902 = n10901 ^ x99 ;
  assign n10633 = n10497 & n10575 ;
  assign n10634 = n10633 ^ n10262 ;
  assign n10903 = n10902 ^ n10634 ;
  assign n10904 = n10902 ^ x100 ;
  assign n10905 = n10903 & n10904 ;
  assign n10906 = n10905 ^ x100 ;
  assign n10631 = n10501 & n10575 ;
  assign n10632 = n10631 ^ n10260 ;
  assign n10907 = n10906 ^ n10632 ;
  assign n10908 = n10906 ^ x101 ;
  assign n10909 = n10907 & n10908 ;
  assign n10910 = n10909 ^ x101 ;
  assign n10629 = n10505 & n10575 ;
  assign n10630 = n10629 ^ n10258 ;
  assign n10911 = n10910 ^ n10630 ;
  assign n10912 = n10910 ^ x102 ;
  assign n10913 = n10911 & n10912 ;
  assign n10914 = n10913 ^ x102 ;
  assign n10627 = n10509 & n10575 ;
  assign n10628 = n10627 ^ n10255 ;
  assign n10915 = n10914 ^ n10628 ;
  assign n10916 = n10914 ^ x103 ;
  assign n10917 = n10915 & n10916 ;
  assign n10918 = n10917 ^ x103 ;
  assign n10625 = n10513 & n10575 ;
  assign n10626 = n10625 ^ n10244 ;
  assign n10919 = n10918 ^ n10626 ;
  assign n10920 = n10918 ^ x104 ;
  assign n10921 = n10919 & n10920 ;
  assign n10922 = n10921 ^ x104 ;
  assign n10623 = n10517 & n10575 ;
  assign n10624 = n10623 ^ n10241 ;
  assign n10923 = n10922 ^ n10624 ;
  assign n10924 = n10922 ^ x105 ;
  assign n10925 = n10923 & n10924 ;
  assign n10926 = n10925 ^ x105 ;
  assign n10621 = n10521 & n10575 ;
  assign n10622 = n10621 ^ n10239 ;
  assign n10927 = n10926 ^ n10622 ;
  assign n10928 = n10926 ^ x106 ;
  assign n10929 = n10927 & n10928 ;
  assign n10930 = n10929 ^ x106 ;
  assign n10931 = n10930 ^ n10614 ;
  assign n10932 = n10931 ^ n10619 ;
  assign n10933 = ~n10620 & n10932 ;
  assign n10934 = n10933 ^ n10619 ;
  assign n10935 = ~n10615 & n10934 ;
  assign n10936 = n10935 ^ x108 ;
  assign n10939 = n10938 ^ n10936 ;
  assign n10940 = n10938 ^ x109 ;
  assign n10941 = n10939 & ~n10940 ;
  assign n10942 = n10941 ^ x109 ;
  assign n10611 = n10537 & n10575 ;
  assign n10612 = n10611 ^ n10231 ;
  assign n10943 = n10942 ^ n10612 ;
  assign n10944 = n10942 ^ x110 ;
  assign n10945 = n10943 & n10944 ;
  assign n10946 = n10945 ^ x110 ;
  assign n10609 = n10541 & n10575 ;
  assign n10610 = n10609 ^ n10229 ;
  assign n10947 = n10946 ^ n10610 ;
  assign n10948 = n10946 ^ x111 ;
  assign n10949 = n10947 & n10948 ;
  assign n10950 = n10949 ^ x111 ;
  assign n10607 = n10545 & n10575 ;
  assign n10608 = n10607 ^ n10227 ;
  assign n10951 = n10950 ^ n10608 ;
  assign n10952 = n10950 ^ x112 ;
  assign n10953 = n10951 & n10952 ;
  assign n10954 = n10953 ^ x112 ;
  assign n10955 = n10954 ^ n10599 ;
  assign n10956 = n10955 ^ n10605 ;
  assign n10957 = ~n10606 & n10956 ;
  assign n10958 = n10957 ^ n10605 ;
  assign n10959 = ~n10600 & n10958 ;
  assign n10960 = n10959 ^ x114 ;
  assign n10961 = n10960 ^ n10581 ;
  assign n10962 = n10961 ^ n10587 ;
  assign n10963 = ~n10588 & n10962 ;
  assign n10964 = n10963 ^ n10587 ;
  assign n10965 = ~n10582 & n10964 ;
  assign n10966 = n10965 ^ x116 ;
  assign n10980 = n10577 ^ x118 ;
  assign n10969 = n10563 ^ x116 ;
  assign n10970 = n10575 & n10969 ;
  assign n10971 = n10970 ^ n10215 ;
  assign n10972 = n10971 ^ n10966 ;
  assign n10982 = n10971 ^ x117 ;
  assign n10983 = ~n10972 & ~n10982 ;
  assign n10981 = n10971 ^ n10577 ;
  assign n10984 = n10983 ^ n10981 ;
  assign n10985 = ~n10980 & ~n10984 ;
  assign n10986 = n10985 ^ x118 ;
  assign n10987 = n10986 ^ n10983 ;
  assign n10988 = n10987 ^ n10986 ;
  assign n10991 = n10986 ^ n10966 ;
  assign n10992 = n10991 ^ n10986 ;
  assign n10993 = n10985 & n10992 ;
  assign n10994 = n10988 & n10993 ;
  assign n10995 = n10994 ^ n10988 ;
  assign n10996 = n10995 ^ n10987 ;
  assign n10997 = n136 & ~n10996 ;
  assign n10999 = n10966 & n10997 ;
  assign n11000 = n10998 & n10999 ;
  assign n11001 = n11000 ^ n10997 ;
  assign n11297 = n10880 & n11001 ;
  assign n11298 = n11297 ^ n10646 ;
  assign n11081 = n10873 & n11001 ;
  assign n11082 = n11081 ^ n10875 ;
  assign n11083 = n11082 ^ x94 ;
  assign n11087 = n11082 ^ x93 ;
  assign n11084 = n10870 & n11001 ;
  assign n11085 = n11084 ^ n10648 ;
  assign n11086 = n11085 ^ n11082 ;
  assign n11088 = n11087 ^ n11086 ;
  assign n11153 = n10747 ^ x10 ;
  assign n11151 = n10713 ^ x65 ;
  assign n11152 = n11001 & n11151 ;
  assign n11154 = n11153 ^ n11152 ;
  assign n11155 = n11154 ^ x66 ;
  assign n11163 = x9 & x65 ;
  assign n11160 = x65 ^ x8 ;
  assign n11156 = x64 ^ x9 ;
  assign n11157 = n11156 ^ x65 ;
  assign n11161 = n11157 ^ n11001 ;
  assign n11162 = ~n11160 & n11161 ;
  assign n11164 = n11163 ^ n11162 ;
  assign n11165 = x64 & n11164 ;
  assign n11166 = n11165 ^ n11163 ;
  assign n11167 = n11166 ^ x65 ;
  assign n11168 = n11167 ^ n11154 ;
  assign n11169 = ~n11155 & n11168 ;
  assign n11170 = n11169 ^ x66 ;
  assign n11171 = n11170 ^ x67 ;
  assign n11176 = n10353 ^ x65 ;
  assign n11177 = n11176 ^ x10 ;
  assign n11180 = x9 & n11177 ;
  assign n11181 = n11180 ^ x10 ;
  assign n11182 = n10747 & ~n11181 ;
  assign n11183 = n11182 ^ x66 ;
  assign n11173 = n10747 ^ n10716 ;
  assign n11174 = n10721 & n11173 ;
  assign n11184 = n11183 ^ n11174 ;
  assign n11185 = n11001 & ~n11184 ;
  assign n11186 = n11185 ^ n10350 ;
  assign n11172 = n10352 & n10575 ;
  assign n11187 = n11186 ^ n11172 ;
  assign n11188 = n11187 ^ n11170 ;
  assign n11189 = n11171 & n11188 ;
  assign n11190 = n11189 ^ x67 ;
  assign n11148 = n10765 ^ x67 ;
  assign n11149 = n11001 & n11148 ;
  assign n11150 = n11149 ^ n10768 ;
  assign n11191 = n11190 ^ n11150 ;
  assign n11192 = n11190 ^ x68 ;
  assign n11193 = n11191 & n11192 ;
  assign n11194 = n11193 ^ x68 ;
  assign n11146 = n10774 & n11001 ;
  assign n11147 = n11146 ^ n10710 ;
  assign n11195 = n11194 ^ n11147 ;
  assign n11196 = n11194 ^ x69 ;
  assign n11197 = n11195 & n11196 ;
  assign n11198 = n11197 ^ x69 ;
  assign n11144 = n10778 & n11001 ;
  assign n11145 = n11144 ^ n10708 ;
  assign n11199 = n11198 ^ n11145 ;
  assign n11200 = n11198 ^ x70 ;
  assign n11201 = n11199 & n11200 ;
  assign n11202 = n11201 ^ x70 ;
  assign n11141 = n10780 ^ x70 ;
  assign n11142 = n11001 & n11141 ;
  assign n11143 = n11142 ^ n10703 ;
  assign n11203 = n11202 ^ n11143 ;
  assign n11204 = n11202 ^ x71 ;
  assign n11205 = n11203 & n11204 ;
  assign n11206 = n11205 ^ x71 ;
  assign n11130 = n10703 ^ x71 ;
  assign n11131 = n11130 ^ n10780 ;
  assign n11132 = n11131 ^ x70 ;
  assign n11133 = n11132 ^ n11130 ;
  assign n11135 = n10780 ^ x71 ;
  assign n11136 = n11135 ^ n11130 ;
  assign n11137 = ~n11133 & ~n11136 ;
  assign n11138 = n11137 ^ n11130 ;
  assign n11139 = n11001 & ~n11138 ;
  assign n11140 = n11139 ^ n10699 ;
  assign n11207 = n11206 ^ n11140 ;
  assign n11208 = n11206 ^ x72 ;
  assign n11209 = n11207 & n11208 ;
  assign n11210 = n11209 ^ x72 ;
  assign n11127 = n10786 ^ x72 ;
  assign n11128 = n11001 & n11127 ;
  assign n11129 = n11128 ^ n10788 ;
  assign n11211 = n11210 ^ n11129 ;
  assign n11212 = n11210 ^ x73 ;
  assign n11213 = n11211 & n11212 ;
  assign n11214 = n11213 ^ x73 ;
  assign n11125 = n10794 & n11001 ;
  assign n11126 = n11125 ^ n10697 ;
  assign n11215 = n11214 ^ n11126 ;
  assign n11216 = n11214 ^ x74 ;
  assign n11217 = n11215 & n11216 ;
  assign n11218 = n11217 ^ x74 ;
  assign n11123 = n10798 & n11001 ;
  assign n11124 = n11123 ^ n10695 ;
  assign n11219 = n11218 ^ n11124 ;
  assign n11220 = n11218 ^ x75 ;
  assign n11221 = n11219 & n11220 ;
  assign n11222 = n11221 ^ x75 ;
  assign n11121 = n10802 & n11001 ;
  assign n11122 = n11121 ^ n10693 ;
  assign n11223 = n11222 ^ n11122 ;
  assign n11224 = n11222 ^ x76 ;
  assign n11225 = n11223 & n11224 ;
  assign n11226 = n11225 ^ x76 ;
  assign n11119 = n10806 & n11001 ;
  assign n11120 = n11119 ^ n10691 ;
  assign n11227 = n11226 ^ n11120 ;
  assign n11228 = n11226 ^ x77 ;
  assign n11229 = n11227 & n11228 ;
  assign n11230 = n11229 ^ x77 ;
  assign n11117 = n10810 & n11001 ;
  assign n11118 = n11117 ^ n10689 ;
  assign n11231 = n11230 ^ n11118 ;
  assign n11232 = n11230 ^ x78 ;
  assign n11233 = n11231 & n11232 ;
  assign n11234 = n11233 ^ x78 ;
  assign n11115 = n10814 & n11001 ;
  assign n11116 = n11115 ^ n10686 ;
  assign n11235 = n11234 ^ n11116 ;
  assign n11236 = n11234 ^ x79 ;
  assign n11237 = n11235 & n11236 ;
  assign n11238 = n11237 ^ x79 ;
  assign n11113 = n10818 & n11001 ;
  assign n11114 = n11113 ^ n10675 ;
  assign n11239 = n11238 ^ n11114 ;
  assign n11240 = n11238 ^ x80 ;
  assign n11241 = n11239 & n11240 ;
  assign n11242 = n11241 ^ x80 ;
  assign n11111 = n10822 & n11001 ;
  assign n11112 = n11111 ^ n10672 ;
  assign n11243 = n11242 ^ n11112 ;
  assign n11244 = n11242 ^ x81 ;
  assign n11245 = n11243 & n11244 ;
  assign n11246 = n11245 ^ x81 ;
  assign n11109 = n10826 & n11001 ;
  assign n11110 = n11109 ^ n10670 ;
  assign n11247 = n11246 ^ n11110 ;
  assign n11248 = n11246 ^ x82 ;
  assign n11249 = n11247 & n11248 ;
  assign n11250 = n11249 ^ x82 ;
  assign n11107 = n10830 & n11001 ;
  assign n11108 = n11107 ^ n10668 ;
  assign n11251 = n11250 ^ n11108 ;
  assign n11252 = n11250 ^ x83 ;
  assign n11253 = n11251 & n11252 ;
  assign n11254 = n11253 ^ x83 ;
  assign n11105 = n10834 & n11001 ;
  assign n11106 = n11105 ^ n10666 ;
  assign n11255 = n11254 ^ n11106 ;
  assign n11256 = n11254 ^ x84 ;
  assign n11257 = n11255 & n11256 ;
  assign n11258 = n11257 ^ x84 ;
  assign n11103 = n10838 & n11001 ;
  assign n11104 = n11103 ^ n10664 ;
  assign n11259 = n11258 ^ n11104 ;
  assign n11260 = n11258 ^ x85 ;
  assign n11261 = n11259 & n11260 ;
  assign n11262 = n11261 ^ x85 ;
  assign n11101 = n10842 & n11001 ;
  assign n11102 = n11101 ^ n10662 ;
  assign n11263 = n11262 ^ n11102 ;
  assign n11264 = n11262 ^ x86 ;
  assign n11265 = n11263 & n11264 ;
  assign n11266 = n11265 ^ x86 ;
  assign n11099 = n10846 & n11001 ;
  assign n11100 = n11099 ^ n10660 ;
  assign n11267 = n11266 ^ n11100 ;
  assign n11268 = n11266 ^ x87 ;
  assign n11269 = n11267 & n11268 ;
  assign n11270 = n11269 ^ x87 ;
  assign n11097 = n10850 & n11001 ;
  assign n11098 = n11097 ^ n10658 ;
  assign n11271 = n11270 ^ n11098 ;
  assign n11272 = n11270 ^ x88 ;
  assign n11273 = n11271 & n11272 ;
  assign n11274 = n11273 ^ x88 ;
  assign n11095 = n10854 & n11001 ;
  assign n11096 = n11095 ^ n10656 ;
  assign n11275 = n11274 ^ n11096 ;
  assign n11276 = n11274 ^ x89 ;
  assign n11277 = n11275 & n11276 ;
  assign n11278 = n11277 ^ x89 ;
  assign n11093 = n10858 & n11001 ;
  assign n11094 = n11093 ^ n10654 ;
  assign n11279 = n11278 ^ n11094 ;
  assign n11280 = n11278 ^ x90 ;
  assign n11281 = n11279 & n11280 ;
  assign n11282 = n11281 ^ x90 ;
  assign n11091 = n10862 & n11001 ;
  assign n11092 = n11091 ^ n10652 ;
  assign n11283 = n11282 ^ n11092 ;
  assign n11284 = n11282 ^ x91 ;
  assign n11285 = n11283 & n11284 ;
  assign n11286 = n11285 ^ x91 ;
  assign n11089 = n10866 & n11001 ;
  assign n11090 = n11089 ^ n10650 ;
  assign n11287 = n11286 ^ n11090 ;
  assign n11288 = n11286 ^ x92 ;
  assign n11289 = n11287 & n11288 ;
  assign n11290 = n11289 ^ x92 ;
  assign n11291 = n11290 ^ n11082 ;
  assign n11292 = n11291 ^ n11087 ;
  assign n11293 = ~n11088 & n11292 ;
  assign n11294 = n11293 ^ n11087 ;
  assign n11295 = ~n11083 & n11294 ;
  assign n11296 = n11295 ^ x94 ;
  assign n11299 = n11298 ^ n11296 ;
  assign n11300 = n11298 ^ x95 ;
  assign n11301 = n11299 & ~n11300 ;
  assign n11302 = n11301 ^ x95 ;
  assign n11079 = n10884 & n11001 ;
  assign n11080 = n11079 ^ n10644 ;
  assign n11303 = n11302 ^ n11080 ;
  assign n11304 = n11302 ^ x96 ;
  assign n11305 = n11303 & n11304 ;
  assign n11306 = n11305 ^ x96 ;
  assign n11077 = n10888 & n11001 ;
  assign n11078 = n11077 ^ n10642 ;
  assign n11307 = n11306 ^ n11078 ;
  assign n11308 = n11306 ^ x97 ;
  assign n11309 = n11307 & n11308 ;
  assign n11310 = n11309 ^ x97 ;
  assign n11075 = n10892 & n11001 ;
  assign n11076 = n11075 ^ n10640 ;
  assign n11311 = n11310 ^ n11076 ;
  assign n11312 = n11310 ^ x98 ;
  assign n11313 = n11311 & n11312 ;
  assign n11314 = n11313 ^ x98 ;
  assign n11073 = n10896 & n11001 ;
  assign n11074 = n11073 ^ n10638 ;
  assign n11315 = n11314 ^ n11074 ;
  assign n11316 = n11314 ^ x99 ;
  assign n11317 = n11315 & n11316 ;
  assign n11318 = n11317 ^ x99 ;
  assign n11071 = n10900 & n11001 ;
  assign n11072 = n11071 ^ n10636 ;
  assign n11319 = n11318 ^ n11072 ;
  assign n11320 = n11318 ^ x100 ;
  assign n11321 = n11319 & n11320 ;
  assign n11322 = n11321 ^ x100 ;
  assign n11069 = n10904 & n11001 ;
  assign n11070 = n11069 ^ n10634 ;
  assign n11323 = n11322 ^ n11070 ;
  assign n11324 = n11322 ^ x101 ;
  assign n11325 = n11323 & n11324 ;
  assign n11326 = n11325 ^ x101 ;
  assign n11067 = n10908 & n11001 ;
  assign n11068 = n11067 ^ n10632 ;
  assign n11327 = n11326 ^ n11068 ;
  assign n11328 = n11326 ^ x102 ;
  assign n11329 = n11327 & n11328 ;
  assign n11330 = n11329 ^ x102 ;
  assign n11065 = n10912 & n11001 ;
  assign n11066 = n11065 ^ n10630 ;
  assign n11331 = n11330 ^ n11066 ;
  assign n11332 = n11330 ^ x103 ;
  assign n11333 = n11331 & n11332 ;
  assign n11334 = n11333 ^ x103 ;
  assign n11063 = n10916 & n11001 ;
  assign n11064 = n11063 ^ n10628 ;
  assign n11335 = n11334 ^ n11064 ;
  assign n11336 = n11334 ^ x104 ;
  assign n11337 = n11335 & n11336 ;
  assign n11338 = n11337 ^ x104 ;
  assign n11061 = n10920 & n11001 ;
  assign n11062 = n11061 ^ n10626 ;
  assign n11339 = n11338 ^ n11062 ;
  assign n11340 = n11338 ^ x105 ;
  assign n11341 = n11339 & n11340 ;
  assign n11342 = n11341 ^ x105 ;
  assign n11059 = n10924 & n11001 ;
  assign n11060 = n11059 ^ n10624 ;
  assign n11343 = n11342 ^ n11060 ;
  assign n11344 = n11342 ^ x106 ;
  assign n11345 = n11343 & n11344 ;
  assign n11346 = n11345 ^ x106 ;
  assign n11347 = n11346 ^ x107 ;
  assign n11348 = n10928 & n11001 ;
  assign n11349 = n11348 ^ n10622 ;
  assign n11350 = n11349 ^ n11346 ;
  assign n11351 = n11347 & n11350 ;
  assign n11352 = n11351 ^ x107 ;
  assign n11354 = n11352 ^ x108 ;
  assign n10967 = n10966 ^ x118 ;
  assign n10578 = x118 ^ x117 ;
  assign n10968 = n10967 ^ n10578 ;
  assign n10975 = n10968 & n10972 ;
  assign n10976 = n10975 ^ n10578 ;
  assign n10977 = n136 & n10976 ;
  assign n10978 = n10577 & ~n10977 ;
  assign n11401 = n10978 ^ n10153 ;
  assign n11402 = ~x119 & ~n11401 ;
  assign n11403 = n11402 ^ n10153 ;
  assign n11013 = n10966 ^ x117 ;
  assign n11014 = n10997 & n11013 ;
  assign n11015 = n11014 ^ n10971 ;
  assign n11017 = n11015 ^ x117 ;
  assign n11002 = n10585 ^ x116 ;
  assign n11003 = n11002 ^ x115 ;
  assign n11004 = n11003 ^ n10960 ;
  assign n11005 = n11004 ^ n11002 ;
  assign n11007 = x116 ^ x115 ;
  assign n11008 = n11007 ^ n11002 ;
  assign n11009 = ~n11005 & ~n11008 ;
  assign n11010 = n11009 ^ n11002 ;
  assign n11011 = n11001 & ~n11010 ;
  assign n11012 = n11011 ^ n10581 ;
  assign n11016 = n11015 ^ n11012 ;
  assign n11018 = n11017 ^ n11016 ;
  assign n11056 = n10930 ^ x107 ;
  assign n11057 = n11001 & n11056 ;
  assign n11058 = n11057 ^ n10617 ;
  assign n11353 = n11352 ^ n11058 ;
  assign n11355 = n11353 & n11354 ;
  assign n11356 = n11355 ^ x108 ;
  assign n11045 = n10617 ^ x108 ;
  assign n11046 = n11045 ^ n10930 ;
  assign n11047 = n11046 ^ x107 ;
  assign n11048 = n11047 ^ n11045 ;
  assign n11050 = n10930 ^ x108 ;
  assign n11051 = n11050 ^ n11045 ;
  assign n11052 = ~n11048 & ~n11051 ;
  assign n11053 = n11052 ^ n11045 ;
  assign n11054 = n11001 & ~n11053 ;
  assign n11055 = n11054 ^ n10614 ;
  assign n11357 = n11356 ^ n11055 ;
  assign n11358 = n11356 ^ x109 ;
  assign n11359 = n11357 & n11358 ;
  assign n11360 = n11359 ^ x109 ;
  assign n11042 = n10936 ^ x109 ;
  assign n11043 = n11001 & n11042 ;
  assign n11044 = n11043 ^ n10938 ;
  assign n11361 = n11360 ^ n11044 ;
  assign n11362 = n11360 ^ x110 ;
  assign n11363 = n11361 & n11362 ;
  assign n11364 = n11363 ^ x110 ;
  assign n11040 = n10944 & n11001 ;
  assign n11041 = n11040 ^ n10612 ;
  assign n11365 = n11364 ^ n11041 ;
  assign n11366 = n11364 ^ x111 ;
  assign n11367 = n11365 & n11366 ;
  assign n11368 = n11367 ^ x111 ;
  assign n11038 = n10948 & n11001 ;
  assign n11039 = n11038 ^ n10610 ;
  assign n11369 = n11368 ^ n11039 ;
  assign n11370 = n11368 ^ x112 ;
  assign n11371 = n11369 & n11370 ;
  assign n11372 = n11371 ^ x112 ;
  assign n11036 = n10952 & n11001 ;
  assign n11037 = n11036 ^ n10608 ;
  assign n11373 = n11372 ^ n11037 ;
  assign n11374 = n11372 ^ x113 ;
  assign n11375 = n11373 & n11374 ;
  assign n11376 = n11375 ^ x113 ;
  assign n11033 = n10954 ^ x113 ;
  assign n11034 = n11001 & n11033 ;
  assign n11035 = n11034 ^ n10603 ;
  assign n11377 = n11376 ^ n11035 ;
  assign n11378 = n11376 ^ x114 ;
  assign n11379 = n11377 & n11378 ;
  assign n11380 = n11379 ^ x114 ;
  assign n11022 = n10603 ^ x114 ;
  assign n11023 = n11022 ^ n10954 ;
  assign n11024 = n11023 ^ x113 ;
  assign n11025 = n11024 ^ n11022 ;
  assign n11027 = n10954 ^ x114 ;
  assign n11028 = n11027 ^ n11022 ;
  assign n11029 = ~n11025 & ~n11028 ;
  assign n11030 = n11029 ^ n11022 ;
  assign n11031 = n11001 & ~n11030 ;
  assign n11032 = n11031 ^ n10599 ;
  assign n11381 = n11380 ^ n11032 ;
  assign n11382 = n11380 ^ x115 ;
  assign n11383 = n11381 & n11382 ;
  assign n11384 = n11383 ^ x115 ;
  assign n11019 = n10960 ^ x115 ;
  assign n11020 = n11001 & n11019 ;
  assign n11021 = n11020 ^ n10585 ;
  assign n11385 = n11384 ^ n11021 ;
  assign n11386 = n11384 ^ x116 ;
  assign n11387 = n11385 & n11386 ;
  assign n11388 = n11387 ^ x116 ;
  assign n11389 = n11388 ^ n11015 ;
  assign n11390 = n11389 ^ n11017 ;
  assign n11391 = ~n11018 & n11390 ;
  assign n11392 = n11391 ^ n11017 ;
  assign n11394 = x119 ^ x118 ;
  assign n11393 = n11015 ^ x119 ;
  assign n11395 = n11394 ^ n11393 ;
  assign n11396 = n11392 & ~n11395 ;
  assign n11397 = n11396 ^ n11394 ;
  assign n11406 = n11397 ^ n135 ;
  assign n11407 = n11403 & ~n11406 ;
  assign n11408 = n11407 ^ x119 ;
  assign n11409 = n135 & ~n11408 ;
  assign n11733 = n11354 & n11409 ;
  assign n11734 = n11733 ^ n11058 ;
  assign n11442 = n11347 & n11409 ;
  assign n11443 = n11442 ^ n11349 ;
  assign n11444 = n11443 ^ x108 ;
  assign n11448 = n11443 ^ x107 ;
  assign n11445 = n11344 & n11409 ;
  assign n11446 = n11445 ^ n11060 ;
  assign n11447 = n11446 ^ n11443 ;
  assign n11449 = n11448 ^ n11447 ;
  assign n11464 = n11308 & n11409 ;
  assign n11465 = n11464 ^ n11078 ;
  assign n11466 = n11465 ^ x98 ;
  assign n11467 = n11304 & n11409 ;
  assign n11468 = n11467 ^ n11080 ;
  assign n11469 = n11468 ^ x97 ;
  assign n11621 = n11240 & n11409 ;
  assign n11622 = n11621 ^ n11114 ;
  assign n11511 = n11236 & n11409 ;
  assign n11512 = n11511 ^ n11116 ;
  assign n11513 = n11512 ^ x80 ;
  assign n11517 = n11512 ^ x79 ;
  assign n11514 = n11232 & n11409 ;
  assign n11515 = n11514 ^ n11118 ;
  assign n11516 = n11515 ^ n11512 ;
  assign n11518 = n11517 ^ n11516 ;
  assign n11529 = n11208 & n11409 ;
  assign n11530 = n11529 ^ n11140 ;
  assign n11531 = n11530 ^ x73 ;
  assign n11532 = n11204 & n11409 ;
  assign n11533 = n11532 ^ n11143 ;
  assign n11534 = n11533 ^ x72 ;
  assign n11575 = n11192 & n11409 ;
  assign n11576 = n11575 ^ n11150 ;
  assign n11569 = n11171 & n11409 ;
  assign n11570 = n11569 ^ n11187 ;
  assign n11562 = n11167 ^ x66 ;
  assign n11563 = n11409 & n11562 ;
  assign n11564 = n11563 ^ n11154 ;
  assign n11556 = x64 & n11001 ;
  assign n11552 = ~x8 & x64 ;
  assign n11553 = n11552 ^ x65 ;
  assign n11554 = n11409 & n11553 ;
  assign n11555 = n11554 ^ x9 ;
  assign n11557 = n11556 ^ n11555 ;
  assign n11544 = x8 & x65 ;
  assign n11539 = x65 ^ x7 ;
  assign n11540 = x64 ^ x8 ;
  assign n11541 = n11540 ^ x65 ;
  assign n11542 = n11541 ^ n11409 ;
  assign n11543 = ~n11539 & n11542 ;
  assign n11545 = n11544 ^ n11543 ;
  assign n11548 = x64 & n11545 ;
  assign n11549 = n11548 ^ n11544 ;
  assign n11550 = n11549 ^ x65 ;
  assign n11558 = n11557 ^ n11550 ;
  assign n11559 = n11557 ^ x66 ;
  assign n11560 = n11558 & ~n11559 ;
  assign n11561 = n11560 ^ x66 ;
  assign n11565 = n11564 ^ n11561 ;
  assign n11566 = n11564 ^ x67 ;
  assign n11567 = n11565 & ~n11566 ;
  assign n11568 = n11567 ^ x67 ;
  assign n11571 = n11570 ^ n11568 ;
  assign n11572 = n11570 ^ x68 ;
  assign n11573 = n11571 & ~n11572 ;
  assign n11574 = n11573 ^ x68 ;
  assign n11577 = n11576 ^ n11574 ;
  assign n11578 = n11576 ^ x69 ;
  assign n11579 = n11577 & ~n11578 ;
  assign n11580 = n11579 ^ x69 ;
  assign n11537 = n11196 & n11409 ;
  assign n11538 = n11537 ^ n11147 ;
  assign n11581 = n11580 ^ n11538 ;
  assign n11582 = n11580 ^ x70 ;
  assign n11583 = n11581 & n11582 ;
  assign n11584 = n11583 ^ x70 ;
  assign n11535 = n11200 & n11409 ;
  assign n11536 = n11535 ^ n11145 ;
  assign n11585 = n11584 ^ n11536 ;
  assign n11586 = n11584 ^ x71 ;
  assign n11587 = n11585 & n11586 ;
  assign n11588 = n11587 ^ x71 ;
  assign n11589 = n11588 ^ n11533 ;
  assign n11590 = ~n11534 & n11589 ;
  assign n11591 = n11590 ^ x72 ;
  assign n11592 = n11591 ^ n11530 ;
  assign n11593 = ~n11531 & n11592 ;
  assign n11594 = n11593 ^ x73 ;
  assign n11527 = n11212 & n11409 ;
  assign n11528 = n11527 ^ n11129 ;
  assign n11595 = n11594 ^ n11528 ;
  assign n11596 = n11594 ^ x74 ;
  assign n11597 = n11595 & n11596 ;
  assign n11598 = n11597 ^ x74 ;
  assign n11525 = n11216 & n11409 ;
  assign n11526 = n11525 ^ n11126 ;
  assign n11599 = n11598 ^ n11526 ;
  assign n11600 = n11598 ^ x75 ;
  assign n11601 = n11599 & n11600 ;
  assign n11602 = n11601 ^ x75 ;
  assign n11523 = n11220 & n11409 ;
  assign n11524 = n11523 ^ n11124 ;
  assign n11603 = n11602 ^ n11524 ;
  assign n11604 = n11602 ^ x76 ;
  assign n11605 = n11603 & n11604 ;
  assign n11606 = n11605 ^ x76 ;
  assign n11521 = n11224 & n11409 ;
  assign n11522 = n11521 ^ n11122 ;
  assign n11607 = n11606 ^ n11522 ;
  assign n11608 = n11606 ^ x77 ;
  assign n11609 = n11607 & n11608 ;
  assign n11610 = n11609 ^ x77 ;
  assign n11519 = n11228 & n11409 ;
  assign n11520 = n11519 ^ n11120 ;
  assign n11611 = n11610 ^ n11520 ;
  assign n11612 = n11610 ^ x78 ;
  assign n11613 = n11611 & n11612 ;
  assign n11614 = n11613 ^ x78 ;
  assign n11615 = n11614 ^ n11512 ;
  assign n11616 = n11615 ^ n11517 ;
  assign n11617 = ~n11518 & n11616 ;
  assign n11618 = n11617 ^ n11517 ;
  assign n11619 = ~n11513 & n11618 ;
  assign n11620 = n11619 ^ x80 ;
  assign n11623 = n11622 ^ n11620 ;
  assign n11624 = n11622 ^ x81 ;
  assign n11625 = n11623 & ~n11624 ;
  assign n11626 = n11625 ^ x81 ;
  assign n11509 = n11244 & n11409 ;
  assign n11510 = n11509 ^ n11112 ;
  assign n11627 = n11626 ^ n11510 ;
  assign n11628 = n11626 ^ x82 ;
  assign n11629 = n11627 & n11628 ;
  assign n11630 = n11629 ^ x82 ;
  assign n11507 = n11248 & n11409 ;
  assign n11508 = n11507 ^ n11110 ;
  assign n11631 = n11630 ^ n11508 ;
  assign n11632 = n11630 ^ x83 ;
  assign n11633 = n11631 & n11632 ;
  assign n11634 = n11633 ^ x83 ;
  assign n11505 = n11252 & n11409 ;
  assign n11506 = n11505 ^ n11108 ;
  assign n11635 = n11634 ^ n11506 ;
  assign n11636 = n11634 ^ x84 ;
  assign n11637 = n11635 & n11636 ;
  assign n11638 = n11637 ^ x84 ;
  assign n11503 = n11256 & n11409 ;
  assign n11504 = n11503 ^ n11106 ;
  assign n11639 = n11638 ^ n11504 ;
  assign n11640 = n11638 ^ x85 ;
  assign n11641 = n11639 & n11640 ;
  assign n11642 = n11641 ^ x85 ;
  assign n11501 = n11260 & n11409 ;
  assign n11502 = n11501 ^ n11104 ;
  assign n11643 = n11642 ^ n11502 ;
  assign n11644 = n11642 ^ x86 ;
  assign n11645 = n11643 & n11644 ;
  assign n11646 = n11645 ^ x86 ;
  assign n11499 = n11264 & n11409 ;
  assign n11500 = n11499 ^ n11102 ;
  assign n11647 = n11646 ^ n11500 ;
  assign n11648 = n11646 ^ x87 ;
  assign n11649 = n11647 & n11648 ;
  assign n11650 = n11649 ^ x87 ;
  assign n11497 = n11268 & n11409 ;
  assign n11498 = n11497 ^ n11100 ;
  assign n11651 = n11650 ^ n11498 ;
  assign n11652 = n11650 ^ x88 ;
  assign n11653 = n11651 & n11652 ;
  assign n11654 = n11653 ^ x88 ;
  assign n11495 = n11272 & n11409 ;
  assign n11496 = n11495 ^ n11098 ;
  assign n11655 = n11654 ^ n11496 ;
  assign n11656 = n11654 ^ x89 ;
  assign n11657 = n11655 & n11656 ;
  assign n11658 = n11657 ^ x89 ;
  assign n11493 = n11276 & n11409 ;
  assign n11494 = n11493 ^ n11096 ;
  assign n11659 = n11658 ^ n11494 ;
  assign n11660 = n11658 ^ x90 ;
  assign n11661 = n11659 & n11660 ;
  assign n11662 = n11661 ^ x90 ;
  assign n11491 = n11280 & n11409 ;
  assign n11492 = n11491 ^ n11094 ;
  assign n11663 = n11662 ^ n11492 ;
  assign n11664 = n11662 ^ x91 ;
  assign n11665 = n11663 & n11664 ;
  assign n11666 = n11665 ^ x91 ;
  assign n11489 = n11284 & n11409 ;
  assign n11490 = n11489 ^ n11092 ;
  assign n11667 = n11666 ^ n11490 ;
  assign n11668 = n11666 ^ x92 ;
  assign n11669 = n11667 & n11668 ;
  assign n11670 = n11669 ^ x92 ;
  assign n11487 = n11288 & n11409 ;
  assign n11488 = n11487 ^ n11090 ;
  assign n11671 = n11670 ^ n11488 ;
  assign n11672 = n11670 ^ x93 ;
  assign n11673 = n11671 & n11672 ;
  assign n11674 = n11673 ^ x93 ;
  assign n11484 = n11290 ^ x93 ;
  assign n11485 = n11409 & n11484 ;
  assign n11486 = n11485 ^ n11085 ;
  assign n11675 = n11674 ^ n11486 ;
  assign n11676 = n11674 ^ x94 ;
  assign n11677 = n11675 & n11676 ;
  assign n11678 = n11677 ^ x94 ;
  assign n11473 = n11085 ^ x94 ;
  assign n11474 = n11473 ^ n11290 ;
  assign n11475 = n11474 ^ x93 ;
  assign n11476 = n11475 ^ n11473 ;
  assign n11477 = n11473 ^ n11085 ;
  assign n11478 = n11477 ^ n11290 ;
  assign n11479 = n11478 ^ n11473 ;
  assign n11480 = ~n11476 & ~n11479 ;
  assign n11481 = n11480 ^ n11473 ;
  assign n11482 = n11409 & ~n11481 ;
  assign n11483 = n11482 ^ n11082 ;
  assign n11679 = n11678 ^ n11483 ;
  assign n11680 = n11678 ^ x95 ;
  assign n11681 = n11679 & n11680 ;
  assign n11682 = n11681 ^ x95 ;
  assign n11470 = n11296 ^ x95 ;
  assign n11471 = n11409 & n11470 ;
  assign n11472 = n11471 ^ n11298 ;
  assign n11683 = n11682 ^ n11472 ;
  assign n11684 = n11682 ^ x96 ;
  assign n11685 = n11683 & n11684 ;
  assign n11686 = n11685 ^ x96 ;
  assign n11687 = n11686 ^ n11468 ;
  assign n11688 = ~n11469 & n11687 ;
  assign n11689 = n11688 ^ x97 ;
  assign n11690 = n11689 ^ n11465 ;
  assign n11691 = ~n11466 & n11690 ;
  assign n11692 = n11691 ^ x98 ;
  assign n11693 = n11692 ^ x99 ;
  assign n11694 = n11312 & n11409 ;
  assign n11695 = n11694 ^ n11076 ;
  assign n11696 = n11695 ^ n11692 ;
  assign n11697 = n11693 & n11696 ;
  assign n11698 = n11697 ^ x99 ;
  assign n11462 = n11316 & n11409 ;
  assign n11463 = n11462 ^ n11074 ;
  assign n11699 = n11698 ^ n11463 ;
  assign n11700 = n11698 ^ x100 ;
  assign n11701 = n11699 & n11700 ;
  assign n11702 = n11701 ^ x100 ;
  assign n11460 = n11320 & n11409 ;
  assign n11461 = n11460 ^ n11072 ;
  assign n11703 = n11702 ^ n11461 ;
  assign n11704 = n11702 ^ x101 ;
  assign n11705 = n11703 & n11704 ;
  assign n11706 = n11705 ^ x101 ;
  assign n11458 = n11324 & n11409 ;
  assign n11459 = n11458 ^ n11070 ;
  assign n11707 = n11706 ^ n11459 ;
  assign n11708 = n11706 ^ x102 ;
  assign n11709 = n11707 & n11708 ;
  assign n11710 = n11709 ^ x102 ;
  assign n11456 = n11328 & n11409 ;
  assign n11457 = n11456 ^ n11068 ;
  assign n11711 = n11710 ^ n11457 ;
  assign n11712 = n11710 ^ x103 ;
  assign n11713 = n11711 & n11712 ;
  assign n11714 = n11713 ^ x103 ;
  assign n11454 = n11332 & n11409 ;
  assign n11455 = n11454 ^ n11066 ;
  assign n11715 = n11714 ^ n11455 ;
  assign n11716 = n11714 ^ x104 ;
  assign n11717 = n11715 & n11716 ;
  assign n11718 = n11717 ^ x104 ;
  assign n11452 = n11336 & n11409 ;
  assign n11453 = n11452 ^ n11064 ;
  assign n11719 = n11718 ^ n11453 ;
  assign n11720 = n11718 ^ x105 ;
  assign n11721 = n11719 & n11720 ;
  assign n11722 = n11721 ^ x105 ;
  assign n11450 = n11340 & n11409 ;
  assign n11451 = n11450 ^ n11062 ;
  assign n11723 = n11722 ^ n11451 ;
  assign n11724 = n11722 ^ x106 ;
  assign n11725 = n11723 & n11724 ;
  assign n11726 = n11725 ^ x106 ;
  assign n11727 = n11726 ^ n11443 ;
  assign n11728 = n11727 ^ n11448 ;
  assign n11729 = ~n11449 & n11728 ;
  assign n11730 = n11729 ^ n11448 ;
  assign n11731 = ~n11444 & n11730 ;
  assign n11732 = n11731 ^ x108 ;
  assign n11735 = n11734 ^ n11732 ;
  assign n11736 = n11734 ^ x109 ;
  assign n11737 = n11735 & ~n11736 ;
  assign n11738 = n11737 ^ x109 ;
  assign n11440 = n11358 & n11409 ;
  assign n11441 = n11440 ^ n11055 ;
  assign n11739 = n11738 ^ n11441 ;
  assign n11740 = n11738 ^ x110 ;
  assign n11741 = n11739 & n11740 ;
  assign n11742 = n11741 ^ x110 ;
  assign n11438 = n11362 & n11409 ;
  assign n11439 = n11438 ^ n11044 ;
  assign n11743 = n11742 ^ n11439 ;
  assign n11744 = n11742 ^ x111 ;
  assign n11745 = n11743 & n11744 ;
  assign n11746 = n11745 ^ x111 ;
  assign n11747 = n11746 ^ x112 ;
  assign n11748 = n11366 & n11409 ;
  assign n11749 = n11748 ^ n11041 ;
  assign n11750 = n11749 ^ n11746 ;
  assign n11751 = n11747 & n11750 ;
  assign n11752 = n11751 ^ x112 ;
  assign n11754 = n11752 ^ x113 ;
  assign n11410 = n11388 ^ x118 ;
  assign n11411 = n11410 ^ n11012 ;
  assign n11412 = n11411 ^ x117 ;
  assign n11413 = n11412 ^ n11410 ;
  assign n11415 = n11012 ^ x118 ;
  assign n11416 = n11415 ^ n11410 ;
  assign n11417 = n11413 & ~n11416 ;
  assign n11418 = n11417 ^ n11410 ;
  assign n11419 = n11409 & n11418 ;
  assign n11420 = n11419 ^ n11015 ;
  assign n11421 = n11420 ^ x119 ;
  assign n11426 = n11420 ^ x118 ;
  assign n11422 = n11388 ^ x117 ;
  assign n11423 = n11409 & n11422 ;
  assign n11424 = n11423 ^ n11012 ;
  assign n11425 = n11424 ^ n11420 ;
  assign n11427 = n11426 ^ n11425 ;
  assign n11436 = n11370 & n11409 ;
  assign n11437 = n11436 ^ n11039 ;
  assign n11753 = n11752 ^ n11437 ;
  assign n11755 = n11753 & n11754 ;
  assign n11756 = n11755 ^ x113 ;
  assign n11434 = n11374 & n11409 ;
  assign n11435 = n11434 ^ n11037 ;
  assign n11757 = n11756 ^ n11435 ;
  assign n11758 = n11756 ^ x114 ;
  assign n11759 = n11757 & n11758 ;
  assign n11760 = n11759 ^ x114 ;
  assign n11432 = n11378 & n11409 ;
  assign n11433 = n11432 ^ n11035 ;
  assign n11761 = n11760 ^ n11433 ;
  assign n11762 = n11760 ^ x115 ;
  assign n11763 = n11761 & n11762 ;
  assign n11764 = n11763 ^ x115 ;
  assign n11430 = n11382 & n11409 ;
  assign n11431 = n11430 ^ n11032 ;
  assign n11765 = n11764 ^ n11431 ;
  assign n11766 = n11764 ^ x116 ;
  assign n11767 = n11765 & n11766 ;
  assign n11768 = n11767 ^ x116 ;
  assign n11428 = n11386 & n11409 ;
  assign n11429 = n11428 ^ n11021 ;
  assign n11769 = n11768 ^ n11429 ;
  assign n11770 = n11768 ^ x117 ;
  assign n11771 = n11769 & n11770 ;
  assign n11772 = n11771 ^ x117 ;
  assign n11773 = n11772 ^ n11420 ;
  assign n11774 = n11773 ^ n11426 ;
  assign n11775 = ~n11427 & n11774 ;
  assign n11776 = n11775 ^ n11426 ;
  assign n11777 = ~n11421 & n11776 ;
  assign n11778 = n11777 ^ x119 ;
  assign n11779 = x120 & n134 ;
  assign n11780 = ~n10577 & n11779 ;
  assign n11781 = n11780 ^ n134 ;
  assign n10979 = n135 & n10978 ;
  assign n11398 = n10979 & n11397 ;
  assign n11399 = n11398 ^ n10978 ;
  assign n11782 = n11399 ^ x120 ;
  assign n11783 = n11782 ^ n11778 ;
  assign n11784 = n11783 ^ n134 ;
  assign n11785 = n11781 & ~n11784 ;
  assign n11786 = n11778 & n11785 ;
  assign n11787 = n11786 ^ n11780 ;
  assign n11788 = n11787 ^ n134 ;
  assign n12149 = n11754 & n11788 ;
  assign n12150 = n12149 ^ n11437 ;
  assign n11808 = n11747 & n11788 ;
  assign n11809 = n11808 ^ n11749 ;
  assign n11810 = n11809 ^ x113 ;
  assign n11814 = n11809 ^ x112 ;
  assign n11811 = n11744 & n11788 ;
  assign n11812 = n11811 ^ n11439 ;
  assign n11813 = n11812 ^ n11809 ;
  assign n11815 = n11814 ^ n11813 ;
  assign n12137 = n11740 & n11788 ;
  assign n12138 = n12137 ^ n11441 ;
  assign n12130 = n11732 ^ x109 ;
  assign n12131 = n11788 & n12130 ;
  assign n12132 = n12131 ^ n11734 ;
  assign n11816 = n11446 ^ x108 ;
  assign n11817 = n11816 ^ n11726 ;
  assign n11818 = n11817 ^ x107 ;
  assign n11819 = n11818 ^ n11816 ;
  assign n11821 = n11726 ^ x108 ;
  assign n11822 = n11821 ^ n11816 ;
  assign n11823 = ~n11819 & ~n11822 ;
  assign n11824 = n11823 ^ n11816 ;
  assign n11825 = n11788 & ~n11824 ;
  assign n11826 = n11825 ^ n11443 ;
  assign n11827 = n11826 ^ x109 ;
  assign n11832 = n11826 ^ x108 ;
  assign n11828 = n11726 ^ x107 ;
  assign n11829 = n11788 & n11828 ;
  assign n11830 = n11829 ^ n11446 ;
  assign n11831 = n11830 ^ n11826 ;
  assign n11833 = n11832 ^ n11831 ;
  assign n11848 = n11693 & n11788 ;
  assign n11849 = n11848 ^ n11695 ;
  assign n11850 = n11849 ^ x100 ;
  assign n11851 = n11689 ^ x98 ;
  assign n11852 = n11788 & n11851 ;
  assign n11853 = n11852 ^ n11465 ;
  assign n11854 = n11853 ^ x99 ;
  assign n11860 = n11680 & n11788 ;
  assign n11861 = n11860 ^ n11483 ;
  assign n11862 = n11861 ^ x96 ;
  assign n11863 = n11676 & n11788 ;
  assign n11864 = n11863 ^ n11486 ;
  assign n11865 = n11864 ^ x95 ;
  assign n11874 = n11652 & n11788 ;
  assign n11875 = n11874 ^ n11498 ;
  assign n11876 = n11875 ^ x89 ;
  assign n12005 = n11608 & n11788 ;
  assign n12006 = n12005 ^ n11522 ;
  assign n11908 = n11604 & n11788 ;
  assign n11909 = n11908 ^ n11524 ;
  assign n11910 = n11909 ^ x77 ;
  assign n11914 = n11909 ^ x76 ;
  assign n11911 = n11600 & n11788 ;
  assign n11912 = n11911 ^ n11526 ;
  assign n11913 = n11912 ^ n11909 ;
  assign n11915 = n11914 ^ n11913 ;
  assign n11943 = x65 & n11788 ;
  assign n11942 = x64 & n11409 ;
  assign n11944 = n11943 ^ n11942 ;
  assign n11945 = n11944 ^ x8 ;
  assign n11940 = x64 & n11788 ;
  assign n11941 = ~x7 & n11940 ;
  assign n11946 = n11945 ^ n11941 ;
  assign n11947 = n11946 ^ x66 ;
  assign n11955 = x7 & x65 ;
  assign n11952 = x65 ^ x6 ;
  assign n11948 = x64 ^ x7 ;
  assign n11949 = n11948 ^ x65 ;
  assign n11953 = n11949 ^ n11788 ;
  assign n11954 = ~n11952 & n11953 ;
  assign n11956 = n11955 ^ n11954 ;
  assign n11957 = x64 & n11956 ;
  assign n11958 = n11957 ^ n11955 ;
  assign n11959 = n11958 ^ x65 ;
  assign n11960 = n11959 ^ n11946 ;
  assign n11961 = ~n11947 & n11960 ;
  assign n11962 = n11961 ^ x66 ;
  assign n11937 = n11550 ^ x66 ;
  assign n11938 = n11788 & n11937 ;
  assign n11939 = n11938 ^ n11557 ;
  assign n11963 = n11962 ^ n11939 ;
  assign n11964 = n11962 ^ x67 ;
  assign n11965 = n11963 & n11964 ;
  assign n11966 = n11965 ^ x67 ;
  assign n11934 = n11561 ^ x67 ;
  assign n11935 = n11788 & n11934 ;
  assign n11936 = n11935 ^ n11564 ;
  assign n11967 = n11966 ^ n11936 ;
  assign n11968 = n11966 ^ x68 ;
  assign n11969 = n11967 & n11968 ;
  assign n11970 = n11969 ^ x68 ;
  assign n11931 = n11568 ^ x68 ;
  assign n11932 = n11788 & n11931 ;
  assign n11933 = n11932 ^ n11570 ;
  assign n11971 = n11970 ^ n11933 ;
  assign n11972 = n11970 ^ x69 ;
  assign n11973 = n11971 & n11972 ;
  assign n11974 = n11973 ^ x69 ;
  assign n11928 = n11574 ^ x69 ;
  assign n11929 = n11788 & n11928 ;
  assign n11930 = n11929 ^ n11576 ;
  assign n11975 = n11974 ^ n11930 ;
  assign n11976 = n11974 ^ x70 ;
  assign n11977 = n11975 & n11976 ;
  assign n11978 = n11977 ^ x70 ;
  assign n11926 = n11582 & n11788 ;
  assign n11927 = n11926 ^ n11538 ;
  assign n11979 = n11978 ^ n11927 ;
  assign n11980 = n11978 ^ x71 ;
  assign n11981 = n11979 & n11980 ;
  assign n11982 = n11981 ^ x71 ;
  assign n11924 = n11586 & n11788 ;
  assign n11925 = n11924 ^ n11536 ;
  assign n11983 = n11982 ^ n11925 ;
  assign n11984 = n11982 ^ x72 ;
  assign n11985 = n11983 & n11984 ;
  assign n11986 = n11985 ^ x72 ;
  assign n11921 = n11588 ^ x72 ;
  assign n11922 = n11788 & n11921 ;
  assign n11923 = n11922 ^ n11533 ;
  assign n11987 = n11986 ^ n11923 ;
  assign n11988 = n11986 ^ x73 ;
  assign n11989 = n11987 & n11988 ;
  assign n11990 = n11989 ^ x73 ;
  assign n11918 = n11591 ^ x73 ;
  assign n11919 = n11788 & n11918 ;
  assign n11920 = n11919 ^ n11530 ;
  assign n11991 = n11990 ^ n11920 ;
  assign n11992 = n11990 ^ x74 ;
  assign n11993 = n11991 & n11992 ;
  assign n11994 = n11993 ^ x74 ;
  assign n11916 = n11596 & n11788 ;
  assign n11917 = n11916 ^ n11528 ;
  assign n11995 = n11994 ^ n11917 ;
  assign n11996 = n11994 ^ x75 ;
  assign n11997 = n11995 & n11996 ;
  assign n11998 = n11997 ^ x75 ;
  assign n11999 = n11998 ^ n11909 ;
  assign n12000 = n11999 ^ n11914 ;
  assign n12001 = ~n11915 & n12000 ;
  assign n12002 = n12001 ^ n11914 ;
  assign n12003 = ~n11910 & n12002 ;
  assign n12004 = n12003 ^ x77 ;
  assign n12007 = n12006 ^ n12004 ;
  assign n12008 = n12006 ^ x78 ;
  assign n12009 = n12007 & ~n12008 ;
  assign n12010 = n12009 ^ x78 ;
  assign n11906 = n11612 & n11788 ;
  assign n11907 = n11906 ^ n11520 ;
  assign n12011 = n12010 ^ n11907 ;
  assign n12012 = n12010 ^ x79 ;
  assign n12013 = n12011 & n12012 ;
  assign n12014 = n12013 ^ x79 ;
  assign n11903 = n11614 ^ x79 ;
  assign n11904 = n11788 & n11903 ;
  assign n11905 = n11904 ^ n11515 ;
  assign n12015 = n12014 ^ n11905 ;
  assign n12016 = n12014 ^ x80 ;
  assign n12017 = n12015 & n12016 ;
  assign n12018 = n12017 ^ x80 ;
  assign n11892 = n11515 ^ x80 ;
  assign n11893 = n11892 ^ n11614 ;
  assign n11894 = n11893 ^ x79 ;
  assign n11895 = n11894 ^ n11892 ;
  assign n11897 = n11614 ^ x80 ;
  assign n11898 = n11897 ^ n11892 ;
  assign n11899 = ~n11895 & ~n11898 ;
  assign n11900 = n11899 ^ n11892 ;
  assign n11901 = n11788 & ~n11900 ;
  assign n11902 = n11901 ^ n11512 ;
  assign n12019 = n12018 ^ n11902 ;
  assign n12020 = n12018 ^ x81 ;
  assign n12021 = n12019 & n12020 ;
  assign n12022 = n12021 ^ x81 ;
  assign n11889 = n11620 ^ x81 ;
  assign n11890 = n11788 & n11889 ;
  assign n11891 = n11890 ^ n11622 ;
  assign n12023 = n12022 ^ n11891 ;
  assign n12024 = n12022 ^ x82 ;
  assign n12025 = n12023 & n12024 ;
  assign n12026 = n12025 ^ x82 ;
  assign n11887 = n11628 & n11788 ;
  assign n11888 = n11887 ^ n11510 ;
  assign n12027 = n12026 ^ n11888 ;
  assign n12028 = n12026 ^ x83 ;
  assign n12029 = n12027 & n12028 ;
  assign n12030 = n12029 ^ x83 ;
  assign n11885 = n11632 & n11788 ;
  assign n11886 = n11885 ^ n11508 ;
  assign n12031 = n12030 ^ n11886 ;
  assign n12032 = n12030 ^ x84 ;
  assign n12033 = n12031 & n12032 ;
  assign n12034 = n12033 ^ x84 ;
  assign n11883 = n11636 & n11788 ;
  assign n11884 = n11883 ^ n11506 ;
  assign n12035 = n12034 ^ n11884 ;
  assign n12036 = n12034 ^ x85 ;
  assign n12037 = n12035 & n12036 ;
  assign n12038 = n12037 ^ x85 ;
  assign n11881 = n11640 & n11788 ;
  assign n11882 = n11881 ^ n11504 ;
  assign n12039 = n12038 ^ n11882 ;
  assign n12040 = n12038 ^ x86 ;
  assign n12041 = n12039 & n12040 ;
  assign n12042 = n12041 ^ x86 ;
  assign n11879 = n11644 & n11788 ;
  assign n11880 = n11879 ^ n11502 ;
  assign n12043 = n12042 ^ n11880 ;
  assign n12044 = n12042 ^ x87 ;
  assign n12045 = n12043 & n12044 ;
  assign n12046 = n12045 ^ x87 ;
  assign n11877 = n11648 & n11788 ;
  assign n11878 = n11877 ^ n11500 ;
  assign n12047 = n12046 ^ n11878 ;
  assign n12048 = n12046 ^ x88 ;
  assign n12049 = n12047 & n12048 ;
  assign n12050 = n12049 ^ x88 ;
  assign n12051 = n12050 ^ n11875 ;
  assign n12052 = ~n11876 & n12051 ;
  assign n12053 = n12052 ^ x89 ;
  assign n12054 = n12053 ^ x90 ;
  assign n12055 = n11656 & n11788 ;
  assign n12056 = n12055 ^ n11496 ;
  assign n12057 = n12056 ^ n12053 ;
  assign n12058 = n12054 & n12057 ;
  assign n12059 = n12058 ^ x90 ;
  assign n11872 = n11660 & n11788 ;
  assign n11873 = n11872 ^ n11494 ;
  assign n12060 = n12059 ^ n11873 ;
  assign n12061 = n12059 ^ x91 ;
  assign n12062 = n12060 & n12061 ;
  assign n12063 = n12062 ^ x91 ;
  assign n11870 = n11664 & n11788 ;
  assign n11871 = n11870 ^ n11492 ;
  assign n12064 = n12063 ^ n11871 ;
  assign n12065 = n12063 ^ x92 ;
  assign n12066 = n12064 & n12065 ;
  assign n12067 = n12066 ^ x92 ;
  assign n11868 = n11668 & n11788 ;
  assign n11869 = n11868 ^ n11490 ;
  assign n12068 = n12067 ^ n11869 ;
  assign n12069 = n12067 ^ x93 ;
  assign n12070 = n12068 & n12069 ;
  assign n12071 = n12070 ^ x93 ;
  assign n11866 = n11672 & n11788 ;
  assign n11867 = n11866 ^ n11488 ;
  assign n12072 = n12071 ^ n11867 ;
  assign n12073 = n12071 ^ x94 ;
  assign n12074 = n12072 & n12073 ;
  assign n12075 = n12074 ^ x94 ;
  assign n12076 = n12075 ^ n11864 ;
  assign n12077 = ~n11865 & n12076 ;
  assign n12078 = n12077 ^ x95 ;
  assign n12079 = n12078 ^ n11861 ;
  assign n12080 = ~n11862 & n12079 ;
  assign n12081 = n12080 ^ x96 ;
  assign n11858 = n11684 & n11788 ;
  assign n11859 = n11858 ^ n11472 ;
  assign n12082 = n12081 ^ n11859 ;
  assign n12083 = n12081 ^ x97 ;
  assign n12084 = n12082 & n12083 ;
  assign n12085 = n12084 ^ x97 ;
  assign n11855 = n11686 ^ x97 ;
  assign n11856 = n11788 & n11855 ;
  assign n11857 = n11856 ^ n11468 ;
  assign n12086 = n12085 ^ n11857 ;
  assign n12087 = n12085 ^ x98 ;
  assign n12088 = n12086 & n12087 ;
  assign n12089 = n12088 ^ x98 ;
  assign n12090 = n12089 ^ n11853 ;
  assign n12091 = ~n11854 & n12090 ;
  assign n12092 = n12091 ^ x99 ;
  assign n12093 = n12092 ^ n11849 ;
  assign n12094 = ~n11850 & n12093 ;
  assign n12095 = n12094 ^ x100 ;
  assign n11846 = n11700 & n11788 ;
  assign n11847 = n11846 ^ n11463 ;
  assign n12096 = n12095 ^ n11847 ;
  assign n12097 = n12095 ^ x101 ;
  assign n12098 = n12096 & n12097 ;
  assign n12099 = n12098 ^ x101 ;
  assign n11844 = n11704 & n11788 ;
  assign n11845 = n11844 ^ n11461 ;
  assign n12100 = n12099 ^ n11845 ;
  assign n12101 = n12099 ^ x102 ;
  assign n12102 = n12100 & n12101 ;
  assign n12103 = n12102 ^ x102 ;
  assign n11842 = n11708 & n11788 ;
  assign n11843 = n11842 ^ n11459 ;
  assign n12104 = n12103 ^ n11843 ;
  assign n12105 = n12103 ^ x103 ;
  assign n12106 = n12104 & n12105 ;
  assign n12107 = n12106 ^ x103 ;
  assign n11840 = n11712 & n11788 ;
  assign n11841 = n11840 ^ n11457 ;
  assign n12108 = n12107 ^ n11841 ;
  assign n12109 = n12107 ^ x104 ;
  assign n12110 = n12108 & n12109 ;
  assign n12111 = n12110 ^ x104 ;
  assign n11838 = n11716 & n11788 ;
  assign n11839 = n11838 ^ n11455 ;
  assign n12112 = n12111 ^ n11839 ;
  assign n12113 = n12111 ^ x105 ;
  assign n12114 = n12112 & n12113 ;
  assign n12115 = n12114 ^ x105 ;
  assign n11836 = n11720 & n11788 ;
  assign n11837 = n11836 ^ n11453 ;
  assign n12116 = n12115 ^ n11837 ;
  assign n12117 = n12115 ^ x106 ;
  assign n12118 = n12116 & n12117 ;
  assign n12119 = n12118 ^ x106 ;
  assign n11834 = n11724 & n11788 ;
  assign n11835 = n11834 ^ n11451 ;
  assign n12120 = n12119 ^ n11835 ;
  assign n12121 = n12119 ^ x107 ;
  assign n12122 = n12120 & n12121 ;
  assign n12123 = n12122 ^ x107 ;
  assign n12124 = n12123 ^ n11826 ;
  assign n12125 = n12124 ^ n11832 ;
  assign n12126 = ~n11833 & n12125 ;
  assign n12127 = n12126 ^ n11832 ;
  assign n12128 = ~n11827 & n12127 ;
  assign n12129 = n12128 ^ x109 ;
  assign n12133 = n12132 ^ n12129 ;
  assign n12134 = n12132 ^ x110 ;
  assign n12135 = n12133 & ~n12134 ;
  assign n12136 = n12135 ^ x110 ;
  assign n12139 = n12138 ^ n12136 ;
  assign n12140 = n12138 ^ x111 ;
  assign n12141 = n12139 & ~n12140 ;
  assign n12142 = n12141 ^ x111 ;
  assign n12143 = n12142 ^ n11809 ;
  assign n12144 = n12143 ^ n11814 ;
  assign n12145 = ~n11815 & n12144 ;
  assign n12146 = n12145 ^ n11814 ;
  assign n12147 = ~n11810 & n12146 ;
  assign n12148 = n12147 ^ x113 ;
  assign n12151 = n12150 ^ n12148 ;
  assign n12152 = n12150 ^ x114 ;
  assign n12153 = n12151 & ~n12152 ;
  assign n12154 = n12153 ^ x114 ;
  assign n11806 = n11758 & n11788 ;
  assign n11807 = n11806 ^ n11435 ;
  assign n12155 = n12154 ^ n11807 ;
  assign n12156 = n12154 ^ x115 ;
  assign n12157 = n12155 & n12156 ;
  assign n12158 = n12157 ^ x115 ;
  assign n11804 = n11762 & n11788 ;
  assign n11805 = n11804 ^ n11433 ;
  assign n12159 = n12158 ^ n11805 ;
  assign n12160 = n12158 ^ x116 ;
  assign n12161 = n12159 & n12160 ;
  assign n12162 = n12161 ^ x116 ;
  assign n11802 = n11766 & n11788 ;
  assign n11803 = n11802 ^ n11431 ;
  assign n12163 = n12162 ^ n11803 ;
  assign n12164 = n12162 ^ x117 ;
  assign n12165 = n12163 & n12164 ;
  assign n12166 = n12165 ^ x117 ;
  assign n11800 = n11770 & n11788 ;
  assign n11801 = n11800 ^ n11429 ;
  assign n12167 = n12166 ^ n11801 ;
  assign n12168 = n12166 ^ x118 ;
  assign n12169 = n12167 & n12168 ;
  assign n12170 = n12169 ^ x118 ;
  assign n12171 = n12170 ^ x119 ;
  assign n12172 = n11772 ^ x118 ;
  assign n12173 = n11788 & n12172 ;
  assign n12174 = n12173 ^ n11424 ;
  assign n12175 = n12174 ^ n12170 ;
  assign n12176 = n12171 & n12175 ;
  assign n12177 = n12176 ^ x119 ;
  assign n11789 = n11424 ^ x119 ;
  assign n11790 = n11789 ^ n11772 ;
  assign n11791 = n11790 ^ x118 ;
  assign n11792 = n11791 ^ n11789 ;
  assign n11794 = n11772 ^ x119 ;
  assign n11795 = n11794 ^ n11789 ;
  assign n11796 = ~n11792 & ~n11795 ;
  assign n11797 = n11796 ^ n11789 ;
  assign n11798 = n11788 & ~n11797 ;
  assign n11799 = n11798 ^ n11420 ;
  assign n12178 = n12177 ^ n11799 ;
  assign n12179 = n12177 ^ x120 ;
  assign n12180 = n12178 & n12179 ;
  assign n12181 = n12180 ^ x120 ;
  assign n12183 = n11778 ^ x120 ;
  assign n12184 = n134 & n11399 ;
  assign n12185 = n12183 & n12184 ;
  assign n12186 = n12185 ^ n11399 ;
  assign n12955 = ~x121 & n12186 ;
  assign n12956 = ~n12181 & n12955 ;
  assign n12189 = n12186 ^ n10978 ;
  assign n12190 = ~x121 & ~n12189 ;
  assign n12191 = n12190 ^ n10978 ;
  assign n12182 = n12181 ^ x121 ;
  assign n12192 = n12182 ^ n133 ;
  assign n12193 = n12191 & ~n12192 ;
  assign n12194 = n12193 ^ x121 ;
  assign n12195 = n133 & ~n12194 ;
  assign n12198 = n12171 & n12195 ;
  assign n12199 = n12198 ^ n12174 ;
  assign n12200 = n12199 ^ x120 ;
  assign n12201 = n12168 & n12195 ;
  assign n12202 = n12201 ^ n11801 ;
  assign n12203 = n12202 ^ x119 ;
  assign n12204 = n12164 & n12195 ;
  assign n12205 = n12204 ^ n11803 ;
  assign n12206 = n12205 ^ x118 ;
  assign n12211 = n12148 ^ x114 ;
  assign n12212 = n12195 & n12211 ;
  assign n12213 = n12212 ^ n12150 ;
  assign n12214 = n12213 ^ x115 ;
  assign n12536 = n12123 ^ x108 ;
  assign n12537 = n12195 & n12536 ;
  assign n12538 = n12537 ^ n11830 ;
  assign n12246 = n12121 & n12195 ;
  assign n12247 = n12246 ^ n11835 ;
  assign n12248 = n12247 ^ x108 ;
  assign n12252 = n12247 ^ x107 ;
  assign n12249 = n12117 & n12195 ;
  assign n12250 = n12249 ^ n11837 ;
  assign n12251 = n12250 ^ n12247 ;
  assign n12253 = n12252 ^ n12251 ;
  assign n12282 = n12069 & n12195 ;
  assign n12283 = n12282 ^ n11869 ;
  assign n12284 = n12283 ^ x94 ;
  assign n12285 = n12065 & n12195 ;
  assign n12286 = n12285 ^ n11871 ;
  assign n12287 = n12286 ^ x93 ;
  assign n12297 = n12044 & n12195 ;
  assign n12298 = n12297 ^ n11880 ;
  assign n12299 = n12298 ^ x88 ;
  assign n12300 = n12040 & n12195 ;
  assign n12301 = n12300 ^ n11882 ;
  assign n12302 = n12301 ^ x87 ;
  assign n12331 = n11998 ^ x76 ;
  assign n12332 = n12195 & n12331 ;
  assign n12333 = n12332 ^ n11912 ;
  assign n12334 = n12333 ^ x77 ;
  assign n12335 = n11996 & n12195 ;
  assign n12336 = n12335 ^ n11917 ;
  assign n12337 = n12336 ^ x76 ;
  assign n12361 = n11940 ^ x7 ;
  assign n12358 = ~x6 & x64 ;
  assign n12359 = n12358 ^ x65 ;
  assign n12360 = n12195 & n12359 ;
  assign n12362 = n12361 ^ n12360 ;
  assign n12363 = n12362 ^ x66 ;
  assign n12365 = x64 & n12195 ;
  assign n12371 = x5 & n12365 ;
  assign n12364 = ~x5 & x64 ;
  assign n12368 = n12364 ^ x65 ;
  assign n12369 = x6 & n12368 ;
  assign n12366 = n12365 ^ n12364 ;
  assign n12367 = ~x65 & ~n12366 ;
  assign n12370 = n12369 ^ n12367 ;
  assign n12372 = n12371 ^ n12370 ;
  assign n12373 = n12372 ^ n12362 ;
  assign n12374 = ~n12363 & ~n12373 ;
  assign n12375 = n12374 ^ x66 ;
  assign n12354 = n11959 ^ x66 ;
  assign n12355 = n12195 & n12354 ;
  assign n12356 = n12355 ^ n11946 ;
  assign n12376 = n12375 ^ n12356 ;
  assign n12377 = n12375 ^ x67 ;
  assign n12378 = n12376 & n12377 ;
  assign n12379 = n12378 ^ x67 ;
  assign n12352 = n11964 & n12195 ;
  assign n12353 = n12352 ^ n11939 ;
  assign n12380 = n12379 ^ n12353 ;
  assign n12381 = n12379 ^ x68 ;
  assign n12382 = n12380 & n12381 ;
  assign n12383 = n12382 ^ x68 ;
  assign n12350 = n11968 & n12195 ;
  assign n12351 = n12350 ^ n11936 ;
  assign n12384 = n12383 ^ n12351 ;
  assign n12385 = n12383 ^ x69 ;
  assign n12386 = n12384 & n12385 ;
  assign n12387 = n12386 ^ x69 ;
  assign n12348 = n11972 & n12195 ;
  assign n12349 = n12348 ^ n11933 ;
  assign n12388 = n12387 ^ n12349 ;
  assign n12389 = n12387 ^ x70 ;
  assign n12390 = n12388 & n12389 ;
  assign n12391 = n12390 ^ x70 ;
  assign n12346 = n11976 & n12195 ;
  assign n12347 = n12346 ^ n11930 ;
  assign n12392 = n12391 ^ n12347 ;
  assign n12393 = n12391 ^ x71 ;
  assign n12394 = n12392 & n12393 ;
  assign n12395 = n12394 ^ x71 ;
  assign n12344 = n11980 & n12195 ;
  assign n12345 = n12344 ^ n11927 ;
  assign n12396 = n12395 ^ n12345 ;
  assign n12397 = n12395 ^ x72 ;
  assign n12398 = n12396 & n12397 ;
  assign n12399 = n12398 ^ x72 ;
  assign n12342 = n11984 & n12195 ;
  assign n12343 = n12342 ^ n11925 ;
  assign n12400 = n12399 ^ n12343 ;
  assign n12401 = n12399 ^ x73 ;
  assign n12402 = n12400 & n12401 ;
  assign n12403 = n12402 ^ x73 ;
  assign n12340 = n11988 & n12195 ;
  assign n12341 = n12340 ^ n11923 ;
  assign n12404 = n12403 ^ n12341 ;
  assign n12405 = n12403 ^ x74 ;
  assign n12406 = n12404 & n12405 ;
  assign n12407 = n12406 ^ x74 ;
  assign n12338 = n11992 & n12195 ;
  assign n12339 = n12338 ^ n11920 ;
  assign n12408 = n12407 ^ n12339 ;
  assign n12409 = n12407 ^ x75 ;
  assign n12410 = n12408 & n12409 ;
  assign n12411 = n12410 ^ x75 ;
  assign n12412 = n12411 ^ n12336 ;
  assign n12413 = ~n12337 & n12412 ;
  assign n12414 = n12413 ^ x76 ;
  assign n12415 = n12414 ^ n12333 ;
  assign n12416 = ~n12334 & n12415 ;
  assign n12417 = n12416 ^ x77 ;
  assign n12320 = n11912 ^ x77 ;
  assign n12321 = n12320 ^ n11998 ;
  assign n12322 = n12321 ^ x76 ;
  assign n12323 = n12322 ^ n12320 ;
  assign n12325 = n11998 ^ x77 ;
  assign n12326 = n12325 ^ n12320 ;
  assign n12327 = ~n12323 & ~n12326 ;
  assign n12328 = n12327 ^ n12320 ;
  assign n12329 = n12195 & ~n12328 ;
  assign n12330 = n12329 ^ n11909 ;
  assign n12418 = n12417 ^ n12330 ;
  assign n12419 = n12417 ^ x78 ;
  assign n12420 = n12418 & n12419 ;
  assign n12421 = n12420 ^ x78 ;
  assign n12317 = n12004 ^ x78 ;
  assign n12318 = n12195 & n12317 ;
  assign n12319 = n12318 ^ n12006 ;
  assign n12422 = n12421 ^ n12319 ;
  assign n12423 = n12421 ^ x79 ;
  assign n12424 = n12422 & n12423 ;
  assign n12425 = n12424 ^ x79 ;
  assign n12315 = n12012 & n12195 ;
  assign n12316 = n12315 ^ n11907 ;
  assign n12426 = n12425 ^ n12316 ;
  assign n12427 = n12425 ^ x80 ;
  assign n12428 = n12426 & n12427 ;
  assign n12429 = n12428 ^ x80 ;
  assign n12313 = n12016 & n12195 ;
  assign n12314 = n12313 ^ n11905 ;
  assign n12430 = n12429 ^ n12314 ;
  assign n12431 = n12429 ^ x81 ;
  assign n12432 = n12430 & n12431 ;
  assign n12433 = n12432 ^ x81 ;
  assign n12311 = n12020 & n12195 ;
  assign n12312 = n12311 ^ n11902 ;
  assign n12434 = n12433 ^ n12312 ;
  assign n12435 = n12433 ^ x82 ;
  assign n12436 = n12434 & n12435 ;
  assign n12437 = n12436 ^ x82 ;
  assign n12309 = n12024 & n12195 ;
  assign n12310 = n12309 ^ n11891 ;
  assign n12438 = n12437 ^ n12310 ;
  assign n12439 = n12437 ^ x83 ;
  assign n12440 = n12438 & n12439 ;
  assign n12441 = n12440 ^ x83 ;
  assign n12307 = n12028 & n12195 ;
  assign n12308 = n12307 ^ n11888 ;
  assign n12442 = n12441 ^ n12308 ;
  assign n12443 = n12441 ^ x84 ;
  assign n12444 = n12442 & n12443 ;
  assign n12445 = n12444 ^ x84 ;
  assign n12305 = n12032 & n12195 ;
  assign n12306 = n12305 ^ n11886 ;
  assign n12446 = n12445 ^ n12306 ;
  assign n12447 = n12445 ^ x85 ;
  assign n12448 = n12446 & n12447 ;
  assign n12449 = n12448 ^ x85 ;
  assign n12303 = n12036 & n12195 ;
  assign n12304 = n12303 ^ n11884 ;
  assign n12450 = n12449 ^ n12304 ;
  assign n12451 = n12449 ^ x86 ;
  assign n12452 = n12450 & n12451 ;
  assign n12453 = n12452 ^ x86 ;
  assign n12454 = n12453 ^ n12301 ;
  assign n12455 = ~n12302 & n12454 ;
  assign n12456 = n12455 ^ x87 ;
  assign n12457 = n12456 ^ n12298 ;
  assign n12458 = ~n12299 & n12457 ;
  assign n12459 = n12458 ^ x88 ;
  assign n12295 = n12048 & n12195 ;
  assign n12296 = n12295 ^ n11878 ;
  assign n12460 = n12459 ^ n12296 ;
  assign n12461 = n12459 ^ x89 ;
  assign n12462 = n12460 & n12461 ;
  assign n12463 = n12462 ^ x89 ;
  assign n12292 = n12050 ^ x89 ;
  assign n12293 = n12195 & n12292 ;
  assign n12294 = n12293 ^ n11875 ;
  assign n12464 = n12463 ^ n12294 ;
  assign n12465 = n12463 ^ x90 ;
  assign n12466 = n12464 & n12465 ;
  assign n12467 = n12466 ^ x90 ;
  assign n12290 = n12054 & n12195 ;
  assign n12291 = n12290 ^ n12056 ;
  assign n12468 = n12467 ^ n12291 ;
  assign n12469 = n12467 ^ x91 ;
  assign n12470 = n12468 & n12469 ;
  assign n12471 = n12470 ^ x91 ;
  assign n12288 = n12061 & n12195 ;
  assign n12289 = n12288 ^ n11873 ;
  assign n12472 = n12471 ^ n12289 ;
  assign n12473 = n12471 ^ x92 ;
  assign n12474 = n12472 & n12473 ;
  assign n12475 = n12474 ^ x92 ;
  assign n12476 = n12475 ^ n12286 ;
  assign n12477 = ~n12287 & n12476 ;
  assign n12478 = n12477 ^ x93 ;
  assign n12479 = n12478 ^ n12283 ;
  assign n12480 = ~n12284 & n12479 ;
  assign n12481 = n12480 ^ x94 ;
  assign n12280 = n12073 & n12195 ;
  assign n12281 = n12280 ^ n11867 ;
  assign n12482 = n12481 ^ n12281 ;
  assign n12483 = n12481 ^ x95 ;
  assign n12484 = n12482 & n12483 ;
  assign n12485 = n12484 ^ x95 ;
  assign n12277 = n12075 ^ x95 ;
  assign n12278 = n12195 & n12277 ;
  assign n12279 = n12278 ^ n11864 ;
  assign n12486 = n12485 ^ n12279 ;
  assign n12487 = n12485 ^ x96 ;
  assign n12488 = n12486 & n12487 ;
  assign n12489 = n12488 ^ x96 ;
  assign n12274 = n12078 ^ x96 ;
  assign n12275 = n12195 & n12274 ;
  assign n12276 = n12275 ^ n11861 ;
  assign n12490 = n12489 ^ n12276 ;
  assign n12491 = n12489 ^ x97 ;
  assign n12492 = n12490 & n12491 ;
  assign n12493 = n12492 ^ x97 ;
  assign n12272 = n12083 & n12195 ;
  assign n12273 = n12272 ^ n11859 ;
  assign n12494 = n12493 ^ n12273 ;
  assign n12495 = n12493 ^ x98 ;
  assign n12496 = n12494 & n12495 ;
  assign n12497 = n12496 ^ x98 ;
  assign n12270 = n12087 & n12195 ;
  assign n12271 = n12270 ^ n11857 ;
  assign n12498 = n12497 ^ n12271 ;
  assign n12499 = n12497 ^ x99 ;
  assign n12500 = n12498 & n12499 ;
  assign n12501 = n12500 ^ x99 ;
  assign n12267 = n12089 ^ x99 ;
  assign n12268 = n12195 & n12267 ;
  assign n12269 = n12268 ^ n11853 ;
  assign n12502 = n12501 ^ n12269 ;
  assign n12503 = n12501 ^ x100 ;
  assign n12504 = n12502 & n12503 ;
  assign n12505 = n12504 ^ x100 ;
  assign n12264 = n12092 ^ x100 ;
  assign n12265 = n12195 & n12264 ;
  assign n12266 = n12265 ^ n11849 ;
  assign n12506 = n12505 ^ n12266 ;
  assign n12507 = n12505 ^ x101 ;
  assign n12508 = n12506 & n12507 ;
  assign n12509 = n12508 ^ x101 ;
  assign n12262 = n12097 & n12195 ;
  assign n12263 = n12262 ^ n11847 ;
  assign n12510 = n12509 ^ n12263 ;
  assign n12511 = n12509 ^ x102 ;
  assign n12512 = n12510 & n12511 ;
  assign n12513 = n12512 ^ x102 ;
  assign n12260 = n12101 & n12195 ;
  assign n12261 = n12260 ^ n11845 ;
  assign n12514 = n12513 ^ n12261 ;
  assign n12515 = n12513 ^ x103 ;
  assign n12516 = n12514 & n12515 ;
  assign n12517 = n12516 ^ x103 ;
  assign n12258 = n12105 & n12195 ;
  assign n12259 = n12258 ^ n11843 ;
  assign n12518 = n12517 ^ n12259 ;
  assign n12519 = n12517 ^ x104 ;
  assign n12520 = n12518 & n12519 ;
  assign n12521 = n12520 ^ x104 ;
  assign n12256 = n12109 & n12195 ;
  assign n12257 = n12256 ^ n11841 ;
  assign n12522 = n12521 ^ n12257 ;
  assign n12523 = n12521 ^ x105 ;
  assign n12524 = n12522 & n12523 ;
  assign n12525 = n12524 ^ x105 ;
  assign n12254 = n12113 & n12195 ;
  assign n12255 = n12254 ^ n11839 ;
  assign n12526 = n12525 ^ n12255 ;
  assign n12527 = n12525 ^ x106 ;
  assign n12528 = n12526 & n12527 ;
  assign n12529 = n12528 ^ x106 ;
  assign n12530 = n12529 ^ n12247 ;
  assign n12531 = n12530 ^ n12252 ;
  assign n12532 = ~n12253 & n12531 ;
  assign n12533 = n12532 ^ n12252 ;
  assign n12534 = ~n12248 & n12533 ;
  assign n12535 = n12534 ^ x108 ;
  assign n12539 = n12538 ^ n12535 ;
  assign n12540 = n12538 ^ x109 ;
  assign n12541 = n12539 & ~n12540 ;
  assign n12542 = n12541 ^ x109 ;
  assign n12235 = n11830 ^ x109 ;
  assign n12236 = n12235 ^ n12123 ;
  assign n12237 = n12236 ^ x108 ;
  assign n12238 = n12237 ^ n12235 ;
  assign n12240 = n12123 ^ x109 ;
  assign n12241 = n12240 ^ n12235 ;
  assign n12242 = ~n12238 & ~n12241 ;
  assign n12243 = n12242 ^ n12235 ;
  assign n12244 = n12195 & ~n12243 ;
  assign n12245 = n12244 ^ n11826 ;
  assign n12543 = n12542 ^ n12245 ;
  assign n12544 = n12542 ^ x110 ;
  assign n12545 = n12543 & n12544 ;
  assign n12546 = n12545 ^ x110 ;
  assign n12232 = n12129 ^ x110 ;
  assign n12233 = n12195 & n12232 ;
  assign n12234 = n12233 ^ n12132 ;
  assign n12547 = n12546 ^ n12234 ;
  assign n12548 = n12546 ^ x111 ;
  assign n12549 = n12547 & n12548 ;
  assign n12550 = n12549 ^ x111 ;
  assign n12229 = n12136 ^ x111 ;
  assign n12230 = n12195 & n12229 ;
  assign n12231 = n12230 ^ n12138 ;
  assign n12551 = n12550 ^ n12231 ;
  assign n12552 = n12550 ^ x112 ;
  assign n12553 = n12551 & n12552 ;
  assign n12554 = n12553 ^ x112 ;
  assign n12226 = n12142 ^ x112 ;
  assign n12227 = n12195 & n12226 ;
  assign n12228 = n12227 ^ n11812 ;
  assign n12555 = n12554 ^ n12228 ;
  assign n12556 = n12554 ^ x113 ;
  assign n12557 = n12555 & n12556 ;
  assign n12558 = n12557 ^ x113 ;
  assign n12215 = n11812 ^ x113 ;
  assign n12216 = n12215 ^ n12142 ;
  assign n12217 = n12216 ^ x112 ;
  assign n12218 = n12217 ^ n12215 ;
  assign n12220 = n12142 ^ x113 ;
  assign n12221 = n12220 ^ n12215 ;
  assign n12222 = ~n12218 & ~n12221 ;
  assign n12223 = n12222 ^ n12215 ;
  assign n12224 = n12195 & ~n12223 ;
  assign n12225 = n12224 ^ n11809 ;
  assign n12559 = n12558 ^ n12225 ;
  assign n12560 = n12558 ^ x114 ;
  assign n12561 = n12559 & n12560 ;
  assign n12562 = n12561 ^ x114 ;
  assign n12563 = n12562 ^ n12213 ;
  assign n12564 = ~n12214 & n12563 ;
  assign n12565 = n12564 ^ x115 ;
  assign n12209 = n12156 & n12195 ;
  assign n12210 = n12209 ^ n11807 ;
  assign n12566 = n12565 ^ n12210 ;
  assign n12567 = n12565 ^ x116 ;
  assign n12568 = n12566 & n12567 ;
  assign n12569 = n12568 ^ x116 ;
  assign n12207 = n12160 & n12195 ;
  assign n12208 = n12207 ^ n11805 ;
  assign n12570 = n12569 ^ n12208 ;
  assign n12571 = n12569 ^ x117 ;
  assign n12572 = n12570 & n12571 ;
  assign n12573 = n12572 ^ x117 ;
  assign n12574 = n12573 ^ n12205 ;
  assign n12575 = ~n12206 & n12574 ;
  assign n12576 = n12575 ^ x118 ;
  assign n12577 = n12576 ^ n12202 ;
  assign n12578 = ~n12203 & n12577 ;
  assign n12579 = n12578 ^ x119 ;
  assign n12580 = n12579 ^ n12199 ;
  assign n12581 = ~n12200 & n12580 ;
  assign n12582 = n12581 ^ x120 ;
  assign n12196 = n12179 & n12195 ;
  assign n12197 = n12196 ^ n11799 ;
  assign n12583 = n12582 ^ n12197 ;
  assign n12584 = n12582 ^ x121 ;
  assign n12585 = n12583 & n12584 ;
  assign n12586 = n12585 ^ x121 ;
  assign n12957 = n12956 ^ n12586 ;
  assign n12958 = n12957 ^ n133 ;
  assign n12959 = n12958 ^ n132 ;
  assign n12960 = n12959 ^ n10978 ;
  assign n12961 = n12960 ^ n12959 ;
  assign n12964 = ~n133 & n12961 ;
  assign n12965 = n12964 ^ n12959 ;
  assign n12966 = ~n12956 & n12965 ;
  assign n12967 = ~n12957 & ~n12966 ;
  assign n12968 = n12966 ^ n12959 ;
  assign n12969 = n12968 ^ n12586 ;
  assign n12970 = n12967 & n12969 ;
  assign n12971 = n12970 ^ n12968 ;
  assign n12972 = n12971 ^ x123 ;
  assign n11400 = x122 & ~n11399 ;
  assign n12187 = n133 & n12186 ;
  assign n12188 = ~n12182 & n12187 ;
  assign n12587 = n132 & ~n12586 ;
  assign n12588 = ~n12188 & n12587 ;
  assign n12591 = n11400 & n12588 ;
  assign n12589 = n12588 ^ n12188 ;
  assign n12592 = n12591 ^ n12589 ;
  assign n12600 = n12560 & n12592 ;
  assign n12601 = n12600 ^ n12225 ;
  assign n12602 = n12601 ^ x115 ;
  assign n12603 = n12556 & n12592 ;
  assign n12604 = n12603 ^ n12228 ;
  assign n12605 = n12604 ^ x114 ;
  assign n12926 = n12548 & n12592 ;
  assign n12927 = n12926 ^ n12234 ;
  assign n12920 = n12544 & n12592 ;
  assign n12921 = n12920 ^ n12245 ;
  assign n12913 = n12535 ^ x109 ;
  assign n12914 = n12592 & n12913 ;
  assign n12915 = n12914 ^ n12538 ;
  assign n12608 = n12250 ^ x108 ;
  assign n12609 = n12608 ^ n12529 ;
  assign n12610 = n12609 ^ x107 ;
  assign n12611 = n12610 ^ n12608 ;
  assign n12613 = n12529 ^ x108 ;
  assign n12614 = n12613 ^ n12608 ;
  assign n12615 = ~n12611 & ~n12614 ;
  assign n12616 = n12615 ^ n12608 ;
  assign n12617 = n12592 & ~n12616 ;
  assign n12618 = n12617 ^ n12247 ;
  assign n12619 = n12618 ^ x109 ;
  assign n12624 = n12618 ^ x108 ;
  assign n12620 = n12529 ^ x107 ;
  assign n12621 = n12592 & n12620 ;
  assign n12622 = n12621 ^ n12250 ;
  assign n12623 = n12622 ^ n12618 ;
  assign n12625 = n12624 ^ n12623 ;
  assign n12638 = n12503 & n12592 ;
  assign n12639 = n12638 ^ n12269 ;
  assign n12640 = n12639 ^ x101 ;
  assign n12641 = n12499 & n12592 ;
  assign n12642 = n12641 ^ n12271 ;
  assign n12643 = n12642 ^ x100 ;
  assign n12854 = n12478 ^ x94 ;
  assign n12855 = n12592 & n12854 ;
  assign n12856 = n12855 ^ n12283 ;
  assign n12847 = n12475 ^ x93 ;
  assign n12848 = n12592 & n12847 ;
  assign n12849 = n12848 ^ n12286 ;
  assign n12841 = n12473 & n12592 ;
  assign n12842 = n12841 ^ n12289 ;
  assign n12652 = n12469 & n12592 ;
  assign n12653 = n12652 ^ n12291 ;
  assign n12654 = n12653 ^ x92 ;
  assign n12658 = n12653 ^ x91 ;
  assign n12655 = n12465 & n12592 ;
  assign n12656 = n12655 ^ n12294 ;
  assign n12657 = n12656 ^ n12653 ;
  assign n12659 = n12658 ^ n12657 ;
  assign n12813 = n12447 & n12592 ;
  assign n12814 = n12813 ^ n12306 ;
  assign n12670 = n12443 & n12592 ;
  assign n12671 = n12670 ^ n12308 ;
  assign n12672 = n12671 ^ x85 ;
  assign n12676 = n12671 ^ x84 ;
  assign n12673 = n12439 & n12592 ;
  assign n12674 = n12673 ^ n12310 ;
  assign n12675 = n12674 ^ n12671 ;
  assign n12677 = n12676 ^ n12675 ;
  assign n12678 = n12435 & n12592 ;
  assign n12679 = n12678 ^ n12312 ;
  assign n12680 = n12679 ^ x83 ;
  assign n12684 = n12679 ^ x82 ;
  assign n12681 = n12431 & n12592 ;
  assign n12682 = n12681 ^ n12314 ;
  assign n12683 = n12682 ^ n12679 ;
  assign n12685 = n12684 ^ n12683 ;
  assign n12686 = n12427 & n12592 ;
  assign n12687 = n12686 ^ n12316 ;
  assign n12688 = n12687 ^ x81 ;
  assign n12689 = n12423 & n12592 ;
  assign n12690 = n12689 ^ n12319 ;
  assign n12691 = n12690 ^ x80 ;
  assign n12704 = n12401 & n12592 ;
  assign n12705 = n12704 ^ n12343 ;
  assign n12706 = n12705 ^ x74 ;
  assign n12707 = n12397 & n12592 ;
  assign n12708 = n12707 ^ n12345 ;
  assign n12709 = n12708 ^ x73 ;
  assign n12727 = x65 & n12592 ;
  assign n12725 = n12371 ^ x6 ;
  assign n12723 = n12592 ^ n12195 ;
  assign n12724 = n12364 & n12723 ;
  assign n12726 = n12725 ^ n12724 ;
  assign n12728 = n12727 ^ n12726 ;
  assign n12729 = n12728 ^ x66 ;
  assign n12735 = x5 & x65 ;
  assign n12730 = x65 ^ x4 ;
  assign n12731 = x64 ^ x5 ;
  assign n12732 = n12731 ^ x65 ;
  assign n12733 = n12732 ^ n12592 ;
  assign n12734 = ~n12730 & n12733 ;
  assign n12736 = n12735 ^ n12734 ;
  assign n12737 = n12732 ^ x65 ;
  assign n12738 = n12737 ^ x5 ;
  assign n12739 = n12736 & n12738 ;
  assign n12740 = n12739 ^ n12735 ;
  assign n12741 = n12740 ^ x65 ;
  assign n12742 = n12741 ^ n12728 ;
  assign n12743 = ~n12729 & n12742 ;
  assign n12744 = n12743 ^ x66 ;
  assign n12720 = n12372 ^ x66 ;
  assign n12721 = n12592 & ~n12720 ;
  assign n12722 = n12721 ^ n12362 ;
  assign n12745 = n12744 ^ n12722 ;
  assign n12746 = n12744 ^ x67 ;
  assign n12747 = n12745 & n12746 ;
  assign n12748 = n12747 ^ x67 ;
  assign n12718 = n12377 & n12592 ;
  assign n12719 = n12718 ^ n12356 ;
  assign n12749 = n12748 ^ n12719 ;
  assign n12750 = n12748 ^ x68 ;
  assign n12751 = n12749 & n12750 ;
  assign n12752 = n12751 ^ x68 ;
  assign n12716 = n12381 & n12592 ;
  assign n12717 = n12716 ^ n12353 ;
  assign n12753 = n12752 ^ n12717 ;
  assign n12754 = n12752 ^ x69 ;
  assign n12755 = n12753 & n12754 ;
  assign n12756 = n12755 ^ x69 ;
  assign n12714 = n12385 & n12592 ;
  assign n12715 = n12714 ^ n12351 ;
  assign n12757 = n12756 ^ n12715 ;
  assign n12758 = n12756 ^ x70 ;
  assign n12759 = n12757 & n12758 ;
  assign n12760 = n12759 ^ x70 ;
  assign n12712 = n12389 & n12592 ;
  assign n12713 = n12712 ^ n12349 ;
  assign n12761 = n12760 ^ n12713 ;
  assign n12762 = n12760 ^ x71 ;
  assign n12763 = n12761 & n12762 ;
  assign n12764 = n12763 ^ x71 ;
  assign n12710 = n12393 & n12592 ;
  assign n12711 = n12710 ^ n12347 ;
  assign n12765 = n12764 ^ n12711 ;
  assign n12766 = n12764 ^ x72 ;
  assign n12767 = n12765 & n12766 ;
  assign n12768 = n12767 ^ x72 ;
  assign n12769 = n12768 ^ n12708 ;
  assign n12770 = ~n12709 & n12769 ;
  assign n12771 = n12770 ^ x73 ;
  assign n12772 = n12771 ^ n12705 ;
  assign n12773 = ~n12706 & n12772 ;
  assign n12774 = n12773 ^ x74 ;
  assign n12702 = n12405 & n12592 ;
  assign n12703 = n12702 ^ n12341 ;
  assign n12775 = n12774 ^ n12703 ;
  assign n12776 = n12774 ^ x75 ;
  assign n12777 = n12775 & n12776 ;
  assign n12778 = n12777 ^ x75 ;
  assign n12700 = n12409 & n12592 ;
  assign n12701 = n12700 ^ n12339 ;
  assign n12779 = n12778 ^ n12701 ;
  assign n12780 = n12778 ^ x76 ;
  assign n12781 = n12779 & n12780 ;
  assign n12782 = n12781 ^ x76 ;
  assign n12697 = n12411 ^ x76 ;
  assign n12698 = n12592 & n12697 ;
  assign n12699 = n12698 ^ n12336 ;
  assign n12783 = n12782 ^ n12699 ;
  assign n12784 = n12782 ^ x77 ;
  assign n12785 = n12783 & n12784 ;
  assign n12786 = n12785 ^ x77 ;
  assign n12694 = n12414 ^ x77 ;
  assign n12695 = n12592 & n12694 ;
  assign n12696 = n12695 ^ n12333 ;
  assign n12787 = n12786 ^ n12696 ;
  assign n12788 = n12786 ^ x78 ;
  assign n12789 = n12787 & n12788 ;
  assign n12790 = n12789 ^ x78 ;
  assign n12692 = n12419 & n12592 ;
  assign n12693 = n12692 ^ n12330 ;
  assign n12791 = n12790 ^ n12693 ;
  assign n12792 = n12790 ^ x79 ;
  assign n12793 = n12791 & n12792 ;
  assign n12794 = n12793 ^ x79 ;
  assign n12795 = n12794 ^ n12690 ;
  assign n12796 = ~n12691 & n12795 ;
  assign n12797 = n12796 ^ x80 ;
  assign n12798 = n12797 ^ n12687 ;
  assign n12799 = ~n12688 & n12798 ;
  assign n12800 = n12799 ^ x81 ;
  assign n12801 = n12800 ^ n12679 ;
  assign n12802 = n12801 ^ n12684 ;
  assign n12803 = ~n12685 & n12802 ;
  assign n12804 = n12803 ^ n12684 ;
  assign n12805 = ~n12680 & n12804 ;
  assign n12806 = n12805 ^ x83 ;
  assign n12807 = n12806 ^ n12671 ;
  assign n12808 = n12807 ^ n12676 ;
  assign n12809 = ~n12677 & n12808 ;
  assign n12810 = n12809 ^ n12676 ;
  assign n12811 = ~n12672 & n12810 ;
  assign n12812 = n12811 ^ x85 ;
  assign n12815 = n12814 ^ n12812 ;
  assign n12816 = n12814 ^ x86 ;
  assign n12817 = n12815 & ~n12816 ;
  assign n12818 = n12817 ^ x86 ;
  assign n12668 = n12451 & n12592 ;
  assign n12669 = n12668 ^ n12304 ;
  assign n12819 = n12818 ^ n12669 ;
  assign n12820 = n12818 ^ x87 ;
  assign n12821 = n12819 & n12820 ;
  assign n12822 = n12821 ^ x87 ;
  assign n12665 = n12453 ^ x87 ;
  assign n12666 = n12592 & n12665 ;
  assign n12667 = n12666 ^ n12301 ;
  assign n12823 = n12822 ^ n12667 ;
  assign n12824 = n12822 ^ x88 ;
  assign n12825 = n12823 & n12824 ;
  assign n12826 = n12825 ^ x88 ;
  assign n12662 = n12456 ^ x88 ;
  assign n12663 = n12592 & n12662 ;
  assign n12664 = n12663 ^ n12298 ;
  assign n12827 = n12826 ^ n12664 ;
  assign n12828 = n12826 ^ x89 ;
  assign n12829 = n12827 & n12828 ;
  assign n12830 = n12829 ^ x89 ;
  assign n12660 = n12461 & n12592 ;
  assign n12661 = n12660 ^ n12296 ;
  assign n12831 = n12830 ^ n12661 ;
  assign n12832 = n12830 ^ x90 ;
  assign n12833 = n12831 & n12832 ;
  assign n12834 = n12833 ^ x90 ;
  assign n12835 = n12834 ^ n12653 ;
  assign n12836 = n12835 ^ n12658 ;
  assign n12837 = ~n12659 & n12836 ;
  assign n12838 = n12837 ^ n12658 ;
  assign n12839 = ~n12654 & n12838 ;
  assign n12840 = n12839 ^ x92 ;
  assign n12843 = n12842 ^ n12840 ;
  assign n12844 = n12842 ^ x93 ;
  assign n12845 = n12843 & ~n12844 ;
  assign n12846 = n12845 ^ x93 ;
  assign n12850 = n12849 ^ n12846 ;
  assign n12851 = n12849 ^ x94 ;
  assign n12852 = n12850 & ~n12851 ;
  assign n12853 = n12852 ^ x94 ;
  assign n12857 = n12856 ^ n12853 ;
  assign n12858 = n12856 ^ x95 ;
  assign n12859 = n12857 & ~n12858 ;
  assign n12860 = n12859 ^ x95 ;
  assign n12650 = n12483 & n12592 ;
  assign n12651 = n12650 ^ n12281 ;
  assign n12861 = n12860 ^ n12651 ;
  assign n12862 = n12860 ^ x96 ;
  assign n12863 = n12861 & n12862 ;
  assign n12864 = n12863 ^ x96 ;
  assign n12648 = n12487 & n12592 ;
  assign n12649 = n12648 ^ n12279 ;
  assign n12865 = n12864 ^ n12649 ;
  assign n12866 = n12864 ^ x97 ;
  assign n12867 = n12865 & n12866 ;
  assign n12868 = n12867 ^ x97 ;
  assign n12646 = n12491 & n12592 ;
  assign n12647 = n12646 ^ n12276 ;
  assign n12869 = n12868 ^ n12647 ;
  assign n12870 = n12868 ^ x98 ;
  assign n12871 = n12869 & n12870 ;
  assign n12872 = n12871 ^ x98 ;
  assign n12644 = n12495 & n12592 ;
  assign n12645 = n12644 ^ n12273 ;
  assign n12873 = n12872 ^ n12645 ;
  assign n12874 = n12872 ^ x99 ;
  assign n12875 = n12873 & n12874 ;
  assign n12876 = n12875 ^ x99 ;
  assign n12877 = n12876 ^ n12642 ;
  assign n12878 = ~n12643 & n12877 ;
  assign n12879 = n12878 ^ x100 ;
  assign n12880 = n12879 ^ n12639 ;
  assign n12881 = ~n12640 & n12880 ;
  assign n12882 = n12881 ^ x101 ;
  assign n12636 = n12507 & n12592 ;
  assign n12637 = n12636 ^ n12266 ;
  assign n12883 = n12882 ^ n12637 ;
  assign n12884 = n12882 ^ x102 ;
  assign n12885 = n12883 & n12884 ;
  assign n12886 = n12885 ^ x102 ;
  assign n12634 = n12511 & n12592 ;
  assign n12635 = n12634 ^ n12263 ;
  assign n12887 = n12886 ^ n12635 ;
  assign n12888 = n12886 ^ x103 ;
  assign n12889 = n12887 & n12888 ;
  assign n12890 = n12889 ^ x103 ;
  assign n12632 = n12515 & n12592 ;
  assign n12633 = n12632 ^ n12261 ;
  assign n12891 = n12890 ^ n12633 ;
  assign n12892 = n12890 ^ x104 ;
  assign n12893 = n12891 & n12892 ;
  assign n12894 = n12893 ^ x104 ;
  assign n12630 = n12519 & n12592 ;
  assign n12631 = n12630 ^ n12259 ;
  assign n12895 = n12894 ^ n12631 ;
  assign n12896 = n12894 ^ x105 ;
  assign n12897 = n12895 & n12896 ;
  assign n12898 = n12897 ^ x105 ;
  assign n12628 = n12523 & n12592 ;
  assign n12629 = n12628 ^ n12257 ;
  assign n12899 = n12898 ^ n12629 ;
  assign n12900 = n12898 ^ x106 ;
  assign n12901 = n12899 & n12900 ;
  assign n12902 = n12901 ^ x106 ;
  assign n12626 = n12527 & n12592 ;
  assign n12627 = n12626 ^ n12255 ;
  assign n12903 = n12902 ^ n12627 ;
  assign n12904 = n12902 ^ x107 ;
  assign n12905 = n12903 & n12904 ;
  assign n12906 = n12905 ^ x107 ;
  assign n12907 = n12906 ^ n12618 ;
  assign n12908 = n12907 ^ n12624 ;
  assign n12909 = ~n12625 & n12908 ;
  assign n12910 = n12909 ^ n12624 ;
  assign n12911 = ~n12619 & n12910 ;
  assign n12912 = n12911 ^ x109 ;
  assign n12916 = n12915 ^ n12912 ;
  assign n12917 = n12915 ^ x110 ;
  assign n12918 = n12916 & ~n12917 ;
  assign n12919 = n12918 ^ x110 ;
  assign n12922 = n12921 ^ n12919 ;
  assign n12923 = n12921 ^ x111 ;
  assign n12924 = n12922 & ~n12923 ;
  assign n12925 = n12924 ^ x111 ;
  assign n12928 = n12927 ^ n12925 ;
  assign n12929 = n12927 ^ x112 ;
  assign n12930 = n12928 & ~n12929 ;
  assign n12931 = n12930 ^ x112 ;
  assign n12606 = n12552 & n12592 ;
  assign n12607 = n12606 ^ n12231 ;
  assign n12932 = n12931 ^ n12607 ;
  assign n12933 = n12931 ^ x113 ;
  assign n12934 = n12932 & n12933 ;
  assign n12935 = n12934 ^ x113 ;
  assign n12936 = n12935 ^ n12604 ;
  assign n12937 = ~n12605 & n12936 ;
  assign n12938 = n12937 ^ x114 ;
  assign n12939 = n12938 ^ n12601 ;
  assign n12940 = ~n12602 & n12939 ;
  assign n12941 = n12940 ^ x115 ;
  assign n12597 = n12562 ^ x115 ;
  assign n12598 = n12592 & n12597 ;
  assign n12599 = n12598 ^ n12213 ;
  assign n12942 = n12941 ^ n12599 ;
  assign n12943 = n12941 ^ x116 ;
  assign n12944 = n12942 & n12943 ;
  assign n12945 = n12944 ^ x116 ;
  assign n12595 = n12567 & n12592 ;
  assign n12596 = n12595 ^ n12210 ;
  assign n12946 = n12945 ^ n12596 ;
  assign n12947 = n12945 ^ x117 ;
  assign n12948 = n12946 & n12947 ;
  assign n12949 = n12948 ^ x117 ;
  assign n12593 = n12571 & n12592 ;
  assign n12594 = n12593 ^ n12208 ;
  assign n12950 = n12949 ^ n12594 ;
  assign n12951 = n12949 ^ x118 ;
  assign n12952 = n12950 & n12951 ;
  assign n12953 = n12952 ^ x118 ;
  assign n12954 = n12953 ^ x119 ;
  assign n12981 = n12573 ^ x118 ;
  assign n12982 = n12592 & n12981 ;
  assign n12983 = n12982 ^ n12205 ;
  assign n12984 = n12983 ^ n12953 ;
  assign n12985 = n12954 & n12984 ;
  assign n12986 = n12985 ^ x119 ;
  assign n12978 = n12576 ^ x119 ;
  assign n12979 = n12592 & n12978 ;
  assign n12980 = n12979 ^ n12202 ;
  assign n12987 = n12986 ^ n12980 ;
  assign n12988 = n12986 ^ x120 ;
  assign n12989 = n12987 & n12988 ;
  assign n12990 = n12989 ^ x120 ;
  assign n12975 = n12579 ^ x120 ;
  assign n12976 = n12592 & n12975 ;
  assign n12977 = n12976 ^ n12199 ;
  assign n12991 = n12990 ^ n12977 ;
  assign n12992 = n12990 ^ x121 ;
  assign n12993 = n12991 & n12992 ;
  assign n12994 = n12993 ^ x121 ;
  assign n12973 = n12584 & n12592 ;
  assign n12974 = n12973 ^ n12197 ;
  assign n12995 = n12994 ^ n12974 ;
  assign n12998 = n12974 ^ x122 ;
  assign n12999 = n12995 & ~n12998 ;
  assign n12996 = x123 ^ x122 ;
  assign n13000 = n12999 ^ n12996 ;
  assign n13003 = ~n12972 & n13000 ;
  assign n13004 = n13003 ^ x123 ;
  assign n13005 = n131 & ~n13004 ;
  assign n13174 = x64 & n13005 ;
  assign n13175 = n13174 ^ x4 ;
  assign n13614 = ~x3 & x65 ;
  assign n13615 = n13175 & ~n13614 ;
  assign n13022 = n12925 ^ x112 ;
  assign n13023 = n13005 & n13022 ;
  assign n13024 = n13023 ^ n12927 ;
  assign n13025 = n13024 ^ x113 ;
  assign n13026 = n12919 ^ x111 ;
  assign n13027 = n13005 & n13026 ;
  assign n13028 = n13027 ^ n12921 ;
  assign n13029 = n13028 ^ x112 ;
  assign n13324 = n12862 & n13005 ;
  assign n13325 = n13324 ^ n12651 ;
  assign n13071 = n12853 ^ x95 ;
  assign n13072 = n13005 & n13071 ;
  assign n13073 = n13072 ^ n12856 ;
  assign n13074 = n13073 ^ x96 ;
  assign n13079 = n13073 ^ x95 ;
  assign n13075 = n12846 ^ x94 ;
  assign n13076 = n13005 & n13075 ;
  assign n13077 = n13076 ^ n12849 ;
  assign n13078 = n13077 ^ n13073 ;
  assign n13080 = n13079 ^ n13078 ;
  assign n13296 = n12828 & n13005 ;
  assign n13297 = n13296 ^ n12664 ;
  assign n13100 = n12824 & n13005 ;
  assign n13101 = n13100 ^ n12667 ;
  assign n13102 = n13101 ^ x89 ;
  assign n13106 = n13101 ^ x88 ;
  assign n13103 = n12820 & n13005 ;
  assign n13104 = n13103 ^ n12669 ;
  assign n13105 = n13104 ^ n13101 ;
  assign n13107 = n13106 ^ n13105 ;
  assign n13240 = n12776 & n13005 ;
  assign n13241 = n13240 ^ n12703 ;
  assign n13153 = n12771 ^ x74 ;
  assign n13154 = n13005 & n13153 ;
  assign n13155 = n13154 ^ n12705 ;
  assign n13156 = n13155 ^ x75 ;
  assign n13161 = n13155 ^ x74 ;
  assign n13157 = n12768 ^ x73 ;
  assign n13158 = n13005 & n13157 ;
  assign n13159 = n13158 ^ n12708 ;
  assign n13160 = n13159 ^ n13155 ;
  assign n13162 = n13161 ^ n13160 ;
  assign n13208 = n12746 & n13005 ;
  assign n13209 = n13208 ^ n12722 ;
  assign n13201 = n12741 ^ x66 ;
  assign n13202 = n13005 & n13201 ;
  assign n13203 = n13202 ^ n12728 ;
  assign n13182 = ~x4 & x65 ;
  assign n13183 = n13182 ^ x64 ;
  assign n13184 = n13005 & ~n13183 ;
  assign n13185 = n13184 ^ n12592 ;
  assign n13193 = n13185 ^ x5 ;
  assign n13194 = n13193 ^ n13005 ;
  assign n13190 = ~x65 & n13005 ;
  assign n13191 = n13190 ^ n13185 ;
  assign n13192 = ~x64 & n13191 ;
  assign n13195 = n13194 ^ n13192 ;
  assign n13180 = x4 & n3646 ;
  assign n13181 = n13005 & n13180 ;
  assign n13196 = n13195 ^ n13181 ;
  assign n13173 = ~x3 & x64 ;
  assign n13176 = n13175 ^ n13173 ;
  assign n13177 = n13175 ^ x65 ;
  assign n13178 = n13176 & ~n13177 ;
  assign n13179 = n13178 ^ x65 ;
  assign n13197 = n13196 ^ n13179 ;
  assign n13198 = n13196 ^ x66 ;
  assign n13199 = n13197 & ~n13198 ;
  assign n13200 = n13199 ^ x66 ;
  assign n13204 = n13203 ^ n13200 ;
  assign n13205 = n13203 ^ x67 ;
  assign n13206 = n13204 & ~n13205 ;
  assign n13207 = n13206 ^ x67 ;
  assign n13210 = n13209 ^ n13207 ;
  assign n13211 = n13209 ^ x68 ;
  assign n13212 = n13210 & ~n13211 ;
  assign n13213 = n13212 ^ x68 ;
  assign n13171 = n12750 & n13005 ;
  assign n13172 = n13171 ^ n12719 ;
  assign n13214 = n13213 ^ n13172 ;
  assign n13215 = n13213 ^ x69 ;
  assign n13216 = n13214 & n13215 ;
  assign n13217 = n13216 ^ x69 ;
  assign n13169 = n12754 & n13005 ;
  assign n13170 = n13169 ^ n12717 ;
  assign n13218 = n13217 ^ n13170 ;
  assign n13219 = n13217 ^ x70 ;
  assign n13220 = n13218 & n13219 ;
  assign n13221 = n13220 ^ x70 ;
  assign n13167 = n12758 & n13005 ;
  assign n13168 = n13167 ^ n12715 ;
  assign n13222 = n13221 ^ n13168 ;
  assign n13223 = n13221 ^ x71 ;
  assign n13224 = n13222 & n13223 ;
  assign n13225 = n13224 ^ x71 ;
  assign n13165 = n12762 & n13005 ;
  assign n13166 = n13165 ^ n12713 ;
  assign n13226 = n13225 ^ n13166 ;
  assign n13227 = n13225 ^ x72 ;
  assign n13228 = n13226 & n13227 ;
  assign n13229 = n13228 ^ x72 ;
  assign n13163 = n12766 & n13005 ;
  assign n13164 = n13163 ^ n12711 ;
  assign n13230 = n13229 ^ n13164 ;
  assign n13231 = n13229 ^ x73 ;
  assign n13232 = n13230 & n13231 ;
  assign n13233 = n13232 ^ x73 ;
  assign n13234 = n13233 ^ n13155 ;
  assign n13235 = n13234 ^ n13161 ;
  assign n13236 = ~n13162 & n13235 ;
  assign n13237 = n13236 ^ n13161 ;
  assign n13238 = ~n13156 & n13237 ;
  assign n13239 = n13238 ^ x75 ;
  assign n13242 = n13241 ^ n13239 ;
  assign n13243 = n13241 ^ x76 ;
  assign n13244 = n13242 & ~n13243 ;
  assign n13245 = n13244 ^ x76 ;
  assign n13151 = n12780 & n13005 ;
  assign n13152 = n13151 ^ n12701 ;
  assign n13246 = n13245 ^ n13152 ;
  assign n13247 = n13245 ^ x77 ;
  assign n13248 = n13246 & n13247 ;
  assign n13249 = n13248 ^ x77 ;
  assign n13149 = n12784 & n13005 ;
  assign n13150 = n13149 ^ n12699 ;
  assign n13250 = n13249 ^ n13150 ;
  assign n13251 = n13249 ^ x78 ;
  assign n13252 = n13250 & n13251 ;
  assign n13253 = n13252 ^ x78 ;
  assign n13147 = n12788 & n13005 ;
  assign n13148 = n13147 ^ n12696 ;
  assign n13254 = n13253 ^ n13148 ;
  assign n13255 = n13253 ^ x79 ;
  assign n13256 = n13254 & n13255 ;
  assign n13257 = n13256 ^ x79 ;
  assign n13145 = n12792 & n13005 ;
  assign n13146 = n13145 ^ n12693 ;
  assign n13258 = n13257 ^ n13146 ;
  assign n13259 = n13257 ^ x80 ;
  assign n13260 = n13258 & n13259 ;
  assign n13261 = n13260 ^ x80 ;
  assign n13142 = n12794 ^ x80 ;
  assign n13143 = n13005 & n13142 ;
  assign n13144 = n13143 ^ n12690 ;
  assign n13262 = n13261 ^ n13144 ;
  assign n13263 = n13261 ^ x81 ;
  assign n13264 = n13262 & n13263 ;
  assign n13265 = n13264 ^ x81 ;
  assign n13139 = n12797 ^ x81 ;
  assign n13140 = n13005 & n13139 ;
  assign n13141 = n13140 ^ n12687 ;
  assign n13266 = n13265 ^ n13141 ;
  assign n13267 = n13265 ^ x82 ;
  assign n13268 = n13266 & n13267 ;
  assign n13269 = n13268 ^ x82 ;
  assign n13136 = n12800 ^ x82 ;
  assign n13137 = n13005 & n13136 ;
  assign n13138 = n13137 ^ n12682 ;
  assign n13270 = n13269 ^ n13138 ;
  assign n13271 = n13269 ^ x83 ;
  assign n13272 = n13270 & n13271 ;
  assign n13273 = n13272 ^ x83 ;
  assign n13125 = n12682 ^ x83 ;
  assign n13126 = n13125 ^ n12800 ;
  assign n13127 = n13126 ^ x82 ;
  assign n13128 = n13127 ^ n13125 ;
  assign n13129 = n13125 ^ n12682 ;
  assign n13130 = n13129 ^ n12800 ;
  assign n13131 = n13130 ^ n13125 ;
  assign n13132 = ~n13128 & ~n13131 ;
  assign n13133 = n13132 ^ n13125 ;
  assign n13134 = n13005 & ~n13133 ;
  assign n13135 = n13134 ^ n12679 ;
  assign n13274 = n13273 ^ n13135 ;
  assign n13275 = n13273 ^ x84 ;
  assign n13276 = n13274 & n13275 ;
  assign n13277 = n13276 ^ x84 ;
  assign n13122 = n12806 ^ x84 ;
  assign n13123 = n13005 & n13122 ;
  assign n13124 = n13123 ^ n12674 ;
  assign n13278 = n13277 ^ n13124 ;
  assign n13279 = n13277 ^ x85 ;
  assign n13280 = n13278 & n13279 ;
  assign n13281 = n13280 ^ x85 ;
  assign n13111 = n12674 ^ x85 ;
  assign n13112 = n13111 ^ n12806 ;
  assign n13113 = n13112 ^ x84 ;
  assign n13114 = n13113 ^ n13111 ;
  assign n13116 = n12806 ^ x85 ;
  assign n13117 = n13116 ^ n13111 ;
  assign n13118 = ~n13114 & ~n13117 ;
  assign n13119 = n13118 ^ n13111 ;
  assign n13120 = n13005 & ~n13119 ;
  assign n13121 = n13120 ^ n12671 ;
  assign n13282 = n13281 ^ n13121 ;
  assign n13283 = n13281 ^ x86 ;
  assign n13284 = n13282 & n13283 ;
  assign n13285 = n13284 ^ x86 ;
  assign n13108 = n12812 ^ x86 ;
  assign n13109 = n13005 & n13108 ;
  assign n13110 = n13109 ^ n12814 ;
  assign n13286 = n13285 ^ n13110 ;
  assign n13287 = n13285 ^ x87 ;
  assign n13288 = n13286 & n13287 ;
  assign n13289 = n13288 ^ x87 ;
  assign n13290 = n13289 ^ n13101 ;
  assign n13291 = n13290 ^ n13106 ;
  assign n13292 = ~n13107 & n13291 ;
  assign n13293 = n13292 ^ n13106 ;
  assign n13294 = ~n13102 & n13293 ;
  assign n13295 = n13294 ^ x89 ;
  assign n13298 = n13297 ^ n13295 ;
  assign n13299 = n13297 ^ x90 ;
  assign n13300 = n13298 & ~n13299 ;
  assign n13301 = n13300 ^ x90 ;
  assign n13098 = n12832 & n13005 ;
  assign n13099 = n13098 ^ n12661 ;
  assign n13302 = n13301 ^ n13099 ;
  assign n13303 = n13301 ^ x91 ;
  assign n13304 = n13302 & n13303 ;
  assign n13305 = n13304 ^ x91 ;
  assign n13095 = n12834 ^ x91 ;
  assign n13096 = n13005 & n13095 ;
  assign n13097 = n13096 ^ n12656 ;
  assign n13306 = n13305 ^ n13097 ;
  assign n13307 = n13305 ^ x92 ;
  assign n13308 = n13306 & n13307 ;
  assign n13309 = n13308 ^ x92 ;
  assign n13084 = n12656 ^ x92 ;
  assign n13085 = n13084 ^ n12834 ;
  assign n13086 = n13085 ^ x91 ;
  assign n13087 = n13086 ^ n13084 ;
  assign n13089 = n12834 ^ x92 ;
  assign n13090 = n13089 ^ n13084 ;
  assign n13091 = ~n13087 & ~n13090 ;
  assign n13092 = n13091 ^ n13084 ;
  assign n13093 = n13005 & ~n13092 ;
  assign n13094 = n13093 ^ n12653 ;
  assign n13310 = n13309 ^ n13094 ;
  assign n13311 = n13309 ^ x93 ;
  assign n13312 = n13310 & n13311 ;
  assign n13313 = n13312 ^ x93 ;
  assign n13081 = n12840 ^ x93 ;
  assign n13082 = n13005 & n13081 ;
  assign n13083 = n13082 ^ n12842 ;
  assign n13314 = n13313 ^ n13083 ;
  assign n13315 = n13313 ^ x94 ;
  assign n13316 = n13314 & n13315 ;
  assign n13317 = n13316 ^ x94 ;
  assign n13318 = n13317 ^ n13073 ;
  assign n13319 = n13318 ^ n13079 ;
  assign n13320 = ~n13080 & n13319 ;
  assign n13321 = n13320 ^ n13079 ;
  assign n13322 = ~n13074 & n13321 ;
  assign n13323 = n13322 ^ x96 ;
  assign n13326 = n13325 ^ n13323 ;
  assign n13327 = n13325 ^ x97 ;
  assign n13328 = n13326 & ~n13327 ;
  assign n13329 = n13328 ^ x97 ;
  assign n13069 = n12866 & n13005 ;
  assign n13070 = n13069 ^ n12649 ;
  assign n13330 = n13329 ^ n13070 ;
  assign n13331 = n13329 ^ x98 ;
  assign n13332 = n13330 & n13331 ;
  assign n13333 = n13332 ^ x98 ;
  assign n13067 = n12870 & n13005 ;
  assign n13068 = n13067 ^ n12647 ;
  assign n13334 = n13333 ^ n13068 ;
  assign n13335 = n13333 ^ x99 ;
  assign n13336 = n13334 & n13335 ;
  assign n13337 = n13336 ^ x99 ;
  assign n13065 = n12874 & n13005 ;
  assign n13066 = n13065 ^ n12645 ;
  assign n13338 = n13337 ^ n13066 ;
  assign n13339 = n13337 ^ x100 ;
  assign n13340 = n13338 & n13339 ;
  assign n13341 = n13340 ^ x100 ;
  assign n13062 = n12876 ^ x100 ;
  assign n13063 = n13005 & n13062 ;
  assign n13064 = n13063 ^ n12642 ;
  assign n13342 = n13341 ^ n13064 ;
  assign n13343 = n13341 ^ x101 ;
  assign n13344 = n13342 & n13343 ;
  assign n13345 = n13344 ^ x101 ;
  assign n13059 = n12879 ^ x101 ;
  assign n13060 = n13005 & n13059 ;
  assign n13061 = n13060 ^ n12639 ;
  assign n13346 = n13345 ^ n13061 ;
  assign n13347 = n13345 ^ x102 ;
  assign n13348 = n13346 & n13347 ;
  assign n13349 = n13348 ^ x102 ;
  assign n13057 = n12884 & n13005 ;
  assign n13058 = n13057 ^ n12637 ;
  assign n13350 = n13349 ^ n13058 ;
  assign n13351 = n13349 ^ x103 ;
  assign n13352 = n13350 & n13351 ;
  assign n13353 = n13352 ^ x103 ;
  assign n13055 = n12888 & n13005 ;
  assign n13056 = n13055 ^ n12635 ;
  assign n13354 = n13353 ^ n13056 ;
  assign n13355 = n13353 ^ x104 ;
  assign n13356 = n13354 & n13355 ;
  assign n13357 = n13356 ^ x104 ;
  assign n13053 = n12892 & n13005 ;
  assign n13054 = n13053 ^ n12633 ;
  assign n13358 = n13357 ^ n13054 ;
  assign n13359 = n13357 ^ x105 ;
  assign n13360 = n13358 & n13359 ;
  assign n13361 = n13360 ^ x105 ;
  assign n13051 = n12896 & n13005 ;
  assign n13052 = n13051 ^ n12631 ;
  assign n13362 = n13361 ^ n13052 ;
  assign n13363 = n13361 ^ x106 ;
  assign n13364 = n13362 & n13363 ;
  assign n13365 = n13364 ^ x106 ;
  assign n13049 = n12900 & n13005 ;
  assign n13050 = n13049 ^ n12629 ;
  assign n13366 = n13365 ^ n13050 ;
  assign n13367 = n13365 ^ x107 ;
  assign n13368 = n13366 & n13367 ;
  assign n13369 = n13368 ^ x107 ;
  assign n13047 = n12904 & n13005 ;
  assign n13048 = n13047 ^ n12627 ;
  assign n13370 = n13369 ^ n13048 ;
  assign n13371 = n13369 ^ x108 ;
  assign n13372 = n13370 & n13371 ;
  assign n13373 = n13372 ^ x108 ;
  assign n13044 = n12906 ^ x108 ;
  assign n13045 = n13005 & n13044 ;
  assign n13046 = n13045 ^ n12622 ;
  assign n13374 = n13373 ^ n13046 ;
  assign n13375 = n13373 ^ x109 ;
  assign n13376 = n13374 & n13375 ;
  assign n13377 = n13376 ^ x109 ;
  assign n13033 = n12622 ^ x109 ;
  assign n13034 = n13033 ^ n12906 ;
  assign n13035 = n13034 ^ x108 ;
  assign n13036 = n13035 ^ n13033 ;
  assign n13038 = n12906 ^ x109 ;
  assign n13039 = n13038 ^ n13033 ;
  assign n13040 = ~n13036 & ~n13039 ;
  assign n13041 = n13040 ^ n13033 ;
  assign n13042 = n13005 & ~n13041 ;
  assign n13043 = n13042 ^ n12618 ;
  assign n13378 = n13377 ^ n13043 ;
  assign n13379 = n13377 ^ x110 ;
  assign n13380 = n13378 & n13379 ;
  assign n13381 = n13380 ^ x110 ;
  assign n13030 = n12912 ^ x110 ;
  assign n13031 = n13005 & n13030 ;
  assign n13032 = n13031 ^ n12915 ;
  assign n13382 = n13381 ^ n13032 ;
  assign n13383 = n13381 ^ x111 ;
  assign n13384 = n13382 & n13383 ;
  assign n13385 = n13384 ^ x111 ;
  assign n13386 = n13385 ^ n13028 ;
  assign n13387 = ~n13029 & n13386 ;
  assign n13388 = n13387 ^ x112 ;
  assign n13389 = n13388 ^ n13024 ;
  assign n13390 = ~n13025 & n13389 ;
  assign n13391 = n13390 ^ x113 ;
  assign n13020 = n12933 & n13005 ;
  assign n13021 = n13020 ^ n12607 ;
  assign n13392 = n13391 ^ n13021 ;
  assign n13393 = n13391 ^ x114 ;
  assign n13394 = n13392 & n13393 ;
  assign n13395 = n13394 ^ x114 ;
  assign n13017 = n12935 ^ x114 ;
  assign n13018 = n13005 & n13017 ;
  assign n13019 = n13018 ^ n12604 ;
  assign n13396 = n13395 ^ n13019 ;
  assign n13397 = n13395 ^ x115 ;
  assign n13398 = n13396 & n13397 ;
  assign n13399 = n13398 ^ x115 ;
  assign n13014 = n12938 ^ x115 ;
  assign n13015 = n13005 & n13014 ;
  assign n13016 = n13015 ^ n12601 ;
  assign n13400 = n13399 ^ n13016 ;
  assign n13401 = n13399 ^ x116 ;
  assign n13402 = n13400 & n13401 ;
  assign n13403 = n13402 ^ x116 ;
  assign n13012 = n12943 & n13005 ;
  assign n13013 = n13012 ^ n12599 ;
  assign n13404 = n13403 ^ n13013 ;
  assign n13405 = n13403 ^ x117 ;
  assign n13406 = n13404 & n13405 ;
  assign n13407 = n13406 ^ x117 ;
  assign n13010 = n12947 & n13005 ;
  assign n13011 = n13010 ^ n12596 ;
  assign n13408 = n13407 ^ n13011 ;
  assign n13409 = n13407 ^ x118 ;
  assign n13410 = n13408 & n13409 ;
  assign n13411 = n13410 ^ x118 ;
  assign n13008 = n12951 & n13005 ;
  assign n13009 = n13008 ^ n12594 ;
  assign n13412 = n13411 ^ n13009 ;
  assign n13413 = n13411 ^ x119 ;
  assign n13414 = n13412 & n13413 ;
  assign n13415 = n13414 ^ x119 ;
  assign n13006 = n12954 & n13005 ;
  assign n13007 = n13006 ^ n12983 ;
  assign n13416 = n13415 ^ n13007 ;
  assign n13417 = n13415 ^ x120 ;
  assign n13418 = n13416 & n13417 ;
  assign n13419 = n13418 ^ x120 ;
  assign n13420 = n13419 ^ x121 ;
  assign n13426 = n12988 & n13005 ;
  assign n13427 = n13426 ^ n12980 ;
  assign n13428 = n13427 ^ n13419 ;
  assign n13429 = n13420 & n13428 ;
  assign n13430 = n13429 ^ x121 ;
  assign n13424 = n12992 & n13005 ;
  assign n13425 = n13424 ^ n12977 ;
  assign n13431 = n13430 ^ n13425 ;
  assign n13432 = n13430 ^ x122 ;
  assign n13433 = n13431 & n13432 ;
  assign n13434 = n13433 ^ x122 ;
  assign n13421 = n12994 ^ x122 ;
  assign n13422 = n13005 & n13421 ;
  assign n13423 = n13422 ^ n12974 ;
  assign n13435 = n13434 ^ n13423 ;
  assign n13436 = n13434 ^ x123 ;
  assign n13437 = n13435 & n13436 ;
  assign n13438 = n13437 ^ x123 ;
  assign n13439 = x124 & n130 ;
  assign n13440 = ~n12186 & n13439 ;
  assign n13441 = n13440 ^ n130 ;
  assign n13442 = n131 & n12971 ;
  assign n13443 = n13000 & n13442 ;
  assign n13444 = n13443 ^ n12971 ;
  assign n13445 = n13444 ^ x124 ;
  assign n13446 = n13445 ^ n13438 ;
  assign n13447 = n13446 ^ n130 ;
  assign n13448 = n13441 & ~n13447 ;
  assign n13449 = n13438 & n13448 ;
  assign n13450 = n13449 ^ n13440 ;
  assign n13451 = n13450 ^ n130 ;
  assign n13624 = n13173 ^ x65 ;
  assign n13625 = n13451 & n13624 ;
  assign n13616 = ~x2 & x64 ;
  assign n13617 = n13451 ^ x3 ;
  assign n13618 = n13617 ^ n13451 ;
  assign n13621 = x65 & n13618 ;
  assign n13622 = n13621 ^ n13617 ;
  assign n13623 = n13616 & ~n13622 ;
  assign n13626 = n13625 ^ n13623 ;
  assign n13627 = n13615 & ~n13626 ;
  assign n13599 = x64 ^ x3 ;
  assign n13600 = n13005 ^ x4 ;
  assign n13601 = n13005 ^ x2 ;
  assign n13602 = n13601 ^ n13005 ;
  assign n13603 = ~n13600 & n13602 ;
  assign n13604 = n13603 ^ n13601 ;
  assign n13608 = ~n191 & n13604 ;
  assign n13609 = n13608 ^ n13600 ;
  assign n13610 = x64 & ~n13609 ;
  assign n13611 = n13610 ^ n13182 ;
  assign n13612 = n13599 & n13611 ;
  assign n13613 = n13451 & n13612 ;
  assign n13628 = n13627 ^ n13613 ;
  assign n13629 = n13175 ^ x2 ;
  assign n13630 = n13629 ^ x65 ;
  assign n13631 = n13630 ^ x3 ;
  assign n13632 = n13631 ^ n13451 ;
  assign n13633 = ~x2 & ~n13632 ;
  assign n13634 = n13633 ^ n13629 ;
  assign n13635 = n13629 ^ n13451 ;
  assign n13636 = n13635 ^ x2 ;
  assign n13637 = ~n13617 & ~n13636 ;
  assign n13638 = n13637 ^ n13629 ;
  assign n13639 = ~n13634 & ~n13638 ;
  assign n13640 = n13639 ^ n13629 ;
  assign n13641 = x64 & ~n13640 ;
  assign n13642 = ~x66 & n13614 ;
  assign n13643 = x64 & n13451 ;
  assign n13644 = n13451 ^ n13175 ;
  assign n13645 = ~n13643 & ~n13644 ;
  assign n13646 = n13642 & n13645 ;
  assign n13647 = n13646 ^ x66 ;
  assign n13648 = ~n13641 & ~n13647 ;
  assign n13649 = ~n13628 & ~n13648 ;
  assign n13650 = n13649 ^ x67 ;
  assign n13651 = n13179 ^ x66 ;
  assign n13652 = n13451 & n13651 ;
  assign n13653 = n13652 ^ n13196 ;
  assign n13654 = n13653 ^ n13649 ;
  assign n13655 = n13650 & n13654 ;
  assign n13656 = n13655 ^ x67 ;
  assign n13657 = n13656 ^ x68 ;
  assign n13658 = n13200 ^ x67 ;
  assign n13659 = n13451 & n13658 ;
  assign n13660 = n13659 ^ n13203 ;
  assign n13661 = n13660 ^ n13656 ;
  assign n13662 = n13657 & n13661 ;
  assign n13663 = n13662 ^ x68 ;
  assign n13665 = n13663 ^ x69 ;
  assign n13886 = n13438 ^ x124 ;
  assign n13887 = n130 & n13444 ;
  assign n13888 = n13886 & n13887 ;
  assign n13889 = n13888 ^ n13444 ;
  assign n13890 = n13889 ^ x125 ;
  assign n13859 = n13401 & n13451 ;
  assign n13860 = n13859 ^ n13016 ;
  assign n13462 = n13397 & n13451 ;
  assign n13463 = n13462 ^ n13019 ;
  assign n13464 = n13463 ^ x116 ;
  assign n13468 = n13463 ^ x115 ;
  assign n13465 = n13393 & n13451 ;
  assign n13466 = n13465 ^ n13021 ;
  assign n13467 = n13466 ^ n13463 ;
  assign n13469 = n13468 ^ n13467 ;
  assign n13807 = n13351 & n13451 ;
  assign n13808 = n13807 ^ n13058 ;
  assign n13492 = n13347 & n13451 ;
  assign n13493 = n13492 ^ n13061 ;
  assign n13494 = n13493 ^ x103 ;
  assign n13498 = n13493 ^ x102 ;
  assign n13495 = n13343 & n13451 ;
  assign n13496 = n13495 ^ n13064 ;
  assign n13497 = n13496 ^ n13493 ;
  assign n13499 = n13498 ^ n13497 ;
  assign n13795 = n13339 & n13451 ;
  assign n13796 = n13795 ^ n13066 ;
  assign n13500 = n13335 & n13451 ;
  assign n13501 = n13500 ^ n13068 ;
  assign n13502 = n13501 ^ x100 ;
  assign n13506 = n13501 ^ x99 ;
  assign n13503 = n13331 & n13451 ;
  assign n13504 = n13503 ^ n13070 ;
  assign n13505 = n13504 ^ n13501 ;
  assign n13507 = n13506 ^ n13505 ;
  assign n13527 = n13307 & n13451 ;
  assign n13528 = n13527 ^ n13097 ;
  assign n13529 = n13528 ^ x93 ;
  assign n13686 = n13231 & n13451 ;
  assign n13687 = n13686 ^ n13164 ;
  assign n13680 = n13227 & n13451 ;
  assign n13681 = n13680 ^ n13166 ;
  assign n13674 = n13223 & n13451 ;
  assign n13675 = n13674 ^ n13168 ;
  assign n13588 = n13219 & n13451 ;
  assign n13589 = n13588 ^ n13170 ;
  assign n13590 = n13589 ^ x71 ;
  assign n13594 = n13589 ^ x70 ;
  assign n13591 = n13215 & n13451 ;
  assign n13592 = n13591 ^ n13172 ;
  assign n13593 = n13592 ^ n13589 ;
  assign n13595 = n13594 ^ n13593 ;
  assign n13596 = n13207 ^ x68 ;
  assign n13597 = n13451 & n13596 ;
  assign n13598 = n13597 ^ n13209 ;
  assign n13664 = n13663 ^ n13598 ;
  assign n13666 = n13664 & n13665 ;
  assign n13667 = n13666 ^ x69 ;
  assign n13668 = n13667 ^ n13589 ;
  assign n13669 = n13668 ^ n13594 ;
  assign n13670 = ~n13595 & n13669 ;
  assign n13671 = n13670 ^ n13594 ;
  assign n13672 = ~n13590 & n13671 ;
  assign n13673 = n13672 ^ x71 ;
  assign n13676 = n13675 ^ n13673 ;
  assign n13677 = n13675 ^ x72 ;
  assign n13678 = n13676 & ~n13677 ;
  assign n13679 = n13678 ^ x72 ;
  assign n13682 = n13681 ^ n13679 ;
  assign n13683 = n13681 ^ x73 ;
  assign n13684 = n13682 & ~n13683 ;
  assign n13685 = n13684 ^ x73 ;
  assign n13688 = n13687 ^ n13685 ;
  assign n13689 = n13687 ^ x74 ;
  assign n13690 = n13688 & ~n13689 ;
  assign n13691 = n13690 ^ x74 ;
  assign n13585 = n13233 ^ x74 ;
  assign n13586 = n13451 & n13585 ;
  assign n13587 = n13586 ^ n13159 ;
  assign n13692 = n13691 ^ n13587 ;
  assign n13693 = n13691 ^ x75 ;
  assign n13694 = n13692 & n13693 ;
  assign n13695 = n13694 ^ x75 ;
  assign n13574 = n13159 ^ x75 ;
  assign n13575 = n13574 ^ n13233 ;
  assign n13576 = n13575 ^ x74 ;
  assign n13577 = n13576 ^ n13574 ;
  assign n13579 = n13233 ^ x75 ;
  assign n13580 = n13579 ^ n13574 ;
  assign n13581 = ~n13577 & ~n13580 ;
  assign n13582 = n13581 ^ n13574 ;
  assign n13583 = n13451 & ~n13582 ;
  assign n13584 = n13583 ^ n13155 ;
  assign n13696 = n13695 ^ n13584 ;
  assign n13697 = n13695 ^ x76 ;
  assign n13698 = n13696 & n13697 ;
  assign n13699 = n13698 ^ x76 ;
  assign n13571 = n13239 ^ x76 ;
  assign n13572 = n13451 & n13571 ;
  assign n13573 = n13572 ^ n13241 ;
  assign n13700 = n13699 ^ n13573 ;
  assign n13701 = n13699 ^ x77 ;
  assign n13702 = n13700 & n13701 ;
  assign n13703 = n13702 ^ x77 ;
  assign n13569 = n13247 & n13451 ;
  assign n13570 = n13569 ^ n13152 ;
  assign n13704 = n13703 ^ n13570 ;
  assign n13705 = n13703 ^ x78 ;
  assign n13706 = n13704 & n13705 ;
  assign n13707 = n13706 ^ x78 ;
  assign n13567 = n13251 & n13451 ;
  assign n13568 = n13567 ^ n13150 ;
  assign n13708 = n13707 ^ n13568 ;
  assign n13709 = n13707 ^ x79 ;
  assign n13710 = n13708 & n13709 ;
  assign n13711 = n13710 ^ x79 ;
  assign n13565 = n13255 & n13451 ;
  assign n13566 = n13565 ^ n13148 ;
  assign n13712 = n13711 ^ n13566 ;
  assign n13713 = n13711 ^ x80 ;
  assign n13714 = n13712 & n13713 ;
  assign n13715 = n13714 ^ x80 ;
  assign n13563 = n13259 & n13451 ;
  assign n13564 = n13563 ^ n13146 ;
  assign n13716 = n13715 ^ n13564 ;
  assign n13717 = n13715 ^ x81 ;
  assign n13718 = n13716 & n13717 ;
  assign n13719 = n13718 ^ x81 ;
  assign n13561 = n13263 & n13451 ;
  assign n13562 = n13561 ^ n13144 ;
  assign n13720 = n13719 ^ n13562 ;
  assign n13721 = n13719 ^ x82 ;
  assign n13722 = n13720 & n13721 ;
  assign n13723 = n13722 ^ x82 ;
  assign n13559 = n13267 & n13451 ;
  assign n13560 = n13559 ^ n13141 ;
  assign n13724 = n13723 ^ n13560 ;
  assign n13725 = n13723 ^ x83 ;
  assign n13726 = n13724 & n13725 ;
  assign n13727 = n13726 ^ x83 ;
  assign n13557 = n13271 & n13451 ;
  assign n13558 = n13557 ^ n13138 ;
  assign n13728 = n13727 ^ n13558 ;
  assign n13729 = n13727 ^ x84 ;
  assign n13730 = n13728 & n13729 ;
  assign n13731 = n13730 ^ x84 ;
  assign n13555 = n13275 & n13451 ;
  assign n13556 = n13555 ^ n13135 ;
  assign n13732 = n13731 ^ n13556 ;
  assign n13733 = n13731 ^ x85 ;
  assign n13734 = n13732 & n13733 ;
  assign n13735 = n13734 ^ x85 ;
  assign n13553 = n13279 & n13451 ;
  assign n13554 = n13553 ^ n13124 ;
  assign n13736 = n13735 ^ n13554 ;
  assign n13737 = n13735 ^ x86 ;
  assign n13738 = n13736 & n13737 ;
  assign n13739 = n13738 ^ x86 ;
  assign n13551 = n13283 & n13451 ;
  assign n13552 = n13551 ^ n13121 ;
  assign n13740 = n13739 ^ n13552 ;
  assign n13741 = n13739 ^ x87 ;
  assign n13742 = n13740 & n13741 ;
  assign n13743 = n13742 ^ x87 ;
  assign n13549 = n13287 & n13451 ;
  assign n13550 = n13549 ^ n13110 ;
  assign n13744 = n13743 ^ n13550 ;
  assign n13745 = n13743 ^ x88 ;
  assign n13746 = n13744 & n13745 ;
  assign n13747 = n13746 ^ x88 ;
  assign n13546 = n13289 ^ x88 ;
  assign n13547 = n13451 & n13546 ;
  assign n13548 = n13547 ^ n13104 ;
  assign n13748 = n13747 ^ n13548 ;
  assign n13749 = n13747 ^ x89 ;
  assign n13750 = n13748 & n13749 ;
  assign n13751 = n13750 ^ x89 ;
  assign n13535 = n13104 ^ x89 ;
  assign n13536 = n13535 ^ n13289 ;
  assign n13537 = n13536 ^ x88 ;
  assign n13538 = n13537 ^ n13535 ;
  assign n13540 = n13289 ^ x89 ;
  assign n13541 = n13540 ^ n13535 ;
  assign n13542 = ~n13538 & ~n13541 ;
  assign n13543 = n13542 ^ n13535 ;
  assign n13544 = n13451 & ~n13543 ;
  assign n13545 = n13544 ^ n13101 ;
  assign n13752 = n13751 ^ n13545 ;
  assign n13753 = n13751 ^ x90 ;
  assign n13754 = n13752 & n13753 ;
  assign n13755 = n13754 ^ x90 ;
  assign n13532 = n13295 ^ x90 ;
  assign n13533 = n13451 & n13532 ;
  assign n13534 = n13533 ^ n13297 ;
  assign n13756 = n13755 ^ n13534 ;
  assign n13757 = n13755 ^ x91 ;
  assign n13758 = n13756 & n13757 ;
  assign n13759 = n13758 ^ x91 ;
  assign n13530 = n13303 & n13451 ;
  assign n13531 = n13530 ^ n13099 ;
  assign n13760 = n13759 ^ n13531 ;
  assign n13761 = n13759 ^ x92 ;
  assign n13762 = n13760 & n13761 ;
  assign n13763 = n13762 ^ x92 ;
  assign n13764 = n13763 ^ n13528 ;
  assign n13765 = ~n13529 & n13764 ;
  assign n13766 = n13765 ^ x93 ;
  assign n13767 = n13766 ^ x94 ;
  assign n13768 = n13311 & n13451 ;
  assign n13769 = n13768 ^ n13094 ;
  assign n13770 = n13769 ^ n13766 ;
  assign n13771 = n13767 & n13770 ;
  assign n13772 = n13771 ^ x94 ;
  assign n13525 = n13315 & n13451 ;
  assign n13526 = n13525 ^ n13083 ;
  assign n13773 = n13772 ^ n13526 ;
  assign n13774 = n13772 ^ x95 ;
  assign n13775 = n13773 & n13774 ;
  assign n13776 = n13775 ^ x95 ;
  assign n13522 = n13317 ^ x95 ;
  assign n13523 = n13451 & n13522 ;
  assign n13524 = n13523 ^ n13077 ;
  assign n13777 = n13776 ^ n13524 ;
  assign n13778 = n13776 ^ x96 ;
  assign n13779 = n13777 & n13778 ;
  assign n13780 = n13779 ^ x96 ;
  assign n13511 = n13077 ^ x96 ;
  assign n13512 = n13511 ^ n13317 ;
  assign n13513 = n13512 ^ x95 ;
  assign n13514 = n13513 ^ n13511 ;
  assign n13516 = n13317 ^ x96 ;
  assign n13517 = n13516 ^ n13511 ;
  assign n13518 = ~n13514 & ~n13517 ;
  assign n13519 = n13518 ^ n13511 ;
  assign n13520 = n13451 & ~n13519 ;
  assign n13521 = n13520 ^ n13073 ;
  assign n13781 = n13780 ^ n13521 ;
  assign n13782 = n13780 ^ x97 ;
  assign n13783 = n13781 & n13782 ;
  assign n13784 = n13783 ^ x97 ;
  assign n13508 = n13323 ^ x97 ;
  assign n13509 = n13451 & n13508 ;
  assign n13510 = n13509 ^ n13325 ;
  assign n13785 = n13784 ^ n13510 ;
  assign n13786 = n13784 ^ x98 ;
  assign n13787 = n13785 & n13786 ;
  assign n13788 = n13787 ^ x98 ;
  assign n13789 = n13788 ^ n13501 ;
  assign n13790 = n13789 ^ n13506 ;
  assign n13791 = ~n13507 & n13790 ;
  assign n13792 = n13791 ^ n13506 ;
  assign n13793 = ~n13502 & n13792 ;
  assign n13794 = n13793 ^ x100 ;
  assign n13797 = n13796 ^ n13794 ;
  assign n13798 = n13796 ^ x101 ;
  assign n13799 = n13797 & ~n13798 ;
  assign n13800 = n13799 ^ x101 ;
  assign n13801 = n13800 ^ n13493 ;
  assign n13802 = n13801 ^ n13498 ;
  assign n13803 = ~n13499 & n13802 ;
  assign n13804 = n13803 ^ n13498 ;
  assign n13805 = ~n13494 & n13804 ;
  assign n13806 = n13805 ^ x103 ;
  assign n13809 = n13808 ^ n13806 ;
  assign n13810 = n13808 ^ x104 ;
  assign n13811 = n13809 & ~n13810 ;
  assign n13812 = n13811 ^ x104 ;
  assign n13490 = n13355 & n13451 ;
  assign n13491 = n13490 ^ n13056 ;
  assign n13813 = n13812 ^ n13491 ;
  assign n13814 = n13812 ^ x105 ;
  assign n13815 = n13813 & n13814 ;
  assign n13816 = n13815 ^ x105 ;
  assign n13488 = n13359 & n13451 ;
  assign n13489 = n13488 ^ n13054 ;
  assign n13817 = n13816 ^ n13489 ;
  assign n13818 = n13816 ^ x106 ;
  assign n13819 = n13817 & n13818 ;
  assign n13820 = n13819 ^ x106 ;
  assign n13486 = n13363 & n13451 ;
  assign n13487 = n13486 ^ n13052 ;
  assign n13821 = n13820 ^ n13487 ;
  assign n13822 = n13820 ^ x107 ;
  assign n13823 = n13821 & n13822 ;
  assign n13824 = n13823 ^ x107 ;
  assign n13484 = n13367 & n13451 ;
  assign n13485 = n13484 ^ n13050 ;
  assign n13825 = n13824 ^ n13485 ;
  assign n13826 = n13824 ^ x108 ;
  assign n13827 = n13825 & n13826 ;
  assign n13828 = n13827 ^ x108 ;
  assign n13482 = n13371 & n13451 ;
  assign n13483 = n13482 ^ n13048 ;
  assign n13829 = n13828 ^ n13483 ;
  assign n13830 = n13828 ^ x109 ;
  assign n13831 = n13829 & n13830 ;
  assign n13832 = n13831 ^ x109 ;
  assign n13480 = n13375 & n13451 ;
  assign n13481 = n13480 ^ n13046 ;
  assign n13833 = n13832 ^ n13481 ;
  assign n13834 = n13832 ^ x110 ;
  assign n13835 = n13833 & n13834 ;
  assign n13836 = n13835 ^ x110 ;
  assign n13478 = n13379 & n13451 ;
  assign n13479 = n13478 ^ n13043 ;
  assign n13837 = n13836 ^ n13479 ;
  assign n13838 = n13836 ^ x111 ;
  assign n13839 = n13837 & n13838 ;
  assign n13840 = n13839 ^ x111 ;
  assign n13476 = n13383 & n13451 ;
  assign n13477 = n13476 ^ n13032 ;
  assign n13841 = n13840 ^ n13477 ;
  assign n13842 = n13840 ^ x112 ;
  assign n13843 = n13841 & n13842 ;
  assign n13844 = n13843 ^ x112 ;
  assign n13473 = n13385 ^ x112 ;
  assign n13474 = n13451 & n13473 ;
  assign n13475 = n13474 ^ n13028 ;
  assign n13845 = n13844 ^ n13475 ;
  assign n13846 = n13844 ^ x113 ;
  assign n13847 = n13845 & n13846 ;
  assign n13848 = n13847 ^ x113 ;
  assign n13470 = n13388 ^ x113 ;
  assign n13471 = n13451 & n13470 ;
  assign n13472 = n13471 ^ n13024 ;
  assign n13849 = n13848 ^ n13472 ;
  assign n13850 = n13848 ^ x114 ;
  assign n13851 = n13849 & n13850 ;
  assign n13852 = n13851 ^ x114 ;
  assign n13853 = n13852 ^ n13463 ;
  assign n13854 = n13853 ^ n13468 ;
  assign n13855 = ~n13469 & n13854 ;
  assign n13856 = n13855 ^ n13468 ;
  assign n13857 = ~n13464 & n13856 ;
  assign n13858 = n13857 ^ x116 ;
  assign n13861 = n13860 ^ n13858 ;
  assign n13862 = n13860 ^ x117 ;
  assign n13863 = n13861 & ~n13862 ;
  assign n13864 = n13863 ^ x117 ;
  assign n13460 = n13405 & n13451 ;
  assign n13461 = n13460 ^ n13013 ;
  assign n13865 = n13864 ^ n13461 ;
  assign n13866 = n13864 ^ x118 ;
  assign n13867 = n13865 & n13866 ;
  assign n13868 = n13867 ^ x118 ;
  assign n13458 = n13409 & n13451 ;
  assign n13459 = n13458 ^ n13011 ;
  assign n13869 = n13868 ^ n13459 ;
  assign n13870 = n13868 ^ x119 ;
  assign n13871 = n13869 & n13870 ;
  assign n13872 = n13871 ^ x119 ;
  assign n13456 = n13413 & n13451 ;
  assign n13457 = n13456 ^ n13009 ;
  assign n13873 = n13872 ^ n13457 ;
  assign n13874 = n13872 ^ x120 ;
  assign n13875 = n13873 & n13874 ;
  assign n13876 = n13875 ^ x120 ;
  assign n13454 = n13417 & n13451 ;
  assign n13455 = n13454 ^ n13007 ;
  assign n13877 = n13876 ^ n13455 ;
  assign n13878 = n13876 ^ x121 ;
  assign n13879 = n13877 & n13878 ;
  assign n13880 = n13879 ^ x121 ;
  assign n13452 = n13420 & n13451 ;
  assign n13453 = n13452 ^ n13427 ;
  assign n13881 = n13880 ^ n13453 ;
  assign n13882 = n13880 ^ x122 ;
  assign n13883 = n13881 & n13882 ;
  assign n13884 = n13883 ^ x122 ;
  assign n13885 = n13884 ^ x123 ;
  assign n13893 = n13432 & n13451 ;
  assign n13894 = n13893 ^ n13425 ;
  assign n13895 = n13894 ^ n13884 ;
  assign n13896 = n13885 & n13895 ;
  assign n13897 = n13896 ^ x123 ;
  assign n13891 = n13436 & n13451 ;
  assign n13892 = n13891 ^ n13423 ;
  assign n13898 = n13897 ^ n13892 ;
  assign n13901 = n13892 ^ x124 ;
  assign n13902 = n13898 & ~n13901 ;
  assign n13899 = x125 ^ x124 ;
  assign n13903 = n13902 ^ n13899 ;
  assign n13906 = ~n13890 & n13903 ;
  assign n13907 = n13906 ^ x125 ;
  assign n13908 = n129 & ~n13907 ;
  assign n14122 = n13665 & n13908 ;
  assign n14123 = n14122 ^ n13598 ;
  assign n14068 = n13657 & n13908 ;
  assign n14069 = n14068 ^ n13660 ;
  assign n14070 = n14069 ^ x69 ;
  assign n14074 = n14069 ^ x68 ;
  assign n14071 = n13650 & n13908 ;
  assign n14072 = n14071 ^ n13653 ;
  assign n14073 = n14072 ^ n14069 ;
  assign n14075 = n14074 ^ n14073 ;
  assign n14078 = n13643 ^ x3 ;
  assign n14076 = n13616 ^ x65 ;
  assign n14077 = n13908 & n14076 ;
  assign n14079 = n14078 ^ n14077 ;
  assign n14080 = n14079 ^ x66 ;
  assign n14088 = x2 & x65 ;
  assign n14085 = x65 ^ x1 ;
  assign n14081 = x64 ^ x2 ;
  assign n14082 = n14081 ^ x65 ;
  assign n14086 = n14082 ^ n13908 ;
  assign n14087 = ~n14085 & n14086 ;
  assign n14089 = n14088 ^ n14087 ;
  assign n14090 = x64 & n14089 ;
  assign n14091 = n14090 ^ n14088 ;
  assign n14092 = n14091 ^ x65 ;
  assign n14093 = n14092 ^ n14079 ;
  assign n14094 = ~n14080 & n14093 ;
  assign n14095 = n14094 ^ x66 ;
  assign n14096 = n14095 ^ x67 ;
  assign n14107 = x3 & x65 ;
  assign n14098 = x65 ^ x2 ;
  assign n14099 = n13599 ^ x65 ;
  assign n14100 = n14099 ^ n13451 ;
  assign n14101 = ~n14098 & n14100 ;
  assign n14108 = n14107 ^ n14101 ;
  assign n14109 = ~x64 & n14108 ;
  assign n14104 = n14101 ^ n6836 ;
  assign n14110 = n14109 ^ n14104 ;
  assign n14111 = n13908 & n14110 ;
  assign n14097 = n13625 ^ n13175 ;
  assign n14112 = n14111 ^ n14097 ;
  assign n14113 = n14112 ^ n14095 ;
  assign n14114 = n14096 & n14113 ;
  assign n14115 = n14114 ^ x67 ;
  assign n14116 = n14115 ^ n14069 ;
  assign n14117 = n14116 ^ n14074 ;
  assign n14118 = ~n14075 & n14117 ;
  assign n14119 = n14118 ^ n14074 ;
  assign n14120 = ~n14070 & n14119 ;
  assign n14121 = n14120 ^ x69 ;
  assign n14124 = n14123 ^ n14121 ;
  assign n14125 = n14123 ^ x70 ;
  assign n14126 = n14124 & ~n14125 ;
  assign n14127 = n14126 ^ x70 ;
  assign n14065 = n13667 ^ x70 ;
  assign n14066 = n13908 & n14065 ;
  assign n14067 = n14066 ^ n13592 ;
  assign n14128 = n14127 ^ n14067 ;
  assign n14129 = n14127 ^ x71 ;
  assign n14130 = n14128 & n14129 ;
  assign n14131 = n14130 ^ x71 ;
  assign n14054 = n13592 ^ x71 ;
  assign n14055 = n14054 ^ n13667 ;
  assign n14056 = n14055 ^ x70 ;
  assign n14057 = n14056 ^ n14054 ;
  assign n14059 = n13667 ^ x71 ;
  assign n14060 = n14059 ^ n14054 ;
  assign n14061 = ~n14057 & ~n14060 ;
  assign n14062 = n14061 ^ n14054 ;
  assign n14063 = n13908 & ~n14062 ;
  assign n14064 = n14063 ^ n13589 ;
  assign n14132 = n14131 ^ n14064 ;
  assign n14133 = n14131 ^ x72 ;
  assign n14134 = n14132 & n14133 ;
  assign n14135 = n14134 ^ x72 ;
  assign n14051 = n13673 ^ x72 ;
  assign n14052 = n13908 & n14051 ;
  assign n14053 = n14052 ^ n13675 ;
  assign n14136 = n14135 ^ n14053 ;
  assign n14137 = n14135 ^ x73 ;
  assign n14138 = n14136 & n14137 ;
  assign n14139 = n14138 ^ x73 ;
  assign n14048 = n13679 ^ x73 ;
  assign n14049 = n13908 & n14048 ;
  assign n14050 = n14049 ^ n13681 ;
  assign n14140 = n14139 ^ n14050 ;
  assign n14141 = n14139 ^ x74 ;
  assign n14142 = n14140 & n14141 ;
  assign n14143 = n14142 ^ x74 ;
  assign n14045 = n13685 ^ x74 ;
  assign n14046 = n13908 & n14045 ;
  assign n14047 = n14046 ^ n13687 ;
  assign n14144 = n14143 ^ n14047 ;
  assign n14145 = n14143 ^ x75 ;
  assign n14146 = n14144 & n14145 ;
  assign n14147 = n14146 ^ x75 ;
  assign n14043 = n13693 & n13908 ;
  assign n14044 = n14043 ^ n13587 ;
  assign n14148 = n14147 ^ n14044 ;
  assign n14149 = n14147 ^ x76 ;
  assign n14150 = n14148 & n14149 ;
  assign n14151 = n14150 ^ x76 ;
  assign n14041 = n13697 & n13908 ;
  assign n14042 = n14041 ^ n13584 ;
  assign n14152 = n14151 ^ n14042 ;
  assign n14153 = n14151 ^ x77 ;
  assign n14154 = n14152 & n14153 ;
  assign n14155 = n14154 ^ x77 ;
  assign n14039 = n13701 & n13908 ;
  assign n14040 = n14039 ^ n13573 ;
  assign n14156 = n14155 ^ n14040 ;
  assign n14157 = n14155 ^ x78 ;
  assign n14158 = n14156 & n14157 ;
  assign n14159 = n14158 ^ x78 ;
  assign n14037 = n13705 & n13908 ;
  assign n14038 = n14037 ^ n13570 ;
  assign n14160 = n14159 ^ n14038 ;
  assign n14161 = n14159 ^ x79 ;
  assign n14162 = n14160 & n14161 ;
  assign n14163 = n14162 ^ x79 ;
  assign n14035 = n13709 & n13908 ;
  assign n14036 = n14035 ^ n13568 ;
  assign n14164 = n14163 ^ n14036 ;
  assign n14165 = n14163 ^ x80 ;
  assign n14166 = n14164 & n14165 ;
  assign n14167 = n14166 ^ x80 ;
  assign n14033 = n13713 & n13908 ;
  assign n14034 = n14033 ^ n13566 ;
  assign n14168 = n14167 ^ n14034 ;
  assign n14169 = n14167 ^ x81 ;
  assign n14170 = n14168 & n14169 ;
  assign n14171 = n14170 ^ x81 ;
  assign n14031 = n13717 & n13908 ;
  assign n14032 = n14031 ^ n13564 ;
  assign n14172 = n14171 ^ n14032 ;
  assign n14173 = n14171 ^ x82 ;
  assign n14174 = n14172 & n14173 ;
  assign n14175 = n14174 ^ x82 ;
  assign n14029 = n13721 & n13908 ;
  assign n14030 = n14029 ^ n13562 ;
  assign n14176 = n14175 ^ n14030 ;
  assign n14177 = n14175 ^ x83 ;
  assign n14178 = n14176 & n14177 ;
  assign n14179 = n14178 ^ x83 ;
  assign n14027 = n13725 & n13908 ;
  assign n14028 = n14027 ^ n13560 ;
  assign n14180 = n14179 ^ n14028 ;
  assign n14181 = n14179 ^ x84 ;
  assign n14182 = n14180 & n14181 ;
  assign n14183 = n14182 ^ x84 ;
  assign n14025 = n13729 & n13908 ;
  assign n14026 = n14025 ^ n13558 ;
  assign n14184 = n14183 ^ n14026 ;
  assign n14185 = n14183 ^ x85 ;
  assign n14186 = n14184 & n14185 ;
  assign n14187 = n14186 ^ x85 ;
  assign n14188 = n14187 ^ x86 ;
  assign n14189 = n13733 & n13908 ;
  assign n14190 = n14189 ^ n13556 ;
  assign n14191 = n14190 ^ n14187 ;
  assign n14192 = n14188 & n14191 ;
  assign n14193 = n14192 ^ x86 ;
  assign n14195 = n14193 ^ x87 ;
  assign n14345 = n129 & n13889 ;
  assign n14346 = n13903 & n14345 ;
  assign n14347 = n14346 ^ n13889 ;
  assign n14348 = n14347 ^ x126 ;
  assign n14349 = n13897 ^ x124 ;
  assign n14350 = n13908 & n14349 ;
  assign n14351 = n14350 ^ n13892 ;
  assign n14322 = n13870 & n13908 ;
  assign n14323 = n14322 ^ n13459 ;
  assign n13917 = n13866 & n13908 ;
  assign n13918 = n13917 ^ n13461 ;
  assign n13919 = n13918 ^ x119 ;
  assign n13924 = n13918 ^ x118 ;
  assign n13920 = n13858 ^ x117 ;
  assign n13921 = n13908 & n13920 ;
  assign n13922 = n13921 ^ n13860 ;
  assign n13923 = n13922 ^ n13918 ;
  assign n13925 = n13924 ^ n13923 ;
  assign n14302 = n13850 & n13908 ;
  assign n14303 = n14302 ^ n13472 ;
  assign n13940 = n13846 & n13908 ;
  assign n13941 = n13940 ^ n13475 ;
  assign n13942 = n13941 ^ x114 ;
  assign n13946 = n13941 ^ x113 ;
  assign n13943 = n13842 & n13908 ;
  assign n13944 = n13943 ^ n13477 ;
  assign n13945 = n13944 ^ n13941 ;
  assign n13947 = n13946 ^ n13945 ;
  assign n13965 = n13496 ^ x103 ;
  assign n13966 = n13965 ^ n13800 ;
  assign n13967 = n13966 ^ x102 ;
  assign n13968 = n13967 ^ n13965 ;
  assign n13970 = n13800 ^ x103 ;
  assign n13971 = n13970 ^ n13965 ;
  assign n13972 = ~n13968 & ~n13971 ;
  assign n13973 = n13972 ^ n13965 ;
  assign n13974 = n13908 & ~n13973 ;
  assign n13975 = n13974 ^ n13493 ;
  assign n13976 = n13975 ^ x104 ;
  assign n13977 = n13800 ^ x102 ;
  assign n13978 = n13908 & n13977 ;
  assign n13979 = n13978 ^ n13496 ;
  assign n13980 = n13979 ^ x103 ;
  assign n14023 = n13737 & n13908 ;
  assign n14024 = n14023 ^ n13554 ;
  assign n14194 = n14193 ^ n14024 ;
  assign n14196 = n14194 & n14195 ;
  assign n14197 = n14196 ^ x87 ;
  assign n14021 = n13741 & n13908 ;
  assign n14022 = n14021 ^ n13552 ;
  assign n14198 = n14197 ^ n14022 ;
  assign n14199 = n14197 ^ x88 ;
  assign n14200 = n14198 & n14199 ;
  assign n14201 = n14200 ^ x88 ;
  assign n14019 = n13745 & n13908 ;
  assign n14020 = n14019 ^ n13550 ;
  assign n14202 = n14201 ^ n14020 ;
  assign n14203 = n14201 ^ x89 ;
  assign n14204 = n14202 & n14203 ;
  assign n14205 = n14204 ^ x89 ;
  assign n14017 = n13749 & n13908 ;
  assign n14018 = n14017 ^ n13548 ;
  assign n14206 = n14205 ^ n14018 ;
  assign n14207 = n14205 ^ x90 ;
  assign n14208 = n14206 & n14207 ;
  assign n14209 = n14208 ^ x90 ;
  assign n14015 = n13753 & n13908 ;
  assign n14016 = n14015 ^ n13545 ;
  assign n14210 = n14209 ^ n14016 ;
  assign n14211 = n14209 ^ x91 ;
  assign n14212 = n14210 & n14211 ;
  assign n14213 = n14212 ^ x91 ;
  assign n14013 = n13757 & n13908 ;
  assign n14014 = n14013 ^ n13534 ;
  assign n14214 = n14213 ^ n14014 ;
  assign n14215 = n14213 ^ x92 ;
  assign n14216 = n14214 & n14215 ;
  assign n14217 = n14216 ^ x92 ;
  assign n14011 = n13761 & n13908 ;
  assign n14012 = n14011 ^ n13531 ;
  assign n14218 = n14217 ^ n14012 ;
  assign n14219 = n14217 ^ x93 ;
  assign n14220 = n14218 & n14219 ;
  assign n14221 = n14220 ^ x93 ;
  assign n14008 = n13763 ^ x93 ;
  assign n14009 = n13908 & n14008 ;
  assign n14010 = n14009 ^ n13528 ;
  assign n14222 = n14221 ^ n14010 ;
  assign n14223 = n14221 ^ x94 ;
  assign n14224 = n14222 & n14223 ;
  assign n14225 = n14224 ^ x94 ;
  assign n14006 = n13767 & n13908 ;
  assign n14007 = n14006 ^ n13769 ;
  assign n14226 = n14225 ^ n14007 ;
  assign n14227 = n14225 ^ x95 ;
  assign n14228 = n14226 & n14227 ;
  assign n14229 = n14228 ^ x95 ;
  assign n14004 = n13774 & n13908 ;
  assign n14005 = n14004 ^ n13526 ;
  assign n14230 = n14229 ^ n14005 ;
  assign n14231 = n14229 ^ x96 ;
  assign n14232 = n14230 & n14231 ;
  assign n14233 = n14232 ^ x96 ;
  assign n14002 = n13778 & n13908 ;
  assign n14003 = n14002 ^ n13524 ;
  assign n14234 = n14233 ^ n14003 ;
  assign n14235 = n14233 ^ x97 ;
  assign n14236 = n14234 & n14235 ;
  assign n14237 = n14236 ^ x97 ;
  assign n14000 = n13782 & n13908 ;
  assign n14001 = n14000 ^ n13521 ;
  assign n14238 = n14237 ^ n14001 ;
  assign n14239 = n14237 ^ x98 ;
  assign n14240 = n14238 & n14239 ;
  assign n14241 = n14240 ^ x98 ;
  assign n13998 = n13786 & n13908 ;
  assign n13999 = n13998 ^ n13510 ;
  assign n14242 = n14241 ^ n13999 ;
  assign n14243 = n14241 ^ x99 ;
  assign n14244 = n14242 & n14243 ;
  assign n14245 = n14244 ^ x99 ;
  assign n13995 = n13788 ^ x99 ;
  assign n13996 = n13908 & n13995 ;
  assign n13997 = n13996 ^ n13504 ;
  assign n14246 = n14245 ^ n13997 ;
  assign n14247 = n14245 ^ x100 ;
  assign n14248 = n14246 & n14247 ;
  assign n14249 = n14248 ^ x100 ;
  assign n13984 = n13504 ^ x100 ;
  assign n13985 = n13984 ^ n13788 ;
  assign n13986 = n13985 ^ x99 ;
  assign n13987 = n13986 ^ n13984 ;
  assign n13989 = n13788 ^ x100 ;
  assign n13990 = n13989 ^ n13984 ;
  assign n13991 = ~n13987 & ~n13990 ;
  assign n13992 = n13991 ^ n13984 ;
  assign n13993 = n13908 & ~n13992 ;
  assign n13994 = n13993 ^ n13501 ;
  assign n14250 = n14249 ^ n13994 ;
  assign n14251 = n14249 ^ x101 ;
  assign n14252 = n14250 & n14251 ;
  assign n14253 = n14252 ^ x101 ;
  assign n13981 = n13794 ^ x101 ;
  assign n13982 = n13908 & n13981 ;
  assign n13983 = n13982 ^ n13796 ;
  assign n14254 = n14253 ^ n13983 ;
  assign n14255 = n14253 ^ x102 ;
  assign n14256 = n14254 & n14255 ;
  assign n14257 = n14256 ^ x102 ;
  assign n14258 = n14257 ^ n13979 ;
  assign n14259 = ~n13980 & n14258 ;
  assign n14260 = n14259 ^ x103 ;
  assign n14261 = n14260 ^ n13975 ;
  assign n14262 = ~n13976 & n14261 ;
  assign n14263 = n14262 ^ x104 ;
  assign n13962 = n13806 ^ x104 ;
  assign n13963 = n13908 & n13962 ;
  assign n13964 = n13963 ^ n13808 ;
  assign n14264 = n14263 ^ n13964 ;
  assign n14265 = n14263 ^ x105 ;
  assign n14266 = n14264 & n14265 ;
  assign n14267 = n14266 ^ x105 ;
  assign n13960 = n13814 & n13908 ;
  assign n13961 = n13960 ^ n13491 ;
  assign n14268 = n14267 ^ n13961 ;
  assign n14269 = n14267 ^ x106 ;
  assign n14270 = n14268 & n14269 ;
  assign n14271 = n14270 ^ x106 ;
  assign n13958 = n13818 & n13908 ;
  assign n13959 = n13958 ^ n13489 ;
  assign n14272 = n14271 ^ n13959 ;
  assign n14273 = n14271 ^ x107 ;
  assign n14274 = n14272 & n14273 ;
  assign n14275 = n14274 ^ x107 ;
  assign n13956 = n13822 & n13908 ;
  assign n13957 = n13956 ^ n13487 ;
  assign n14276 = n14275 ^ n13957 ;
  assign n14277 = n14275 ^ x108 ;
  assign n14278 = n14276 & n14277 ;
  assign n14279 = n14278 ^ x108 ;
  assign n13954 = n13826 & n13908 ;
  assign n13955 = n13954 ^ n13485 ;
  assign n14280 = n14279 ^ n13955 ;
  assign n14281 = n14279 ^ x109 ;
  assign n14282 = n14280 & n14281 ;
  assign n14283 = n14282 ^ x109 ;
  assign n13952 = n13830 & n13908 ;
  assign n13953 = n13952 ^ n13483 ;
  assign n14284 = n14283 ^ n13953 ;
  assign n14285 = n14283 ^ x110 ;
  assign n14286 = n14284 & n14285 ;
  assign n14287 = n14286 ^ x110 ;
  assign n13950 = n13834 & n13908 ;
  assign n13951 = n13950 ^ n13481 ;
  assign n14288 = n14287 ^ n13951 ;
  assign n14289 = n14287 ^ x111 ;
  assign n14290 = n14288 & n14289 ;
  assign n14291 = n14290 ^ x111 ;
  assign n13948 = n13838 & n13908 ;
  assign n13949 = n13948 ^ n13479 ;
  assign n14292 = n14291 ^ n13949 ;
  assign n14293 = n14291 ^ x112 ;
  assign n14294 = n14292 & n14293 ;
  assign n14295 = n14294 ^ x112 ;
  assign n14296 = n14295 ^ n13941 ;
  assign n14297 = n14296 ^ n13946 ;
  assign n14298 = ~n13947 & n14297 ;
  assign n14299 = n14298 ^ n13946 ;
  assign n14300 = ~n13942 & n14299 ;
  assign n14301 = n14300 ^ x114 ;
  assign n14304 = n14303 ^ n14301 ;
  assign n14305 = n14303 ^ x115 ;
  assign n14306 = n14304 & ~n14305 ;
  assign n14307 = n14306 ^ x115 ;
  assign n13937 = n13852 ^ x115 ;
  assign n13938 = n13908 & n13937 ;
  assign n13939 = n13938 ^ n13466 ;
  assign n14308 = n14307 ^ n13939 ;
  assign n14309 = n14307 ^ x116 ;
  assign n14310 = n14308 & n14309 ;
  assign n14311 = n14310 ^ x116 ;
  assign n13926 = n13466 ^ x116 ;
  assign n13927 = n13926 ^ n13852 ;
  assign n13928 = n13927 ^ x115 ;
  assign n13929 = n13928 ^ n13926 ;
  assign n13931 = n13852 ^ x116 ;
  assign n13932 = n13931 ^ n13926 ;
  assign n13933 = ~n13929 & ~n13932 ;
  assign n13934 = n13933 ^ n13926 ;
  assign n13935 = n13908 & ~n13934 ;
  assign n13936 = n13935 ^ n13463 ;
  assign n14312 = n14311 ^ n13936 ;
  assign n14313 = n14311 ^ x117 ;
  assign n14314 = n14312 & n14313 ;
  assign n14315 = n14314 ^ x117 ;
  assign n14316 = n14315 ^ n13918 ;
  assign n14317 = n14316 ^ n13924 ;
  assign n14318 = ~n13925 & n14317 ;
  assign n14319 = n14318 ^ n13924 ;
  assign n14320 = ~n13919 & n14319 ;
  assign n14321 = n14320 ^ x119 ;
  assign n14324 = n14323 ^ n14321 ;
  assign n14325 = n14323 ^ x120 ;
  assign n14326 = n14324 & ~n14325 ;
  assign n14327 = n14326 ^ x120 ;
  assign n13915 = n13874 & n13908 ;
  assign n13916 = n13915 ^ n13457 ;
  assign n14328 = n14327 ^ n13916 ;
  assign n14329 = n14327 ^ x121 ;
  assign n14330 = n14328 & n14329 ;
  assign n14331 = n14330 ^ x121 ;
  assign n13913 = n13878 & n13908 ;
  assign n13914 = n13913 ^ n13455 ;
  assign n14332 = n14331 ^ n13914 ;
  assign n14333 = n14331 ^ x122 ;
  assign n14334 = n14332 & n14333 ;
  assign n14335 = n14334 ^ x122 ;
  assign n13911 = n13882 & n13908 ;
  assign n13912 = n13911 ^ n13453 ;
  assign n14336 = n14335 ^ n13912 ;
  assign n14337 = n14335 ^ x123 ;
  assign n14338 = n14336 & n14337 ;
  assign n14339 = n14338 ^ x123 ;
  assign n13909 = n13885 & n13908 ;
  assign n13910 = n13909 ^ n13894 ;
  assign n14340 = n14339 ^ n13910 ;
  assign n14341 = n14339 ^ x124 ;
  assign n14342 = n14340 & n14341 ;
  assign n14343 = n14342 ^ x124 ;
  assign n14352 = n14351 ^ n14343 ;
  assign n14355 = n14351 ^ x125 ;
  assign n14356 = n14352 & ~n14355 ;
  assign n14353 = x126 ^ x125 ;
  assign n14357 = n14356 ^ n14353 ;
  assign n14360 = ~n14348 & n14357 ;
  assign n14361 = n14360 ^ x126 ;
  assign n14362 = ~x127 & ~n14361 ;
  assign n14628 = n14195 & n14362 ;
  assign n14629 = n14628 ^ n14024 ;
  assign n14463 = n14188 & n14362 ;
  assign n14464 = n14463 ^ n14190 ;
  assign n14465 = n14464 ^ x87 ;
  assign n14469 = n14464 ^ x86 ;
  assign n14466 = n14185 & n14362 ;
  assign n14467 = n14466 ^ n14026 ;
  assign n14468 = n14467 ^ n14464 ;
  assign n14470 = n14469 ^ n14468 ;
  assign n14588 = n14153 & n14362 ;
  assign n14589 = n14588 ^ n14042 ;
  assign n14485 = n14149 & n14362 ;
  assign n14486 = n14485 ^ n14044 ;
  assign n14487 = n14486 ^ x77 ;
  assign n14491 = n14486 ^ x76 ;
  assign n14488 = n14145 & n14362 ;
  assign n14489 = n14488 ^ n14047 ;
  assign n14490 = n14489 ^ n14486 ;
  assign n14492 = n14491 ^ n14490 ;
  assign n14499 = n14129 & n14362 ;
  assign n14500 = n14499 ^ n14067 ;
  assign n14501 = n14500 ^ x72 ;
  assign n14502 = n14121 ^ x70 ;
  assign n14503 = n14362 & n14502 ;
  assign n14504 = n14503 ^ n14123 ;
  assign n14505 = n14504 ^ x71 ;
  assign n14550 = n14096 & n14362 ;
  assign n14551 = n14550 ^ n14112 ;
  assign n14543 = n14092 ^ x66 ;
  assign n14544 = n14362 & n14543 ;
  assign n14545 = n14544 ^ n14079 ;
  assign n14537 = x64 & n13908 ;
  assign n14533 = ~x1 & x64 ;
  assign n14534 = n14533 ^ x65 ;
  assign n14535 = n14362 & n14534 ;
  assign n14536 = n14535 ^ x2 ;
  assign n14538 = n14537 ^ n14536 ;
  assign n14527 = x1 & x65 ;
  assign n14524 = x65 ^ x0 ;
  assign n14520 = x64 ^ x1 ;
  assign n14521 = n14520 ^ x65 ;
  assign n14525 = n14521 ^ n14362 ;
  assign n14526 = ~n14524 & n14525 ;
  assign n14528 = n14527 ^ n14526 ;
  assign n14529 = x64 & n14528 ;
  assign n14530 = n14529 ^ n14527 ;
  assign n14531 = n14530 ^ x65 ;
  assign n14539 = n14538 ^ n14531 ;
  assign n14540 = n14538 ^ x66 ;
  assign n14541 = n14539 & ~n14540 ;
  assign n14542 = n14541 ^ x66 ;
  assign n14546 = n14545 ^ n14542 ;
  assign n14547 = n14545 ^ x67 ;
  assign n14548 = n14546 & ~n14547 ;
  assign n14549 = n14548 ^ x67 ;
  assign n14552 = n14551 ^ n14549 ;
  assign n14553 = n14551 ^ x68 ;
  assign n14554 = n14552 & ~n14553 ;
  assign n14555 = n14554 ^ x68 ;
  assign n14517 = n14115 ^ x68 ;
  assign n14518 = n14362 & n14517 ;
  assign n14519 = n14518 ^ n14072 ;
  assign n14556 = n14555 ^ n14519 ;
  assign n14557 = n14555 ^ x69 ;
  assign n14558 = n14556 & n14557 ;
  assign n14559 = n14558 ^ x69 ;
  assign n14506 = n14072 ^ x69 ;
  assign n14507 = n14506 ^ n14115 ;
  assign n14508 = n14507 ^ x68 ;
  assign n14509 = n14508 ^ n14506 ;
  assign n14511 = n14115 ^ x69 ;
  assign n14512 = n14511 ^ n14506 ;
  assign n14513 = ~n14509 & ~n14512 ;
  assign n14514 = n14513 ^ n14506 ;
  assign n14515 = n14362 & ~n14514 ;
  assign n14516 = n14515 ^ n14069 ;
  assign n14560 = n14559 ^ n14516 ;
  assign n14561 = n14559 ^ x70 ;
  assign n14562 = n14560 & n14561 ;
  assign n14563 = n14562 ^ x70 ;
  assign n14564 = n14563 ^ n14504 ;
  assign n14565 = ~n14505 & n14564 ;
  assign n14566 = n14565 ^ x71 ;
  assign n14567 = n14566 ^ n14500 ;
  assign n14568 = ~n14501 & n14567 ;
  assign n14569 = n14568 ^ x72 ;
  assign n14497 = n14133 & n14362 ;
  assign n14498 = n14497 ^ n14064 ;
  assign n14570 = n14569 ^ n14498 ;
  assign n14571 = n14569 ^ x73 ;
  assign n14572 = n14570 & n14571 ;
  assign n14573 = n14572 ^ x73 ;
  assign n14495 = n14137 & n14362 ;
  assign n14496 = n14495 ^ n14053 ;
  assign n14574 = n14573 ^ n14496 ;
  assign n14575 = n14573 ^ x74 ;
  assign n14576 = n14574 & n14575 ;
  assign n14577 = n14576 ^ x74 ;
  assign n14493 = n14141 & n14362 ;
  assign n14494 = n14493 ^ n14050 ;
  assign n14578 = n14577 ^ n14494 ;
  assign n14579 = n14577 ^ x75 ;
  assign n14580 = n14578 & n14579 ;
  assign n14581 = n14580 ^ x75 ;
  assign n14582 = n14581 ^ n14486 ;
  assign n14583 = n14582 ^ n14491 ;
  assign n14584 = ~n14492 & n14583 ;
  assign n14585 = n14584 ^ n14491 ;
  assign n14586 = ~n14487 & n14585 ;
  assign n14587 = n14586 ^ x77 ;
  assign n14590 = n14589 ^ n14587 ;
  assign n14591 = n14589 ^ x78 ;
  assign n14592 = n14590 & ~n14591 ;
  assign n14593 = n14592 ^ x78 ;
  assign n14483 = n14157 & n14362 ;
  assign n14484 = n14483 ^ n14040 ;
  assign n14594 = n14593 ^ n14484 ;
  assign n14595 = n14593 ^ x79 ;
  assign n14596 = n14594 & n14595 ;
  assign n14597 = n14596 ^ x79 ;
  assign n14481 = n14161 & n14362 ;
  assign n14482 = n14481 ^ n14038 ;
  assign n14598 = n14597 ^ n14482 ;
  assign n14599 = n14597 ^ x80 ;
  assign n14600 = n14598 & n14599 ;
  assign n14601 = n14600 ^ x80 ;
  assign n14479 = n14165 & n14362 ;
  assign n14480 = n14479 ^ n14036 ;
  assign n14602 = n14601 ^ n14480 ;
  assign n14603 = n14601 ^ x81 ;
  assign n14604 = n14602 & n14603 ;
  assign n14605 = n14604 ^ x81 ;
  assign n14477 = n14169 & n14362 ;
  assign n14478 = n14477 ^ n14034 ;
  assign n14606 = n14605 ^ n14478 ;
  assign n14607 = n14605 ^ x82 ;
  assign n14608 = n14606 & n14607 ;
  assign n14609 = n14608 ^ x82 ;
  assign n14475 = n14173 & n14362 ;
  assign n14476 = n14475 ^ n14032 ;
  assign n14610 = n14609 ^ n14476 ;
  assign n14611 = n14609 ^ x83 ;
  assign n14612 = n14610 & n14611 ;
  assign n14613 = n14612 ^ x83 ;
  assign n14473 = n14177 & n14362 ;
  assign n14474 = n14473 ^ n14030 ;
  assign n14614 = n14613 ^ n14474 ;
  assign n14615 = n14613 ^ x84 ;
  assign n14616 = n14614 & n14615 ;
  assign n14617 = n14616 ^ x84 ;
  assign n14471 = n14181 & n14362 ;
  assign n14472 = n14471 ^ n14028 ;
  assign n14618 = n14617 ^ n14472 ;
  assign n14619 = n14617 ^ x85 ;
  assign n14620 = n14618 & n14619 ;
  assign n14621 = n14620 ^ x85 ;
  assign n14622 = n14621 ^ n14464 ;
  assign n14623 = n14622 ^ n14469 ;
  assign n14624 = ~n14470 & n14623 ;
  assign n14625 = n14624 ^ n14469 ;
  assign n14626 = ~n14465 & n14625 ;
  assign n14627 = n14626 ^ x87 ;
  assign n14630 = n14629 ^ n14627 ;
  assign n14631 = n14629 ^ x88 ;
  assign n14632 = n14630 & ~n14631 ;
  assign n14633 = n14632 ^ x88 ;
  assign n14461 = n14199 & n14362 ;
  assign n14462 = n14461 ^ n14022 ;
  assign n14634 = n14633 ^ n14462 ;
  assign n14635 = n14633 ^ x89 ;
  assign n14636 = n14634 & n14635 ;
  assign n14637 = n14636 ^ x89 ;
  assign n14459 = n14203 & n14362 ;
  assign n14460 = n14459 ^ n14020 ;
  assign n14638 = n14637 ^ n14460 ;
  assign n14639 = n14637 ^ x90 ;
  assign n14640 = n14638 & n14639 ;
  assign n14641 = n14640 ^ x90 ;
  assign n14457 = n14207 & n14362 ;
  assign n14458 = n14457 ^ n14018 ;
  assign n14642 = n14641 ^ n14458 ;
  assign n14643 = n14641 ^ x91 ;
  assign n14644 = n14642 & n14643 ;
  assign n14645 = n14644 ^ x91 ;
  assign n14455 = n14211 & n14362 ;
  assign n14456 = n14455 ^ n14016 ;
  assign n14646 = n14645 ^ n14456 ;
  assign n14647 = n14645 ^ x92 ;
  assign n14648 = n14646 & n14647 ;
  assign n14649 = n14648 ^ x92 ;
  assign n14453 = n14215 & n14362 ;
  assign n14454 = n14453 ^ n14014 ;
  assign n14650 = n14649 ^ n14454 ;
  assign n14651 = n14649 ^ x93 ;
  assign n14652 = n14650 & n14651 ;
  assign n14653 = n14652 ^ x93 ;
  assign n14451 = n14219 & n14362 ;
  assign n14452 = n14451 ^ n14012 ;
  assign n14654 = n14653 ^ n14452 ;
  assign n14655 = n14653 ^ x94 ;
  assign n14656 = n14654 & n14655 ;
  assign n14657 = n14656 ^ x94 ;
  assign n14449 = n14223 & n14362 ;
  assign n14450 = n14449 ^ n14010 ;
  assign n14658 = n14657 ^ n14450 ;
  assign n14659 = n14657 ^ x95 ;
  assign n14660 = n14658 & n14659 ;
  assign n14661 = n14660 ^ x95 ;
  assign n14447 = n14227 & n14362 ;
  assign n14448 = n14447 ^ n14007 ;
  assign n14662 = n14661 ^ n14448 ;
  assign n14663 = n14661 ^ x96 ;
  assign n14664 = n14662 & n14663 ;
  assign n14665 = n14664 ^ x96 ;
  assign n14445 = n14231 & n14362 ;
  assign n14446 = n14445 ^ n14005 ;
  assign n14666 = n14665 ^ n14446 ;
  assign n14667 = n14665 ^ x97 ;
  assign n14668 = n14666 & n14667 ;
  assign n14669 = n14668 ^ x97 ;
  assign n14443 = n14235 & n14362 ;
  assign n14444 = n14443 ^ n14003 ;
  assign n14670 = n14669 ^ n14444 ;
  assign n14671 = n14669 ^ x98 ;
  assign n14672 = n14670 & n14671 ;
  assign n14673 = n14672 ^ x98 ;
  assign n14441 = n14239 & n14362 ;
  assign n14442 = n14441 ^ n14001 ;
  assign n14674 = n14673 ^ n14442 ;
  assign n14675 = n14673 ^ x99 ;
  assign n14676 = n14674 & n14675 ;
  assign n14677 = n14676 ^ x99 ;
  assign n14439 = n14243 & n14362 ;
  assign n14440 = n14439 ^ n13999 ;
  assign n14678 = n14677 ^ n14440 ;
  assign n14679 = n14677 ^ x100 ;
  assign n14680 = n14678 & n14679 ;
  assign n14681 = n14680 ^ x100 ;
  assign n14437 = n14247 & n14362 ;
  assign n14438 = n14437 ^ n13997 ;
  assign n14682 = n14681 ^ n14438 ;
  assign n14683 = n14681 ^ x101 ;
  assign n14684 = n14682 & n14683 ;
  assign n14685 = n14684 ^ x101 ;
  assign n14435 = n14251 & n14362 ;
  assign n14436 = n14435 ^ n13994 ;
  assign n14686 = n14685 ^ n14436 ;
  assign n14687 = n14685 ^ x102 ;
  assign n14688 = n14686 & n14687 ;
  assign n14689 = n14688 ^ x102 ;
  assign n14433 = n14255 & n14362 ;
  assign n14434 = n14433 ^ n13983 ;
  assign n14690 = n14689 ^ n14434 ;
  assign n14691 = n14689 ^ x103 ;
  assign n14692 = n14690 & n14691 ;
  assign n14693 = n14692 ^ x103 ;
  assign n14430 = n14257 ^ x103 ;
  assign n14431 = n14362 & n14430 ;
  assign n14432 = n14431 ^ n13979 ;
  assign n14694 = n14693 ^ n14432 ;
  assign n14695 = n14693 ^ x104 ;
  assign n14696 = n14694 & n14695 ;
  assign n14697 = n14696 ^ x104 ;
  assign n14427 = n14260 ^ x104 ;
  assign n14428 = n14362 & n14427 ;
  assign n14429 = n14428 ^ n13975 ;
  assign n14698 = n14697 ^ n14429 ;
  assign n14699 = n14697 ^ x105 ;
  assign n14700 = n14698 & n14699 ;
  assign n14701 = n14700 ^ x105 ;
  assign n14425 = n14265 & n14362 ;
  assign n14426 = n14425 ^ n13964 ;
  assign n14702 = n14701 ^ n14426 ;
  assign n14703 = n14701 ^ x106 ;
  assign n14704 = n14702 & n14703 ;
  assign n14705 = n14704 ^ x106 ;
  assign n14423 = n14269 & n14362 ;
  assign n14424 = n14423 ^ n13961 ;
  assign n14706 = n14705 ^ n14424 ;
  assign n14707 = n14705 ^ x107 ;
  assign n14708 = n14706 & n14707 ;
  assign n14709 = n14708 ^ x107 ;
  assign n14421 = n14273 & n14362 ;
  assign n14422 = n14421 ^ n13959 ;
  assign n14710 = n14709 ^ n14422 ;
  assign n14711 = n14709 ^ x108 ;
  assign n14712 = n14710 & n14711 ;
  assign n14713 = n14712 ^ x108 ;
  assign n14419 = n14277 & n14362 ;
  assign n14420 = n14419 ^ n13957 ;
  assign n14714 = n14713 ^ n14420 ;
  assign n14715 = n14713 ^ x109 ;
  assign n14716 = n14714 & n14715 ;
  assign n14717 = n14716 ^ x109 ;
  assign n14417 = n14281 & n14362 ;
  assign n14418 = n14417 ^ n13955 ;
  assign n14718 = n14717 ^ n14418 ;
  assign n14719 = n14717 ^ x110 ;
  assign n14720 = n14718 & n14719 ;
  assign n14721 = n14720 ^ x110 ;
  assign n14415 = n14285 & n14362 ;
  assign n14416 = n14415 ^ n13953 ;
  assign n14722 = n14721 ^ n14416 ;
  assign n14723 = n14721 ^ x111 ;
  assign n14724 = n14722 & n14723 ;
  assign n14725 = n14724 ^ x111 ;
  assign n14413 = n14289 & n14362 ;
  assign n14414 = n14413 ^ n13951 ;
  assign n14726 = n14725 ^ n14414 ;
  assign n14727 = n14725 ^ x112 ;
  assign n14728 = n14726 & n14727 ;
  assign n14729 = n14728 ^ x112 ;
  assign n14411 = n14293 & n14362 ;
  assign n14412 = n14411 ^ n13949 ;
  assign n14730 = n14729 ^ n14412 ;
  assign n14731 = n14729 ^ x113 ;
  assign n14732 = n14730 & n14731 ;
  assign n14733 = n14732 ^ x113 ;
  assign n14408 = n14295 ^ x113 ;
  assign n14409 = n14362 & n14408 ;
  assign n14410 = n14409 ^ n13944 ;
  assign n14734 = n14733 ^ n14410 ;
  assign n14735 = n14733 ^ x114 ;
  assign n14736 = n14734 & n14735 ;
  assign n14737 = n14736 ^ x114 ;
  assign n14397 = n13944 ^ x114 ;
  assign n14398 = n14397 ^ n14295 ;
  assign n14399 = n14398 ^ x113 ;
  assign n14400 = n14399 ^ n14397 ;
  assign n14402 = n14295 ^ x114 ;
  assign n14403 = n14402 ^ n14397 ;
  assign n14404 = ~n14400 & ~n14403 ;
  assign n14405 = n14404 ^ n14397 ;
  assign n14406 = n14362 & ~n14405 ;
  assign n14407 = n14406 ^ n13941 ;
  assign n14738 = n14737 ^ n14407 ;
  assign n14739 = n14737 ^ x115 ;
  assign n14740 = n14738 & n14739 ;
  assign n14741 = n14740 ^ x115 ;
  assign n14394 = n14301 ^ x115 ;
  assign n14395 = n14362 & n14394 ;
  assign n14396 = n14395 ^ n14303 ;
  assign n14742 = n14741 ^ n14396 ;
  assign n14743 = n14741 ^ x116 ;
  assign n14744 = n14742 & n14743 ;
  assign n14745 = n14744 ^ x116 ;
  assign n14392 = n14309 & n14362 ;
  assign n14393 = n14392 ^ n13939 ;
  assign n14746 = n14745 ^ n14393 ;
  assign n14747 = n14745 ^ x117 ;
  assign n14748 = n14746 & n14747 ;
  assign n14749 = n14748 ^ x117 ;
  assign n14390 = n14313 & n14362 ;
  assign n14391 = n14390 ^ n13936 ;
  assign n14750 = n14749 ^ n14391 ;
  assign n14751 = n14749 ^ x118 ;
  assign n14752 = n14750 & n14751 ;
  assign n14753 = n14752 ^ x118 ;
  assign n14387 = n14315 ^ x118 ;
  assign n14388 = n14362 & n14387 ;
  assign n14389 = n14388 ^ n13922 ;
  assign n14754 = n14753 ^ n14389 ;
  assign n14755 = n14753 ^ x119 ;
  assign n14756 = n14754 & n14755 ;
  assign n14757 = n14756 ^ x119 ;
  assign n14376 = n13922 ^ x119 ;
  assign n14377 = n14376 ^ n14315 ;
  assign n14378 = n14377 ^ x118 ;
  assign n14379 = n14378 ^ n14376 ;
  assign n14381 = n14315 ^ x119 ;
  assign n14382 = n14381 ^ n14376 ;
  assign n14383 = ~n14379 & ~n14382 ;
  assign n14384 = n14383 ^ n14376 ;
  assign n14385 = n14362 & ~n14384 ;
  assign n14386 = n14385 ^ n13918 ;
  assign n14758 = n14757 ^ n14386 ;
  assign n14759 = n14757 ^ x120 ;
  assign n14760 = n14758 & n14759 ;
  assign n14761 = n14760 ^ x120 ;
  assign n14373 = n14321 ^ x120 ;
  assign n14374 = n14362 & n14373 ;
  assign n14375 = n14374 ^ n14323 ;
  assign n14762 = n14761 ^ n14375 ;
  assign n14763 = n14761 ^ x121 ;
  assign n14764 = n14762 & n14763 ;
  assign n14765 = n14764 ^ x121 ;
  assign n14371 = n14329 & n14362 ;
  assign n14372 = n14371 ^ n13916 ;
  assign n14766 = n14765 ^ n14372 ;
  assign n14767 = n14765 ^ x122 ;
  assign n14768 = n14766 & n14767 ;
  assign n14769 = n14768 ^ x122 ;
  assign n14369 = n14333 & n14362 ;
  assign n14370 = n14369 ^ n13914 ;
  assign n14770 = n14769 ^ n14370 ;
  assign n14771 = n14769 ^ x123 ;
  assign n14772 = n14770 & n14771 ;
  assign n14773 = n14772 ^ x123 ;
  assign n14367 = n14337 & n14362 ;
  assign n14368 = n14367 ^ n13912 ;
  assign n14774 = n14773 ^ n14368 ;
  assign n14775 = n14773 ^ x124 ;
  assign n14776 = n14774 & n14775 ;
  assign n14777 = n14776 ^ x124 ;
  assign n14365 = n14341 & n14362 ;
  assign n14366 = n14365 ^ n13910 ;
  assign n14778 = n14777 ^ n14366 ;
  assign n14779 = n14777 ^ x125 ;
  assign n14780 = n14778 & n14779 ;
  assign n14781 = n14780 ^ x125 ;
  assign n14344 = n14343 ^ x125 ;
  assign n14363 = n14344 & n14362 ;
  assign n14364 = n14363 ^ n14351 ;
  assign n14782 = n14781 ^ n14364 ;
  assign n14783 = n14781 ^ x126 ;
  assign n14784 = n14782 & n14783 ;
  assign n14785 = n14784 ^ x126 ;
  assign n14786 = n14785 ^ x127 ;
  assign n14789 = n14347 & ~n14357 ;
  assign n14790 = n14789 ^ n12971 ;
  assign n14791 = n14785 & ~n14790 ;
  assign n14792 = n14791 ^ n12971 ;
  assign n14793 = n14786 & ~n14792 ;
  assign n14794 = n14793 ^ n14785 ;
  assign n14795 = n251 ^ n208 ;
  assign n14796 = ~x65 & ~x66 ;
  assign n14797 = n189 & n14796 ;
  assign n14798 = ~x63 & x64 ;
  assign n14799 = n14797 & n14798 ;
  assign n14800 = n14799 ^ n14797 ;
  assign n14801 = x64 & ~n14794 ;
  assign n14802 = n14801 ^ x0 ;
  assign n14808 = x64 & n14362 ;
  assign n14804 = ~x0 & x64 ;
  assign n14805 = n14804 ^ x65 ;
  assign n14806 = ~n14794 & n14805 ;
  assign n14807 = n14806 ^ x1 ;
  assign n14809 = n14808 ^ n14807 ;
  assign n14810 = n14531 ^ x66 ;
  assign n14811 = ~n14794 & n14810 ;
  assign n14812 = n14811 ^ n14538 ;
  assign n14813 = n14542 ^ x67 ;
  assign n14814 = ~n14794 & n14813 ;
  assign n14815 = n14814 ^ n14545 ;
  assign n14816 = n14549 ^ x68 ;
  assign n14817 = ~n14794 & n14816 ;
  assign n14818 = n14817 ^ n14551 ;
  assign n14819 = n14557 & ~n14794 ;
  assign n14820 = n14819 ^ n14519 ;
  assign n14821 = n14561 & ~n14794 ;
  assign n14822 = n14821 ^ n14516 ;
  assign n14823 = n14563 ^ x71 ;
  assign n14824 = ~n14794 & n14823 ;
  assign n14825 = n14824 ^ n14504 ;
  assign n14826 = n14566 ^ x72 ;
  assign n14827 = ~n14794 & n14826 ;
  assign n14828 = n14827 ^ n14500 ;
  assign n14829 = n14571 & ~n14794 ;
  assign n14830 = n14829 ^ n14498 ;
  assign n14831 = n14575 & ~n14794 ;
  assign n14832 = n14831 ^ n14496 ;
  assign n14833 = n14579 & ~n14794 ;
  assign n14834 = n14833 ^ n14494 ;
  assign n14835 = n14581 ^ x76 ;
  assign n14836 = ~n14794 & n14835 ;
  assign n14837 = n14836 ^ n14489 ;
  assign n14838 = n14489 ^ x77 ;
  assign n14839 = n14838 ^ n14581 ;
  assign n14840 = n14839 ^ x76 ;
  assign n14841 = n14840 ^ n14838 ;
  assign n14843 = n14581 ^ x77 ;
  assign n14844 = n14843 ^ n14838 ;
  assign n14845 = ~n14841 & ~n14844 ;
  assign n14846 = n14845 ^ n14838 ;
  assign n14847 = ~n14794 & ~n14846 ;
  assign n14848 = n14847 ^ n14486 ;
  assign n14849 = n14587 ^ x78 ;
  assign n14850 = ~n14794 & n14849 ;
  assign n14851 = n14850 ^ n14589 ;
  assign n14852 = n14595 & ~n14794 ;
  assign n14853 = n14852 ^ n14484 ;
  assign n14854 = n14599 & ~n14794 ;
  assign n14855 = n14854 ^ n14482 ;
  assign n14856 = n14603 & ~n14794 ;
  assign n14857 = n14856 ^ n14480 ;
  assign n14858 = n14607 & ~n14794 ;
  assign n14859 = n14858 ^ n14478 ;
  assign n14860 = n14611 & ~n14794 ;
  assign n14861 = n14860 ^ n14476 ;
  assign n14862 = n14615 & ~n14794 ;
  assign n14863 = n14862 ^ n14474 ;
  assign n14864 = n14619 & ~n14794 ;
  assign n14865 = n14864 ^ n14472 ;
  assign n14866 = n14621 ^ x86 ;
  assign n14867 = ~n14794 & n14866 ;
  assign n14868 = n14867 ^ n14467 ;
  assign n14869 = n14467 ^ x87 ;
  assign n14870 = n14869 ^ n14621 ;
  assign n14871 = n14870 ^ x86 ;
  assign n14872 = n14871 ^ n14869 ;
  assign n14874 = n14621 ^ x87 ;
  assign n14875 = n14874 ^ n14869 ;
  assign n14876 = ~n14872 & ~n14875 ;
  assign n14877 = n14876 ^ n14869 ;
  assign n14878 = ~n14794 & ~n14877 ;
  assign n14879 = n14878 ^ n14464 ;
  assign n14880 = n14627 ^ x88 ;
  assign n14881 = ~n14794 & n14880 ;
  assign n14882 = n14881 ^ n14629 ;
  assign n14883 = n14635 & ~n14794 ;
  assign n14884 = n14883 ^ n14462 ;
  assign n14885 = n14639 & ~n14794 ;
  assign n14886 = n14885 ^ n14460 ;
  assign n14887 = n14643 & ~n14794 ;
  assign n14888 = n14887 ^ n14458 ;
  assign n14889 = n14647 & ~n14794 ;
  assign n14890 = n14889 ^ n14456 ;
  assign n14891 = n14651 & ~n14794 ;
  assign n14892 = n14891 ^ n14454 ;
  assign n14893 = n14655 & ~n14794 ;
  assign n14894 = n14893 ^ n14452 ;
  assign n14895 = n14659 & ~n14794 ;
  assign n14896 = n14895 ^ n14450 ;
  assign n14897 = n14663 & ~n14794 ;
  assign n14898 = n14897 ^ n14448 ;
  assign n14899 = n14667 & ~n14794 ;
  assign n14900 = n14899 ^ n14446 ;
  assign n14901 = n14671 & ~n14794 ;
  assign n14902 = n14901 ^ n14444 ;
  assign n14903 = n14675 & ~n14794 ;
  assign n14904 = n14903 ^ n14442 ;
  assign n14905 = n14679 & ~n14794 ;
  assign n14906 = n14905 ^ n14440 ;
  assign n14907 = n14683 & ~n14794 ;
  assign n14908 = n14907 ^ n14438 ;
  assign n14909 = n14687 & ~n14794 ;
  assign n14910 = n14909 ^ n14436 ;
  assign n14911 = n14691 & ~n14794 ;
  assign n14912 = n14911 ^ n14434 ;
  assign n14913 = n14695 & ~n14794 ;
  assign n14914 = n14913 ^ n14432 ;
  assign n14915 = n14699 & ~n14794 ;
  assign n14916 = n14915 ^ n14429 ;
  assign n14917 = n14703 & ~n14794 ;
  assign n14918 = n14917 ^ n14426 ;
  assign n14919 = n14707 & ~n14794 ;
  assign n14920 = n14919 ^ n14424 ;
  assign n14921 = n14711 & ~n14794 ;
  assign n14922 = n14921 ^ n14422 ;
  assign n14923 = n14715 & ~n14794 ;
  assign n14924 = n14923 ^ n14420 ;
  assign n14925 = n14719 & ~n14794 ;
  assign n14926 = n14925 ^ n14418 ;
  assign n14927 = n14723 & ~n14794 ;
  assign n14928 = n14927 ^ n14416 ;
  assign n14929 = n14727 & ~n14794 ;
  assign n14930 = n14929 ^ n14414 ;
  assign n14931 = n14731 & ~n14794 ;
  assign n14932 = n14931 ^ n14412 ;
  assign n14933 = n14735 & ~n14794 ;
  assign n14934 = n14933 ^ n14410 ;
  assign n14935 = n14739 & ~n14794 ;
  assign n14936 = n14935 ^ n14407 ;
  assign n14937 = n14743 & ~n14794 ;
  assign n14938 = n14937 ^ n14396 ;
  assign n14939 = n14747 & ~n14794 ;
  assign n14940 = n14939 ^ n14393 ;
  assign n14941 = n14751 & ~n14794 ;
  assign n14942 = n14941 ^ n14391 ;
  assign n14943 = n14755 & ~n14794 ;
  assign n14944 = n14943 ^ n14389 ;
  assign n14945 = n14759 & ~n14794 ;
  assign n14946 = n14945 ^ n14386 ;
  assign n14947 = n14763 & ~n14794 ;
  assign n14948 = n14947 ^ n14375 ;
  assign n14949 = n14767 & ~n14794 ;
  assign n14950 = n14949 ^ n14372 ;
  assign n14951 = n14771 & ~n14794 ;
  assign n14952 = n14951 ^ n14370 ;
  assign n14953 = n14775 & ~n14794 ;
  assign n14954 = n14953 ^ n14368 ;
  assign n14955 = n14779 & ~n14794 ;
  assign n14956 = n14955 ^ n14366 ;
  assign n14957 = n14783 & ~n14794 ;
  assign n14958 = n14957 ^ n14364 ;
  assign n14959 = n14347 & ~n14786 ;
  assign n14960 = ~n14785 & n14959 ;
  assign n14961 = n14357 & n14960 ;
  assign n14962 = n14961 ^ n14959 ;
  assign y0 = ~n14794 ;
  assign y1 = n14362 ;
  assign y2 = n13908 ;
  assign y3 = n13451 ;
  assign y4 = n13005 ;
  assign y5 = n12592 ;
  assign y6 = n12195 ;
  assign y7 = n11788 ;
  assign y8 = n11409 ;
  assign y9 = n11001 ;
  assign y10 = n10575 ;
  assign y11 = n10212 ;
  assign y12 = n9788 ;
  assign y13 = n9428 ;
  assign y14 = n9045 ;
  assign y15 = n8707 ;
  assign y16 = n8357 ;
  assign y17 = n8026 ;
  assign y18 = n7696 ;
  assign y19 = n7360 ;
  assign y20 = n7028 ;
  assign y21 = n6697 ;
  assign y22 = n6379 ;
  assign y23 = n6087 ;
  assign y24 = n5811 ;
  assign y25 = n5536 ;
  assign y26 = n5246 ;
  assign y27 = n4950 ;
  assign y28 = n4679 ;
  assign y29 = n4447 ;
  assign y30 = n4227 ;
  assign y31 = n3999 ;
  assign y32 = n3771 ;
  assign y33 = n3559 ;
  assign y34 = n3323 ;
  assign y35 = n3113 ;
  assign y36 = n2927 ;
  assign y37 = n2742 ;
  assign y38 = n2557 ;
  assign y39 = n2384 ;
  assign y40 = n2229 ;
  assign y41 = n2065 ;
  assign y42 = n1914 ;
  assign y43 = n1779 ;
  assign y44 = n1639 ;
  assign y45 = n1502 ;
  assign y46 = n1386 ;
  assign y47 = n1266 ;
  assign y48 = n1159 ;
  assign y49 = n1065 ;
  assign y50 = n966 ;
  assign y51 = n879 ;
  assign y52 = n792 ;
  assign y53 = n711 ;
  assign y54 = n626 ;
  assign y55 = n546 ;
  assign y56 = n480 ;
  assign y57 = n423 ;
  assign y58 = n372 ;
  assign y59 = n330 ;
  assign y60 = n285 ;
  assign y61 = n241 ;
  assign y62 = n14795 ;
  assign y63 = n14800 ;
  assign y64 = n14802 ;
  assign y65 = n14809 ;
  assign y66 = n14812 ;
  assign y67 = n14815 ;
  assign y68 = n14818 ;
  assign y69 = n14820 ;
  assign y70 = n14822 ;
  assign y71 = n14825 ;
  assign y72 = n14828 ;
  assign y73 = n14830 ;
  assign y74 = n14832 ;
  assign y75 = n14834 ;
  assign y76 = n14837 ;
  assign y77 = n14848 ;
  assign y78 = n14851 ;
  assign y79 = n14853 ;
  assign y80 = n14855 ;
  assign y81 = n14857 ;
  assign y82 = n14859 ;
  assign y83 = n14861 ;
  assign y84 = n14863 ;
  assign y85 = n14865 ;
  assign y86 = n14868 ;
  assign y87 = n14879 ;
  assign y88 = n14882 ;
  assign y89 = n14884 ;
  assign y90 = n14886 ;
  assign y91 = n14888 ;
  assign y92 = n14890 ;
  assign y93 = n14892 ;
  assign y94 = n14894 ;
  assign y95 = n14896 ;
  assign y96 = n14898 ;
  assign y97 = n14900 ;
  assign y98 = n14902 ;
  assign y99 = n14904 ;
  assign y100 = n14906 ;
  assign y101 = n14908 ;
  assign y102 = n14910 ;
  assign y103 = n14912 ;
  assign y104 = n14914 ;
  assign y105 = n14916 ;
  assign y106 = n14918 ;
  assign y107 = n14920 ;
  assign y108 = n14922 ;
  assign y109 = n14924 ;
  assign y110 = n14926 ;
  assign y111 = n14928 ;
  assign y112 = n14930 ;
  assign y113 = n14932 ;
  assign y114 = n14934 ;
  assign y115 = n14936 ;
  assign y116 = n14938 ;
  assign y117 = n14940 ;
  assign y118 = n14942 ;
  assign y119 = n14944 ;
  assign y120 = n14946 ;
  assign y121 = n14948 ;
  assign y122 = n14950 ;
  assign y123 = n14952 ;
  assign y124 = n14954 ;
  assign y125 = n14956 ;
  assign y126 = n14958 ;
  assign y127 = n14962 ;
endmodule
