module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528, n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552, n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677, n_5678, n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705, n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713, n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743, n_5744, n_5745, n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772, n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789, n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907, n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983, n_5984, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208, n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263, n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311, n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319, n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359, n_6360, n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408, n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416, n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424, n_6425, n_6426, n_6427, n_6428, n_6429, n_6430, n_6431, n_6432, n_6433, n_6434, n_6435, n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443, n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457, n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, n_6465, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472, n_6473, n_6474, n_6475, n_6476, n_6477, n_6478, n_6479, n_6480, n_6481, n_6482, n_6483, n_6484, n_6485, n_6486, n_6487, n_6488, n_6489, n_6490, n_6491, n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504, n_6505, n_6506, n_6507, n_6508, n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524, n_6525, n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540, n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556, n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564, n_6565, n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572, n_6573, n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592, n_6593, n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608, n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617, n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704, n_6705, n_6706, n_6707, n_6708, n_6709, n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723, n_6724, n_6725, n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740, n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748, n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764, n_6765, n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772, n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788, n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796, n_6797, n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804, n_6805, n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812, n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820, n_6821, n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828, n_6829, n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6839, n_6840, n_6841, n_6842, n_6843, n_6844, n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853, n_6854, n_6855, n_6856, n_6857, n_6858, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864, n_6865, n_6866, n_6867, n_6868, n_6869, n_6870, n_6871, n_6872, n_6873, n_6874, n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881, n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888, n_6889, n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6898, n_6899, n_6900, n_6901, n_6902, n_6903, n_6904, n_6905, n_6906, n_6907, n_6908, n_6909, n_6910, n_6911, n_6912, n_6913, n_6914, n_6915, n_6916, n_6917, n_6918, n_6919, n_6920, n_6921, n_6922, n_6923, n_6924, n_6925, n_6926, n_6927, n_6928, n_6929, n_6930, n_6931, n_6932, n_6933, n_6934, n_6935, n_6936, n_6937, n_6938, n_6939, n_6940, n_6941, n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948, n_6949, n_6950, n_6951, n_6952, n_6953, n_6954, n_6955, n_6956, n_6957, n_6958, n_6959, n_6960, n_6961, n_6962, n_6963, n_6964, n_6965, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971, n_6972, n_6973, n_6974, n_6975, n_6976, n_6977, n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, n_7003, n_7004, n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012, n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020, n_7021, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030, n_7031, n_7032, n_7033, n_7034, n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041, n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7056, n_7057, n_7058, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065, n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073, n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081, n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089, n_7090, n_7091, n_7092, n_7093, n_7094, n_7095, n_7096, n_7097, n_7098, n_7099, n_7100, n_7101, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108, n_7109, n_7110, n_7111, n_7112, n_7113, n_7114, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129, n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136, n_7137, n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145, n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153, n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7160, n_7161, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172, n_7173, n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181, n_7182, n_7183, n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198, n_7199, n_7200, n_7201, n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212, n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220, n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228, n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236, n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7256, n_7257, n_7258, n_7259, n_7260, n_7261, n_7262, n_7263, n_7264, n_7265, n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273, n_7274, n_7275, n_7276, n_7277, n_7278, n_7279, n_7280, n_7281, n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288, n_7289, n_7290, n_7291, n_7292, n_7293, n_7294, n_7295, n_7296, n_7297, n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304, n_7305, n_7306, n_7307, n_7308, n_7309, n_7310, n_7311, n_7312, n_7313, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332, n_7333, n_7334, n_7335, n_7336, n_7337, n_7338, n_7339, n_7340, n_7341, n_7342, n_7343, n_7344, n_7345, n_7346, n_7347, n_7348, n_7349, n_7350, n_7351, n_7352, n_7353, n_7354, n_7355, n_7356, n_7357, n_7358, n_7359, n_7360, n_7361, n_7362, n_7363, n_7364, n_7365, n_7366, n_7367, n_7368, n_7369, n_7370, n_7371, n_7372, n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, n_7380, n_7381, n_7382, n_7383, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389, n_7390, n_7391, n_7392, n_7393, n_7394, n_7395, n_7396, n_7397, n_7398, n_7399, n_7400, n_7401, n_7402, n_7403, n_7404, n_7405, n_7406, n_7407, n_7408, n_7409, n_7410, n_7411, n_7412, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7421, n_7422, n_7423, n_7424, n_7425, n_7426, n_7427, n_7428, n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7435, n_7436, n_7437, n_7438, n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7446, n_7447, n_7448, n_7449, n_7450, n_7451, n_7452, n_7453, n_7454, n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461, n_7462, n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469, n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502, n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518, n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541, n_7542, n_7543, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552, n_7553, n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565, n_7566, n_7567, n_7568, n_7569, n_7570, n_7571, n_7572, n_7573, n_7574, n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7584, n_7585, n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596, n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603, n_7604, n_7605, n_7606, n_7607, n_7608, n_7609, n_7610, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625, n_7626, n_7627, n_7628, n_7629, n_7630, n_7631, n_7632, n_7633, n_7634, n_7635, n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643, n_7644, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650, n_7651, n_7652, n_7653, n_7654, n_7655, n_7656, n_7657, n_7658, n_7659, n_7660, n_7661, n_7662, n_7663, n_7664, n_7665, n_7666, n_7667, n_7668, n_7669, n_7670, n_7671, n_7672, n_7673, n_7674, n_7675, n_7676, n_7677, n_7678, n_7679, n_7680, n_7681, n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688, n_7689, n_7690, n_7691, n_7692, n_7693, n_7694, n_7695, n_7696, n_7697, n_7698, n_7699, n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, n_7706, n_7707, n_7708, n_7709, n_7710, n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717, n_7718, n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726, n_7727, n_7728, n_7729, n_7730, n_7731, n_7732, n_7733, n_7734, n_7735, n_7736, n_7737, n_7738, n_7739, n_7740, n_7741, n_7742, n_7743, n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750, n_7751, n_7752, n_7753, n_7754, n_7755, n_7756, n_7757, n_7758, n_7759, n_7760, n_7761, n_7762, n_7763, n_7764, n_7765, n_7766, n_7767, n_7768, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781, n_7782, n_7783, n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7806, n_7807, n_7808, n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816, n_7817, n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824, n_7825, n_7826, n_7827, n_7828, n_7829, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835, n_7836, n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7843, n_7844, n_7845, n_7846, n_7847, n_7848, n_7849, n_7850, n_7851, n_7852, n_7853, n_7854, n_7855, n_7856, n_7857, n_7858, n_7859, n_7860, n_7861, n_7862, n_7863, n_7864, n_7865, n_7866, n_7867, n_7868, n_7869, n_7870, n_7871, n_7872, n_7873, n_7874, n_7875, n_7876, n_7877, n_7878, n_7879, n_7880, n_7881, n_7882, n_7883, n_7884, n_7885, n_7886, n_7887, n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, n_7895, n_7896, n_7897, n_7898, n_7899, n_7900, n_7901, n_7902, n_7903, n_7904, n_7905, n_7906, n_7907, n_7908, n_7909, n_7910, n_7911, n_7912, n_7913, n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920, n_7921, n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928, n_7929, n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937, n_7938, n_7939, n_7940, n_7941, n_7942, n_7943, n_7944, n_7945, n_7946, n_7947, n_7948, n_7949, n_7950, n_7951, n_7952, n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960, n_7961, n_7962, n_7963, n_7964, n_7965, n_7966, n_7967, n_7968, n_7969, n_7970, n_7971, n_7972, n_7973, n_7974, n_7975, n_7976, n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991, n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999, n_8000, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007, n_8008, n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016, n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025, n_8026, n_8027, n_8028, n_8029, n_8030, n_8031, n_8032, n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, n_8039, n_8040, n_8041, n_8042, n_8043, n_8044, n_8045, n_8046, n_8047, n_8048, n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055, n_8056, n_8057, n_8058, n_8059, n_8060, n_8061, n_8062, n_8063, n_8064, n_8065, n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072, n_8073, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080, n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088, n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096, n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104, n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112, n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120, n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128, n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136, n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144, n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152, n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160, n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168, n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176, n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184, n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192, n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200, n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208, n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216, n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224, n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232, n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240, n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248, n_8249, n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256, n_8257, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272, n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280, n_8281, n_8282, n_8283, n_8284, n_8285, n_8286, n_8287, n_8288, n_8289, n_8290, n_8291, n_8292, n_8293, n_8294, n_8295, n_8296, n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304, n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320, n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328, n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354, n_8355, n_8356, n_8357, n_8358, n_8359, n_8360, n_8361, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367, n_8368, n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376, n_8377, n_8378, n_8379, n_8380, n_8381, n_8382, n_8383, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389, n_8390, n_8391, n_8392, n_8393, n_8394, n_8395, n_8396, n_8397, n_8398, n_8399, n_8400, n_8401, n_8402, n_8403, n_8404, n_8405, n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416, n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424, n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432, n_8433, n_8434, n_8435, n_8436, n_8437, n_8438, n_8439, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448, n_8449, n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456, n_8457, n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464, n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472, n_8473, n_8474, n_8475, n_8476, n_8477, n_8478, n_8479, n_8480, n_8481, n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488, n_8489, n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496, n_8497, n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, n_8504, n_8505, n_8506, n_8507, n_8508, n_8509, n_8510, n_8511, n_8512, n_8513, n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528, n_8529, n_8530, n_8531, n_8532, n_8533, n_8534, n_8535, n_8536, n_8537, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544, n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552, n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560, n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568, n_8569, n_8570, n_8571, n_8572, n_8573, n_8574, n_8575, n_8576, n_8577, n_8578, n_8579, n_8580, n_8581, n_8582, n_8583, n_8584, n_8585, n_8586, n_8587, n_8588, n_8589, n_8590, n_8591, n_8592, n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600, n_8601, n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613, n_8614, n_8615, n_8616, n_8617, n_8618, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8625, n_8626, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632, n_8633, n_8634, n_8635, n_8636, n_8637, n_8638, n_8639, n_8640, n_8641, n_8642, n_8643, n_8644, n_8645, n_8646, n_8647, n_8648, n_8649, n_8650, n_8651, n_8652, n_8653, n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8660, n_8661, n_8662, n_8663, n_8664, n_8665, n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, n_8672, n_8673, n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681, n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689, n_8690, n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697, n_8698, n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705, n_8706, n_8707, n_8708, n_8709, n_8710, n_8711, n_8712, n_8713, n_8714, n_8715, n_8716, n_8717, n_8718, n_8719, n_8720, n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727, n_8728, n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735, n_8736, n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743, n_8744, n_8745, n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8752, n_8753, n_8754, n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761, n_8762, n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769, n_8770, n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777, n_8778, n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786, n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793, n_8794, n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802, n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8809, n_8810, n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817, n_8818, n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, n_8825, n_8826, n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833, n_8834, n_8835, n_8836, n_8837, n_8838, n_8839, n_8840, n_8841, n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8848, n_8849, n_8850, n_8851, n_8852, n_8853, n_8854, n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861, n_8862, n_8863, n_8864, n_8865, n_8866, n_8867, n_8868, n_8869, n_8870, n_8871, n_8872, n_8873, n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881, n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889, n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897, n_8898, n_8899, n_8900, n_8901, n_8902, n_8903, n_8904, n_8905, n_8906, n_8907, n_8908, n_8909, n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916, n_8917, n_8918, n_8919, n_8920, n_8921, n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928, n_8929, n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936, n_8937, n_8938, n_8939, n_8940, n_8941, n_8942, n_8943, n_8944, n_8945, n_8946, n_8947, n_8948, n_8949, n_8950, n_8951, n_8952, n_8953, n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960, n_8961, n_8962, n_8963, n_8964, n_8965, n_8966, n_8967, n_8968, n_8969, n_8970, n_8971, n_8972, n_8973, n_8974, n_8975, n_8976, n_8977, n_8978, n_8979, n_8980, n_8981, n_8982, n_8983, n_8984, n_8985, n_8986, n_8987, n_8988, n_8989, n_8990, n_8991, n_8992, n_8993, n_8994, n_8995, n_8996, n_8997, n_8998, n_8999, n_9000, n_9001, n_9002, n_9003, n_9004, n_9005, n_9006, n_9007, n_9008, n_9009, n_9010, n_9011, n_9012, n_9013, n_9014, n_9015, n_9016, n_9017, n_9018, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024, n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032, n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040, n_9041, n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048, n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056, n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9064, n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071, n_9072, n_9073, n_9074, n_9075, n_9076, n_9077, n_9078, n_9079, n_9080, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087, n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095, n_9096, n_9097, n_9098, n_9099, n_9100, n_9101, n_9102, n_9103, n_9104, n_9105, n_9106, n_9107, n_9108, n_9109, n_9110, n_9111, n_9112, n_9113, n_9114, n_9115, n_9116, n_9117, n_9118, n_9119, n_9120, n_9121, n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128, n_9129, n_9130, n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137, n_9138, n_9139, n_9140, n_9141, n_9142, n_9143, n_9144, n_9145, n_9146, n_9147, n_9148, n_9149, n_9150, n_9151, n_9152, n_9153, n_9154, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160, n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9168, n_9169, n_9170, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176, n_9177, n_9178, n_9179, n_9180, n_9181, n_9182, n_9183, n_9184, n_9185, n_9186, n_9187, n_9188, n_9189, n_9190, n_9191, n_9192, n_9193, n_9194, n_9195, n_9196, n_9197, n_9198, n_9199, n_9200, n_9201, n_9202, n_9203, n_9204, n_9205, n_9206, n_9207, n_9208, n_9209, n_9210, n_9211, n_9212, n_9213, n_9214, n_9215, n_9216, n_9217, n_9218, n_9219, n_9220, n_9221, n_9222, n_9223, n_9224, n_9225, n_9226, n_9227, n_9228, n_9229, n_9230, n_9231, n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9239, n_9240, n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9247, n_9248, n_9249, n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256, n_9257, n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265, n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, n_9273, n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281, n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288, n_9289, n_9290, n_9291, n_9292, n_9293, n_9294, n_9295, n_9296, n_9297, n_9298, n_9299, n_9300, n_9301, n_9302, n_9303, n_9304, n_9305, n_9306, n_9307, n_9308, n_9309, n_9310, n_9311, n_9312, n_9313, n_9314, n_9315, n_9316, n_9317, n_9318, n_9319, n_9320, n_9321, n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9328, n_9329, n_9330, n_9331, n_9332, n_9333, n_9334, n_9335, n_9336, n_9337, n_9338, n_9339, n_9340, n_9341, n_9342, n_9343, n_9344, n_9345, n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353, n_9354, n_9355, n_9356, n_9357, n_9358, n_9359, n_9360, n_9361, n_9362, n_9363, n_9364, n_9365, n_9366, n_9367, n_9368, n_9369, n_9370, n_9371, n_9372, n_9373, n_9374, n_9375, n_9376, n_9377, n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9384, n_9385, n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396, n_9397, n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405, n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413, n_9414, n_9415, n_9416, n_9417, n_9418, n_9419, n_9420, n_9421, n_9422, n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430, n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438, n_9439, n_9440, n_9441, n_9442, n_9443, n_9444, n_9445, n_9446, n_9447, n_9448, n_9449, n_9450, n_9451, n_9452, n_9453, n_9454, n_9455, n_9456, n_9457, n_9458, n_9459, n_9460, n_9461, n_9462, n_9463, n_9464, n_9465, n_9466, n_9467, n_9468, n_9469, n_9470, n_9471, n_9472, n_9473, n_9474, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480, n_9481, n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489, n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496, n_9497, n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504, n_9505, n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512, n_9513, n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520, n_9521, n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, n_9528, n_9529, n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536, n_9537, n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545, n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552, n_9553, n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561, n_9562, n_9563, n_9564, n_9565, n_9566, n_9567, n_9568, n_9569, n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576, n_9577, n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584, n_9585, n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, n_9596, n_9597, n_9598, n_9599, n_9600, n_9601, n_9602, n_9603, n_9604, n_9605, n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612, n_9613, n_9614, n_9615, n_9616, n_9617, n_9618, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624, n_9625, n_9626, n_9627, n_9628, n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635, n_9636, n_9637, n_9638, n_9639, n_9640, n_9641, n_9642, n_9643, n_9644, n_9645, n_9646, n_9647, n_9648, n_9649, n_9650, n_9651, n_9652, n_9653, n_9654, n_9655, n_9656, n_9657, n_9658, n_9659, n_9660, n_9661, n_9662, n_9663, n_9664, n_9665, n_9666, n_9667, n_9668, n_9669, n_9670, n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677, n_9678, n_9679, n_9680, n_9681, n_9682, n_9683, n_9684, n_9685, n_9686, n_9687, n_9688, n_9689, n_9690, n_9691, n_9692, n_9693, n_9694, n_9695, n_9696, n_9697, n_9698, n_9699, n_9700, n_9701, n_9702, n_9703, n_9704, n_9705, n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712, n_9713, n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720, n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728, n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736, n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744, n_9745, n_9746, n_9747, n_9748, n_9749, n_9750, n_9751, n_9752, n_9753, n_9754, n_9755, n_9756, n_9757, n_9758, n_9759, n_9760, n_9761, n_9762, n_9763, n_9764, n_9765, n_9766, n_9767, n_9768, n_9769, n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776, n_9777, n_9778, n_9779, n_9780, n_9781, n_9782, n_9783, n_9784, n_9785, n_9786, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792, n_9793, n_9794, n_9795, n_9796, n_9797, n_9798, n_9799, n_9800, n_9801, n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808, n_9809, n_9810, n_9811, n_9812, n_9813, n_9814, n_9815, n_9816, n_9817, n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_9825, n_9826, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832, n_9833, n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848, n_9849, n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856, n_9857, n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864, n_9865, n_9866, n_9867, n_9868, n_9869, n_9870, n_9871, n_9872, n_9873, n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880, n_9881, n_9882, n_9883, n_9884, n_9885, n_9886, n_9887, n_9888, n_9889, n_9890, n_9891, n_9892, n_9893, n_9894, n_9895, n_9896, n_9897, n_9898, n_9899, n_9900, n_9901, n_9902, n_9903, n_9904, n_9905, n_9906, n_9907, n_9908, n_9909, n_9910, n_9911, n_9912, n_9913, n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920, n_9921, n_9922, n_9923, n_9924, n_9925, n_9926, n_9927, n_9928, n_9929, n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937, n_9938, n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945, n_9946, n_9947, n_9948, n_9949, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955, n_9956, n_9957, n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964, n_9965, n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972, n_9973, n_9974, n_9975, n_9976, n_9977, n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984, n_9985, n_9986, n_9987, n_9988, n_9989, n_9990, n_9991, n_9992, n_9993, n_9994, n_9995, n_9996, n_9997, n_9998, n_9999, n_10000, n_10001, n_10002, n_10003, n_10004, n_10005, n_10006, n_10007, n_10008, n_10009, n_10010, n_10011, n_10012, n_10013, n_10014, n_10015, n_10016, n_10017, n_10018, n_10019, n_10020, n_10021, n_10022, n_10023, n_10024, n_10025, n_10026, n_10027, n_10028, n_10029, n_10030, n_10031, n_10032, n_10033, n_10034, n_10035, n_10036, n_10037, n_10038, n_10039, n_10040, n_10041, n_10042, n_10043, n_10044, n_10045, n_10046, n_10047, n_10048, n_10049, n_10050, n_10051, n_10052, n_10053, n_10054, n_10055, n_10056, n_10057, n_10058, n_10059, n_10060, n_10061, n_10062, n_10063, n_10064, n_10065, n_10066, n_10067, n_10068, n_10069, n_10070, n_10071, n_10072, n_10073, n_10074, n_10075, n_10076, n_10077, n_10078, n_10079, n_10080, n_10081, n_10082, n_10083, n_10084, n_10085, n_10086, n_10087, n_10088, n_10089, n_10090, n_10091, n_10092, n_10093, n_10094, n_10095, n_10096, n_10097, n_10098, n_10099, n_10100, n_10101, n_10102, n_10103, n_10104, n_10105, n_10106, n_10107, n_10108, n_10109, n_10110, n_10111, n_10112, n_10113, n_10114, n_10115, n_10116, n_10117, n_10118, n_10119, n_10120, n_10121, n_10122, n_10123, n_10124, n_10125, n_10126, n_10127, n_10128, n_10129, n_10130, n_10131, n_10132, n_10133, n_10134, n_10135, n_10136, n_10137, n_10138, n_10139, n_10140, n_10141, n_10142, n_10143, n_10144, n_10145, n_10146, n_10147, n_10148, n_10149, n_10150, n_10151, n_10152, n_10153, n_10154, n_10155, n_10156, n_10157, n_10158, n_10159, n_10160, n_10161, n_10162, n_10163, n_10164, n_10165, n_10166, n_10167, n_10168, n_10169, n_10170, n_10171, n_10172, n_10173, n_10174, n_10175, n_10176, n_10177, n_10178, n_10179, n_10180, n_10181, n_10182, n_10183, n_10184, n_10185, n_10186, n_10187, n_10188, n_10189, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195, n_10196, n_10197, n_10198, n_10199, n_10200, n_10201, n_10202, n_10203, n_10204, n_10205, n_10206, n_10207, n_10208, n_10209, n_10210, n_10211, n_10212, n_10213, n_10214, n_10215, n_10216, n_10217, n_10218, n_10219, n_10220, n_10221, n_10222, n_10223, n_10224, n_10225, n_10226, n_10227, n_10228, n_10229, n_10230, n_10231, n_10232, n_10233, n_10234, n_10235, n_10236, n_10237, n_10238, n_10239, n_10240, n_10241, n_10242, n_10243, n_10244, n_10245, n_10246, n_10247, n_10248, n_10249, n_10250, n_10251, n_10252, n_10253, n_10254, n_10255, n_10256, n_10257, n_10258, n_10259, n_10260, n_10261, n_10262, n_10263, n_10264, n_10265, n_10266, n_10267, n_10268, n_10269, n_10270, n_10271, n_10272, n_10273, n_10274, n_10275, n_10276, n_10277, n_10278, n_10279, n_10280, n_10281, n_10282, n_10283, n_10284, n_10285, n_10286, n_10287, n_10288, n_10289, n_10290, n_10291, n_10292, n_10293, n_10294, n_10295, n_10296, n_10297, n_10298, n_10299, n_10300, n_10301, n_10302, n_10303, n_10304, n_10305, n_10306, n_10307, n_10308, n_10309, n_10310, n_10311, n_10312, n_10313, n_10314, n_10315, n_10316, n_10317, n_10318, n_10319, n_10320, n_10321, n_10322, n_10323, n_10324, n_10325, n_10326, n_10327, n_10328, n_10329, n_10330, n_10331, n_10332, n_10333, n_10334, n_10335, n_10336, n_10337, n_10338, n_10339, n_10340, n_10341, n_10342, n_10343, n_10344, n_10345, n_10346, n_10347, n_10348, n_10349, n_10350, n_10351, n_10352, n_10353, n_10354, n_10355, n_10356, n_10357, n_10358, n_10359, n_10360, n_10361, n_10362, n_10363, n_10364, n_10365, n_10366, n_10367, n_10368, n_10369, n_10370, n_10371, n_10372, n_10373, n_10374, n_10375, n_10376, n_10377, n_10378, n_10379, n_10380, n_10381, n_10382, n_10383, n_10384, n_10385, n_10386, n_10387, n_10388, n_10389, n_10390, n_10391, n_10392, n_10393, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399, n_10400, n_10401, n_10402, n_10403, n_10404, n_10405, n_10406, n_10407, n_10408, n_10409, n_10410, n_10411, n_10412, n_10413, n_10414, n_10415, n_10416, n_10417, n_10418, n_10419, n_10420, n_10421, n_10422, n_10423, n_10424, n_10425, n_10426, n_10427, n_10428, n_10429, n_10430, n_10431, n_10432, n_10433, n_10434, n_10435, n_10436, n_10437, n_10438, n_10439, n_10440, n_10441, n_10442, n_10443, n_10444, n_10445, n_10446, n_10447, n_10448, n_10449, n_10450, n_10451, n_10452, n_10453, n_10454, n_10455, n_10456, n_10457, n_10458, n_10459, n_10460, n_10461, n_10462, n_10463, n_10464, n_10465, n_10466, n_10467, n_10468, n_10469, n_10470, n_10471, n_10472, n_10473, n_10474, n_10475, n_10476, n_10477, n_10478, n_10479, n_10480, n_10481, n_10482, n_10483, n_10484, n_10485, n_10486, n_10487, n_10488, n_10489, n_10490, n_10491, n_10492, n_10493, n_10494, n_10495, n_10496, n_10497, n_10498, n_10499, n_10500, n_10501, n_10502, n_10503, n_10504, n_10505, n_10506, n_10507, n_10508, n_10509, n_10510, n_10511, n_10512, n_10513, n_10514, n_10515, n_10516, n_10517, n_10518, n_10519, n_10520, n_10521, n_10522, n_10523, n_10524, n_10525, n_10526, n_10527, n_10528, n_10529, n_10530, n_10531, n_10532, n_10533, n_10534, n_10535, n_10536, n_10537, n_10538, n_10539, n_10540, n_10541, n_10542, n_10543, n_10544, n_10545, n_10546, n_10547, n_10548, n_10549, n_10550, n_10551, n_10552, n_10553, n_10554, n_10555, n_10556, n_10557, n_10558, n_10559, n_10560, n_10561, n_10562, n_10563, n_10564, n_10565, n_10566, n_10567, n_10568, n_10569, n_10570, n_10571, n_10572, n_10573, n_10574, n_10575, n_10576, n_10577, n_10578, n_10579, n_10580, n_10581, n_10582, n_10583, n_10584, n_10585, n_10586, n_10587, n_10588, n_10589, n_10590, n_10591, n_10592, n_10593, n_10594, n_10595, n_10596, n_10597, n_10598, n_10599, n_10600, n_10601, n_10602, n_10603, n_10604, n_10605, n_10606, n_10607, n_10608, n_10609, n_10610, n_10611, n_10612, n_10613, n_10614, n_10615, n_10616, n_10617, n_10618, n_10619, n_10620, n_10621, n_10622, n_10623, n_10624, n_10625, n_10626, n_10627, n_10628, n_10629, n_10630, n_10631, n_10632, n_10633, n_10634, n_10635, n_10636, n_10637, n_10638, n_10639, n_10640, n_10641, n_10642, n_10643, n_10644, n_10645, n_10646, n_10647, n_10648, n_10649, n_10650, n_10651, n_10652, n_10653, n_10654, n_10655, n_10656, n_10657, n_10658, n_10659, n_10660, n_10661, n_10662, n_10663, n_10664, n_10665, n_10666, n_10667, n_10668, n_10669, n_10670, n_10671, n_10672, n_10673, n_10674, n_10675, n_10676, n_10677, n_10678, n_10679, n_10680, n_10681, n_10682, n_10683, n_10684, n_10685, n_10686, n_10687, n_10688, n_10689, n_10690, n_10691, n_10692, n_10693, n_10694, n_10695, n_10696, n_10697, n_10698, n_10699, n_10700, n_10701, n_10702, n_10703, n_10704, n_10705, n_10706, n_10707, n_10708, n_10709, n_10710, n_10711, n_10712, n_10713, n_10714, n_10715, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721, n_10722, n_10723, n_10724, n_10725, n_10726, n_10727, n_10728, n_10729, n_10730, n_10731, n_10732, n_10733, n_10734, n_10735, n_10736, n_10737, n_10738, n_10739, n_10740, n_10741, n_10742, n_10743, n_10744, n_10745, n_10746, n_10747, n_10748, n_10749, n_10750, n_10751, n_10752, n_10753, n_10754, n_10755, n_10756, n_10757, n_10758, n_10759, n_10760, n_10761, n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768, n_10769, n_10770, n_10771, n_10772, n_10773, n_10774, n_10775, n_10776, n_10777, n_10778, n_10779, n_10780, n_10781, n_10782, n_10783, n_10784, n_10785, n_10786, n_10787, n_10788, n_10789, n_10790, n_10791, n_10792, n_10793, n_10794, n_10795, n_10796, n_10797, n_10798, n_10799, n_10800, n_10801, n_10802, n_10803, n_10804, n_10805, n_10806, n_10807, n_10808, n_10809, n_10810, n_10811, n_10812, n_10813, n_10814, n_10815, n_10816, n_10817, n_10818, n_10819, n_10820, n_10821, n_10822, n_10823, n_10824, n_10825, n_10826, n_10827, n_10828, n_10829, n_10830, n_10831, n_10832, n_10833, n_10834, n_10835, n_10836, n_10837, n_10838, n_10839, n_10840, n_10841, n_10842, n_10843, n_10844, n_10845, n_10846, n_10847, n_10848, n_10849, n_10850, n_10851, n_10852, n_10853, n_10854, n_10855, n_10856, n_10857, n_10858, n_10859, n_10860, n_10861, n_10862, n_10863, n_10864, n_10865, n_10866, n_10867, n_10868, n_10869, n_10870, n_10871, n_10872, n_10873, n_10874, n_10875, n_10876, n_10877, n_10878, n_10879, n_10880, n_10881, n_10882, n_10883, n_10884, n_10885, n_10886, n_10887, n_10888, n_10889, n_10890, n_10891, n_10892, n_10893, n_10894, n_10895, n_10896, n_10897, n_10898, n_10899, n_10900, n_10901, n_10902, n_10903, n_10904, n_10905, n_10906, n_10907, n_10908, n_10909, n_10910, n_10911, n_10912, n_10913, n_10914, n_10915, n_10916, n_10917, n_10918, n_10919, n_10920, n_10921, n_10922, n_10923, n_10924, n_10925, n_10926, n_10927, n_10928, n_10929, n_10930, n_10931, n_10932, n_10933, n_10934, n_10935, n_10936, n_10937, n_10938, n_10939, n_10940, n_10941, n_10942, n_10943, n_10944, n_10945, n_10946, n_10947, n_10948, n_10949, n_10950, n_10951, n_10952, n_10953, n_10954, n_10955, n_10956, n_10957, n_10958, n_10959, n_10960, n_10961, n_10962, n_10963, n_10964, n_10965, n_10966, n_10967, n_10968, n_10969, n_10970, n_10971, n_10972, n_10973, n_10974, n_10975, n_10976, n_10977, n_10978, n_10979, n_10980, n_10981, n_10982, n_10983, n_10984, n_10985, n_10986, n_10987, n_10988, n_10989, n_10990, n_10991, n_10992, n_10993, n_10994, n_10995, n_10996, n_10997, n_10998, n_10999, n_11000, n_11001, n_11002, n_11003, n_11004, n_11005, n_11006, n_11007, n_11008, n_11009, n_11010, n_11011, n_11012, n_11013, n_11014, n_11015, n_11016, n_11017, n_11018, n_11019, n_11020, n_11021, n_11022, n_11023, n_11024, n_11025, n_11026, n_11027, n_11028, n_11029, n_11030, n_11031, n_11032, n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, n_11039, n_11040, n_11041, n_11042, n_11043, n_11044, n_11045, n_11046, n_11047, n_11048, n_11049, n_11050, n_11051, n_11052, n_11053, n_11054, n_11055, n_11056, n_11057, n_11058, n_11059, n_11060, n_11061, n_11062, n_11063, n_11064, n_11065, n_11066, n_11067, n_11068, n_11069, n_11070, n_11071, n_11072, n_11073, n_11074, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080, n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087, n_11088, n_11089, n_11090, n_11091, n_11092, n_11093, n_11094, n_11095, n_11096, n_11097, n_11098, n_11099, n_11100, n_11101, n_11102, n_11103, n_11104, n_11105, n_11106, n_11107, n_11108, n_11109, n_11110, n_11111, n_11112, n_11113, n_11114, n_11115, n_11116, n_11117, n_11118, n_11119, n_11120, n_11121, n_11122, n_11123, n_11124, n_11125, n_11126, n_11127, n_11128, n_11129, n_11130, n_11131, n_11132, n_11133, n_11134, n_11135, n_11136, n_11137, n_11138, n_11139, n_11140, n_11141, n_11142, n_11143, n_11144, n_11145, n_11146, n_11147, n_11148, n_11149, n_11150, n_11151, n_11152, n_11153, n_11154, n_11155, n_11156, n_11157, n_11158, n_11159, n_11160, n_11161, n_11162, n_11163, n_11164, n_11165, n_11166, n_11167, n_11168, n_11169, n_11170, n_11171, n_11172, n_11173, n_11174, n_11175, n_11176, n_11177, n_11178, n_11179, n_11180, n_11181, n_11182, n_11183, n_11184, n_11185, n_11186, n_11187, n_11188, n_11189, n_11190, n_11191, n_11192, n_11193, n_11194, n_11195, n_11196, n_11197, n_11198, n_11199, n_11200, n_11201, n_11202, n_11203, n_11204, n_11205, n_11206, n_11207, n_11208, n_11209, n_11210, n_11211, n_11212, n_11213, n_11214, n_11215, n_11216, n_11217, n_11218, n_11219, n_11220, n_11221, n_11222, n_11223, n_11224, n_11225, n_11226, n_11227, n_11228, n_11229, n_11230, n_11231, n_11232, n_11233, n_11234, n_11235, n_11236, n_11237, n_11238, n_11239, n_11240, n_11241, n_11242, n_11243, n_11244, n_11245, n_11246, n_11247, n_11248, n_11249, n_11250, n_11251, n_11252, n_11253, n_11254, n_11255, n_11256, n_11257, n_11258, n_11259, n_11260, n_11261, n_11262, n_11263, n_11264, n_11265, n_11266, n_11267, n_11268, n_11269, n_11270, n_11271, n_11272, n_11273, n_11274, n_11275, n_11276, n_11277, n_11278, n_11279, n_11280, n_11281, n_11282, n_11283, n_11284, n_11285, n_11286, n_11287, n_11288, n_11289, n_11290, n_11291, n_11292, n_11293, n_11294, n_11295, n_11296, n_11297, n_11298, n_11299, n_11300, n_11301, n_11302, n_11303, n_11304, n_11305, n_11306, n_11307, n_11308, n_11309, n_11310, n_11311, n_11312, n_11313, n_11314, n_11315, n_11316, n_11317, n_11318, n_11319, n_11320, n_11321, n_11322, n_11323, n_11324, n_11325, n_11326, n_11327, n_11328, n_11329, n_11330, n_11331, n_11332, n_11333, n_11334, n_11335, n_11336, n_11337, n_11338, n_11339, n_11340, n_11341, n_11342, n_11343, n_11344, n_11345, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351, n_11352, n_11353, n_11354, n_11355, n_11356, n_11357, n_11358, n_11359, n_11360, n_11361, n_11362, n_11363, n_11364, n_11365, n_11366, n_11367, n_11368, n_11369, n_11370, n_11371, n_11372, n_11373, n_11374, n_11375, n_11376, n_11377, n_11378, n_11379, n_11380, n_11381, n_11382, n_11383, n_11384, n_11385, n_11386, n_11387, n_11388, n_11389, n_11390, n_11391, n_11392, n_11393, n_11394, n_11395, n_11396, n_11397, n_11398, n_11399, n_11400, n_11401, n_11402, n_11403, n_11404, n_11405, n_11406, n_11407, n_11408, n_11409, n_11410, n_11411, n_11412, n_11413, n_11414, n_11415, n_11416, n_11417, n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424, n_11425, n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432, n_11433, n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440, n_11441, n_11442, n_11443, n_11444, n_11445, n_11446, n_11447, n_11448, n_11449, n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11456, n_11457, n_11458, n_11459, n_11460, n_11461, n_11462, n_11463, n_11464, n_11465, n_11466, n_11467, n_11468, n_11469, n_11470, n_11471, n_11472, n_11473, n_11474, n_11475, n_11476, n_11477, n_11478, n_11479, n_11480, n_11481, n_11482, n_11483, n_11484, n_11485, n_11486, n_11487, n_11488, n_11489, n_11490, n_11491, n_11492, n_11493, n_11494, n_11495, n_11496, n_11497, n_11498, n_11499, n_11500, n_11501, n_11502, n_11503, n_11504, n_11505, n_11506, n_11507, n_11508, n_11509, n_11510, n_11511, n_11512, n_11513, n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520, n_11521, n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528, n_11529, n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536, n_11537, n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544, n_11545, n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552, n_11553, n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560, n_11561, n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568, n_11569, n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576, n_11577, n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584, n_11585, n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592, n_11593, n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600, n_11601, n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11608, n_11609, n_11610, n_11611, n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618, n_11619, n_11620, n_11621, n_11622, n_11623, n_11624, n_11625, n_11626, n_11627, n_11628, n_11629, n_11630, n_11631, n_11632, n_11633, n_11634, n_11635, n_11636, n_11637, n_11638, n_11639, n_11640, n_11641, n_11642, n_11643, n_11644, n_11645, n_11646, n_11647, n_11648, n_11649, n_11650, n_11651, n_11652, n_11653, n_11654, n_11655, n_11656, n_11657, n_11658, n_11659, n_11660, n_11661, n_11662, n_11663, n_11664, n_11665, n_11666, n_11667, n_11668, n_11669, n_11670, n_11671, n_11672, n_11673, n_11674, n_11675, n_11676, n_11677, n_11678, n_11679, n_11680, n_11681, n_11682, n_11683, n_11684, n_11685, n_11686, n_11687, n_11688, n_11689, n_11690, n_11691, n_11692, n_11693, n_11694, n_11695, n_11696, n_11697, n_11698, n_11699, n_11700, n_11701, n_11702, n_11703, n_11704, n_11705, n_11706, n_11707, n_11708, n_11709, n_11710, n_11711, n_11712, n_11713, n_11714, n_11715, n_11716, n_11717, n_11718, n_11719, n_11720, n_11721, n_11722, n_11723, n_11724, n_11725, n_11726, n_11727, n_11728, n_11729, n_11730, n_11731, n_11732, n_11733, n_11734, n_11735, n_11736, n_11737, n_11738, n_11739, n_11740, n_11741, n_11742, n_11743, n_11744, n_11745, n_11746, n_11747, n_11748, n_11749, n_11750, n_11751, n_11752, n_11753, n_11754, n_11755, n_11756, n_11757, n_11758, n_11759, n_11760, n_11761, n_11762, n_11763, n_11764, n_11765, n_11766, n_11767, n_11768, n_11769, n_11770, n_11771, n_11772, n_11773, n_11774, n_11775, n_11776, n_11777, n_11778, n_11779, n_11780, n_11781, n_11782, n_11783, n_11784, n_11785, n_11786, n_11787, n_11788, n_11789, n_11790, n_11791, n_11792, n_11793, n_11794, n_11795, n_11796, n_11797, n_11798, n_11799, n_11800, n_11801, n_11802, n_11803, n_11804, n_11805, n_11806, n_11807, n_11808, n_11809, n_11810, n_11811, n_11812, n_11813, n_11814, n_11815, n_11816, n_11817, n_11818, n_11819, n_11820, n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827, n_11828, n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835, n_11836, n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843, n_11844, n_11845, n_11846, n_11847, n_11848, n_11849, n_11850, n_11851, n_11852, n_11853, n_11854, n_11855, n_11856, n_11857, n_11858, n_11859, n_11860, n_11861, n_11862, n_11863, n_11864, n_11865, n_11866, n_11867, n_11868, n_11869, n_11870, n_11871, n_11872, n_11873, n_11874, n_11875, n_11876, n_11877, n_11878, n_11879, n_11880, n_11881, n_11882, n_11883, n_11884, n_11885, n_11886, n_11887, n_11888, n_11889, n_11890, n_11891, n_11892, n_11893, n_11894, n_11895, n_11896, n_11897, n_11898, n_11899, n_11900, n_11901, n_11902, n_11903, n_11904, n_11905, n_11906, n_11907, n_11908, n_11909, n_11910, n_11911, n_11912, n_11913, n_11914, n_11915, n_11916, n_11917, n_11918, n_11919, n_11920, n_11921, n_11922, n_11923, n_11924, n_11925, n_11926, n_11927, n_11928, n_11929, n_11930, n_11931, n_11932, n_11933, n_11934, n_11935, n_11936, n_11937, n_11938, n_11939, n_11940, n_11941, n_11942, n_11943, n_11944, n_11945, n_11946, n_11947, n_11948, n_11949, n_11950, n_11951, n_11952, n_11953, n_11954, n_11955, n_11956, n_11957, n_11958, n_11959, n_11960, n_11961, n_11962, n_11963, n_11964, n_11965, n_11966, n_11967, n_11968, n_11969, n_11970, n_11971, n_11972, n_11973, n_11974, n_11975, n_11976, n_11977, n_11978, n_11979, n_11980, n_11981, n_11982, n_11983, n_11984, n_11985, n_11986, n_11987, n_11988, n_11989, n_11990, n_11991, n_11992, n_11993, n_11994, n_11995, n_11996, n_11997, n_11998, n_11999, n_12000, n_12001, n_12002, n_12003, n_12004, n_12005, n_12006, n_12007, n_12008, n_12009, n_12010, n_12011, n_12012, n_12013, n_12014, n_12015, n_12016, n_12017, n_12018, n_12019, n_12020, n_12021, n_12022, n_12023, n_12024, n_12025, n_12026, n_12027, n_12028, n_12029, n_12030, n_12031, n_12032, n_12033, n_12034, n_12035, n_12036, n_12037, n_12038, n_12039, n_12040, n_12041, n_12042, n_12043, n_12044, n_12045, n_12046, n_12047, n_12048, n_12049, n_12050, n_12051, n_12052, n_12053, n_12054, n_12055, n_12056, n_12057, n_12058, n_12059, n_12060, n_12061, n_12062, n_12063, n_12064, n_12065, n_12066, n_12067, n_12068, n_12069, n_12070, n_12071, n_12072, n_12073, n_12074, n_12075, n_12076, n_12077, n_12078, n_12079, n_12080, n_12081, n_12082, n_12083, n_12084, n_12085, n_12086, n_12087, n_12088, n_12089, n_12090, n_12091, n_12092, n_12093, n_12094, n_12095, n_12096, n_12097, n_12098, n_12099, n_12100, n_12101, n_12102, n_12103, n_12104, n_12105, n_12106, n_12107, n_12108, n_12109, n_12110, n_12111, n_12112, n_12113, n_12114, n_12115, n_12116, n_12117, n_12118, n_12119, n_12120, n_12121, n_12122, n_12123, n_12124, n_12125, n_12126, n_12127, n_12128, n_12129, n_12130, n_12131, n_12132, n_12133, n_12134, n_12135, n_12136, n_12137, n_12138, n_12139, n_12140, n_12141, n_12142, n_12143, n_12144, n_12145, n_12146, n_12147, n_12148, n_12149, n_12150, n_12151, n_12152, n_12153, n_12154, n_12155, n_12156, n_12157, n_12158, n_12159, n_12160, n_12161, n_12162, n_12163, n_12164, n_12165, n_12166, n_12167, n_12168, n_12169, n_12170, n_12171, n_12172, n_12173, n_12174, n_12175, n_12176, n_12177, n_12178, n_12179, n_12180, n_12181, n_12182, n_12183, n_12184, n_12185, n_12186, n_12187, n_12188, n_12189, n_12190, n_12191, n_12192, n_12193, n_12194, n_12195, n_12196, n_12197, n_12198, n_12199, n_12200, n_12201, n_12202, n_12203, n_12204, n_12205, n_12206, n_12207, n_12208, n_12209, n_12210, n_12211, n_12212, n_12213, n_12214, n_12215, n_12216, n_12217, n_12218, n_12219, n_12220, n_12221, n_12222, n_12223, n_12224, n_12225, n_12226, n_12227, n_12228, n_12229, n_12230, n_12231, n_12232, n_12233, n_12234, n_12235, n_12236, n_12237, n_12238, n_12239, n_12240, n_12241, n_12242, n_12243, n_12244, n_12245, n_12246, n_12247, n_12248, n_12249, n_12250, n_12251, n_12252, n_12253, n_12254, n_12255, n_12256, n_12257, n_12258, n_12259, n_12260, n_12261, n_12262, n_12263, n_12264, n_12265, n_12266, n_12267, n_12268, n_12269, n_12270, n_12271, n_12272, n_12273, n_12274, n_12275, n_12276, n_12277, n_12278, n_12279, n_12280, n_12281, n_12282, n_12283, n_12284, n_12285, n_12286, n_12287, n_12288, n_12289, n_12290, n_12291, n_12292, n_12293, n_12294, n_12295, n_12296, n_12297, n_12298, n_12299, n_12300, n_12301, n_12302, n_12303, n_12304, n_12305, n_12306, n_12307, n_12308, n_12309, n_12310, n_12311, n_12312, n_12313, n_12314, n_12315, n_12316, n_12317, n_12318, n_12319, n_12320, n_12321, n_12322, n_12323, n_12324, n_12325, n_12326, n_12327, n_12328, n_12329, n_12330, n_12331, n_12332, n_12333, n_12334, n_12335, n_12336, n_12337, n_12338, n_12339, n_12340, n_12341, n_12342, n_12343, n_12344, n_12345, n_12346, n_12347, n_12348, n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355, n_12356, n_12357, n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364, n_12365, n_12366, n_12367, n_12368, n_12369, n_12370, n_12371, n_12372, n_12373, n_12374, n_12375, n_12376, n_12377, n_12378, n_12379, n_12380, n_12381, n_12382, n_12383, n_12384, n_12385, n_12386, n_12387, n_12388, n_12389, n_12390, n_12391, n_12392, n_12393, n_12394, n_12395, n_12396, n_12397, n_12398, n_12399, n_12400, n_12401, n_12402, n_12403, n_12404, n_12405, n_12406, n_12407, n_12408, n_12409, n_12410, n_12411, n_12412, n_12413, n_12414, n_12415, n_12416, n_12417, n_12418, n_12419, n_12420, n_12421, n_12422, n_12423, n_12424, n_12425, n_12426, n_12427, n_12428, n_12429, n_12430, n_12431, n_12432, n_12433, n_12434, n_12435, n_12436, n_12437, n_12438, n_12439, n_12440, n_12441, n_12442, n_12443, n_12444, n_12445, n_12446, n_12447, n_12448, n_12449, n_12450, n_12451, n_12452, n_12453, n_12454, n_12455, n_12456, n_12457, n_12458, n_12459, n_12460, n_12461, n_12462, n_12463, n_12464, n_12465, n_12466, n_12467, n_12468, n_12469, n_12470, n_12471, n_12472, n_12473, n_12474, n_12475, n_12476, n_12477, n_12478, n_12479, n_12480, n_12481, n_12482, n_12483, n_12484, n_12485, n_12486, n_12487, n_12488, n_12489, n_12490, n_12491, n_12492, n_12493, n_12494, n_12495, n_12496, n_12497, n_12498, n_12499, n_12500, n_12501, n_12502, n_12503, n_12504, n_12505, n_12506, n_12507, n_12508, n_12509, n_12510, n_12511, n_12512, n_12513, n_12514, n_12515, n_12516, n_12517, n_12518, n_12519, n_12520, n_12521, n_12522, n_12523, n_12524, n_12525, n_12526, n_12527, n_12528, n_12529, n_12530, n_12531, n_12532, n_12533, n_12534, n_12535, n_12536, n_12537, n_12538, n_12539, n_12540, n_12541, n_12542, n_12543, n_12544, n_12545, n_12546, n_12547, n_12548, n_12549, n_12550, n_12551, n_12552, n_12553, n_12554, n_12555, n_12556, n_12557, n_12558, n_12559, n_12560, n_12561, n_12562, n_12563, n_12564, n_12565, n_12566, n_12567, n_12568, n_12569, n_12570, n_12571, n_12572, n_12573, n_12574, n_12575, n_12576, n_12577, n_12578, n_12579, n_12580, n_12581, n_12582, n_12583, n_12584, n_12585, n_12586, n_12587, n_12588, n_12589, n_12590, n_12591, n_12592, n_12593, n_12594, n_12595, n_12596, n_12597, n_12598, n_12599, n_12600, n_12601, n_12602, n_12603, n_12604, n_12605, n_12606, n_12607, n_12608, n_12609, n_12610, n_12611, n_12612, n_12613, n_12614, n_12615, n_12616, n_12617, n_12618, n_12619, n_12620, n_12621, n_12622, n_12623, n_12624, n_12625, n_12626, n_12627, n_12628, n_12629, n_12630, n_12631, n_12632, n_12633, n_12634, n_12635, n_12636, n_12637, n_12638, n_12639, n_12640, n_12641, n_12642, n_12643, n_12644, n_12645, n_12646, n_12647, n_12648, n_12649, n_12650, n_12651, n_12652, n_12653, n_12654, n_12655, n_12656, n_12657, n_12658, n_12659, n_12660, n_12661, n_12662, n_12663, n_12664, n_12665, n_12666, n_12667, n_12668, n_12669, n_12670, n_12671, n_12672, n_12673, n_12674, n_12675, n_12676, n_12677, n_12678, n_12679, n_12680, n_12681, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687, n_12688, n_12689, n_12690, n_12691, n_12692, n_12693, n_12694, n_12695, n_12696, n_12697, n_12698, n_12699, n_12700, n_12701, n_12702, n_12703, n_12704, n_12705, n_12706, n_12707, n_12708, n_12709, n_12710, n_12711, n_12712, n_12713, n_12714, n_12715, n_12716, n_12717, n_12718, n_12719, n_12720, n_12721, n_12722, n_12723, n_12724, n_12725, n_12726, n_12727, n_12728, n_12729, n_12730, n_12731, n_12732, n_12733, n_12734, n_12735, n_12736, n_12737, n_12738, n_12739, n_12740, n_12741, n_12742, n_12743, n_12744, n_12745, n_12746, n_12747, n_12748, n_12749, n_12750, n_12751, n_12752, n_12753, n_12754, n_12755, n_12756, n_12757, n_12758, n_12759, n_12760, n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767, n_12768, n_12769, n_12770, n_12771, n_12772, n_12773, n_12774, n_12775, n_12776, n_12777, n_12778, n_12779, n_12780, n_12781, n_12782, n_12783, n_12784, n_12785, n_12786, n_12787, n_12788, n_12789, n_12790, n_12791, n_12792, n_12793, n_12794, n_12795, n_12796, n_12797, n_12798, n_12799, n_12800, n_12801, n_12802, n_12803, n_12804, n_12805, n_12806, n_12807, n_12808, n_12809, n_12810, n_12811, n_12812, n_12813, n_12814, n_12815, n_12816, n_12817, n_12818, n_12819, n_12820, n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827, n_12828, n_12829, n_12830, n_12831, n_12832, n_12833, n_12834, n_12835, n_12836, n_12837, n_12838, n_12839, n_12840, n_12841, n_12842, n_12843, n_12844, n_12845, n_12846, n_12847, n_12848, n_12849, n_12850, n_12851, n_12852, n_12853, n_12854, n_12855, n_12856, n_12857, n_12858, n_12859, n_12860, n_12861, n_12862, n_12863, n_12864, n_12865, n_12866, n_12867, n_12868, n_12869, n_12870, n_12871, n_12872, n_12873, n_12874, n_12875, n_12876, n_12877, n_12878, n_12879, n_12880, n_12881, n_12882, n_12883, n_12884, n_12885, n_12886, n_12887, n_12888, n_12889, n_12890, n_12891, n_12892, n_12893, n_12894, n_12895, n_12896, n_12897, n_12898, n_12899, n_12900, n_12901, n_12902, n_12903, n_12904, n_12905, n_12906, n_12907, n_12908, n_12909, n_12910, n_12911, n_12912, n_12913, n_12914, n_12915, n_12916, n_12917, n_12918, n_12919, n_12920, n_12921, n_12922, n_12923, n_12924, n_12925, n_12926, n_12927, n_12928, n_12929, n_12930, n_12931, n_12932, n_12933, n_12934, n_12935, n_12936, n_12937, n_12938, n_12939, n_12940, n_12941, n_12942, n_12943, n_12944, n_12945, n_12946, n_12947, n_12948, n_12949, n_12950, n_12951, n_12952, n_12953, n_12954, n_12955, n_12956, n_12957, n_12958, n_12959, n_12960, n_12961, n_12962, n_12963, n_12964, n_12965, n_12966, n_12967, n_12968, n_12969, n_12970, n_12971, n_12972, n_12973, n_12974, n_12975, n_12976, n_12977, n_12978, n_12979, n_12980, n_12981, n_12982, n_12983, n_12984, n_12985, n_12986, n_12987, n_12988, n_12989, n_12990, n_12991, n_12992, n_12993, n_12994, n_12995, n_12996, n_12997, n_12998, n_12999, n_13000, n_13001, n_13002, n_13003, n_13004, n_13005, n_13006, n_13007, n_13008, n_13009, n_13010, n_13011, n_13012, n_13013, n_13014, n_13015, n_13016, n_13017, n_13018, n_13019, n_13020, n_13021, n_13022, n_13023, n_13024, n_13025, n_13026, n_13027, n_13028, n_13029, n_13030, n_13031, n_13032, n_13033, n_13034, n_13035, n_13036, n_13037, n_13038, n_13039, n_13040, n_13041, n_13042, n_13043, n_13044, n_13045, n_13046, n_13047, n_13048, n_13049, n_13050, n_13051, n_13052, n_13053, n_13054, n_13055, n_13056, n_13057, n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064, n_13065, n_13066, n_13067, n_13068, n_13069, n_13070, n_13071, n_13072, n_13073, n_13074, n_13075, n_13076, n_13077, n_13078, n_13079, n_13080, n_13081, n_13082, n_13083, n_13084, n_13085, n_13086, n_13087, n_13088, n_13089, n_13090, n_13091, n_13092, n_13093, n_13094, n_13095, n_13096, n_13097, n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104, n_13105, n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13112, n_13113, n_13114, n_13115, n_13116, n_13117, n_13118, n_13119, n_13120, n_13121, n_13122, n_13123, n_13124, n_13125, n_13126, n_13127, n_13128, n_13129, n_13130, n_13131, n_13132, n_13133, n_13134, n_13135, n_13136, n_13137, n_13138, n_13139, n_13140, n_13141, n_13142, n_13143, n_13144, n_13145, n_13146, n_13147, n_13148, n_13149, n_13150, n_13151, n_13152, n_13153, n_13154, n_13155, n_13156, n_13157, n_13158, n_13159, n_13160, n_13161, n_13162, n_13163, n_13164, n_13165, n_13166, n_13167, n_13168, n_13169, n_13170, n_13171, n_13172, n_13173, n_13174, n_13175, n_13176, n_13177, n_13178, n_13179, n_13180, n_13181, n_13182, n_13183, n_13184, n_13185, n_13186, n_13187, n_13188, n_13189, n_13190, n_13191, n_13192, n_13193, n_13194, n_13195, n_13196, n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203, n_13204, n_13205, n_13206, n_13207, n_13208, n_13209, n_13210, n_13211, n_13212, n_13213, n_13214, n_13215, n_13216, n_13217, n_13218, n_13219, n_13220, n_13221, n_13222, n_13223, n_13224, n_13225, n_13226, n_13227, n_13228, n_13229, n_13230, n_13231, n_13232, n_13233, n_13234, n_13235, n_13236, n_13237, n_13238, n_13239, n_13240, n_13241, n_13242, n_13243, n_13244, n_13245, n_13246, n_13247, n_13248, n_13249, n_13250, n_13251, n_13252, n_13253, n_13254, n_13255, n_13256, n_13257, n_13258, n_13259, n_13260, n_13261, n_13262, n_13263, n_13264, n_13265, n_13266, n_13267, n_13268, n_13269, n_13270, n_13271, n_13272, n_13273, n_13274, n_13275, n_13276, n_13277, n_13278, n_13279, n_13280, n_13281, n_13282, n_13283, n_13284, n_13285, n_13286, n_13287, n_13288, n_13289, n_13290, n_13291, n_13292, n_13293, n_13294, n_13295, n_13296, n_13297, n_13298, n_13299, n_13300, n_13301, n_13302, n_13303, n_13304, n_13305, n_13306, n_13307, n_13308, n_13309, n_13310, n_13311, n_13312, n_13313, n_13314, n_13315, n_13316, n_13317, n_13318, n_13319, n_13320, n_13321, n_13322, n_13323, n_13324, n_13325, n_13326, n_13327, n_13328, n_13329, n_13330, n_13331, n_13332, n_13333, n_13334, n_13335, n_13336, n_13337, n_13338, n_13339, n_13340, n_13341, n_13342, n_13343, n_13344, n_13345, n_13346, n_13347, n_13348, n_13349, n_13350, n_13351, n_13352, n_13353, n_13354, n_13355, n_13356, n_13357, n_13358, n_13359, n_13360, n_13361, n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368, n_13369, n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376, n_13377, n_13378, n_13379, n_13380, n_13381, n_13382, n_13383, n_13384, n_13385, n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392, n_13393, n_13394, n_13395, n_13396, n_13397, n_13398, n_13399, n_13400, n_13401, n_13402, n_13403, n_13404, n_13405, n_13406, n_13407, n_13408, n_13409, n_13410, n_13411, n_13412, n_13413, n_13414, n_13415, n_13416, n_13417, n_13418, n_13419, n_13420, n_13421, n_13422, n_13423, n_13424, n_13425, n_13426, n_13427, n_13428, n_13429, n_13430, n_13431, n_13432, n_13433, n_13434, n_13435, n_13436, n_13437, n_13438, n_13439, n_13440, n_13441, n_13442, n_13443, n_13444, n_13445, n_13446, n_13447, n_13448, n_13449, n_13450, n_13451, n_13452, n_13453, n_13454, n_13455, n_13456, n_13457, n_13458, n_13459, n_13460, n_13461, n_13462, n_13463, n_13464, n_13465, n_13466, n_13467, n_13468, n_13469, n_13470, n_13471, n_13472, n_13473, n_13474, n_13475, n_13476, n_13477, n_13478, n_13479, n_13480, n_13481, n_13482, n_13483, n_13484, n_13485, n_13486, n_13487, n_13488, n_13489, n_13490, n_13491, n_13492, n_13493, n_13494, n_13495, n_13496, n_13497, n_13498, n_13499, n_13500, n_13501, n_13502, n_13503, n_13504, n_13505, n_13506, n_13507, n_13508, n_13509, n_13510, n_13511, n_13512, n_13513, n_13514, n_13515, n_13516, n_13517, n_13518, n_13519, n_13520, n_13521, n_13522, n_13523, n_13524, n_13525, n_13526, n_13527, n_13528, n_13529, n_13530, n_13531, n_13532, n_13533, n_13534, n_13535, n_13536, n_13537, n_13538, n_13539, n_13540, n_13541, n_13542, n_13543, n_13544, n_13545, n_13546, n_13547, n_13548, n_13549, n_13550, n_13551, n_13552, n_13553, n_13554, n_13555, n_13556, n_13557, n_13558, n_13559, n_13560, n_13561, n_13562, n_13563, n_13564, n_13565, n_13566, n_13567, n_13568, n_13569, n_13570, n_13571, n_13572, n_13573, n_13574, n_13575, n_13576, n_13577, n_13578, n_13579, n_13580, n_13581, n_13582, n_13583, n_13584, n_13585, n_13586, n_13587, n_13588, n_13589, n_13590, n_13591, n_13592, n_13593, n_13594, n_13595, n_13596, n_13597, n_13598, n_13599, n_13600, n_13601, n_13602, n_13603, n_13604, n_13605, n_13606, n_13607, n_13608, n_13609, n_13610, n_13611, n_13612, n_13613, n_13614, n_13615, n_13616, n_13617, n_13618, n_13619, n_13620, n_13621, n_13622, n_13623, n_13624, n_13625, n_13626, n_13627, n_13628, n_13629, n_13630, n_13631, n_13632, n_13633, n_13634, n_13635, n_13636, n_13637, n_13638, n_13639, n_13640, n_13641, n_13642, n_13643, n_13644, n_13645, n_13646, n_13647, n_13648, n_13649, n_13650, n_13651, n_13652, n_13653, n_13654, n_13655, n_13656, n_13657, n_13658, n_13659, n_13660, n_13661, n_13662, n_13663, n_13664, n_13665, n_13666, n_13667, n_13668, n_13669, n_13670, n_13671, n_13672, n_13673, n_13674, n_13675, n_13676, n_13677, n_13678, n_13679, n_13680, n_13681, n_13682, n_13683, n_13684, n_13685, n_13686, n_13687, n_13688, n_13689, n_13690, n_13691, n_13692, n_13693, n_13694, n_13695, n_13696, n_13697, n_13698, n_13699, n_13700, n_13701, n_13702, n_13703, n_13704, n_13705, n_13706, n_13707, n_13708, n_13709, n_13710, n_13711, n_13712, n_13713, n_13714, n_13715, n_13716, n_13717, n_13718, n_13719, n_13720, n_13721, n_13722, n_13723, n_13724, n_13725, n_13726, n_13727, n_13728, n_13729, n_13730, n_13731, n_13732, n_13733, n_13734, n_13735, n_13736, n_13737, n_13738, n_13739, n_13740, n_13741, n_13742, n_13743, n_13744, n_13745, n_13746, n_13747, n_13748, n_13749, n_13750, n_13751, n_13752, n_13753, n_13754, n_13755, n_13756, n_13757, n_13758, n_13759, n_13760, n_13761, n_13762, n_13763, n_13764, n_13765, n_13766, n_13767, n_13768, n_13769, n_13770, n_13771, n_13772, n_13773, n_13774, n_13775, n_13776, n_13777, n_13778, n_13779, n_13780, n_13781, n_13782, n_13783, n_13784, n_13785, n_13786, n_13787, n_13788, n_13789, n_13790, n_13791, n_13792, n_13793, n_13794, n_13795, n_13796, n_13797, n_13798, n_13799, n_13800, n_13801, n_13802, n_13803, n_13804, n_13805, n_13806, n_13807, n_13808, n_13809, n_13810, n_13811, n_13812, n_13813, n_13814, n_13815, n_13816, n_13817, n_13818, n_13819, n_13820, n_13821, n_13822, n_13823, n_13824, n_13825, n_13826, n_13827, n_13828, n_13829, n_13830, n_13831, n_13832, n_13833, n_13834, n_13835, n_13836, n_13837, n_13838, n_13839, n_13840, n_13841, n_13842, n_13843, n_13844, n_13845, n_13846, n_13847, n_13848, n_13849, n_13850, n_13851, n_13852, n_13853, n_13854, n_13855, n_13856, n_13857, n_13858, n_13859, n_13860, n_13861, n_13862, n_13863, n_13864, n_13865, n_13866, n_13867, n_13868, n_13869, n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13876, n_13877, n_13878, n_13879, n_13880, n_13881, n_13882, n_13883, n_13884, n_13885, n_13886, n_13887, n_13888, n_13889, n_13890, n_13891, n_13892, n_13893, n_13894, n_13895, n_13896, n_13897, n_13898, n_13899, n_13900, n_13901, n_13902, n_13903, n_13904, n_13905, n_13906, n_13907, n_13908, n_13909, n_13910, n_13911, n_13912, n_13913, n_13914, n_13915, n_13916, n_13917, n_13918, n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925, n_13926, n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933, n_13934, n_13935, n_13936, n_13937, n_13938, n_13939, n_13940, n_13941, n_13942, n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949, n_13950, n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957, n_13958, n_13959, n_13960, n_13961, n_13962, n_13963, n_13964, n_13965, n_13966, n_13967, n_13968, n_13969, n_13970, n_13971, n_13972, n_13973, n_13974, n_13975, n_13976, n_13977, n_13978, n_13979, n_13980, n_13981, n_13982, n_13983, n_13984, n_13985, n_13986, n_13987, n_13988, n_13989, n_13990, n_13991, n_13992, n_13993, n_13994, n_13995, n_13996, n_13997, n_13998, n_13999, n_14000, n_14001, n_14002, n_14003, n_14004, n_14005, n_14006, n_14007, n_14008, n_14009, n_14010, n_14011, n_14012, n_14013, n_14014, n_14015, n_14016, n_14017, n_14018, n_14019, n_14020, n_14021, n_14022, n_14023, n_14024, n_14025, n_14026, n_14027, n_14028, n_14029, n_14030, n_14031, n_14032, n_14033, n_14034, n_14035, n_14036, n_14037, n_14038, n_14039, n_14040, n_14041, n_14042, n_14043, n_14044, n_14045, n_14046, n_14047, n_14048, n_14049, n_14050, n_14051, n_14052, n_14053, n_14054, n_14055, n_14056, n_14057, n_14058, n_14059, n_14060, n_14061, n_14062, n_14063, n_14064, n_14065, n_14066, n_14067, n_14068, n_14069, n_14070, n_14071, n_14072, n_14073, n_14074, n_14075, n_14076, n_14077, n_14078, n_14079, n_14080, n_14081, n_14082, n_14083, n_14084, n_14085, n_14086, n_14087, n_14088, n_14089, n_14090, n_14091, n_14092, n_14093, n_14094, n_14095, n_14096, n_14097, n_14098, n_14099, n_14100, n_14101, n_14102, n_14103, n_14104, n_14105, n_14106, n_14107, n_14108, n_14109, n_14110, n_14111, n_14112, n_14113, n_14114, n_14115, n_14116, n_14117, n_14118, n_14119, n_14120, n_14121, n_14122, n_14123, n_14124, n_14125, n_14126, n_14127, n_14128, n_14129, n_14130, n_14131, n_14132, n_14133, n_14134, n_14135, n_14136, n_14137, n_14138, n_14139, n_14140, n_14141, n_14142, n_14143, n_14144, n_14145, n_14146, n_14147, n_14148, n_14149, n_14150, n_14151, n_14152, n_14153, n_14154, n_14155, n_14156, n_14157, n_14158, n_14159, n_14160, n_14161, n_14162, n_14163, n_14164, n_14165, n_14166, n_14167, n_14168, n_14169, n_14170, n_14171, n_14172, n_14173, n_14174, n_14175, n_14176, n_14177, n_14178, n_14179, n_14180, n_14181, n_14182, n_14183, n_14184, n_14185, n_14186, n_14187, n_14188, n_14189, n_14190, n_14191, n_14192, n_14193, n_14194, n_14195, n_14196, n_14197, n_14198, n_14199, n_14200, n_14201, n_14202, n_14203, n_14204, n_14205, n_14206, n_14207, n_14208, n_14209, n_14210, n_14211, n_14212, n_14213, n_14214, n_14215, n_14216, n_14217, n_14218, n_14219, n_14220, n_14221, n_14222, n_14223, n_14224, n_14225, n_14226, n_14227, n_14228, n_14229, n_14230, n_14231, n_14232, n_14233, n_14234, n_14235, n_14236, n_14237, n_14238, n_14239, n_14240, n_14241, n_14242, n_14243, n_14244, n_14245, n_14246, n_14247, n_14248, n_14249, n_14250, n_14251, n_14252, n_14253, n_14254, n_14255, n_14256, n_14257, n_14258, n_14259, n_14260, n_14261, n_14262, n_14263, n_14264, n_14265, n_14266, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272, n_14273, n_14274, n_14275, n_14276, n_14277, n_14278, n_14279, n_14280, n_14281, n_14282, n_14283, n_14284, n_14285, n_14286, n_14287, n_14288, n_14289, n_14290, n_14291, n_14292, n_14293, n_14294, n_14295, n_14296, n_14297, n_14298, n_14299, n_14300, n_14301, n_14302, n_14303, n_14304, n_14305, n_14306, n_14307, n_14308, n_14309, n_14310, n_14311, n_14312, n_14313, n_14314, n_14315, n_14316, n_14317, n_14318, n_14319, n_14320, n_14321, n_14322, n_14323, n_14324, n_14325, n_14326, n_14327, n_14328, n_14329, n_14330, n_14331, n_14332, n_14333, n_14334, n_14335, n_14336, n_14337, n_14338, n_14339, n_14340, n_14341, n_14342, n_14343, n_14344, n_14345, n_14346, n_14347, n_14348, n_14349, n_14350, n_14351, n_14352, n_14353, n_14354, n_14355, n_14356, n_14357, n_14358, n_14359, n_14360, n_14361, n_14362, n_14363, n_14364, n_14365, n_14366, n_14367, n_14368, n_14369, n_14370, n_14371, n_14372, n_14373, n_14374, n_14375, n_14376, n_14377, n_14378, n_14379, n_14380, n_14381, n_14382, n_14383, n_14384, n_14385, n_14386, n_14387, n_14388, n_14389, n_14390, n_14391, n_14392, n_14393, n_14394, n_14395, n_14396, n_14397, n_14398, n_14399, n_14400, n_14401, n_14402, n_14403, n_14404, n_14405, n_14406, n_14407, n_14408, n_14409, n_14410, n_14411, n_14412, n_14413, n_14414, n_14415, n_14416, n_14417, n_14418, n_14419, n_14420, n_14421, n_14422, n_14423, n_14424, n_14425, n_14426, n_14427, n_14428, n_14429, n_14430, n_14431, n_14432, n_14433, n_14434, n_14435, n_14436, n_14437, n_14438, n_14439, n_14440, n_14441, n_14442, n_14443, n_14444, n_14445, n_14446, n_14447, n_14448, n_14449, n_14450, n_14451, n_14452, n_14453, n_14454, n_14455, n_14456, n_14457, n_14458, n_14459, n_14460, n_14461, n_14462, n_14463, n_14464, n_14465, n_14466, n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, n_14473, n_14474, n_14475, n_14476, n_14477, n_14478, n_14479, n_14480, n_14481, n_14482, n_14483, n_14484, n_14485, n_14486, n_14487, n_14488, n_14489, n_14490, n_14491, n_14492, n_14493, n_14494, n_14495, n_14496, n_14497, n_14498, n_14499, n_14500, n_14501, n_14502, n_14503, n_14504, n_14505, n_14506, n_14507, n_14508, n_14509, n_14510, n_14511, n_14512, n_14513, n_14514, n_14515, n_14516, n_14517, n_14518, n_14519, n_14520, n_14521, n_14522, n_14523, n_14524, n_14525, n_14526, n_14527, n_14528, n_14529, n_14530, n_14531, n_14532, n_14533, n_14534, n_14535, n_14536, n_14537, n_14538, n_14539, n_14540, n_14541, n_14542, n_14543, n_14544, n_14545, n_14546, n_14547, n_14548, n_14549, n_14550, n_14551, n_14552, n_14553, n_14554, n_14555, n_14556, n_14557, n_14558, n_14559, n_14560, n_14561, n_14562, n_14563, n_14564, n_14565, n_14566, n_14567, n_14568, n_14569, n_14570, n_14571, n_14572, n_14573, n_14574, n_14575, n_14576, n_14577, n_14578, n_14579, n_14580, n_14581, n_14582, n_14583, n_14584, n_14585, n_14586, n_14587, n_14588, n_14589, n_14590, n_14591, n_14592, n_14593, n_14594, n_14595, n_14596, n_14597, n_14598, n_14599, n_14600, n_14601, n_14602, n_14603, n_14604, n_14605, n_14606, n_14607, n_14608, n_14609, n_14610, n_14611, n_14612, n_14613, n_14614, n_14615, n_14616, n_14617, n_14618, n_14619, n_14620, n_14621, n_14622, n_14623, n_14624, n_14625, n_14626, n_14627, n_14628, n_14629, n_14630, n_14631, n_14632, n_14633, n_14634, n_14635, n_14636, n_14637, n_14638, n_14639, n_14640, n_14641, n_14642, n_14643, n_14644, n_14645, n_14646, n_14647, n_14648, n_14649, n_14650, n_14651, n_14652, n_14653, n_14654, n_14655, n_14656, n_14657, n_14658, n_14659, n_14660, n_14661, n_14662, n_14663, n_14664, n_14665, n_14666, n_14667, n_14668, n_14669, n_14670, n_14671, n_14672, n_14673, n_14674, n_14675, n_14676, n_14677, n_14678, n_14679, n_14680, n_14681, n_14682, n_14683, n_14684, n_14685, n_14686, n_14687, n_14688, n_14689, n_14690, n_14691, n_14692, n_14693, n_14694, n_14695, n_14696, n_14697, n_14698, n_14699, n_14700, n_14701, n_14702, n_14703, n_14704, n_14705, n_14706, n_14707, n_14708, n_14709, n_14710, n_14711, n_14712, n_14713, n_14714, n_14715, n_14716, n_14717, n_14718, n_14719, n_14720, n_14721, n_14722, n_14723, n_14724, n_14725, n_14726, n_14727, n_14728, n_14729, n_14730, n_14731, n_14732, n_14733, n_14734, n_14735, n_14736, n_14737, n_14738, n_14739, n_14740, n_14741, n_14742, n_14743, n_14744, n_14745, n_14746, n_14747, n_14748, n_14749, n_14750, n_14751, n_14752, n_14753, n_14754, n_14755, n_14756, n_14757, n_14758, n_14759, n_14760, n_14761, n_14762, n_14763, n_14764, n_14765, n_14766, n_14767, n_14768, n_14769, n_14770, n_14771, n_14772, n_14773, n_14774, n_14775, n_14776, n_14777, n_14778, n_14779, n_14780, n_14781, n_14782, n_14783, n_14784, n_14785, n_14786, n_14787, n_14788, n_14789, n_14790, n_14791, n_14792, n_14793, n_14794, n_14795, n_14796, n_14797, n_14798, n_14799, n_14800, n_14801, n_14802, n_14803, n_14804, n_14805, n_14806, n_14807, n_14808, n_14809, n_14810, n_14811, n_14812, n_14813, n_14814, n_14815, n_14816, n_14817, n_14818, n_14819, n_14820, n_14821, n_14822, n_14823, n_14824, n_14825, n_14826, n_14827, n_14828, n_14829, n_14830, n_14831, n_14832, n_14833, n_14834, n_14835, n_14836, n_14837, n_14838, n_14839, n_14840, n_14841, n_14842, n_14843, n_14844, n_14845, n_14846, n_14847, n_14848, n_14849, n_14850, n_14851, n_14852, n_14853, n_14854, n_14855, n_14856, n_14857, n_14858, n_14859, n_14860, n_14861, n_14862, n_14863, n_14864, n_14865, n_14866, n_14867, n_14868, n_14869, n_14870, n_14871, n_14872, n_14873, n_14874, n_14875, n_14876, n_14877, n_14878, n_14879, n_14880, n_14881, n_14882, n_14883, n_14884, n_14885, n_14886, n_14887, n_14888, n_14889, n_14890, n_14891, n_14892, n_14893, n_14894, n_14895, n_14896, n_14897, n_14898, n_14899, n_14900, n_14901, n_14902, n_14903, n_14904, n_14905, n_14906, n_14907, n_14908, n_14909, n_14910, n_14911, n_14912, n_14913, n_14914, n_14915, n_14916, n_14917, n_14918, n_14919, n_14920, n_14921, n_14922, n_14923, n_14924, n_14925, n_14926, n_14927, n_14928, n_14929, n_14930, n_14931, n_14932, n_14933, n_14934, n_14935, n_14936, n_14937, n_14938, n_14939, n_14940, n_14941, n_14942, n_14943, n_14944, n_14945, n_14946, n_14947, n_14948, n_14949, n_14950, n_14951, n_14952, n_14953, n_14954, n_14955, n_14956, n_14957, n_14958, n_14959, n_14960, n_14961, n_14962, n_14963, n_14964, n_14965, n_14966, n_14967, n_14968, n_14969, n_14970, n_14971, n_14972, n_14973, n_14974, n_14975, n_14976, n_14977, n_14978, n_14979, n_14980, n_14981, n_14982, n_14983, n_14984, n_14985, n_14986, n_14987, n_14988, n_14989, n_14990, n_14991, n_14992, n_14993, n_14994, n_14995, n_14996, n_14997, n_14998, n_14999, n_15000, n_15001, n_15002, n_15003, n_15004, n_15005, n_15006, n_15007, n_15008, n_15009, n_15010, n_15011, n_15012, n_15013, n_15014, n_15015, n_15016, n_15017, n_15018, n_15019, n_15020, n_15021, n_15022, n_15023, n_15024, n_15025, n_15026, n_15027, n_15028, n_15029, n_15030, n_15031, n_15032, n_15033, n_15034, n_15035, n_15036, n_15037, n_15038, n_15039, n_15040, n_15041, n_15042, n_15043, n_15044, n_15045, n_15046, n_15047, n_15048, n_15049, n_15050, n_15051, n_15052, n_15053, n_15054, n_15055, n_15056, n_15057, n_15058, n_15059, n_15060, n_15061, n_15062, n_15063, n_15064, n_15065, n_15066, n_15067, n_15068, n_15069, n_15070, n_15071, n_15072, n_15073, n_15074, n_15075, n_15076, n_15077, n_15078, n_15079, n_15080, n_15081, n_15082, n_15083, n_15084, n_15085, n_15086, n_15087, n_15088, n_15089, n_15090, n_15091, n_15092, n_15093, n_15094, n_15095, n_15096, n_15097, n_15098, n_15099, n_15100, n_15101, n_15102, n_15103, n_15104, n_15105, n_15106, n_15107, n_15108, n_15109, n_15110, n_15111, n_15112, n_15113, n_15114, n_15115, n_15116, n_15117, n_15118, n_15119, n_15120, n_15121, n_15122, n_15123, n_15124, n_15125, n_15126, n_15127, n_15128, n_15129, n_15130, n_15131, n_15132, n_15133, n_15134, n_15135, n_15136, n_15137, n_15138, n_15139, n_15140, n_15141, n_15142, n_15143, n_15144, n_15145, n_15146, n_15147, n_15148, n_15149, n_15150, n_15151, n_15152, n_15153, n_15154, n_15155, n_15156, n_15157, n_15158, n_15159, n_15160, n_15161, n_15162, n_15163, n_15164, n_15165, n_15166, n_15167, n_15168, n_15169, n_15170, n_15171, n_15172, n_15173, n_15174, n_15175, n_15176, n_15177, n_15178, n_15179, n_15180, n_15181, n_15182, n_15183, n_15184, n_15185, n_15186, n_15187, n_15188, n_15189, n_15190, n_15191, n_15192, n_15193, n_15194, n_15195, n_15196, n_15197, n_15198, n_15199, n_15200, n_15201, n_15202, n_15203, n_15204, n_15205, n_15206, n_15207, n_15208, n_15209, n_15210, n_15211, n_15212, n_15213, n_15214, n_15215, n_15216, n_15217, n_15218, n_15219, n_15220, n_15221, n_15222, n_15223, n_15224, n_15225, n_15226, n_15227, n_15228, n_15229, n_15230, n_15231, n_15232, n_15233, n_15234, n_15235, n_15236, n_15237, n_15238, n_15239, n_15240, n_15241, n_15242, n_15243, n_15244, n_15245, n_15246, n_15247, n_15248, n_15249, n_15250, n_15251, n_15252, n_15253, n_15254, n_15255, n_15256, n_15257, n_15258, n_15259, n_15260, n_15261, n_15262, n_15263, n_15264, n_15265, n_15266, n_15267, n_15268, n_15269, n_15270, n_15271, n_15272, n_15273, n_15274, n_15275, n_15276, n_15277, n_15278, n_15279, n_15280, n_15281, n_15282, n_15283, n_15284, n_15285, n_15286, n_15287, n_15288, n_15289, n_15290, n_15291, n_15292, n_15293, n_15294, n_15295, n_15296, n_15297, n_15298, n_15299, n_15300, n_15301, n_15302, n_15303, n_15304, n_15305, n_15306, n_15307, n_15308, n_15309, n_15310, n_15311, n_15312, n_15313, n_15314, n_15315, n_15316, n_15317, n_15318, n_15319, n_15320, n_15321, n_15322, n_15323, n_15324, n_15325, n_15326, n_15327, n_15328, n_15329, n_15330, n_15331, n_15332, n_15333, n_15334, n_15335, n_15336, n_15337, n_15338, n_15339, n_15340, n_15341, n_15342, n_15343, n_15344, n_15345, n_15346, n_15347, n_15348, n_15349, n_15350, n_15351, n_15352, n_15353, n_15354, n_15355, n_15356, n_15357, n_15358, n_15359, n_15360, n_15361, n_15362, n_15363, n_15364, n_15365, n_15366, n_15367, n_15368, n_15369, n_15370, n_15371, n_15372, n_15373, n_15374, n_15375, n_15376, n_15377, n_15378, n_15379, n_15380, n_15381, n_15382, n_15383, n_15384, n_15385, n_15386, n_15387, n_15388, n_15389, n_15390, n_15391, n_15392, n_15393, n_15394, n_15395, n_15396, n_15397, n_15398, n_15399, n_15400, n_15401, n_15402, n_15403, n_15404, n_15405, n_15406, n_15407, n_15408, n_15409, n_15410, n_15411, n_15412, n_15413, n_15414, n_15415, n_15416, n_15417, n_15418, n_15419, n_15420, n_15421, n_15422, n_15423, n_15424, n_15425, n_15426, n_15427, n_15428, n_15429, n_15430, n_15431, n_15432, n_15433, n_15434, n_15435, n_15436, n_15437, n_15438, n_15439, n_15440, n_15441, n_15442, n_15443, n_15444, n_15445, n_15446, n_15447, n_15448, n_15449, n_15450, n_15451, n_15452, n_15453, n_15454, n_15455, n_15456, n_15457, n_15458, n_15459, n_15460, n_15461, n_15462, n_15463, n_15464, n_15465, n_15466, n_15467, n_15468, n_15469, n_15470, n_15471, n_15472, n_15473, n_15474, n_15475, n_15476, n_15477, n_15478, n_15479, n_15480, n_15481, n_15482, n_15483, n_15484, n_15485, n_15486, n_15487, n_15488, n_15489, n_15490, n_15491, n_15492, n_15493, n_15494, n_15495, n_15496, n_15497, n_15498, n_15499, n_15500, n_15501, n_15502, n_15503, n_15504, n_15505, n_15506, n_15507, n_15508, n_15509, n_15510, n_15511, n_15512, n_15513, n_15514, n_15515, n_15516, n_15517, n_15518, n_15519, n_15520, n_15521, n_15522, n_15523, n_15524, n_15525, n_15526, n_15527, n_15528, n_15529, n_15530, n_15531, n_15532, n_15533, n_15534, n_15535, n_15536, n_15537, n_15538, n_15539, n_15540, n_15541, n_15542, n_15543, n_15544, n_15545, n_15546, n_15547, n_15548, n_15549, n_15550, n_15551, n_15552, n_15553, n_15554, n_15555, n_15556, n_15557, n_15558, n_15559, n_15560, n_15561, n_15562, n_15563, n_15564, n_15565, n_15566, n_15567, n_15568, n_15569, n_15570, n_15571, n_15572, n_15573, n_15574, n_15575, n_15576, n_15577, n_15578, n_15579, n_15580, n_15581, n_15582, n_15583, n_15584, n_15585, n_15586, n_15587, n_15588, n_15589, n_15590, n_15591, n_15592, n_15593, n_15594, n_15595, n_15596, n_15597, n_15598, n_15599, n_15600, n_15601, n_15602, n_15603, n_15604, n_15605, n_15606, n_15607, n_15608, n_15609, n_15610, n_15611, n_15612, n_15613, n_15614, n_15615, n_15616, n_15617, n_15618, n_15619, n_15620, n_15621, n_15622, n_15623, n_15624, n_15625, n_15626, n_15627, n_15628, n_15629, n_15630, n_15631, n_15632, n_15633, n_15634, n_15635, n_15636, n_15637, n_15638, n_15639, n_15640, n_15641, n_15642, n_15643, n_15644, n_15645, n_15646, n_15647, n_15648, n_15649, n_15650, n_15651, n_15652, n_15653, n_15654, n_15655, n_15656, n_15657, n_15658, n_15659, n_15660, n_15661, n_15662, n_15663, n_15664, n_15665, n_15666, n_15667, n_15668, n_15669, n_15670, n_15671, n_15672, n_15673, n_15674, n_15675, n_15676, n_15677, n_15678, n_15679, n_15680, n_15681, n_15682, n_15683, n_15684, n_15685, n_15686, n_15687, n_15688, n_15689, n_15690, n_15691, n_15692, n_15693, n_15694, n_15695, n_15696, n_15697, n_15698, n_15699, n_15700, n_15701, n_15702, n_15703, n_15704, n_15705, n_15706, n_15707, n_15708, n_15709, n_15710, n_15711, n_15712, n_15713, n_15714, n_15715, n_15716, n_15717, n_15718, n_15719, n_15720, n_15721, n_15722, n_15723, n_15724, n_15725, n_15726, n_15727, n_15728, n_15729, n_15730, n_15731, n_15732, n_15733, n_15734, n_15735, n_15736, n_15737, n_15738, n_15739, n_15740, n_15741, n_15742, n_15743, n_15744, n_15745, n_15746, n_15747, n_15748, n_15749, n_15750, n_15751, n_15752, n_15753, n_15754, n_15755, n_15756, n_15757, n_15758, n_15759, n_15760, n_15761, n_15762, n_15763, n_15764, n_15765, n_15766, n_15767, n_15768, n_15769, n_15770, n_15771, n_15772, n_15773, n_15774, n_15775, n_15776, n_15777, n_15778, n_15779, n_15780, n_15781, n_15782, n_15783, n_15784, n_15785, n_15786, n_15787, n_15788, n_15789, n_15790, n_15791, n_15792, n_15793, n_15794, n_15795, n_15796, n_15797, n_15798, n_15799, n_15800, n_15801, n_15802, n_15803, n_15804, n_15805, n_15806, n_15807, n_15808, n_15809, n_15810, n_15811, n_15812, n_15813, n_15814, n_15815, n_15816, n_15817, n_15818, n_15819, n_15820, n_15821, n_15822, n_15823, n_15824, n_15825, n_15826, n_15827, n_15828, n_15829, n_15830, n_15831, n_15832, n_15833, n_15834, n_15835, n_15836, n_15837, n_15838, n_15839, n_15840, n_15841, n_15842, n_15843, n_15844, n_15845, n_15846, n_15847, n_15848, n_15849, n_15850, n_15851, n_15852, n_15853, n_15854, n_15855, n_15856, n_15857, n_15858, n_15859, n_15860, n_15861, n_15862, n_15863, n_15864, n_15865, n_15866, n_15867, n_15868, n_15869, n_15870, n_15871, n_15872, n_15873, n_15874, n_15875, n_15876, n_15877, n_15878, n_15879, n_15880, n_15881, n_15882, n_15883, n_15884, n_15885, n_15886, n_15887, n_15888, n_15889, n_15890, n_15891, n_15892, n_15893, n_15894, n_15895, n_15896, n_15897, n_15898, n_15899, n_15900, n_15901, n_15902, n_15903, n_15904, n_15905, n_15906, n_15907, n_15908, n_15909, n_15910, n_15911, n_15912, n_15913, n_15914, n_15915, n_15916, n_15917, n_15918, n_15919, n_15920, n_15921, n_15922, n_15923, n_15924, n_15925, n_15926, n_15927, n_15928, n_15929, n_15930, n_15931, n_15932, n_15933, n_15934, n_15935, n_15936, n_15937, n_15938, n_15939, n_15940, n_15941, n_15942, n_15943, n_15944, n_15945, n_15946, n_15947, n_15948, n_15949, n_15950, n_15951, n_15952, n_15953, n_15954, n_15955, n_15956, n_15957, n_15958, n_15959, n_15960, n_15961, n_15962, n_15963, n_15964, n_15965, n_15966, n_15967, n_15968, n_15969, n_15970, n_15971, n_15972, n_15973, n_15974, n_15975, n_15976, n_15977, n_15978, n_15979, n_15980, n_15981, n_15982, n_15983, n_15984, n_15985, n_15986, n_15987, n_15988, n_15989, n_15990, n_15991, n_15992, n_15993, n_15994, n_15995, n_15996, n_15997, n_15998, n_15999, n_16000, n_16001, n_16002, n_16003, n_16004, n_16005, n_16006, n_16007, n_16008, n_16009, n_16010, n_16011, n_16012, n_16013, n_16014, n_16015, n_16016, n_16017, n_16018, n_16019, n_16020, n_16021, n_16022, n_16023, n_16024, n_16025, n_16026, n_16027, n_16028, n_16029, n_16030, n_16031, n_16032, n_16033, n_16034, n_16035, n_16036, n_16037, n_16038, n_16039, n_16040, n_16041, n_16042, n_16043, n_16044, n_16045, n_16046, n_16047, n_16048, n_16049, n_16050, n_16051, n_16052, n_16053, n_16054, n_16055, n_16056, n_16057, n_16058, n_16059, n_16060, n_16061, n_16062, n_16063, n_16064, n_16065, n_16066, n_16067, n_16068, n_16069, n_16070, n_16071, n_16072, n_16073, n_16074, n_16075, n_16076, n_16077, n_16078, n_16079, n_16080, n_16081, n_16082, n_16083, n_16084, n_16085, n_16086, n_16087, n_16088, n_16089, n_16090, n_16091, n_16092, n_16093, n_16094, n_16095, n_16096, n_16097, n_16098, n_16099, n_16100, n_16101, n_16102, n_16103, n_16104, n_16105, n_16106, n_16107, n_16108, n_16109, n_16110, n_16111, n_16112, n_16113, n_16114, n_16115, n_16116, n_16117, n_16118, n_16119, n_16120, n_16121, n_16122, n_16123, n_16124, n_16125, n_16126, n_16127, n_16128, n_16129, n_16130, n_16131, n_16132, n_16133, n_16134, n_16135, n_16136, n_16137, n_16138, n_16139, n_16140, n_16141, n_16142, n_16143, n_16144, n_16145, n_16146, n_16147, n_16148, n_16149, n_16150, n_16151, n_16152, n_16153, n_16154, n_16155, n_16156, n_16157, n_16158, n_16159, n_16160, n_16161, n_16162, n_16163, n_16164, n_16165, n_16166, n_16167, n_16168, n_16169, n_16170, n_16171, n_16172, n_16173, n_16174, n_16175, n_16176, n_16177, n_16178, n_16179, n_16180, n_16181, n_16182, n_16183, n_16184, n_16185, n_16186, n_16187, n_16188, n_16189, n_16190, n_16191, n_16192, n_16193, n_16194, n_16195, n_16196, n_16197, n_16198, n_16199, n_16200, n_16201, n_16202, n_16203, n_16204, n_16205, n_16206, n_16207, n_16208, n_16209, n_16210, n_16211, n_16212, n_16213, n_16214, n_16215, n_16216, n_16217, n_16218, n_16219, n_16220, n_16221, n_16222, n_16223, n_16224, n_16225, n_16226, n_16227, n_16228, n_16229, n_16230, n_16231, n_16232, n_16233, n_16234, n_16235, n_16236, n_16237, n_16238, n_16239, n_16240, n_16241, n_16242, n_16243, n_16244, n_16245, n_16246, n_16247, n_16248, n_16249, n_16250, n_16251, n_16252, n_16253, n_16254, n_16255, n_16256, n_16257, n_16258, n_16259, n_16260, n_16261, n_16262, n_16263, n_16264, n_16265, n_16266, n_16267, n_16268, n_16269, n_16270, n_16271, n_16272, n_16273, n_16274, n_16275, n_16276, n_16277, n_16278, n_16279, n_16280, n_16281, n_16282, n_16283, n_16284, n_16285, n_16286, n_16287, n_16288, n_16289, n_16290, n_16291, n_16292, n_16293, n_16294, n_16295, n_16296, n_16297, n_16298, n_16299, n_16300, n_16301, n_16302, n_16303, n_16304, n_16305, n_16306, n_16307, n_16308, n_16309, n_16310, n_16311, n_16312, n_16313, n_16314, n_16315, n_16316, n_16317, n_16318, n_16319, n_16320, n_16321, n_16322, n_16323, n_16324, n_16325, n_16326, n_16327, n_16328, n_16329, n_16330, n_16331, n_16332, n_16333, n_16334, n_16335, n_16336, n_16337, n_16338, n_16339, n_16340, n_16341, n_16342, n_16343, n_16344, n_16345, n_16346, n_16347, n_16348, n_16349, n_16350, n_16351, n_16352, n_16353, n_16354, n_16355, n_16356, n_16357, n_16358, n_16359, n_16360, n_16361, n_16362, n_16363, n_16364, n_16365, n_16366, n_16367, n_16368, n_16369, n_16370, n_16371, n_16372, n_16373, n_16374, n_16375, n_16376, n_16377, n_16378, n_16379, n_16380, n_16381, n_16382, n_16383, n_16384, n_16385, n_16386, n_16387, n_16388, n_16389, n_16390, n_16391, n_16392, n_16393, n_16394, n_16395, n_16396, n_16397, n_16398, n_16399, n_16400, n_16401, n_16402, n_16403, n_16404, n_16405, n_16406, n_16407, n_16408, n_16409, n_16410, n_16411, n_16412, n_16413, n_16414, n_16415, n_16416, n_16417, n_16418, n_16419, n_16420, n_16421, n_16422, n_16423, n_16424, n_16425, n_16426, n_16427, n_16428, n_16429, n_16430, n_16431, n_16432, n_16433, n_16434, n_16435, n_16436, n_16437, n_16438, n_16439, n_16440, n_16441, n_16442, n_16443, n_16444, n_16445, n_16446, n_16447, n_16448, n_16449, n_16450, n_16451, n_16452, n_16453, n_16454, n_16455, n_16456, n_16457, n_16458, n_16459, n_16460, n_16461, n_16462, n_16463, n_16464, n_16465, n_16466, n_16467, n_16468, n_16469, n_16470, n_16471, n_16472, n_16473, n_16474, n_16475, n_16476, n_16477, n_16478, n_16479, n_16480, n_16481, n_16482, n_16483, n_16484, n_16485, n_16486, n_16487, n_16488, n_16489, n_16490, n_16491, n_16492, n_16493, n_16494, n_16495, n_16496, n_16497, n_16498, n_16499, n_16500, n_16501, n_16502, n_16503, n_16504, n_16505, n_16506, n_16507, n_16508, n_16509, n_16510, n_16511, n_16512, n_16513, n_16514, n_16515, n_16516, n_16517, n_16518, n_16519, n_16520, n_16521, n_16522, n_16523, n_16524, n_16525, n_16526, n_16527, n_16528, n_16529, n_16530, n_16531, n_16532, n_16533, n_16534, n_16535, n_16536, n_16537, n_16538, n_16539, n_16540, n_16541, n_16542, n_16543, n_16544, n_16545, n_16546, n_16547, n_16548, n_16549, n_16550, n_16551, n_16552, n_16553, n_16554, n_16555, n_16556, n_16557, n_16558, n_16559, n_16560, n_16561, n_16562, n_16563, n_16564, n_16565, n_16566, n_16567, n_16568, n_16569, n_16570, n_16571, n_16572, n_16573, n_16574, n_16575, n_16576, n_16577, n_16578, n_16579, n_16580, n_16581, n_16582, n_16583, n_16584, n_16585, n_16586, n_16587, n_16588, n_16589, n_16590, n_16591, n_16592, n_16593, n_16594, n_16595, n_16596, n_16597, n_16598, n_16599, n_16600, n_16601, n_16602, n_16603, n_16604, n_16605, n_16606, n_16607, n_16608, n_16609, n_16610, n_16611, n_16612, n_16613, n_16614, n_16615, n_16616, n_16617, n_16618, n_16619, n_16620, n_16621, n_16622, n_16623, n_16624, n_16625, n_16626, n_16627, n_16628, n_16629, n_16630, n_16631, n_16632, n_16633, n_16634, n_16635, n_16636, n_16637, n_16638, n_16639, n_16640, n_16641, n_16642, n_16643, n_16644, n_16645, n_16646, n_16647, n_16648, n_16649, n_16650, n_16651, n_16652, n_16653, n_16654, n_16655, n_16656, n_16657, n_16658, n_16659, n_16660, n_16661, n_16662, n_16663, n_16664, n_16665, n_16666, n_16667, n_16668, n_16669, n_16670, n_16671, n_16672, n_16673, n_16674, n_16675, n_16676, n_16677, n_16678, n_16679, n_16680, n_16681, n_16682, n_16683, n_16684, n_16685, n_16686, n_16687, n_16688, n_16689, n_16690, n_16691, n_16692, n_16693, n_16694, n_16695, n_16696, n_16697, n_16698, n_16699, n_16700, n_16701, n_16702, n_16703, n_16704, n_16705, n_16706, n_16707, n_16708, n_16709, n_16710, n_16711, n_16712, n_16713, n_16714, n_16715, n_16716, n_16717, n_16718, n_16719, n_16720, n_16721, n_16722, n_16723, n_16724, n_16725, n_16726, n_16727, n_16728, n_16729, n_16730, n_16731, n_16732, n_16733, n_16734, n_16735, n_16736, n_16737, n_16738, n_16739, n_16740, n_16741, n_16742, n_16743, n_16744, n_16745, n_16746, n_16747, n_16748, n_16749, n_16750, n_16751, n_16752, n_16753, n_16754, n_16755, n_16756, n_16757, n_16758, n_16759, n_16760, n_16761, n_16762, n_16763, n_16764, n_16765, n_16766, n_16767, n_16768, n_16769, n_16770, n_16771, n_16772, n_16773, n_16774, n_16775, n_16776, n_16777, n_16778, n_16779, n_16780, n_16781, n_16782, n_16783, n_16784, n_16785, n_16786, n_16787, n_16788, n_16789, n_16790, n_16791, n_16792, n_16793, n_16794, n_16795, n_16796, n_16797, n_16798, n_16799, n_16800, n_16801, n_16802, n_16803, n_16804, n_16805, n_16806, n_16807, n_16808, n_16809, n_16810, n_16811, n_16812, n_16813, n_16814, n_16815, n_16816, n_16817, n_16818, n_16819, n_16820, n_16821, n_16822, n_16823, n_16824, n_16825, n_16826, n_16827, n_16828, n_16829, n_16830, n_16831, n_16832, n_16833, n_16834, n_16835, n_16836, n_16837, n_16838, n_16839, n_16840, n_16841, n_16842, n_16843, n_16844, n_16845, n_16846, n_16847, n_16848, n_16849, n_16850, n_16851, n_16852, n_16853, n_16854, n_16855, n_16856, n_16857, n_16858, n_16859, n_16860, n_16861, n_16862, n_16863, n_16864, n_16865, n_16866, n_16867, n_16868, n_16869, n_16870, n_16871, n_16872, n_16873, n_16874, n_16875, n_16876, n_16877, n_16878, n_16879, n_16880, n_16881, n_16882, n_16883, n_16884, n_16885, n_16886, n_16887, n_16888, n_16889, n_16890, n_16891, n_16892, n_16893, n_16894, n_16895, n_16896, n_16897, n_16898, n_16899, n_16900, n_16901, n_16902, n_16903, n_16904, n_16905, n_16906, n_16907, n_16908, n_16909, n_16910, n_16911, n_16912, n_16913, n_16914, n_16915, n_16916, n_16917, n_16918, n_16919, n_16920, n_16921, n_16922, n_16923, n_16924, n_16925, n_16926, n_16927, n_16928, n_16929, n_16930, n_16931, n_16932, n_16933, n_16934, n_16935, n_16936, n_16937, n_16938, n_16939, n_16940, n_16941, n_16942, n_16943, n_16944, n_16945, n_16946, n_16947, n_16948, n_16949, n_16950, n_16951, n_16952, n_16953, n_16954, n_16955, n_16956, n_16957, n_16958, n_16959, n_16960, n_16961, n_16962, n_16963, n_16964, n_16965, n_16966, n_16967, n_16968, n_16969, n_16970, n_16971, n_16972, n_16973, n_16974, n_16975, n_16976, n_16977, n_16978, n_16979, n_16980, n_16981, n_16982, n_16983, n_16984, n_16985, n_16986, n_16987, n_16988, n_16989, n_16990, n_16991, n_16992, n_16993, n_16994, n_16995, n_16996, n_16997, n_16998, n_16999, n_17000, n_17001, n_17002, n_17003, n_17004, n_17005, n_17006, n_17007, n_17008, n_17009, n_17010, n_17011, n_17012, n_17013, n_17014, n_17015, n_17016, n_17017, n_17018, n_17019, n_17020, n_17021, n_17022, n_17023, n_17024, n_17025, n_17026, n_17027, n_17028, n_17029, n_17030, n_17031, n_17032, n_17033, n_17034, n_17035, n_17036, n_17037, n_17038, n_17039, n_17040, n_17041, n_17042, n_17043, n_17044, n_17045, n_17046, n_17047, n_17048, n_17049, n_17050, n_17051, n_17052, n_17053, n_17054, n_17055, n_17056, n_17057, n_17058, n_17059, n_17060, n_17061, n_17062, n_17063, n_17064, n_17065, n_17066, n_17067, n_17068, n_17069, n_17070, n_17071, n_17072, n_17073, n_17074, n_17075, n_17076, n_17077, n_17078, n_17079, n_17080, n_17081, n_17082, n_17083, n_17084, n_17085, n_17086, n_17087, n_17088, n_17089, n_17090, n_17091, n_17092, n_17093, n_17094, n_17095, n_17096, n_17097, n_17098, n_17099, n_17100, n_17101, n_17102, n_17103, n_17104, n_17105, n_17106, n_17107, n_17108, n_17109, n_17110, n_17111, n_17112, n_17113, n_17114, n_17115, n_17116, n_17117, n_17118, n_17119, n_17120, n_17121, n_17122, n_17123, n_17124, n_17125, n_17126, n_17127, n_17128, n_17129, n_17130, n_17131, n_17132, n_17133, n_17134, n_17135, n_17136, n_17137, n_17138, n_17139, n_17140, n_17141, n_17142, n_17143, n_17144, n_17145, n_17146, n_17147, n_17148, n_17149, n_17150, n_17151, n_17152, n_17153, n_17154, n_17155, n_17156, n_17157, n_17158, n_17159, n_17160, n_17161, n_17162, n_17163, n_17164, n_17165, n_17166, n_17167, n_17168, n_17169, n_17170, n_17171, n_17172, n_17173, n_17174, n_17175, n_17176, n_17177, n_17178, n_17179, n_17180, n_17181, n_17182, n_17183, n_17184, n_17185, n_17186, n_17187, n_17188, n_17189, n_17190, n_17191, n_17192, n_17193, n_17194, n_17195, n_17196, n_17197, n_17198, n_17199, n_17200, n_17201, n_17202, n_17203, n_17204, n_17205, n_17206, n_17207, n_17208, n_17209, n_17210, n_17211, n_17212, n_17213, n_17214, n_17215, n_17216, n_17217, n_17218, n_17219, n_17220, n_17221, n_17222, n_17223, n_17224, n_17225, n_17226, n_17227, n_17228, n_17229, n_17230, n_17231, n_17232, n_17233, n_17234, n_17235, n_17236, n_17237, n_17238, n_17239, n_17240, n_17241, n_17242, n_17243, n_17244, n_17245, n_17246, n_17247, n_17248, n_17249, n_17250, n_17251, n_17252, n_17253, n_17254, n_17255, n_17256, n_17257, n_17258, n_17259, n_17260, n_17261, n_17262, n_17263, n_17264, n_17265, n_17266, n_17267, n_17268, n_17269, n_17270, n_17271, n_17272, n_17273, n_17274, n_17275, n_17276, n_17277, n_17278, n_17279, n_17280, n_17281, n_17282, n_17283, n_17284, n_17285, n_17286, n_17287, n_17288, n_17289, n_17290, n_17291, n_17292, n_17293, n_17294, n_17295, n_17296, n_17297, n_17298, n_17299, n_17300, n_17301, n_17302, n_17303, n_17304, n_17305, n_17306, n_17307, n_17308, n_17309, n_17310, n_17311, n_17312, n_17313, n_17314, n_17315, n_17316, n_17317, n_17318, n_17319, n_17320, n_17321, n_17322, n_17323, n_17324, n_17325, n_17326, n_17327, n_17328, n_17329, n_17330, n_17331, n_17332, n_17333, n_17334, n_17335, n_17336, n_17337, n_17338, n_17339, n_17340, n_17341, n_17342, n_17343, n_17344, n_17345, n_17346, n_17347, n_17348, n_17349, n_17350, n_17351, n_17352, n_17353, n_17354, n_17355, n_17356, n_17357, n_17358, n_17359, n_17360, n_17361, n_17362, n_17363, n_17364, n_17365, n_17366, n_17367, n_17368, n_17369, n_17370, n_17371, n_17372, n_17373, n_17374, n_17375, n_17376, n_17377, n_17378, n_17379, n_17380, n_17381, n_17382, n_17383, n_17384, n_17385, n_17386, n_17387, n_17388, n_17389, n_17390, n_17391, n_17392, n_17393, n_17394, n_17395, n_17396, n_17397, n_17398, n_17399, n_17400, n_17401, n_17402, n_17403, n_17404, n_17405, n_17406, n_17407, n_17408, n_17409, n_17410, n_17411, n_17412, n_17413, n_17414, n_17415, n_17416, n_17417, n_17418, n_17419, n_17420, n_17421, n_17422, n_17423, n_17424, n_17425, n_17426, n_17427, n_17428, n_17429, n_17430, n_17431, n_17432, n_17433, n_17434, n_17435, n_17436, n_17437, n_17438, n_17439, n_17440, n_17441, n_17442, n_17443, n_17444, n_17445, n_17446, n_17447, n_17448, n_17449, n_17450, n_17451, n_17452, n_17453, n_17454, n_17455, n_17456, n_17457, n_17458, n_17459, n_17460, n_17461, n_17462, n_17463, n_17464, n_17465, n_17466, n_17467, n_17468, n_17469, n_17470, n_17471, n_17472, n_17473, n_17474, n_17475, n_17476, n_17477, n_17478, n_17479, n_17480, n_17481, n_17482, n_17483, n_17484, n_17485, n_17486, n_17487, n_17488, n_17489, n_17490, n_17491, n_17492, n_17493, n_17494, n_17495, n_17496, n_17497, n_17498, n_17499, n_17500, n_17501, n_17502, n_17503, n_17504, n_17505, n_17506, n_17507, n_17508, n_17509, n_17510, n_17511, n_17512, n_17513, n_17514, n_17515, n_17516, n_17517, n_17518, n_17519, n_17520, n_17521, n_17522, n_17523, n_17524, n_17525, n_17526, n_17527, n_17528, n_17529, n_17530, n_17531, n_17532, n_17533, n_17534, n_17535, n_17536, n_17537, n_17538, n_17539, n_17540, n_17541, n_17542, n_17543, n_17544, n_17545, n_17546, n_17547, n_17548, n_17549, n_17550, n_17551, n_17552, n_17553, n_17554, n_17555, n_17556, n_17557, n_17558, n_17559, n_17560, n_17561, n_17562, n_17563, n_17564, n_17565, n_17566, n_17567, n_17568, n_17569, n_17570, n_17571, n_17572, n_17573, n_17574, n_17575, n_17576, n_17577, n_17578, n_17579, n_17580, n_17581, n_17582, n_17583, n_17584, n_17585, n_17586, n_17587, n_17588, n_17589, n_17590, n_17591, n_17592, n_17593, n_17594, n_17595, n_17596, n_17597, n_17598, n_17599, n_17600, n_17601, n_17602, n_17603, n_17604, n_17605, n_17606, n_17607, n_17608, n_17609, n_17610, n_17611, n_17612, n_17613, n_17614, n_17615, n_17616, n_17617, n_17618, n_17619, n_17620, n_17621, n_17622, n_17623, n_17624, n_17625, n_17626, n_17627, n_17628, n_17629, n_17630, n_17631, n_17632, n_17633, n_17634, n_17635, n_17636, n_17637, n_17638, n_17639, n_17640, n_17641, n_17642, n_17643, n_17644, n_17645, n_17646, n_17647, n_17648, n_17649, n_17650, n_17651, n_17652, n_17653, n_17654, n_17655, n_17656, n_17657, n_17658, n_17659, n_17660, n_17661, n_17662, n_17663, n_17664, n_17665, n_17666, n_17667, n_17668, n_17669, n_17670, n_17671, n_17672, n_17673, n_17674, n_17675, n_17676, n_17677, n_17678, n_17679, n_17680, n_17681, n_17682, n_17683, n_17684, n_17685, n_17686, n_17687, n_17688, n_17689, n_17690, n_17691, n_17692, n_17693, n_17694, n_17695, n_17696, n_17697, n_17698, n_17699, n_17700, n_17701, n_17702, n_17703, n_17704, n_17705, n_17706, n_17707, n_17708, n_17709, n_17710, n_17711, n_17712, n_17713, n_17714, n_17715, n_17716, n_17717, n_17718, n_17719, n_17720, n_17721, n_17722, n_17723, n_17724, n_17725, n_17726, n_17727, n_17728, n_17729, n_17730, n_17731, n_17732, n_17733, n_17734, n_17735, n_17736, n_17737, n_17738, n_17739, n_17740, n_17741, n_17742, n_17743, n_17744, n_17745, n_17746, n_17747, n_17748, n_17749, n_17750, n_17751, n_17752, n_17753, n_17754, n_17755, n_17756, n_17757, n_17758, n_17759, n_17760, n_17761, n_17762, n_17763, n_17764, n_17765, n_17766, n_17767, n_17768, n_17769, n_17770, n_17771, n_17772, n_17773, n_17774, n_17775, n_17776, n_17777, n_17778, n_17779, n_17780, n_17781, n_17782, n_17783, n_17784, n_17785, n_17786, n_17787, n_17788, n_17789, n_17790, n_17791, n_17792, n_17793, n_17794, n_17795, n_17796, n_17797, n_17798, n_17799, n_17800, n_17801, n_17802, n_17803, n_17804, n_17805, n_17806, n_17807, n_17808, n_17809, n_17810, n_17811, n_17812, n_17813, n_17814, n_17815, n_17816, n_17817, n_17818, n_17819, n_17820, n_17821, n_17822, n_17823, n_17824, n_17825, n_17826, n_17827, n_17828, n_17829, n_17830, n_17831, n_17832, n_17833, n_17834, n_17835, n_17836, n_17837, n_17838, n_17839, n_17840, n_17841, n_17842, n_17843, n_17844, n_17845, n_17846, n_17847, n_17848, n_17849, n_17850, n_17851, n_17852, n_17853, n_17854, n_17855, n_17856, n_17857, n_17858, n_17859, n_17860, n_17861, n_17862, n_17863, n_17864, n_17865, n_17866, n_17867, n_17868, n_17869, n_17870, n_17871, n_17872, n_17873, n_17874, n_17875, n_17876, n_17877, n_17878, n_17879, n_17880, n_17881, n_17882, n_17883, n_17884, n_17885, n_17886, n_17887, n_17888, n_17889, n_17890, n_17891, n_17892, n_17893, n_17894, n_17895, n_17896, n_17897, n_17898, n_17899, n_17900, n_17901, n_17902, n_17903, n_17904, n_17905, n_17906, n_17907, n_17908, n_17909, n_17910, n_17911, n_17912, n_17913, n_17914, n_17915, n_17916, n_17917, n_17918, n_17919, n_17920, n_17921, n_17922, n_17923, n_17924, n_17925, n_17926, n_17927, n_17928, n_17929, n_17930, n_17931, n_17932, n_17933, n_17934, n_17935, n_17936, n_17937, n_17938, n_17939, n_17940, n_17941, n_17942, n_17943, n_17944, n_17945, n_17946, n_17947, n_17948, n_17949, n_17950, n_17951, n_17952, n_17953, n_17954, n_17955, n_17956, n_17957, n_17958, n_17959, n_17960, n_17961, n_17962, n_17963, n_17964, n_17965, n_17966, n_17967, n_17968, n_17969, n_17970, n_17971, n_17972, n_17973, n_17974, n_17975, n_17976, n_17977, n_17978, n_17979, n_17980, n_17981, n_17982, n_17983, n_17984, n_17985, n_17986, n_17987, n_17988, n_17989, n_17990, n_17991, n_17992, n_17993, n_17994, n_17995, n_17996, n_17997, n_17998, n_17999, n_18000, n_18001, n_18002, n_18003, n_18004, n_18005, n_18006, n_18007, n_18008, n_18009, n_18010, n_18011, n_18012, n_18013, n_18014, n_18015, n_18016, n_18017, n_18018, n_18019, n_18020, n_18021, n_18022, n_18023, n_18024, n_18025, n_18026, n_18027, n_18028, n_18029, n_18030, n_18031, n_18032, n_18033, n_18034, n_18035, n_18036, n_18037, n_18038, n_18039, n_18040, n_18041, n_18042, n_18043, n_18044, n_18045, n_18046, n_18047, n_18048, n_18049, n_18050, n_18051, n_18052, n_18053, n_18054, n_18055, n_18056, n_18057, n_18058, n_18059, n_18060, n_18061, n_18062, n_18063, n_18064, n_18065, n_18066, n_18067, n_18068, n_18069, n_18070, n_18071, n_18072, n_18073, n_18074, n_18075, n_18076, n_18077, n_18078, n_18079, n_18080, n_18081, n_18082, n_18083, n_18084, n_18085, n_18086, n_18087, n_18088, n_18089, n_18090, n_18091, n_18092, n_18093, n_18094, n_18095, n_18096, n_18097, n_18098, n_18099, n_18100, n_18101, n_18102, n_18103, n_18104, n_18105, n_18106, n_18107, n_18108, n_18109, n_18110, n_18111, n_18112, n_18113, n_18114, n_18115, n_18116, n_18117, n_18118, n_18119, n_18120, n_18121, n_18122, n_18123, n_18124, n_18125, n_18126, n_18127, n_18128, n_18129, n_18130, n_18131, n_18132, n_18133, n_18134, n_18135, n_18136, n_18137, n_18138, n_18139, n_18140, n_18141, n_18142, n_18143, n_18144, n_18145, n_18146, n_18147, n_18148, n_18149, n_18150, n_18151, n_18152, n_18153, n_18154, n_18155, n_18156, n_18157, n_18158, n_18159, n_18160, n_18161, n_18162, n_18163, n_18164, n_18165, n_18166, n_18167, n_18168, n_18169, n_18170, n_18171, n_18172, n_18173, n_18174, n_18175, n_18176, n_18177, n_18178, n_18179, n_18180, n_18181, n_18182, n_18183, n_18184, n_18185, n_18186, n_18187, n_18188, n_18189, n_18190, n_18191, n_18192, n_18193, n_18194, n_18195, n_18196, n_18197, n_18198, n_18199, n_18200, n_18201, n_18202, n_18203, n_18204, n_18205, n_18206, n_18207, n_18208, n_18209, n_18210, n_18211, n_18212, n_18213, n_18214, n_18215, n_18216, n_18217, n_18218, n_18219, n_18220, n_18221, n_18222, n_18223, n_18224, n_18225, n_18226, n_18227, n_18228, n_18229, n_18230, n_18231, n_18232, n_18233, n_18234, n_18235, n_18236, n_18237, n_18238, n_18239, n_18240, n_18241, n_18242, n_18243, n_18244, n_18245, n_18246, n_18247, n_18248, n_18249, n_18250, n_18251, n_18252, n_18253, n_18254, n_18255, n_18256, n_18257, n_18258, n_18259, n_18260, n_18261, n_18262, n_18263, n_18264, n_18265, n_18266, n_18267, n_18268, n_18269, n_18270, n_18271, n_18272, n_18273, n_18274, n_18275, n_18276, n_18277, n_18278, n_18279, n_18280, n_18281, n_18282, n_18283, n_18284, n_18285, n_18286, n_18287, n_18288, n_18289, n_18290, n_18291, n_18292, n_18293, n_18294, n_18295, n_18296, n_18297, n_18298, n_18299, n_18300, n_18301, n_18302, n_18303, n_18304, n_18305, n_18306, n_18307, n_18308, n_18309, n_18310, n_18311, n_18312, n_18313, n_18314, n_18315, n_18316, n_18317, n_18318, n_18319, n_18320, n_18321, n_18322, n_18323, n_18324, n_18325, n_18326, n_18327, n_18328, n_18329, n_18330, n_18331, n_18332, n_18333, n_18334, n_18335, n_18336, n_18337, n_18338, n_18339, n_18340, n_18341, n_18342, n_18343, n_18344, n_18345, n_18346, n_18347, n_18348, n_18349, n_18350, n_18351, n_18352, n_18353, n_18354, n_18355, n_18356, n_18357, n_18358, n_18359, n_18360, n_18361, n_18362, n_18363, n_18364, n_18365, n_18366, n_18367, n_18368, n_18369, n_18370, n_18371, n_18372, n_18373, n_18374, n_18375, n_18376, n_18377, n_18378, n_18379, n_18380, n_18381, n_18382, n_18383, n_18384, n_18385, n_18386, n_18387, n_18388, n_18389, n_18390, n_18391, n_18392, n_18393, n_18394, n_18395, n_18396, n_18397, n_18398, n_18399, n_18400, n_18401, n_18402, n_18403, n_18404, n_18405, n_18406, n_18407, n_18408, n_18409, n_18410, n_18411, n_18412, n_18413, n_18414, n_18415, n_18416, n_18417, n_18418, n_18419, n_18420, n_18421, n_18422, n_18423, n_18424, n_18425, n_18426, n_18427, n_18428, n_18429, n_18430, n_18431, n_18432, n_18433, n_18434, n_18435, n_18436, n_18437, n_18438, n_18439, n_18440, n_18441, n_18442, n_18443, n_18444, n_18445, n_18446, n_18447, n_18448, n_18449, n_18450, n_18451, n_18452, n_18453, n_18454, n_18455, n_18456, n_18457, n_18458, n_18459, n_18460, n_18461, n_18462, n_18463, n_18464, n_18465, n_18466, n_18467, n_18468, n_18469, n_18470, n_18471, n_18472, n_18473, n_18474, n_18475, n_18476, n_18477, n_18478, n_18479, n_18480, n_18481, n_18482, n_18483, n_18484, n_18485, n_18486, n_18487, n_18488, n_18489, n_18490, n_18491, n_18492, n_18493, n_18494, n_18495, n_18496, n_18497, n_18498, n_18499, n_18500, n_18501, n_18502, n_18503, n_18504, n_18505, n_18506, n_18507, n_18508, n_18509, n_18510, n_18511, n_18512, n_18513, n_18514, n_18515, n_18516, n_18517, n_18518, n_18519, n_18520, n_18521, n_18522, n_18523, n_18524, n_18525, n_18526, n_18527, n_18528, n_18529, n_18530, n_18531, n_18532, n_18533, n_18534, n_18535, n_18536, n_18537, n_18538, n_18539, n_18540, n_18541, n_18542, n_18543, n_18544, n_18545, n_18546, n_18547, n_18548, n_18549, n_18550, n_18551, n_18552, n_18553, n_18554, n_18555, n_18556, n_18557, n_18558, n_18559, n_18560, n_18561, n_18562, n_18563, n_18564, n_18565, n_18566, n_18567, n_18568, n_18569, n_18570, n_18571, n_18572, n_18573, n_18574, n_18575, n_18576, n_18577, n_18578, n_18579, n_18580, n_18581, n_18582, n_18583, n_18584, n_18585, n_18586, n_18587, n_18588, n_18589, n_18590, n_18591, n_18592, n_18593, n_18594, n_18595, n_18596, n_18597, n_18598, n_18599, n_18600, n_18601, n_18602, n_18603, n_18604, n_18605, n_18606, n_18607, n_18608, n_18609, n_18610, n_18611, n_18612, n_18613, n_18614, n_18615, n_18616, n_18617, n_18618, n_18619, n_18620, n_18621, n_18622, n_18623, n_18624, n_18625, n_18626, n_18627, n_18628, n_18629, n_18630, n_18631, n_18632, n_18633, n_18634, n_18635, n_18636, n_18637, n_18638, n_18639, n_18640, n_18641, n_18642, n_18643, n_18644, n_18645, n_18646, n_18647, n_18648, n_18649, n_18650, n_18651, n_18652, n_18653, n_18654, n_18655, n_18656, n_18657, n_18658, n_18659, n_18660, n_18661, n_18662, n_18663, n_18664, n_18665, n_18666, n_18667, n_18668, n_18669, n_18670, n_18671, n_18672, n_18673, n_18674, n_18675, n_18676, n_18677, n_18678, n_18679, n_18680, n_18681, n_18682, n_18683, n_18684, n_18685, n_18686, n_18687, n_18688, n_18689, n_18690, n_18691, n_18692, n_18693, n_18694, n_18695, n_18696, n_18697, n_18698, n_18699, n_18700, n_18701, n_18702, n_18703, n_18704, n_18705, n_18706, n_18707, n_18708, n_18709, n_18710, n_18711, n_18712, n_18713, n_18714, n_18715, n_18716, n_18717, n_18718, n_18719, n_18720, n_18721, n_18722, n_18723, n_18724, n_18725, n_18726, n_18727, n_18728, n_18729, n_18730, n_18731, n_18732, n_18733, n_18734, n_18735, n_18736, n_18737, n_18738, n_18739, n_18740, n_18741, n_18742, n_18743, n_18744, n_18745, n_18746, n_18747, n_18748, n_18749, n_18750, n_18751, n_18752, n_18753, n_18754, n_18755, n_18756, n_18757, n_18758, n_18759, n_18760, n_18761, n_18762, n_18763, n_18764, n_18765, n_18766, n_18767, n_18768, n_18769, n_18770, n_18771, n_18772, n_18773, n_18774, n_18775, n_18776, n_18777, n_18778, n_18779, n_18780, n_18781, n_18782, n_18783, n_18784, n_18785, n_18786, n_18787, n_18788, n_18789, n_18790, n_18791, n_18792, n_18793, n_18794, n_18795, n_18796, n_18797, n_18798, n_18799, n_18800, n_18801, n_18802, n_18803, n_18804, n_18805, n_18806, n_18807, n_18808, n_18809, n_18810, n_18811, n_18812, n_18813, n_18814, n_18815, n_18816, n_18817, n_18818, n_18819, n_18820, n_18821, n_18822, n_18823, n_18824, n_18825, n_18826, n_18827, n_18828, n_18829, n_18830, n_18831, n_18832, n_18833, n_18834, n_18835, n_18836, n_18837, n_18838, n_18839, n_18840, n_18841, n_18842, n_18843, n_18844, n_18845, n_18846, n_18847, n_18848, n_18849, n_18850, n_18851, n_18852, n_18853, n_18854, n_18855, n_18856, n_18857, n_18858, n_18859, n_18860, n_18861, n_18862, n_18863, n_18864, n_18865, n_18866, n_18867, n_18868, n_18869, n_18870, n_18871, n_18872, n_18873, n_18874, n_18875, n_18876, n_18877, n_18878, n_18879, n_18880, n_18881, n_18882, n_18883, n_18884, n_18885, n_18886, n_18887, n_18888, n_18889, n_18890, n_18891, n_18892, n_18893, n_18894, n_18895, n_18896, n_18897, n_18898, n_18899, n_18900, n_18901, n_18902, n_18903, n_18904, n_18905, n_18906, n_18907, n_18908, n_18909, n_18910, n_18911, n_18912, n_18913, n_18914, n_18915, n_18916, n_18917, n_18918, n_18919, n_18920, n_18921, n_18922, n_18923, n_18924, n_18925, n_18926, n_18927, n_18928, n_18929, n_18930, n_18931, n_18932, n_18933, n_18934, n_18935, n_18936, n_18937, n_18938, n_18939, n_18940, n_18941, n_18942, n_18943, n_18944, n_18945, n_18946, n_18947, n_18948, n_18949, n_18950, n_18951, n_18952, n_18953, n_18954, n_18955, n_18956, n_18957, n_18958, n_18959, n_18960, n_18961, n_18962, n_18963, n_18964, n_18965, n_18966, n_18967, n_18968, n_18969, n_18970, n_18971, n_18972, n_18973, n_18974, n_18975, n_18976, n_18977, n_18978, n_18979, n_18980, n_18981, n_18982, n_18983, n_18984, n_18985, n_18986, n_18987, n_18988, n_18989, n_18990, n_18991, n_18992, n_18993, n_18994, n_18995, n_18996, n_18997, n_18998, n_18999, n_19000, n_19001, n_19002, n_19003, n_19004, n_19005, n_19006, n_19007, n_19008, n_19009, n_19010, n_19011, n_19012, n_19013, n_19014, n_19015, n_19016, n_19017, n_19018, n_19019, n_19020, n_19021, n_19022, n_19023, n_19024, n_19025, n_19026, n_19027, n_19028, n_19029, n_19030, n_19031, n_19032, n_19033, n_19034, n_19035, n_19036, n_19037, n_19038, n_19039, n_19040, n_19041, n_19042, n_19043, n_19044, n_19045, n_19046, n_19047, n_19048, n_19049, n_19050, n_19051, n_19052, n_19053, n_19054, n_19055, n_19056, n_19057, n_19058, n_19059, n_19060, n_19061, n_19062, n_19063, n_19064, n_19065, n_19066, n_19067, n_19068, n_19069, n_19070, n_19071, n_19072, n_19073, n_19074, n_19075, n_19076, n_19077, n_19078, n_19079, n_19080, n_19081, n_19082, n_19083, n_19084, n_19085, n_19086, n_19087, n_19088, n_19089, n_19090, n_19091, n_19092, n_19093, n_19094, n_19095, n_19096, n_19097, n_19098, n_19099, n_19100, n_19101, n_19102, n_19103, n_19104, n_19105, n_19106, n_19107, n_19108, n_19109, n_19110, n_19111, n_19112, n_19113, n_19114, n_19115, n_19116, n_19117, n_19118, n_19119, n_19120, n_19121, n_19122, n_19123, n_19124, n_19125, n_19126, n_19127, n_19128, n_19129, n_19130, n_19131, n_19132, n_19133, n_19134, n_19135, n_19136, n_19137, n_19138, n_19139, n_19140, n_19141, n_19142, n_19143, n_19144, n_19145, n_19146, n_19147, n_19148, n_19149, n_19150, n_19151, n_19152, n_19153, n_19154, n_19155, n_19156, n_19157, n_19158, n_19159, n_19160, n_19161, n_19162, n_19163, n_19164, n_19165, n_19166, n_19167, n_19168, n_19169, n_19170, n_19171, n_19172, n_19173, n_19174, n_19175, n_19176, n_19177, n_19178, n_19179, n_19180, n_19181, n_19182, n_19183, n_19184, n_19185, n_19186, n_19187, n_19188, n_19189, n_19190, n_19191, n_19192, n_19193, n_19194, n_19195, n_19196, n_19197, n_19198, n_19199, n_19200, n_19201, n_19202, n_19203, n_19204, n_19205, n_19206, n_19207, n_19208, n_19209, n_19210, n_19211, n_19212, n_19213, n_19214, n_19215, n_19216, n_19217, n_19218, n_19219, n_19220, n_19221, n_19222, n_19223, n_19224, n_19225, n_19226, n_19227, n_19228, n_19229, n_19230, n_19231, n_19232, n_19233, n_19234, n_19235, n_19236, n_19237, n_19238, n_19239, n_19240, n_19241, n_19242, n_19243, n_19244, n_19245, n_19246, n_19247, n_19248, n_19249, n_19250, n_19251, n_19252, n_19253, n_19254, n_19255, n_19256, n_19257, n_19258, n_19259, n_19260, n_19261, n_19262, n_19263, n_19264, n_19265, n_19266, n_19267, n_19268, n_19269, n_19270, n_19271, n_19272, n_19273, n_19274, n_19275, n_19276, n_19277, n_19278, n_19279, n_19280, n_19281, n_19282, n_19283, n_19284, n_19285, n_19286, n_19287, n_19288, n_19289, n_19290, n_19291, n_19292, n_19293, n_19294, n_19295, n_19296, n_19297, n_19298, n_19299, n_19300, n_19301, n_19302, n_19303, n_19304, n_19305, n_19306, n_19307, n_19308, n_19309, n_19310, n_19311, n_19312, n_19313, n_19314, n_19315, n_19316, n_19317, n_19318, n_19319, n_19320, n_19321, n_19322, n_19323, n_19324, n_19325, n_19326, n_19327, n_19328, n_19329, n_19330, n_19331, n_19332, n_19333, n_19334, n_19335, n_19336, n_19337, n_19338, n_19339, n_19340, n_19341, n_19342, n_19343, n_19344, n_19345, n_19346, n_19347, n_19348, n_19349, n_19350, n_19351, n_19352, n_19353, n_19354, n_19355, n_19356, n_19357, n_19358, n_19359, n_19360, n_19361, n_19362, n_19363, n_19364, n_19365, n_19366, n_19367, n_19368, n_19369, n_19370, n_19371, n_19372, n_19373, n_19374, n_19375, n_19376, n_19377, n_19378, n_19379, n_19380, n_19381, n_19382, n_19383, n_19384, n_19385, n_19386, n_19387, n_19388, n_19389, n_19390, n_19391, n_19392, n_19393, n_19394, n_19395, n_19396, n_19397, n_19398, n_19399, n_19400, n_19401, n_19402, n_19403, n_19404, n_19405, n_19406, n_19407, n_19408, n_19409, n_19410, n_19411, n_19412, n_19413, n_19414, n_19415, n_19416, n_19417, n_19418, n_19419, n_19420, n_19421, n_19422, n_19423, n_19424, n_19425, n_19426, n_19427, n_19428, n_19429, n_19430, n_19431, n_19432, n_19433, n_19434, n_19435, n_19436, n_19437, n_19438, n_19439, n_19440, n_19441, n_19442, n_19443, n_19444, n_19445, n_19446, n_19447, n_19448, n_19449, n_19450, n_19451, n_19452, n_19453, n_19454, n_19455, n_19456, n_19457, n_19458, n_19459, n_19460, n_19461, n_19462, n_19463, n_19464, n_19465, n_19466, n_19467, n_19468, n_19469, n_19470, n_19471, n_19472, n_19473, n_19474, n_19475, n_19476, n_19477, n_19478, n_19479, n_19480, n_19481, n_19482, n_19483, n_19484, n_19485, n_19486, n_19487, n_19488, n_19489, n_19490, n_19491, n_19492, n_19493, n_19494, n_19495, n_19496, n_19497, n_19498, n_19499, n_19500, n_19501, n_19502, n_19503, n_19504, n_19505, n_19506, n_19507, n_19508, n_19509, n_19510, n_19511, n_19512, n_19513, n_19514, n_19515, n_19516, n_19517, n_19518, n_19519, n_19520, n_19521, n_19522, n_19523, n_19524, n_19525, n_19526, n_19527, n_19528, n_19529, n_19530, n_19531, n_19532, n_19533, n_19534, n_19535, n_19536, n_19537, n_19538, n_19539, n_19540, n_19541, n_19542, n_19543, n_19544, n_19545, n_19546, n_19547, n_19548, n_19549, n_19550, n_19551, n_19552, n_19553, n_19554, n_19555, n_19556, n_19557, n_19558, n_19559, n_19560, n_19561, n_19562, n_19563, n_19564, n_19565, n_19566, n_19567, n_19568, n_19569, n_19570, n_19571, n_19572, n_19573, n_19574, n_19575, n_19576, n_19577, n_19578, n_19579, n_19580, n_19581, n_19582, n_19583, n_19584, n_19585, n_19586, n_19587, n_19588, n_19589, n_19590, n_19591, n_19592, n_19593, n_19594, n_19595, n_19596, n_19597, n_19598, n_19599, n_19600, n_19601, n_19602, n_19603, n_19604, n_19605, n_19606, n_19607, n_19608, n_19609, n_19610, n_19611, n_19612, n_19613, n_19614, n_19615, n_19616, n_19617, n_19618, n_19619, n_19620, n_19621, n_19622, n_19623, n_19624, n_19625, n_19626, n_19627, n_19628, n_19629, n_19630, n_19631, n_19632, n_19633, n_19634, n_19635, n_19636, n_19637, n_19638, n_19639, n_19640, n_19641, n_19642, n_19643, n_19644, n_19645, n_19646, n_19647, n_19648, n_19649, n_19650, n_19651, n_19652, n_19653, n_19654, n_19655, n_19656, n_19657, n_19658, n_19659, n_19660, n_19661, n_19662, n_19663, n_19664, n_19665, n_19666, n_19667, n_19668, n_19669, n_19670, n_19671, n_19672, n_19673, n_19674, n_19675, n_19676, n_19677, n_19678, n_19679, n_19680, n_19681, n_19682, n_19683, n_19684, n_19685, n_19686, n_19687, n_19688, n_19689, n_19690, n_19691, n_19692, n_19693, n_19694, n_19695, n_19696, n_19697, n_19698, n_19699, n_19700, n_19701, n_19702, n_19703, n_19704, n_19705, n_19706, n_19707, n_19708, n_19709, n_19710, n_19711, n_19712, n_19713, n_19714, n_19715, n_19716, n_19717, n_19718, n_19719, n_19720, n_19721, n_19722, n_19723, n_19724, n_19725, n_19726, n_19727, n_19728, n_19729, n_19730, n_19731, n_19732, n_19733, n_19734, n_19735, n_19736, n_19737, n_19738, n_19739, n_19740, n_19741, n_19742, n_19743, n_19744, n_19745, n_19746, n_19747, n_19748, n_19749, n_19750, n_19751, n_19752, n_19753, n_19754, n_19755, n_19756, n_19757, n_19758, n_19759, n_19760, n_19761, n_19762, n_19763, n_19764, n_19765, n_19766, n_19767, n_19768, n_19769, n_19770, n_19771, n_19772, n_19773, n_19774, n_19775, n_19776, n_19777, n_19778, n_19779, n_19780, n_19781, n_19782, n_19783, n_19784, n_19785, n_19786, n_19787, n_19788, n_19789, n_19790, n_19791, n_19792, n_19793, n_19794, n_19795, n_19796, n_19797, n_19798, n_19799, n_19800, n_19801, n_19802, n_19803, n_19804, n_19805, n_19806, n_19807, n_19808, n_19809, n_19810, n_19811, n_19812, n_19813, n_19814, n_19815, n_19816, n_19817, n_19818, n_19819, n_19820, n_19821, n_19822, n_19823, n_19824, n_19825, n_19826, n_19827, n_19828, n_19829, n_19830, n_19831, n_19832, n_19833, n_19834, n_19835, n_19836, n_19837, n_19838, n_19839, n_19840, n_19841, n_19842, n_19843, n_19844, n_19845, n_19846, n_19847, n_19848, n_19849, n_19850, n_19851, n_19852, n_19853, n_19854, n_19855, n_19856, n_19857, n_19858, n_19859, n_19860, n_19861, n_19862, n_19863, n_19864, n_19865, n_19866, n_19867, n_19868, n_19869, n_19870, n_19871, n_19872, n_19873, n_19874, n_19875, n_19876, n_19877, n_19878, n_19879, n_19880, n_19881, n_19882, n_19883, n_19884, n_19885, n_19886, n_19887, n_19888, n_19889, n_19890, n_19891, n_19892, n_19893, n_19894, n_19895, n_19896, n_19897, n_19898, n_19899, n_19900, n_19901, n_19902, n_19903, n_19904, n_19905, n_19906, n_19907, n_19908, n_19909, n_19910, n_19911, n_19912, n_19913, n_19914, n_19915, n_19916, n_19917, n_19918, n_19919, n_19920, n_19921, n_19922, n_19923, n_19924, n_19925, n_19926, n_19927, n_19928, n_19929, n_19930, n_19931, n_19932, n_19933, n_19934, n_19935, n_19936, n_19937, n_19938, n_19939, n_19940, n_19941, n_19942, n_19943, n_19944, n_19945, n_19946, n_19947, n_19948, n_19949, n_19950, n_19951, n_19952, n_19953, n_19954, n_19955, n_19956, n_19957, n_19958, n_19959, n_19960, n_19961, n_19962, n_19963, n_19964, n_19965, n_19966, n_19967, n_19968, n_19969, n_19970, n_19971, n_19972, n_19973, n_19974, n_19975, n_19976, n_19977, n_19978, n_19979, n_19980, n_19981, n_19982, n_19983, n_19984, n_19985, n_19986, n_19987, n_19988, n_19989, n_19990, n_19991, n_19992, n_19993, n_19994, n_19995, n_19996, n_19997, n_19998, n_19999, n_20000, n_20001, n_20002, n_20003, n_20004, n_20005, n_20006, n_20007, n_20008, n_20009, n_20010, n_20011, n_20012, n_20013, n_20014, n_20015, n_20016, n_20017, n_20018, n_20019, n_20020, n_20021, n_20022, n_20023, n_20024, n_20025, n_20026, n_20027, n_20028, n_20029, n_20030, n_20031, n_20032, n_20033, n_20034, n_20035, n_20036, n_20037, n_20038, n_20039, n_20040, n_20041, n_20042, n_20043, n_20044, n_20045, n_20046, n_20047, n_20048, n_20049, n_20050, n_20051, n_20052, n_20053, n_20054, n_20055, n_20056, n_20057, n_20058, n_20059, n_20060, n_20061, n_20062, n_20063, n_20064, n_20065, n_20066, n_20067, n_20068, n_20069, n_20070, n_20071, n_20072, n_20073, n_20074, n_20075, n_20076, n_20077, n_20078, n_20079, n_20080, n_20081, n_20082, n_20083, n_20084, n_20085, n_20086, n_20087, n_20088, n_20089, n_20090, n_20091, n_20092, n_20093, n_20094, n_20095, n_20096, n_20097, n_20098, n_20099, n_20100, n_20101, n_20102, n_20103, n_20104, n_20105, n_20106, n_20107, n_20108, n_20109, n_20110, n_20111, n_20112, n_20113, n_20114, n_20115, n_20116, n_20117, n_20118, n_20119, n_20120, n_20121, n_20122, n_20123, n_20124, n_20125, n_20126, n_20127, n_20128, n_20129, n_20130, n_20131, n_20132, n_20133, n_20134, n_20135, n_20136, n_20137, n_20138, n_20139, n_20140, n_20141, n_20142, n_20143, n_20144, n_20145, n_20146, n_20147, n_20148, n_20149, n_20150, n_20151, n_20152, n_20153, n_20154, n_20155, n_20156, n_20157, n_20158, n_20159, n_20160, n_20161, n_20162, n_20163, n_20164, n_20165, n_20166, n_20167, n_20168, n_20169, n_20170, n_20171, n_20172, n_20173, n_20174, n_20175, n_20176, n_20177, n_20178, n_20179, n_20180, n_20181, n_20182, n_20183, n_20184, n_20185, n_20186, n_20187, n_20188, n_20189, n_20190, n_20191, n_20192, n_20193, n_20194, n_20195, n_20196, n_20197, n_20198, n_20199, n_20200, n_20201, n_20202, n_20203, n_20204, n_20205, n_20206, n_20207, n_20208, n_20209, n_20210, n_20211, n_20212, n_20213, n_20214, n_20215, n_20216, n_20217, n_20218, n_20219, n_20220, n_20221, n_20222, n_20223, n_20224, n_20225, n_20226, n_20227, n_20228, n_20229, n_20230, n_20231, n_20232, n_20233, n_20234, n_20235, n_20236, n_20237, n_20238, n_20239, n_20240, n_20241, n_20242, n_20243, n_20244, n_20245, n_20246, n_20247, n_20248, n_20249, n_20250, n_20251, n_20252, n_20253, n_20254, n_20255, n_20256, n_20257, n_20258, n_20259, n_20260, n_20261, n_20262, n_20263, n_20264, n_20265, n_20266, n_20267, n_20268, n_20269, n_20270, n_20271, n_20272, n_20273, n_20274, n_20275, n_20276, n_20277, n_20278, n_20279, n_20280, n_20281, n_20282, n_20283, n_20284, n_20285, n_20286, n_20287, n_20288, n_20289, n_20290, n_20291, n_20292, n_20293, n_20294, n_20295, n_20296, n_20297, n_20298, n_20299, n_20300, n_20301, n_20302, n_20303, n_20304, n_20305, n_20306, n_20307, n_20308, n_20309, n_20310, n_20311, n_20312, n_20313, n_20314, n_20315, n_20316, n_20317, n_20318, n_20319, n_20320, n_20321, n_20322, n_20323, n_20324, n_20325, n_20326, n_20327, n_20328, n_20329, n_20330, n_20331, n_20332, n_20333, n_20334, n_20335, n_20336, n_20337, n_20338, n_20339, n_20340, n_20341, n_20342, n_20343, n_20344, n_20345, n_20346, n_20347, n_20348, n_20349, n_20350, n_20351, n_20352, n_20353, n_20354, n_20355, n_20356, n_20357, n_20358, n_20359, n_20360, n_20361, n_20362, n_20363, n_20364, n_20365, n_20366, n_20367, n_20368, n_20369, n_20370, n_20371, n_20372, n_20373, n_20374, n_20375, n_20376, n_20377, n_20378, n_20379, n_20380, n_20381, n_20382, n_20383, n_20384, n_20385, n_20386, n_20387, n_20388, n_20389, n_20390, n_20391, n_20392, n_20393, n_20394, n_20395, n_20396, n_20397, n_20398, n_20399, n_20400, n_20401, n_20402, n_20403, n_20404, n_20405, n_20406, n_20407, n_20408, n_20409, n_20410, n_20411, n_20412, n_20413, n_20414, n_20415, n_20416, n_20417, n_20418, n_20419, n_20420, n_20421, n_20422, n_20423, n_20424, n_20425, n_20426, n_20427, n_20428, n_20429, n_20430, n_20431, n_20432, n_20433, n_20434, n_20435, n_20436, n_20437, n_20438, n_20439, n_20440, n_20441, n_20442, n_20443, n_20444, n_20445, n_20446, n_20447, n_20448, n_20449, n_20450, n_20451, n_20452, n_20453, n_20454, n_20455, n_20456, n_20457, n_20458, n_20459, n_20460, n_20461, n_20462, n_20463, n_20464, n_20465, n_20466, n_20467, n_20468, n_20469, n_20470, n_20471, n_20472, n_20473, n_20474, n_20475, n_20476, n_20477, n_20478, n_20479, n_20480, n_20481, n_20482, n_20483, n_20484, n_20485, n_20486, n_20487, n_20488, n_20489, n_20490, n_20491, n_20492, n_20493, n_20494, n_20495, n_20496, n_20497, n_20498, n_20499, n_20500, n_20501, n_20502, n_20503, n_20504, n_20505, n_20506, n_20507, n_20508, n_20509, n_20510, n_20511, n_20512, n_20513, n_20514, n_20515, n_20516, n_20517, n_20518, n_20519, n_20520, n_20521, n_20522, n_20523, n_20524, n_20525, n_20526, n_20527, n_20528, n_20529, n_20530, n_20531, n_20532, n_20533, n_20534, n_20535, n_20536, n_20537, n_20538, n_20539, n_20540, n_20541, n_20542, n_20543, n_20544, n_20545, n_20546, n_20547, n_20548, n_20549, n_20550, n_20551, n_20552, n_20553, n_20554, n_20555, n_20556, n_20557, n_20558, n_20559, n_20560, n_20561, n_20562, n_20563, n_20564, n_20565, n_20566, n_20567, n_20568, n_20569, n_20570, n_20571, n_20572, n_20573, n_20574, n_20575, n_20576, n_20577, n_20578, n_20579, n_20580, n_20581, n_20582, n_20583, n_20584, n_20585, n_20586, n_20587, n_20588, n_20589, n_20590, n_20591, n_20592, n_20593, n_20594, n_20595, n_20596, n_20597, n_20598, n_20599, n_20600, n_20601, n_20602, n_20603, n_20604, n_20605, n_20606, n_20607, n_20608, n_20609, n_20610, n_20611, n_20612, n_20613, n_20614, n_20615, n_20616, n_20617, n_20618, n_20619, n_20620, n_20621, n_20622, n_20623, n_20624, n_20625, n_20626, n_20627, n_20628, n_20629, n_20630, n_20631, n_20632, n_20633, n_20634, n_20635, n_20636, n_20637, n_20638, n_20639, n_20640, n_20641, n_20642, n_20643, n_20644, n_20645, n_20646, n_20647, n_20648, n_20649, n_20650, n_20651, n_20652, n_20653, n_20654, n_20655, n_20656, n_20657, n_20658, n_20659, n_20660, n_20661, n_20662, n_20663, n_20664, n_20665, n_20666, n_20667, n_20668, n_20669, n_20670, n_20671, n_20672, n_20673, n_20674, n_20675, n_20676, n_20677, n_20678, n_20679, n_20680, n_20681, n_20682, n_20683, n_20684, n_20685, n_20686, n_20687, n_20688, n_20689, n_20690, n_20691, n_20692, n_20693, n_20694, n_20695, n_20696, n_20697, n_20698, n_20699, n_20700, n_20701, n_20702, n_20703, n_20704, n_20705, n_20706, n_20707, n_20708, n_20709, n_20710, n_20711, n_20712, n_20713, n_20714, n_20715, n_20716, n_20717, n_20718, n_20719, n_20720, n_20721, n_20722, n_20723, n_20724, n_20725, n_20726, n_20727, n_20728, n_20729, n_20730, n_20731, n_20732, n_20733, n_20734, n_20735, n_20736, n_20737, n_20738, n_20739, n_20740, n_20741, n_20742, n_20743, n_20744, n_20745, n_20746, n_20747, n_20748, n_20749, n_20750, n_20751, n_20752, n_20753, n_20754, n_20755, n_20756, n_20757, n_20758, n_20759, n_20760, n_20761, n_20762, n_20763, n_20764, n_20765, n_20766, n_20767, n_20768, n_20769, n_20770, n_20771, n_20772, n_20773, n_20774, n_20775, n_20776, n_20777, n_20778, n_20779, n_20780, n_20781, n_20782, n_20783, n_20784, n_20785, n_20786, n_20787, n_20788, n_20789, n_20790, n_20791, n_20792, n_20793, n_20794, n_20795, n_20796, n_20797, n_20798, n_20799, n_20800, n_20801, n_20802, n_20803, n_20804, n_20805, n_20806, n_20807, n_20808, n_20809, n_20810, n_20811, n_20812, n_20813, n_20814, n_20815, n_20816, n_20817, n_20818, n_20819, n_20820, n_20821, n_20822, n_20823, n_20824, n_20825, n_20826, n_20827, n_20828, n_20829, n_20830, n_20831, n_20832, n_20833, n_20834, n_20835, n_20836, n_20837, n_20838, n_20839, n_20840, n_20841, n_20842, n_20843, n_20844, n_20845, n_20846, n_20847, n_20848, n_20849, n_20850, n_20851, n_20852, n_20853, n_20854, n_20855, n_20856, n_20857, n_20858, n_20859, n_20860, n_20861, n_20862, n_20863, n_20864, n_20865, n_20866, n_20867, n_20868, n_20869, n_20870, n_20871, n_20872, n_20873, n_20874, n_20875, n_20876, n_20877, n_20878, n_20879, n_20880, n_20881, n_20882, n_20883, n_20884, n_20885, n_20886, n_20887, n_20888, n_20889, n_20890, n_20891, n_20892, n_20893, n_20894, n_20895, n_20896, n_20897, n_20898, n_20899, n_20900, n_20901, n_20902, n_20903, n_20904, n_20905, n_20906, n_20907, n_20908, n_20909, n_20910, n_20911, n_20912, n_20913, n_20914, n_20915, n_20916, n_20917, n_20918, n_20919, n_20920, n_20921, n_20922, n_20923, n_20924, n_20925, n_20926, n_20927, n_20928, n_20929, n_20930, n_20931, n_20932, n_20933, n_20934, n_20935, n_20936, n_20937, n_20938, n_20939, n_20940, n_20941, n_20942, n_20943, n_20944, n_20945, n_20946, n_20947, n_20948, n_20949, n_20950, n_20951, n_20952, n_20953, n_20954, n_20955, n_20956, n_20957, n_20958, n_20959, n_20960, n_20961, n_20962, n_20963, n_20964, n_20965, n_20966, n_20967, n_20968, n_20969, n_20970, n_20971, n_20972, n_20973, n_20974, n_20975, n_20976, n_20977, n_20978, n_20979, n_20980, n_20981, n_20982, n_20983, n_20984, n_20985, n_20986, n_20987, n_20988, n_20989, n_20990, n_20991, n_20992, n_20993, n_20994, n_20995, n_20996, n_20997, n_20998, n_20999, n_21000, n_21001, n_21002, n_21003, n_21004, n_21005, n_21006, n_21007, n_21008, n_21009, n_21010, n_21011, n_21012, n_21013, n_21014, n_21015, n_21016, n_21017, n_21018, n_21019, n_21020, n_21021, n_21022, n_21023, n_21024, n_21025, n_21026, n_21027, n_21028, n_21029, n_21030, n_21031, n_21032, n_21033, n_21034, n_21035, n_21036, n_21037, n_21038, n_21039, n_21040, n_21041, n_21042, n_21043, n_21044, n_21045, n_21046, n_21047, n_21048, n_21049, n_21050, n_21051, n_21052, n_21053, n_21054, n_21055, n_21056, n_21057, n_21058, n_21059, n_21060, n_21061, n_21062, n_21063, n_21064, n_21065, n_21066, n_21067, n_21068, n_21069, n_21070, n_21071, n_21072, n_21073, n_21074, n_21075, n_21076, n_21077, n_21078, n_21079, n_21080, n_21081, n_21082, n_21083, n_21084, n_21085, n_21086, n_21087, n_21088, n_21089, n_21090, n_21091, n_21092, n_21093, n_21094, n_21095, n_21096, n_21097, n_21098, n_21099, n_21100, n_21101, n_21102, n_21103, n_21104, n_21105, n_21106, n_21107, n_21108, n_21109, n_21110, n_21111, n_21112, n_21113, n_21114, n_21115, n_21116, n_21117, n_21118, n_21119, n_21120, n_21121, n_21122, n_21123, n_21124, n_21125, n_21126, n_21127, n_21128, n_21129, n_21130, n_21131, n_21132, n_21133, n_21134, n_21135, n_21136, n_21137, n_21138, n_21139, n_21140, n_21141, n_21142, n_21143, n_21144, n_21145, n_21146, n_21147, n_21148, n_21149, n_21150, n_21151, n_21152, n_21153, n_21154, n_21155, n_21156, n_21157, n_21158, n_21159, n_21160, n_21161, n_21162, n_21163, n_21164, n_21165, n_21166, n_21167, n_21168, n_21169, n_21170, n_21171, n_21172, n_21173, n_21174, n_21175, n_21176, n_21177, n_21178, n_21179, n_21180, n_21181, n_21182, n_21183, n_21184, n_21185, n_21186, n_21187, n_21188, n_21189, n_21190, n_21191, n_21192, n_21193, n_21194, n_21195, n_21196, n_21197, n_21198, n_21199, n_21200, n_21201, n_21202, n_21203, n_21204, n_21205, n_21206, n_21207, n_21208, n_21209, n_21210, n_21211, n_21212, n_21213, n_21214, n_21215, n_21216, n_21217, n_21218, n_21219, n_21220, n_21221, n_21222, n_21223, n_21224, n_21225, n_21226, n_21227, n_21228, n_21229, n_21230, n_21231, n_21232, n_21233, n_21234, n_21235, n_21236, n_21237, n_21238, n_21239, n_21240, n_21241, n_21242, n_21243, n_21244, n_21245, n_21246, n_21247, n_21248, n_21249, n_21250, n_21251, n_21252, n_21253, n_21254, n_21255, n_21256, n_21257, n_21258, n_21259, n_21260, n_21261, n_21262, n_21263, n_21264, n_21265, n_21266, n_21267, n_21268, n_21269, n_21270, n_21271, n_21272, n_21273, n_21274, n_21275, n_21276, n_21277, n_21278, n_21279, n_21280, n_21281, n_21282, n_21283, n_21284, n_21285, n_21286, n_21287, n_21288, n_21289, n_21290, n_21291, n_21292, n_21293, n_21294, n_21295, n_21296, n_21297, n_21298, n_21299, n_21300, n_21301, n_21302, n_21303, n_21304, n_21305, n_21306, n_21307, n_21308, n_21309, n_21310, n_21311, n_21312, n_21313, n_21314, n_21315, n_21316, n_21317, n_21318, n_21319, n_21320, n_21321, n_21322, n_21323, n_21324, n_21325, n_21326, n_21327, n_21328, n_21329, n_21330, n_21331, n_21332, n_21333, n_21334, n_21335, n_21336, n_21337, n_21338, n_21339, n_21340, n_21341, n_21342, n_21343, n_21344, n_21345, n_21346, n_21347, n_21348, n_21349, n_21350, n_21351, n_21352, n_21353, n_21354, n_21355, n_21356, n_21357, n_21358, n_21359, n_21360, n_21361, n_21362, n_21363, n_21364, n_21365, n_21366, n_21367, n_21368, n_21369, n_21370, n_21371, n_21372, n_21373, n_21374, n_21375, n_21376, n_21377, n_21378, n_21379, n_21380, n_21381, n_21382, n_21383, n_21384, n_21385, n_21386, n_21387, n_21388, n_21389, n_21390, n_21391, n_21392, n_21393, n_21394, n_21395, n_21396, n_21397, n_21398, n_21399, n_21400, n_21401, n_21402, n_21403, n_21404, n_21405, n_21406, n_21407, n_21408, n_21409, n_21410, n_21411, n_21412, n_21413, n_21414, n_21415, n_21416, n_21417, n_21418, n_21419, n_21420, n_21421, n_21422, n_21423, n_21424, n_21425, n_21426, n_21427, n_21428, n_21429, n_21430, n_21431, n_21432, n_21433, n_21434, n_21435, n_21436, n_21437, n_21438, n_21439, n_21440, n_21441, n_21442, n_21443, n_21444, n_21445, n_21446, n_21447, n_21448, n_21449, n_21450, n_21451, n_21452, n_21453, n_21454, n_21455, n_21456, n_21457, n_21458, n_21459, n_21460, n_21461, n_21462, n_21463, n_21464, n_21465, n_21466, n_21467, n_21468, n_21469, n_21470, n_21471, n_21472, n_21473, n_21474, n_21475, n_21476, n_21477, n_21478, n_21479, n_21480, n_21481, n_21482, n_21483, n_21484, n_21485, n_21486, n_21487, n_21488, n_21489, n_21490, n_21491, n_21492, n_21493, n_21494, n_21495, n_21496, n_21497, n_21498, n_21499, n_21500, n_21501, n_21502, n_21503, n_21504, n_21505, n_21506, n_21507, n_21508, n_21509, n_21510, n_21511, n_21512, n_21513, n_21514, n_21515, n_21516, n_21517, n_21518, n_21519, n_21520, n_21521, n_21522, n_21523, n_21524, n_21525, n_21526, n_21527, n_21528, n_21529, n_21530, n_21531, n_21532, n_21533, n_21534, n_21535, n_21536, n_21537, n_21538, n_21539, n_21540, n_21541, n_21542, n_21543, n_21544, n_21545, n_21546, n_21547, n_21548, n_21549, n_21550, n_21551, n_21552, n_21553, n_21554, n_21555, n_21556, n_21557, n_21558, n_21559, n_21560, n_21561, n_21562, n_21563, n_21564, n_21565, n_21566, n_21567, n_21568, n_21569, n_21570, n_21571, n_21572, n_21573, n_21574, n_21575, n_21576, n_21577, n_21578, n_21579, n_21580, n_21581, n_21582, n_21583, n_21584, n_21585, n_21586, n_21587, n_21588, n_21589, n_21590, n_21591, n_21592, n_21593, n_21594, n_21595, n_21596, n_21597, n_21598, n_21599, n_21600, n_21601, n_21602, n_21603, n_21604, n_21605, n_21606, n_21607, n_21608, n_21609, n_21610, n_21611, n_21612, n_21613, n_21614, n_21615, n_21616, n_21617, n_21618, n_21619, n_21620, n_21621, n_21622, n_21623, n_21624, n_21625, n_21626, n_21627, n_21628, n_21629, n_21630, n_21631, n_21632, n_21633, n_21634, n_21635, n_21636, n_21637, n_21638, n_21639, n_21640, n_21641, n_21642, n_21643, n_21644, n_21645, n_21646, n_21647, n_21648, n_21649, n_21650, n_21651, n_21652, n_21653, n_21654, n_21655, n_21656, n_21657, n_21658, n_21659, n_21660, n_21661, n_21662, n_21663, n_21664, n_21665, n_21666, n_21667, n_21668, n_21669, n_21670, n_21671, n_21672, n_21673, n_21674, n_21675, n_21676, n_21677, n_21678, n_21679, n_21680, n_21681, n_21682, n_21683, n_21684, n_21685, n_21686, n_21687, n_21688, n_21689, n_21690, n_21691, n_21692, n_21693, n_21694, n_21695, n_21696, n_21697, n_21698, n_21699, n_21700, n_21701, n_21702, n_21703, n_21704, n_21705, n_21706, n_21707, n_21708, n_21709, n_21710, n_21711, n_21712, n_21713, n_21714, n_21715, n_21716, n_21717, n_21718, n_21719, n_21720, n_21721, n_21722, n_21723, n_21724, n_21725, n_21726, n_21727, n_21728, n_21729, n_21730, n_21731, n_21732, n_21733, n_21734, n_21735, n_21736, n_21737, n_21738, n_21739, n_21740, n_21741, n_21742, n_21743, n_21744, n_21745, n_21746, n_21747, n_21748, n_21749, n_21750, n_21751, n_21752, n_21753, n_21754, n_21755, n_21756, n_21757, n_21758, n_21759, n_21760, n_21761, n_21762, n_21763, n_21764, n_21765, n_21766, n_21767, n_21768, n_21769, n_21770, n_21771, n_21772, n_21773, n_21774, n_21775, n_21776, n_21777, n_21778, n_21779, n_21780, n_21781, n_21782, n_21783, n_21784, n_21785, n_21786, n_21787, n_21788, n_21789, n_21790, n_21791, n_21792, n_21793, n_21794, n_21795, n_21796, n_21797, n_21798, n_21799, n_21800, n_21801, n_21802, n_21803, n_21804, n_21805, n_21806, n_21807, n_21808, n_21809, n_21810, n_21811, n_21812, n_21813, n_21814, n_21815, n_21816, n_21817, n_21818, n_21819, n_21820, n_21821, n_21822, n_21823, n_21824, n_21825, n_21826, n_21827, n_21828, n_21829, n_21830, n_21831, n_21832, n_21833, n_21834, n_21835, n_21836, n_21837, n_21838, n_21839, n_21840, n_21841, n_21842, n_21843, n_21844, n_21845, n_21846, n_21847, n_21848, n_21849, n_21850, n_21851, n_21852, n_21853, n_21854, n_21855, n_21856, n_21857, n_21858, n_21859, n_21860, n_21861, n_21862, n_21863, n_21864, n_21865, n_21866, n_21867, n_21868, n_21869, n_21870, n_21871, n_21872, n_21873, n_21874, n_21875, n_21876, n_21877, n_21878, n_21879, n_21880, n_21881, n_21882, n_21883, n_21884, n_21885, n_21886, n_21887, n_21888, n_21889, n_21890, n_21891, n_21892, n_21893, n_21894, n_21895, n_21896, n_21897, n_21898, n_21899, n_21900, n_21901, n_21902, n_21903, n_21904, n_21905, n_21906, n_21907, n_21908, n_21909, n_21910, n_21911, n_21912, n_21913, n_21914, n_21915, n_21916, n_21917, n_21918, n_21919, n_21920, n_21921, n_21922, n_21923, n_21924, n_21925, n_21926, n_21927, n_21928, n_21929, n_21930, n_21931, n_21932, n_21933, n_21934, n_21935, n_21936, n_21937, n_21938, n_21939, n_21940, n_21941, n_21942, n_21943, n_21944, n_21945, n_21946, n_21947, n_21948, n_21949, n_21950, n_21951, n_21952, n_21953, n_21954, n_21955, n_21956, n_21957, n_21958, n_21959, n_21960, n_21961, n_21962, n_21963, n_21964, n_21965, n_21966, n_21967, n_21968, n_21969, n_21970, n_21971, n_21972, n_21973, n_21974, n_21975, n_21976, n_21977, n_21978, n_21979, n_21980, n_21981, n_21982, n_21983, n_21984, n_21985, n_21986, n_21987, n_21988, n_21989, n_21990, n_21991, n_21992, n_21993, n_21994, n_21995, n_21996, n_21997, n_21998, n_21999, n_22000, n_22001, n_22002, n_22003, n_22004, n_22005, n_22006, n_22007, n_22008, n_22009, n_22010, n_22011, n_22012, n_22013, n_22014, n_22015, n_22016, n_22017, n_22018, n_22019, n_22020, n_22021, n_22022, n_22023, n_22024, n_22025, n_22026, n_22027, n_22028, n_22029, n_22030, n_22031, n_22032, n_22033, n_22034, n_22035, n_22036, n_22037, n_22038, n_22039, n_22040, n_22041, n_22042, n_22043, n_22044, n_22045, n_22046, n_22047, n_22048, n_22049, n_22050, n_22051, n_22052, n_22053, n_22054, n_22055, n_22056, n_22057, n_22058, n_22059, n_22060, n_22061, n_22062, n_22063, n_22064, n_22065, n_22066, n_22067, n_22068, n_22069, n_22070, n_22071, n_22072, n_22073, n_22074, n_22075, n_22076, n_22077, n_22078, n_22079, n_22080, n_22081, n_22082, n_22083, n_22084, n_22085, n_22086, n_22087, n_22088, n_22089, n_22090, n_22091, n_22092, n_22093, n_22094, n_22095, n_22096, n_22097, n_22098, n_22099, n_22100, n_22101, n_22102, n_22103, n_22104, n_22105, n_22106, n_22107, n_22108, n_22109, n_22110, n_22111, n_22112, n_22113, n_22114, n_22115, n_22116, n_22117, n_22118, n_22119, n_22120, n_22121, n_22122, n_22123, n_22124, n_22125, n_22126, n_22127, n_22128, n_22129, n_22130, n_22131, n_22132, n_22133, n_22134, n_22135, n_22136, n_22137, n_22138, n_22139, n_22140, n_22141, n_22142, n_22143, n_22144, n_22145, n_22146, n_22147, n_22148, n_22149, n_22150, n_22151, n_22152, n_22153, n_22154, n_22155, n_22156, n_22157, n_22158, n_22159, n_22160, n_22161, n_22162, n_22163, n_22164, n_22165, n_22166, n_22167, n_22168, n_22169, n_22170, n_22171, n_22172, n_22173, n_22174, n_22175, n_22176, n_22177, n_22178, n_22179, n_22180, n_22181, n_22182, n_22183, n_22184, n_22185, n_22186, n_22187, n_22188, n_22189, n_22190, n_22191, n_22192, n_22193, n_22194, n_22195, n_22196, n_22197, n_22198, n_22199, n_22200, n_22201, n_22202, n_22203, n_22204, n_22205, n_22206, n_22207, n_22208, n_22209, n_22210, n_22211, n_22212, n_22213, n_22214, n_22215, n_22216, n_22217, n_22218, n_22219, n_22220, n_22221, n_22222, n_22223, n_22224, n_22225, n_22226, n_22227, n_22228, n_22229, n_22230, n_22231, n_22232, n_22233, n_22234, n_22235, n_22236, n_22237, n_22238, n_22239, n_22240, n_22241, n_22242, n_22243, n_22244, n_22245, n_22246, n_22247, n_22248, n_22249, n_22250, n_22251, n_22252, n_22253, n_22254, n_22255, n_22256, n_22257, n_22258, n_22259, n_22260, n_22261, n_22262, n_22263, n_22264, n_22265, n_22266, n_22267, n_22268, n_22269, n_22270, n_22271, n_22272, n_22273, n_22274, n_22275, n_22276, n_22277, n_22278, n_22279, n_22280, n_22281, n_22282, n_22283, n_22284, n_22285, n_22286, n_22287, n_22288, n_22289, n_22290, n_22291, n_22292, n_22293, n_22294, n_22295, n_22296, n_22297, n_22298, n_22299, n_22300, n_22301, n_22302, n_22303, n_22304, n_22305, n_22306, n_22307, n_22308, n_22309, n_22310, n_22311, n_22312, n_22313, n_22314, n_22315, n_22316, n_22317, n_22318, n_22319, n_22320, n_22321, n_22322, n_22323, n_22324, n_22325, n_22326, n_22327, n_22328, n_22329, n_22330, n_22331, n_22332, n_22333, n_22334, n_22335, n_22336, n_22337, n_22338, n_22339, n_22340, n_22341, n_22342, n_22343, n_22344, n_22345, n_22346, n_22347, n_22348, n_22349, n_22350, n_22351, n_22352, n_22353, n_22354, n_22355, n_22356, n_22357, n_22358, n_22359, n_22360, n_22361, n_22362, n_22363, n_22364, n_22365, n_22366, n_22367, n_22368, n_22369, n_22370, n_22371, n_22372, n_22373, n_22374, n_22375, n_22376, n_22377, n_22378, n_22379, n_22380, n_22381, n_22382, n_22383, n_22384, n_22385, n_22386, n_22387, n_22388, n_22389, n_22390, n_22391, n_22392, n_22393, n_22394, n_22395, n_22396, n_22397, n_22398, n_22399, n_22400, n_22401, n_22402, n_22403, n_22404, n_22405, n_22406, n_22407, n_22408, n_22409, n_22410, n_22411, n_22412, n_22413, n_22414, n_22415, n_22416, n_22417, n_22418, n_22419, n_22420, n_22421, n_22422, n_22423, n_22424, n_22425, n_22426, n_22427, n_22428, n_22429, n_22430, n_22431, n_22432, n_22433, n_22434, n_22435, n_22436, n_22437, n_22438, n_22439, n_22440, n_22441, n_22442, n_22443, n_22444, n_22445, n_22446, n_22447, n_22448, n_22449, n_22450, n_22451, n_22452, n_22453, n_22454, n_22455, n_22456, n_22457, n_22458, n_22459, n_22460, n_22461, n_22462, n_22463, n_22464, n_22465, n_22466, n_22467, n_22468, n_22469, n_22470, n_22471, n_22472, n_22473, n_22474, n_22475, n_22476, n_22477, n_22478, n_22479, n_22480, n_22481, n_22482, n_22483, n_22484, n_22485, n_22486, n_22487, n_22488, n_22489, n_22490, n_22491, n_22492, n_22493, n_22494, n_22495, n_22496, n_22497, n_22498, n_22499, n_22500, n_22501, n_22502, n_22503, n_22504, n_22505, n_22506, n_22507, n_22508, n_22509, n_22510, n_22511, n_22512, n_22513, n_22514, n_22515, n_22516, n_22517, n_22518, n_22519, n_22520, n_22521, n_22522, n_22523, n_22524, n_22525, n_22526, n_22527, n_22528, n_22529, n_22530, n_22531, n_22532, n_22533, n_22534, n_22535, n_22536, n_22537, n_22538, n_22539, n_22540, n_22541, n_22542, n_22543, n_22544, n_22545, n_22546, n_22547, n_22548, n_22549, n_22550, n_22551, n_22552, n_22553, n_22554, n_22555, n_22556, n_22557, n_22558, n_22559, n_22560, n_22561, n_22562, n_22563, n_22564, n_22565, n_22566, n_22567, n_22568, n_22569, n_22570, n_22571, n_22572, n_22573, n_22574, n_22575, n_22576, n_22577, n_22578, n_22579, n_22580, n_22581, n_22582, n_22583, n_22584, n_22585, n_22586, n_22587, n_22588, n_22589, n_22590, n_22591, n_22592, n_22593, n_22594, n_22595, n_22596, n_22597, n_22598, n_22599, n_22600, n_22601, n_22602, n_22603, n_22604, n_22605, n_22606, n_22607, n_22608, n_22609, n_22610, n_22611, n_22612, n_22613, n_22614, n_22615, n_22616, n_22617, n_22618, n_22619, n_22620, n_22621, n_22622, n_22623, n_22624, n_22625, n_22626, n_22627, n_22628, n_22629, n_22630, n_22631, n_22632, n_22633, n_22634, n_22635, n_22636, n_22637, n_22638, n_22639, n_22640, n_22641, n_22642, n_22643, n_22644, n_22645, n_22646, n_22647, n_22648, n_22649, n_22650, n_22651, n_22652, n_22653, n_22654, n_22655, n_22656, n_22657, n_22658, n_22659, n_22660, n_22661, n_22662, n_22663, n_22664, n_22665, n_22666, n_22667, n_22668, n_22669, n_22670, n_22671, n_22672, n_22673, n_22674, n_22675, n_22676, n_22677, n_22678, n_22679, n_22680, n_22681, n_22682, n_22683, n_22684, n_22685, n_22686, n_22687, n_22688, n_22689, n_22690, n_22691, n_22692, n_22693, n_22694, n_22695, n_22696, n_22697, n_22698, n_22699, n_22700, n_22701, n_22702, n_22703, n_22704, n_22705, n_22706, n_22707, n_22708, n_22709, n_22710, n_22711, n_22712, n_22713, n_22714, n_22715, n_22716, n_22717, n_22718, n_22719, n_22720, n_22721, n_22722, n_22723, n_22724, n_22725, n_22726, n_22727, n_22728, n_22729, n_22730, n_22731, n_22732, n_22733, n_22734, n_22735, n_22736, n_22737, n_22738, n_22739, n_22740, n_22741, n_22742, n_22743, n_22744, n_22745, n_22746, n_22747, n_22748, n_22749, n_22750, n_22751, n_22752, n_22753, n_22754, n_22755, n_22756, n_22757, n_22758, n_22759, n_22760, n_22761, n_22762, n_22763, n_22764, n_22765, n_22766, n_22767, n_22768, n_22769, n_22770, n_22771, n_22772, n_22773, n_22774, n_22775, n_22776, n_22777, n_22778, n_22779, n_22780, n_22781, n_22782, n_22783, n_22784, n_22785, n_22786, n_22787, n_22788, n_22789, n_22790, n_22791, n_22792, n_22793, n_22794, n_22795, n_22796, n_22797, n_22798, n_22799, n_22800, n_22801, n_22802, n_22803, n_22804, n_22805, n_22806, n_22807, n_22808, n_22809, n_22810, n_22811, n_22812, n_22813, n_22814, n_22815, n_22816, n_22817, n_22818, n_22819, n_22820, n_22821, n_22822, n_22823, n_22824, n_22825, n_22826, n_22827, n_22828, n_22829, n_22830, n_22831, n_22832, n_22833, n_22834, n_22835, n_22836, n_22837, n_22838, n_22839, n_22840, n_22841, n_22842, n_22843, n_22844, n_22845, n_22846, n_22847, n_22848, n_22849, n_22850, n_22851, n_22852, n_22853, n_22854, n_22855, n_22856, n_22857, n_22858, n_22859, n_22860, n_22861, n_22862, n_22863, n_22864, n_22865, n_22866, n_22867, n_22868, n_22869, n_22870, n_22871, n_22872, n_22873, n_22874, n_22875, n_22876, n_22877, n_22878, n_22879, n_22880, n_22881, n_22882, n_22883, n_22884, n_22885, n_22886, n_22887, n_22888, n_22889, n_22890, n_22891, n_22892, n_22893, n_22894, n_22895, n_22896, n_22897, n_22898, n_22899, n_22900, n_22901, n_22902, n_22903, n_22904, n_22905, n_22906, n_22907, n_22908, n_22909, n_22910, n_22911, n_22912, n_22913, n_22914, n_22915, n_22916, n_22917, n_22918, n_22919, n_22920, n_22921, n_22922, n_22923, n_22924, n_22925, n_22926, n_22927, n_22928, n_22929, n_22930, n_22931, n_22932, n_22933, n_22934, n_22935, n_22936, n_22937, n_22938, n_22939, n_22940, n_22941, n_22942, n_22943, n_22944, n_22945, n_22946, n_22947, n_22948, n_22949, n_22950, n_22951, n_22952, n_22953, n_22954, n_22955, n_22956, n_22957, n_22958, n_22959, n_22960, n_22961, n_22962, n_22963, n_22964, n_22965, n_22966, n_22967, n_22968, n_22969, n_22970, n_22971, n_22972, n_22973, n_22974, n_22975, n_22976, n_22977, n_22978, n_22979, n_22980, n_22981, n_22982, n_22983, n_22984, n_22985, n_22986, n_22987, n_22988, n_22989, n_22990, n_22991, n_22992, n_22993, n_22994, n_22995, n_22996, n_22997, n_22998, n_22999, n_23000, n_23001, n_23002, n_23003, n_23004, n_23005, n_23006, n_23007, n_23008, n_23009, n_23010, n_23011, n_23012, n_23013, n_23014, n_23015, n_23016, n_23017, n_23018, n_23019, n_23020, n_23021, n_23022, n_23023, n_23024, n_23025, n_23026, n_23027, n_23028, n_23029, n_23030, n_23031, n_23032, n_23033, n_23034, n_23035, n_23036, n_23037, n_23038, n_23039, n_23040, n_23041, n_23042, n_23043, n_23044, n_23045, n_23046, n_23047, n_23048, n_23049, n_23050, n_23051, n_23052, n_23053, n_23054, n_23055, n_23056, n_23057, n_23058, n_23059, n_23060, n_23061, n_23062, n_23063, n_23064, n_23065, n_23066, n_23067, n_23068, n_23069, n_23070, n_23071, n_23072, n_23073, n_23074, n_23075, n_23076, n_23077, n_23078, n_23079, n_23080, n_23081, n_23082, n_23083, n_23084, n_23085, n_23086, n_23087, n_23088, n_23089, n_23090, n_23091, n_23092, n_23093, n_23094, n_23095, n_23096, n_23097, n_23098, n_23099, n_23100, n_23101, n_23102, n_23103, n_23104, n_23105, n_23106, n_23107, n_23108, n_23109, n_23110, n_23111, n_23112, n_23113, n_23114, n_23115, n_23116, n_23117, n_23118, n_23119, n_23120, n_23121, n_23122, n_23123, n_23124, n_23125, n_23126, n_23127, n_23128, n_23129, n_23130, n_23131, n_23132, n_23133, n_23134, n_23135, n_23136, n_23137, n_23138, n_23139, n_23140, n_23141, n_23142, n_23143, n_23144, n_23145, n_23146, n_23147, n_23148, n_23149, n_23150, n_23151, n_23152, n_23153, n_23154, n_23155, n_23156, n_23157, n_23158, n_23159, n_23160, n_23161, n_23162, n_23163, n_23164, n_23165, n_23166, n_23167, n_23168, n_23169, n_23170, n_23171, n_23172, n_23173, n_23174, n_23175, n_23176, n_23177, n_23178, n_23179, n_23180, n_23181, n_23182, n_23183, n_23184, n_23185, n_23186, n_23187, n_23188, n_23189, n_23190, n_23191, n_23192, n_23193, n_23194, n_23195, n_23196, n_23197, n_23198, n_23199, n_23200, n_23201, n_23202, n_23203, n_23204, n_23205, n_23206, n_23207, n_23208, n_23209, n_23210, n_23211, n_23212, n_23213, n_23214, n_23215, n_23216, n_23217, n_23218, n_23219, n_23220, n_23221, n_23222, n_23223, n_23224, n_23225, n_23226, n_23227, n_23228, n_23229, n_23230, n_23231, n_23232, n_23233, n_23234, n_23235, n_23236, n_23237, n_23238, n_23239, n_23240, n_23241, n_23242, n_23243, n_23244, n_23245, n_23246, n_23247, n_23248, n_23249, n_23250, n_23251, n_23252, n_23253, n_23254, n_23255, n_23256, n_23257, n_23258, n_23259, n_23260, n_23261, n_23262, n_23263, n_23264, n_23265, n_23266, n_23267, n_23268, n_23269, n_23270, n_23271, n_23272, n_23273, n_23274, n_23275, n_23276, n_23277, n_23278, n_23279, n_23280, n_23281, n_23282, n_23283, n_23284, n_23285, n_23286, n_23287, n_23288, n_23289, n_23290, n_23291, n_23292, n_23293, n_23294, n_23295, n_23296, n_23297, n_23298, n_23299, n_23300, n_23301, n_23302, n_23303, n_23304, n_23305, n_23306, n_23307, n_23308, n_23309, n_23310, n_23311, n_23312, n_23313, n_23314, n_23315, n_23316, n_23317, n_23318, n_23319, n_23320, n_23321, n_23322, n_23323, n_23324, n_23325, n_23326, n_23327, n_23328, n_23329, n_23330, n_23331, n_23332, n_23333, n_23334, n_23335, n_23336, n_23337, n_23338, n_23339, n_23340, n_23341, n_23342, n_23343, n_23344, n_23345, n_23346, n_23347, n_23348, n_23349, n_23350, n_23351, n_23352, n_23353, n_23354, n_23355, n_23356, n_23357, n_23358, n_23359, n_23360, n_23361, n_23362, n_23363, n_23364, n_23365, n_23366, n_23367, n_23368, n_23369, n_23370, n_23371, n_23372, n_23373, n_23374, n_23375, n_23376, n_23377, n_23378, n_23379, n_23380, n_23381, n_23382, n_23383, n_23384, n_23385, n_23386, n_23387, n_23388, n_23389, n_23390, n_23391, n_23392, n_23393, n_23394, n_23395, n_23396, n_23397, n_23398, n_23399, n_23400, n_23401, n_23402, n_23403, n_23404, n_23405, n_23406, n_23407, n_23408, n_23409, n_23410, n_23411, n_23412, n_23413, n_23414, n_23415, n_23416, n_23417, n_23418, n_23419, n_23420, n_23421, n_23422, n_23423, n_23424, n_23425, n_23426, n_23427, n_23428, n_23429, n_23430, n_23431, n_23432, n_23433, n_23434, n_23435, n_23436, n_23437, n_23438, n_23439, n_23440, n_23441, n_23442, n_23443, n_23444, n_23445, n_23446, n_23447, n_23448, n_23449, n_23450, n_23451, n_23452, n_23453, n_23454, n_23455, n_23456, n_23457, n_23458, n_23459, n_23460, n_23461, n_23462, n_23463, n_23464, n_23465, n_23466, n_23467, n_23468, n_23469, n_23470, n_23471, n_23472, n_23473, n_23474, n_23475, n_23476, n_23477, n_23478, n_23479, n_23480, n_23481, n_23482, n_23483, n_23484, n_23485, n_23486, n_23487, n_23488, n_23489, n_23490, n_23491, n_23492, n_23493, n_23494, n_23495, n_23496, n_23497, n_23498, n_23499, n_23500, n_23501, n_23502, n_23503, n_23504, n_23505, n_23506, n_23507, n_23508, n_23509, n_23510, n_23511, n_23512, n_23513, n_23514, n_23515, n_23516, n_23517, n_23518, n_23519, n_23520, n_23521, n_23522, n_23523, n_23524, n_23525, n_23526, n_23527, n_23528, n_23529, n_23530, n_23531, n_23532, n_23533, n_23534, n_23535, n_23536, n_23537, n_23538, n_23539, n_23540, n_23541, n_23542, n_23543, n_23544, n_23545, n_23546, n_23547, n_23548, n_23549, n_23550, n_23551, n_23552, n_23553, n_23554, n_23555, n_23556, n_23557, n_23558, n_23559, n_23560, n_23561, n_23562, n_23563, n_23564, n_23565, n_23566, n_23567, n_23568, n_23569, n_23570, n_23571, n_23572, n_23573, n_23574, n_23575, n_23576, n_23577, n_23578, n_23579, n_23580, n_23581, n_23582, n_23583, n_23584, n_23585, n_23586, n_23587, n_23588, n_23589, n_23590, n_23591, n_23592, n_23593, n_23594, n_23595, n_23596, n_23597, n_23598, n_23599, n_23600, n_23601, n_23602, n_23603, n_23604, n_23605, n_23606, n_23607, n_23608, n_23609, n_23610, n_23611, n_23612, n_23613, n_23614, n_23615, n_23616, n_23617, n_23618, n_23619, n_23620, n_23621, n_23622, n_23623, n_23624, n_23625, n_23626, n_23627, n_23628, n_23629, n_23630, n_23631, n_23632, n_23633, n_23634, n_23635, n_23636, n_23637, n_23638, n_23639, n_23640, n_23641, n_23642, n_23643, n_23644, n_23645, n_23646, n_23647, n_23648, n_23649, n_23650, n_23651, n_23652, n_23653, n_23654, n_23655, n_23656, n_23657, n_23658, n_23659, n_23660, n_23661, n_23662, n_23663, n_23664, n_23665, n_23666, n_23667, n_23668, n_23669, n_23670, n_23671, n_23672, n_23673, n_23674, n_23675, n_23676, n_23677, n_23678, n_23679, n_23680, n_23681, n_23682, n_23683, n_23684, n_23685, n_23686, n_23687, n_23688, n_23689, n_23690, n_23691, n_23692, n_23693, n_23694, n_23695, n_23696, n_23697, n_23698, n_23699, n_23700, n_23701, n_23702, n_23703, n_23704, n_23705, n_23706, n_23707, n_23708, n_23709, n_23710, n_23711, n_23712, n_23713, n_23714, n_23715, n_23716, n_23717, n_23718, n_23719, n_23720, n_23721, n_23722, n_23723, n_23724, n_23725, n_23726, n_23727, n_23728, n_23729, n_23730, n_23731, n_23732, n_23733, n_23734, n_23735, n_23736, n_23737, n_23738, n_23739, n_23740, n_23741, n_23742, n_23743, n_23744, n_23745, n_23746, n_23747, n_23748, n_23749, n_23750, n_23751, n_23752, n_23753, n_23754, n_23755, n_23756, n_23757, n_23758, n_23759, n_23760, n_23761, n_23762, n_23763, n_23764, n_23765, n_23766, n_23767, n_23768, n_23769, n_23770, n_23771, n_23772, n_23773, n_23774, n_23775, n_23776, n_23777, n_23778, n_23779, n_23780, n_23781, n_23782, n_23783, n_23784, n_23785, n_23786, n_23787, n_23788, n_23789, n_23790, n_23791, n_23792, n_23793, n_23794, n_23795, n_23796, n_23797, n_23798, n_23799, n_23800, n_23801, n_23802, n_23803, n_23804, n_23805, n_23806, n_23807, n_23808, n_23809, n_23810, n_23811, n_23812, n_23813, n_23814, n_23815, n_23816, n_23817, n_23818, n_23819, n_23820, n_23821, n_23822, n_23823, n_23824, n_23825, n_23826, n_23827, n_23828, n_23829, n_23830, n_23831, n_23832, n_23833, n_23834, n_23835, n_23836, n_23837, n_23838, n_23839, n_23840, n_23841, n_23842, n_23843, n_23844, n_23845, n_23846, n_23847, n_23848, n_23849, n_23850, n_23851, n_23852, n_23853, n_23854, n_23855, n_23856, n_23857, n_23858, n_23859, n_23860, n_23861, n_23862, n_23863, n_23864, n_23865, n_23866, n_23867, n_23868, n_23869, n_23870, n_23871, n_23872, n_23873, n_23874, n_23875, n_23876, n_23877, n_23878, n_23879, n_23880, n_23881, n_23882, n_23883, n_23884, n_23885, n_23886, n_23887, n_23888, n_23889, n_23890, n_23891, n_23892, n_23893, n_23894, n_23895, n_23896, n_23897, n_23898, n_23899, n_23900, n_23901, n_23902, n_23903, n_23904, n_23905, n_23906, n_23907, n_23908, n_23909, n_23910, n_23911, n_23912, n_23913, n_23914, n_23915, n_23916, n_23917, n_23918, n_23919, n_23920, n_23921, n_23922, n_23923, n_23924, n_23925, n_23926, n_23927, n_23928, n_23929, n_23930, n_23931, n_23932, n_23933, n_23934, n_23935, n_23936, n_23937, n_23938, n_23939, n_23940, n_23941, n_23942, n_23943, n_23944, n_23945, n_23946, n_23947, n_23948, n_23949, n_23950, n_23951, n_23952, n_23953, n_23954, n_23955, n_23956, n_23957, n_23958, n_23959, n_23960, n_23961, n_23962, n_23963, n_23964, n_23965, n_23966, n_23967, n_23968, n_23969, n_23970, n_23971, n_23972, n_23973, n_23974, n_23975, n_23976, n_23977, n_23978, n_23979, n_23980, n_23981, n_23982, n_23983, n_23984, n_23985, n_23986, n_23987, n_23988, n_23989, n_23990, n_23991, n_23992, n_23993, n_23994, n_23995, n_23996, n_23997, n_23998, n_23999, n_24000, n_24001, n_24002, n_24003, n_24004, n_24005, n_24006, n_24007, n_24008, n_24009, n_24010, n_24011, n_24012, n_24013, n_24014, n_24015, n_24016, n_24017, n_24018, n_24019, n_24020, n_24021, n_24022, n_24023, n_24024, n_24025, n_24026, n_24027, n_24028, n_24029, n_24030, n_24031, n_24032, n_24033, n_24034, n_24035, n_24036, n_24037, n_24038, n_24039, n_24040, n_24041, n_24042, n_24043, n_24044, n_24045, n_24046, n_24047, n_24048, n_24049, n_24050, n_24051, n_24052, n_24053, n_24054, n_24055, n_24056, n_24057, n_24058, n_24059, n_24060, n_24061, n_24062, n_24063, n_24064, n_24065, n_24066, n_24067, n_24068, n_24069, n_24070, n_24071, n_24072, n_24073, n_24074, n_24075, n_24076, n_24077, n_24078, n_24079, n_24080, n_24081, n_24082, n_24083, n_24084, n_24085, n_24086, n_24087, n_24088, n_24089, n_24090, n_24091, n_24092, n_24093, n_24094, n_24095, n_24096, n_24097, n_24098, n_24099, n_24100, n_24101, n_24102, n_24103, n_24104, n_24105, n_24106, n_24107, n_24108, n_24109, n_24110, n_24111, n_24112, n_24113, n_24114, n_24115, n_24116, n_24117, n_24118, n_24119, n_24120, n_24121, n_24122, n_24123, n_24124, n_24125, n_24126, n_24127, n_24128, n_24129, n_24130, n_24131, n_24132, n_24133, n_24134, n_24135, n_24136, n_24137, n_24138, n_24139, n_24140, n_24141, n_24142, n_24143, n_24144, n_24145, n_24146, n_24147, n_24148, n_24149, n_24150, n_24151, n_24152, n_24153, n_24154, n_24155, n_24156, n_24157, n_24158, n_24159, n_24160, n_24161, n_24162, n_24163, n_24164, n_24165, n_24166, n_24167, n_24168, n_24169, n_24170, n_24171, n_24172, n_24173, n_24174, n_24175, n_24176, n_24177, n_24178, n_24179, n_24180, n_24181, n_24182, n_24183, n_24184, n_24185, n_24186, n_24187, n_24188, n_24189, n_24190, n_24191, n_24192, n_24193, n_24194, n_24195, n_24196, n_24197, n_24198, n_24199, n_24200, n_24201, n_24202, n_24203, n_24204, n_24205, n_24206, n_24207, n_24208, n_24209, n_24210, n_24211, n_24212, n_24213, n_24214, n_24215, n_24216, n_24217, n_24218, n_24219, n_24220, n_24221, n_24222, n_24223, n_24224, n_24225, n_24226, n_24227, n_24228, n_24229, n_24230, n_24231, n_24232, n_24233, n_24234, n_24235, n_24236, n_24237, n_24238, n_24239, n_24240, n_24241, n_24242, n_24243, n_24244, n_24245, n_24246, n_24247, n_24248, n_24249, n_24250, n_24251, n_24252, n_24253, n_24254, n_24255, n_24256, n_24257, n_24258, n_24259, n_24260, n_24261, n_24262, n_24263, n_24264, n_24265, n_24266, n_24267, n_24268, n_24269, n_24270, n_24271, n_24272, n_24273, n_24274, n_24275, n_24276, n_24277, n_24278, n_24279, n_24280, n_24281, n_24282, n_24283, n_24284, n_24285, n_24286, n_24287, n_24288, n_24289, n_24290, n_24291, n_24292, n_24293, n_24294, n_24295, n_24296, n_24297, n_24298, n_24299, n_24300, n_24301, n_24302, n_24303, n_24304, n_24305, n_24306, n_24307, n_24308, n_24309, n_24310, n_24311, n_24312, n_24313, n_24314, n_24315, n_24316, n_24317, n_24318, n_24319, n_24320, n_24321, n_24322, n_24323, n_24324, n_24325, n_24326, n_24327, n_24328, n_24329, n_24330, n_24331, n_24332, n_24333, n_24334, n_24335, n_24336, n_24337, n_24338, n_24339, n_24340, n_24341, n_24342, n_24343, n_24344, n_24345, n_24346, n_24347, n_24348, n_24349, n_24350, n_24351, n_24352, n_24353, n_24354, n_24355, n_24356, n_24357, n_24358, n_24359, n_24360, n_24361, n_24362, n_24363, n_24364, n_24365, n_24366, n_24367, n_24368, n_24369, n_24370, n_24371, n_24372, n_24373, n_24374, n_24375, n_24376, n_24377, n_24378, n_24379, n_24380, n_24381, n_24382, n_24383, n_24384, n_24385, n_24386, n_24387, n_24388, n_24389, n_24390, n_24391, n_24392, n_24393, n_24394, n_24395, n_24396, n_24397, n_24398, n_24399, n_24400, n_24401, n_24402, n_24403, n_24404, n_24405, n_24406, n_24407, n_24408, n_24409, n_24410, n_24411, n_24412, n_24413, n_24414, n_24415, n_24416, n_24417, n_24418, n_24419, n_24420, n_24421, n_24422, n_24423, n_24424, n_24425, n_24426, n_24427, n_24428, n_24429, n_24430, n_24431, n_24432, n_24433, n_24434, n_24435, n_24436, n_24437, n_24438, n_24439, n_24440, n_24441, n_24442, n_24443, n_24444, n_24445, n_24446, n_24447, n_24448, n_24449, n_24450, n_24451, n_24452, n_24453, n_24454, n_24455, n_24456, n_24457, n_24458, n_24459, n_24460, n_24461, n_24462, n_24463, n_24464, n_24465, n_24466, n_24467, n_24468, n_24469, n_24470, n_24471, n_24472, n_24473, n_24474, n_24475, n_24476, n_24477, n_24478, n_24479, n_24480, n_24481, n_24482, n_24483, n_24484, n_24485, n_24486, n_24487, n_24488, n_24489, n_24490, n_24491, n_24492, n_24493, n_24494, n_24495, n_24496, n_24497, n_24498, n_24499, n_24500, n_24501, n_24502, n_24503, n_24504, n_24505, n_24506, n_24507, n_24508, n_24509, n_24510, n_24511, n_24512, n_24513, n_24514, n_24515, n_24516, n_24517, n_24518, n_24519, n_24520, n_24521, n_24522, n_24523, n_24524, n_24525, n_24526, n_24527, n_24528, n_24529, n_24530, n_24531, n_24532, n_24533, n_24534, n_24535, n_24536, n_24537, n_24538, n_24539, n_24540, n_24541, n_24542, n_24543, n_24544, n_24545, n_24546, n_24547, n_24548, n_24549, n_24550, n_24551, n_24552, n_24553, n_24554, n_24555, n_24556, n_24557, n_24558, n_24559, n_24560, n_24561, n_24562, n_24563, n_24564, n_24565, n_24566, n_24567, n_24568, n_24569, n_24570, n_24571, n_24572, n_24573, n_24574, n_24575, n_24576, n_24577, n_24578, n_24579, n_24580, n_24581, n_24582, n_24583, n_24584, n_24585, n_24586, n_24587, n_24588, n_24589, n_24590, n_24591, n_24592, n_24593, n_24594, n_24595, n_24596, n_24597, n_24598, n_24599, n_24600, n_24601, n_24602, n_24603, n_24604, n_24605, n_24606, n_24607, n_24608, n_24609, n_24610, n_24611, n_24612, n_24613, n_24614, n_24615, n_24616, n_24617, n_24618, n_24619, n_24620, n_24621, n_24622, n_24623, n_24624, n_24625, n_24626, n_24627, n_24628, n_24629, n_24630, n_24631, n_24632, n_24633, n_24634, n_24635, n_24636, n_24637, n_24638, n_24639, n_24640, n_24641, n_24642, n_24643, n_24644, n_24645, n_24646, n_24647, n_24648, n_24649, n_24650, n_24651, n_24652, n_24653, n_24654, n_24655, n_24656, n_24657, n_24658, n_24659, n_24660, n_24661, n_24662, n_24663, n_24664, n_24665, n_24666, n_24667, n_24668, n_24669, n_24670, n_24671, n_24672, n_24673, n_24674, n_24675, n_24676, n_24677, n_24678, n_24679, n_24680, n_24681, n_24682, n_24683, n_24684, n_24685, n_24686, n_24687, n_24688, n_24689, n_24690, n_24691, n_24692, n_24693, n_24694, n_24695, n_24696, n_24697, n_24698, n_24699, n_24700, n_24701, n_24702, n_24703, n_24704, n_24705, n_24706, n_24707, n_24708, n_24709, n_24710, n_24711, n_24712, n_24713, n_24714, n_24715, n_24716, n_24717, n_24718, n_24719, n_24720, n_24721, n_24722, n_24723, n_24724, n_24725, n_24726, n_24727, n_24728, n_24729, n_24730, n_24731, n_24732, n_24733, n_24734, n_24735, n_24736, n_24737, n_24738, n_24739, n_24740, n_24741, n_24742, n_24743, n_24744, n_24745, n_24746, n_24747, n_24748, n_24749, n_24750, n_24751, n_24752, n_24753, n_24754, n_24755, n_24756, n_24757, n_24758, n_24759, n_24760, n_24761, n_24762, n_24763, n_24764, n_24765, n_24766, n_24767, n_24768, n_24769, n_24770, n_24771, n_24772, n_24773, n_24774, n_24775, n_24776, n_24777, n_24778, n_24779, n_24780, n_24781, n_24782, n_24783, n_24784, n_24785, n_24786, n_24787, n_24788, n_24789, n_24790, n_24791, n_24792, n_24793, n_24794, n_24795, n_24796, n_24797, n_24798, n_24799, n_24800, n_24801, n_24802, n_24803, n_24804, n_24805, n_24806, n_24807, n_24808, n_24809, n_24810, n_24811, n_24812, n_24813, n_24814, n_24815, n_24816, n_24817, n_24818, n_24819, n_24820, n_24821, n_24822, n_24823, n_24824, n_24825, n_24826, n_24827, n_24828, n_24829, n_24830, n_24831, n_24832, n_24833, n_24834, n_24835, n_24836, n_24837, n_24838, n_24839, n_24840, n_24841, n_24842, n_24843, n_24844, n_24845, n_24846, n_24847, n_24848, n_24849, n_24850, n_24851, n_24852, n_24853, n_24854, n_24855, n_24856, n_24857, n_24858, n_24859, n_24860, n_24861, n_24862, n_24863, n_24864, n_24865, n_24866, n_24867, n_24868, n_24869, n_24870, n_24871, n_24872, n_24873, n_24874, n_24875, n_24876, n_24877, n_24878, n_24879, n_24880, n_24881, n_24882, n_24883, n_24884, n_24885, n_24886, n_24887, n_24888, n_24889, n_24890, n_24891, n_24892, n_24893, n_24894, n_24895, n_24896, n_24897, n_24898, n_24899, n_24900, n_24901, n_24902, n_24903, n_24904, n_24905, n_24906, n_24907, n_24908, n_24909, n_24910, n_24911, n_24912, n_24913, n_24914, n_24915, n_24916, n_24917, n_24918, n_24919, n_24920, n_24921, n_24922, n_24923, n_24924, n_24925, n_24926, n_24927, n_24928, n_24929, n_24930, n_24931, n_24932, n_24933, n_24934, n_24935, n_24936, n_24937, n_24938, n_24939, n_24940, n_24941, n_24942, n_24943, n_24944, n_24945, n_24946, n_24947, n_24948, n_24949, n_24950, n_24951, n_24952, n_24953, n_24954, n_24955, n_24956, n_24957, n_24958, n_24959, n_24960, n_24961, n_24962, n_24963, n_24964, n_24965, n_24966, n_24967, n_24968, n_24969, n_24970, n_24971, n_24972, n_24973, n_24974, n_24975, n_24976, n_24977, n_24978, n_24979, n_24980, n_24981, n_24982, n_24983, n_24984, n_24985, n_24986, n_24987, n_24988, n_24989, n_24990, n_24991, n_24992, n_24993, n_24994, n_24995, n_24996, n_24997, n_24998, n_24999, n_25000, n_25001, n_25002, n_25003, n_25004, n_25005, n_25006, n_25007, n_25008, n_25009, n_25010, n_25011, n_25012, n_25013, n_25014, n_25015, n_25016, n_25017, n_25018, n_25019, n_25020, n_25021, n_25022, n_25023, n_25024, n_25025, n_25026, n_25027, n_25028, n_25029, n_25030, n_25031, n_25032, n_25033, n_25034, n_25035, n_25036, n_25037, n_25038, n_25039, n_25040, n_25041, n_25042, n_25043, n_25044, n_25045, n_25046, n_25047, n_25048, n_25049, n_25050, n_25051, n_25052, n_25053, n_25054, n_25055, n_25056, n_25057, n_25058, n_25059, n_25060, n_25061, n_25062, n_25063, n_25064, n_25065, n_25066, n_25067, n_25068, n_25069, n_25070, n_25071, n_25072, n_25073, n_25074, n_25075, n_25076, n_25077, n_25078, n_25079, n_25080, n_25081, n_25082, n_25083, n_25084, n_25085, n_25086, n_25087, n_25088, n_25089, n_25090, n_25091, n_25092, n_25093, n_25094, n_25095, n_25096, n_25097, n_25098, n_25099, n_25100, n_25101, n_25102, n_25103, n_25104, n_25105, n_25106, n_25107, n_25108, n_25109, n_25110, n_25111, n_25112, n_25113, n_25114, n_25115, n_25116, n_25117, n_25118, n_25119, n_25120, n_25121, n_25122, n_25123, n_25124, n_25125, n_25126, n_25127, n_25128, n_25129, n_25130, n_25131, n_25132, n_25133, n_25134, n_25135, n_25136, n_25137, n_25138, n_25139, n_25140, n_25141, n_25142, n_25143, n_25144, n_25145, n_25146, n_25147, n_25148, n_25149, n_25150, n_25151, n_25152, n_25153, n_25154, n_25155, n_25156, n_25157, n_25158, n_25159, n_25160, n_25161, n_25162, n_25163, n_25164, n_25165, n_25166, n_25167, n_25168, n_25169, n_25170, n_25171, n_25172, n_25173, n_25174, n_25175, n_25176, n_25177, n_25178, n_25179, n_25180, n_25181, n_25182, n_25183, n_25184, n_25185, n_25186, n_25187, n_25188, n_25189, n_25190, n_25191, n_25192, n_25193, n_25194, n_25195, n_25196, n_25197, n_25198, n_25199, n_25200, n_25201, n_25202, n_25203, n_25204, n_25205, n_25206, n_25207, n_25208, n_25209, n_25210, n_25211, n_25212, n_25213, n_25214, n_25215, n_25216, n_25217, n_25218, n_25219, n_25220, n_25221, n_25222, n_25223, n_25224, n_25225, n_25226, n_25227, n_25228, n_25229, n_25230, n_25231, n_25232, n_25233, n_25234, n_25235, n_25236, n_25237, n_25238, n_25239, n_25240, n_25241, n_25242, n_25243, n_25244, n_25245, n_25246, n_25247, n_25248, n_25249, n_25250, n_25251, n_25252, n_25253, n_25254, n_25255, n_25256, n_25257, n_25258, n_25259, n_25260, n_25261, n_25262, n_25263, n_25264, n_25265, n_25266, n_25267, n_25268, n_25269, n_25270, n_25271, n_25272, n_25273, n_25274, n_25275, n_25276, n_25277, n_25278, n_25279, n_25280, n_25281, n_25282, n_25283, n_25284, n_25285, n_25286, n_25287, n_25288, n_25289, n_25290, n_25291, n_25292, n_25293, n_25294, n_25295, n_25296, n_25297, n_25298, n_25299, n_25300, n_25301, n_25302, n_25303, n_25304, n_25305, n_25306, n_25307, n_25308, n_25309, n_25310, n_25311, n_25312, n_25313, n_25314, n_25315, n_25316, n_25317, n_25318, n_25319, n_25320, n_25321, n_25322, n_25323, n_25324, n_25325, n_25326, n_25327, n_25328, n_25329, n_25330, n_25331, n_25332, n_25333, n_25334, n_25335, n_25336, n_25337, n_25338, n_25339, n_25340, n_25341, n_25342, n_25343, n_25344, n_25345, n_25346, n_25347, n_25348, n_25349, n_25350, n_25351, n_25352, n_25353, n_25354, n_25355, n_25356, n_25357, n_25358, n_25359, n_25360, n_25361, n_25362, n_25363, n_25364, n_25365, n_25366, n_25367, n_25368, n_25369, n_25370, n_25371, n_25372, n_25373, n_25374, n_25375, n_25376, n_25377, n_25378, n_25379, n_25380, n_25381, n_25382, n_25383, n_25384, n_25385, n_25386, n_25387, n_25388, n_25389, n_25390, n_25391, n_25392, n_25393, n_25394, n_25395, n_25396, n_25397, n_25398, n_25399, n_25400, n_25401, n_25402, n_25403, n_25404, n_25405, n_25406, n_25407, n_25408, n_25409, n_25410, n_25411, n_25412, n_25413, n_25414, n_25415, n_25416, n_25417, n_25418, n_25419, n_25420, n_25421, n_25422, n_25423, n_25424, n_25425, n_25426, n_25427, n_25428, n_25429, n_25430, n_25431, n_25432, n_25433, n_25434, n_25435, n_25436, n_25437, n_25438, n_25439, n_25440, n_25441, n_25442, n_25443, n_25444, n_25445, n_25446, n_25447, n_25448, n_25449, n_25450, n_25451, n_25452, n_25453, n_25454, n_25455, n_25456, n_25457, n_25458, n_25459, n_25460, n_25461, n_25462, n_25463, n_25464, n_25465, n_25466, n_25467, n_25468, n_25469, n_25470, n_25471, n_25472, n_25473, n_25474, n_25475, n_25476, n_25477, n_25478, n_25479, n_25480, n_25481, n_25482, n_25483, n_25484, n_25485, n_25486, n_25487, n_25488, n_25489, n_25490, n_25491, n_25492, n_25493, n_25494, n_25495, n_25496, n_25497, n_25498, n_25499, n_25500, n_25501, n_25502, n_25503, n_25504, n_25505, n_25506, n_25507, n_25508, n_25509, n_25510, n_25511, n_25512, n_25513, n_25514, n_25515, n_25516, n_25517, n_25518, n_25519, n_25520, n_25521, n_25522, n_25523, n_25524, n_25525, n_25526, n_25527, n_25528, n_25529, n_25530, n_25531, n_25532, n_25533, n_25534, n_25535, n_25536, n_25537, n_25538, n_25539, n_25540, n_25541, n_25542, n_25543, n_25544, n_25545, n_25546, n_25547, n_25548, n_25549, n_25550, n_25551, n_25552, n_25553, n_25554, n_25555, n_25556, n_25557, n_25558, n_25559, n_25560, n_25561, n_25562, n_25563, n_25564, n_25565, n_25566, n_25567, n_25568, n_25569, n_25570, n_25571, n_25572, n_25573, n_25574, n_25575, n_25576, n_25577, n_25578, n_25579, n_25580, n_25581, n_25582, n_25583, n_25584, n_25585, n_25586, n_25587, n_25588, n_25589, n_25590, n_25591, n_25592, n_25593, n_25594, n_25595, n_25596, n_25597, n_25598, n_25599, n_25600, n_25601, n_25602, n_25603, n_25604, n_25605, n_25606, n_25607, n_25608, n_25609, n_25610, n_25611, n_25612, n_25613, n_25614, n_25615, n_25616, n_25617, n_25618, n_25619, n_25620, n_25621, n_25622, n_25623, n_25624, n_25625, n_25626, n_25627, n_25628, n_25629, n_25630, n_25631, n_25632, n_25633, n_25634, n_25635, n_25636, n_25637, n_25638, n_25639, n_25640, n_25641, n_25642, n_25643, n_25644, n_25645, n_25646, n_25647, n_25648, n_25649, n_25650, n_25651, n_25652, n_25653, n_25654, n_25655, n_25656, n_25657, n_25658, n_25659, n_25660, n_25661, n_25662, n_25663, n_25664, n_25665, n_25666, n_25667, n_25668, n_25669, n_25670, n_25671, n_25672, n_25673, n_25674, n_25675, n_25676, n_25677, n_25678, n_25679, n_25680, n_25681, n_25682, n_25683, n_25684, n_25685, n_25686, n_25687, n_25688, n_25689, n_25690, n_25691, n_25692, n_25693, n_25694, n_25695, n_25696, n_25697, n_25698, n_25699, n_25700, n_25701, n_25702, n_25703, n_25704, n_25705, n_25706, n_25707, n_25708, n_25709, n_25710, n_25711, n_25712, n_25713, n_25714, n_25715, n_25716, n_25717, n_25718, n_25719, n_25720, n_25721, n_25722, n_25723, n_25724, n_25725, n_25726, n_25727, n_25728, n_25729, n_25730, n_25731, n_25732, n_25733, n_25734, n_25735, n_25736, n_25737, n_25738, n_25739, n_25740, n_25741, n_25742, n_25743, n_25744, n_25745, n_25746, n_25747, n_25748, n_25749, n_25750, n_25751, n_25752, n_25753, n_25754, n_25755, n_25756, n_25757, n_25758, n_25759, n_25760, n_25761, n_25762, n_25763, n_25764, n_25765, n_25766, n_25767, n_25768, n_25769, n_25770, n_25771, n_25772, n_25773, n_25774, n_25775, n_25776, n_25777, n_25778, n_25779, n_25780, n_25781, n_25782, n_25783, n_25784, n_25785, n_25786, n_25787, n_25788, n_25789, n_25790, n_25791, n_25792, n_25793, n_25794, n_25795, n_25796, n_25797, n_25798, n_25799, n_25800, n_25801, n_25802, n_25803, n_25804, n_25805, n_25806, n_25807, n_25808, n_25809, n_25810, n_25811, n_25812, n_25813, n_25814, n_25815, n_25816, n_25817, n_25818, n_25819, n_25820, n_25821, n_25822, n_25823, n_25824, n_25825, n_25826, n_25827, n_25828, n_25829, n_25830, n_25831, n_25832, n_25833, n_25834, n_25835, n_25836, n_25837, n_25838, n_25839, n_25840, n_25841, n_25842, n_25843, n_25844, n_25845, n_25846, n_25847, n_25848, n_25849, n_25850, n_25851, n_25852, n_25853, n_25854, n_25855, n_25856, n_25857, n_25858, n_25859, n_25860, n_25861, n_25862, n_25863, n_25864, n_25865, n_25866, n_25867, n_25868, n_25869, n_25870, n_25871, n_25872, n_25873, n_25874, n_25875, n_25876, n_25877, n_25878, n_25879, n_25880, n_25881, n_25882, n_25883, n_25884, n_25885, n_25886, n_25887, n_25888, n_25889, n_25890, n_25891, n_25892, n_25893, n_25894, n_25895, n_25896, n_25897, n_25898, n_25899, n_25900, n_25901, n_25902, n_25903, n_25904, n_25905, n_25906, n_25907, n_25908, n_25909, n_25910, n_25911, n_25912, n_25913, n_25914, n_25915, n_25916, n_25917, n_25918, n_25919, n_25920, n_25921, n_25922, n_25923, n_25924, n_25925, n_25926, n_25927, n_25928, n_25929, n_25930, n_25931, n_25932, n_25933, n_25934, n_25935, n_25936, n_25937, n_25938, n_25939, n_25940, n_25941, n_25942, n_25943, n_25944, n_25945, n_25946, n_25947, n_25948, n_25949, n_25950, n_25951, n_25952, n_25953, n_25954, n_25955, n_25956, n_25957, n_25958, n_25959, n_25960, n_25961, n_25962, n_25963, n_25964, n_25965, n_25966, n_25967, n_25968, n_25969, n_25970, n_25971, n_25972, n_25973, n_25974, n_25975, n_25976, n_25977, n_25978, n_25979, n_25980, n_25981, n_25982, n_25983, n_25984, n_25985, n_25986, n_25987, n_25988, n_25989, n_25990, n_25991, n_25992, n_25993, n_25994, n_25995, n_25996, n_25997, n_25998, n_25999, n_26000, n_26001, n_26002, n_26003, n_26004, n_26005, n_26006, n_26007, n_26008, n_26009, n_26010, n_26011, n_26012, n_26013, n_26014, n_26015, n_26016, n_26017, n_26018, n_26019, n_26020, n_26021, n_26022, n_26023, n_26024, n_26025, n_26026, n_26027, n_26028, n_26029, n_26030, n_26031, n_26032, n_26033, n_26034, n_26035, n_26036, n_26037, n_26038, n_26039, n_26040, n_26041, n_26042, n_26043, n_26044, n_26045, n_26046, n_26047, n_26048, n_26049, n_26050, n_26051, n_26052, n_26053, n_26054, n_26055, n_26056, n_26057, n_26058, n_26059, n_26060, n_26061, n_26062, n_26063, n_26064, n_26065, n_26066, n_26067, n_26068, n_26069, n_26070, n_26071, n_26072, n_26073, n_26074, n_26075, n_26076, n_26077, n_26078, n_26079, n_26080, n_26081, n_26082, n_26083, n_26084, n_26085, n_26086, n_26087, n_26088, n_26089, n_26090, n_26091, n_26092, n_26093, n_26094, n_26095, n_26096, n_26097, n_26098, n_26099, n_26100, n_26101, n_26102, n_26103, n_26104, n_26105, n_26106, n_26107, n_26108, n_26109, n_26110, n_26111, n_26112, n_26113, n_26114, n_26115, n_26116, n_26117, n_26118, n_26119, n_26120, n_26121, n_26122, n_26123, n_26124, n_26125, n_26126, n_26127, n_26128, n_26129, n_26130, n_26131, n_26132, n_26133, n_26134, n_26135, n_26136, n_26137, n_26138, n_26139, n_26140, n_26141, n_26142, n_26143, n_26144, n_26145, n_26146, n_26147, n_26148, n_26149, n_26150, n_26151, n_26152, n_26153, n_26154, n_26155, n_26156, n_26157, n_26158, n_26159, n_26160, n_26161, n_26162, n_26163, n_26164, n_26165, n_26166, n_26167, n_26168, n_26169, n_26170, n_26171, n_26172, n_26173, n_26174, n_26175, n_26176, n_26177, n_26178, n_26179, n_26180, n_26181, n_26182, n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189, n_26190, n_26191, n_26192, n_26193, n_26194, n_26195, n_26196, n_26197, n_26198, n_26199, n_26200, n_26201, n_26202, n_26203, n_26204, n_26205, n_26206, n_26207, n_26208, n_26209, n_26210, n_26211, n_26212, n_26213, n_26214, n_26215, n_26216, n_26217, n_26218, n_26219, n_26220, n_26221, n_26222, n_26223, n_26224, n_26225, n_26226, n_26227, n_26228, n_26229, n_26230, n_26231, n_26232, n_26233, n_26234, n_26235, n_26236, n_26237, n_26238, n_26239, n_26240, n_26241, n_26242, n_26243, n_26244, n_26245, n_26246, n_26247, n_26248, n_26249, n_26250, n_26251, n_26252, n_26253, n_26254, n_26255, n_26256, n_26257, n_26258, n_26259, n_26260, n_26261, n_26262, n_26263, n_26264, n_26265, n_26266, n_26267, n_26268, n_26269, n_26270, n_26271, n_26272, n_26273, n_26274, n_26275, n_26276, n_26277, n_26278, n_26279, n_26280, n_26281, n_26282, n_26283, n_26284, n_26285, n_26286, n_26287, n_26288, n_26289, n_26290, n_26291, n_26292, n_26293, n_26294, n_26295, n_26296, n_26297, n_26298, n_26299, n_26300, n_26301, n_26302, n_26303, n_26304, n_26305, n_26306, n_26307, n_26308, n_26309, n_26310, n_26311, n_26312, n_26313, n_26314, n_26315, n_26316, n_26317, n_26318, n_26319, n_26320, n_26321, n_26322, n_26323, n_26324, n_26325, n_26326, n_26327, n_26328, n_26329, n_26330, n_26331, n_26332, n_26333, n_26334, n_26335, n_26336, n_26337, n_26338, n_26339, n_26340, n_26341, n_26342, n_26343, n_26344, n_26345, n_26346, n_26347, n_26348, n_26349, n_26350, n_26351, n_26352, n_26353, n_26354, n_26355, n_26356, n_26357, n_26358, n_26359, n_26360, n_26361, n_26362, n_26363, n_26364, n_26365, n_26366, n_26367, n_26368, n_26369, n_26370, n_26371, n_26372, n_26373, n_26374, n_26375, n_26376, n_26377, n_26378, n_26379, n_26380, n_26381, n_26382, n_26383, n_26384, n_26385, n_26386, n_26387, n_26388, n_26389, n_26390, n_26391, n_26392, n_26393, n_26394, n_26395, n_26396, n_26397, n_26398, n_26399, n_26400, n_26401, n_26402, n_26403, n_26404, n_26405, n_26406, n_26407, n_26408, n_26409, n_26410, n_26411, n_26412, n_26413, n_26414, n_26415, n_26416, n_26417, n_26418, n_26419, n_26420, n_26421, n_26422, n_26423, n_26424, n_26425, n_26426, n_26427, n_26428, n_26429, n_26430, n_26431, n_26432, n_26433, n_26434, n_26435, n_26436, n_26437, n_26438, n_26439, n_26440, n_26441, n_26442, n_26443, n_26444, n_26445, n_26446, n_26447, n_26448, n_26449, n_26450, n_26451, n_26452, n_26453, n_26454, n_26455, n_26456, n_26457, n_26458, n_26459, n_26460, n_26461, n_26462, n_26463, n_26464, n_26465, n_26466, n_26467, n_26468, n_26469, n_26470, n_26471, n_26472, n_26473, n_26474, n_26475, n_26476, n_26477, n_26478, n_26479, n_26480, n_26481, n_26482, n_26483, n_26484, n_26485, n_26486, n_26487, n_26488, n_26489, n_26490, n_26491, n_26492, n_26493, n_26494, n_26495, n_26496, n_26497, n_26498, n_26499, n_26500, n_26501, n_26502, n_26503, n_26504, n_26505, n_26506, n_26507, n_26508, n_26509, n_26510, n_26511, n_26512, n_26513, n_26514, n_26515, n_26516, n_26517, n_26518, n_26519, n_26520, n_26521, n_26522, n_26523, n_26524, n_26525, n_26526, n_26527, n_26528, n_26529, n_26530, n_26531, n_26532, n_26533, n_26534, n_26535, n_26536, n_26537, n_26538, n_26539, n_26540, n_26541, n_26542, n_26543, n_26544, n_26545, n_26546, n_26547, n_26548, n_26549, n_26550, n_26551, n_26552, n_26553, n_26554, n_26555, n_26556, n_26557, n_26558, n_26559, n_26560, n_26561, n_26562, n_26563, n_26564, n_26565, n_26566, n_26567, n_26568, n_26569, n_26570, n_26571, n_26572, n_26573, n_26574, n_26575, n_26576, n_26577, n_26578, n_26579, n_26580, n_26581, n_26582, n_26583, n_26584, n_26585, n_26586, n_26587, n_26588, n_26589, n_26590, n_26591, n_26592, n_26593, n_26594, n_26595, n_26596, n_26597, n_26598, n_26599, n_26600, n_26601, n_26602, n_26603, n_26604, n_26605, n_26606, n_26607, n_26608, n_26609, n_26610, n_26611, n_26612, n_26613, n_26614, n_26615, n_26616, n_26617, n_26618, n_26619, n_26620, n_26621, n_26622, n_26623, n_26624, n_26625, n_26626, n_26627, n_26628, n_26629, n_26630, n_26631, n_26632, n_26633, n_26634, n_26635, n_26636, n_26637, n_26638, n_26639, n_26640, n_26641, n_26642, n_26643, n_26644, n_26645, n_26646, n_26647, n_26648, n_26649, n_26650, n_26651, n_26652, n_26653, n_26654, n_26655, n_26656, n_26657, n_26658, n_26659, n_26660, n_26661, n_26662, n_26663, n_26664, n_26665, n_26666, n_26667, n_26668, n_26669, n_26670, n_26671, n_26672, n_26673, n_26674, n_26675, n_26676, n_26677, n_26678, n_26679, n_26680, n_26681, n_26682, n_26683, n_26684, n_26685, n_26686, n_26687, n_26688, n_26689, n_26690, n_26691, n_26692, n_26693, n_26694, n_26695, n_26696, n_26697, n_26698, n_26699, n_26700, n_26701, n_26702, n_26703, n_26704, n_26705, n_26706, n_26707, n_26708, n_26709, n_26710, n_26711, n_26712, n_26713, n_26714, n_26715, n_26716, n_26717, n_26718, n_26719, n_26720, n_26721, n_26722, n_26723, n_26724, n_26725, n_26726, n_26727, n_26728, n_26729, n_26730, n_26731, n_26732, n_26733, n_26734, n_26735, n_26736, n_26737, n_26738, n_26739, n_26740, n_26741, n_26742, n_26743, n_26744, n_26745, n_26746, n_26747, n_26748, n_26749, n_26750, n_26751, n_26752, n_26753, n_26754, n_26755, n_26756, n_26757, n_26758, n_26759, n_26760, n_26761, n_26762, n_26763, n_26764, n_26765, n_26766, n_26767, n_26768, n_26769, n_26770, n_26771, n_26772, n_26773, n_26774, n_26775, n_26776, n_26777, n_26778, n_26779, n_26780, n_26781, n_26782, n_26783, n_26784, n_26785, n_26786, n_26787, n_26788, n_26789, n_26790, n_26791, n_26792, n_26793, n_26794, n_26795, n_26796, n_26797, n_26798, n_26799, n_26800, n_26801, n_26802, n_26803, n_26804, n_26805, n_26806, n_26807, n_26808, n_26809, n_26810, n_26811, n_26812, n_26813, n_26814, n_26815, n_26816, n_26817, n_26818, n_26819, n_26820, n_26821, n_26822, n_26823, n_26824, n_26825, n_26826, n_26827, n_26828, n_26829, n_26830, n_26831, n_26832, n_26833, n_26834, n_26835, n_26836, n_26837, n_26838, n_26839, n_26840, n_26841, n_26842, n_26843, n_26844, n_26845, n_26846, n_26847, n_26848, n_26849, n_26850, n_26851, n_26852, n_26853, n_26854, n_26855, n_26856, n_26857, n_26858, n_26859, n_26860, n_26861, n_26862, n_26863, n_26864, n_26865, n_26866, n_26867, n_26868, n_26869, n_26870, n_26871, n_26872, n_26873, n_26874, n_26875, n_26876, n_26877, n_26878, n_26879, n_26880, n_26881, n_26882, n_26883, n_26884, n_26885, n_26886, n_26887, n_26888, n_26889, n_26890, n_26891, n_26892, n_26893, n_26894, n_26895, n_26896, n_26897, n_26898, n_26899, n_26900, n_26901, n_26902, n_26903, n_26904, n_26905, n_26906, n_26907, n_26908, n_26909, n_26910, n_26911, n_26912, n_26913, n_26914, n_26915, n_26916, n_26917, n_26918, n_26919, n_26920, n_26921, n_26922, n_26923, n_26924, n_26925, n_26926, n_26927, n_26928, n_26929, n_26930, n_26931, n_26932, n_26933, n_26934, n_26935, n_26936, n_26937, n_26938, n_26939, n_26940, n_26941, n_26942, n_26943, n_26944, n_26945, n_26946, n_26947, n_26948, n_26949, n_26950, n_26951, n_26952, n_26953, n_26954, n_26955, n_26956, n_26957, n_26958, n_26959, n_26960, n_26961, n_26962, n_26963, n_26964, n_26965, n_26966, n_26967, n_26968, n_26969, n_26970, n_26971, n_26972, n_26973, n_26974, n_26975, n_26976, n_26977, n_26978, n_26979, n_26980, n_26981, n_26982, n_26983, n_26984, n_26985, n_26986, n_26987, n_26988, n_26989, n_26990, n_26991, n_26992, n_26993, n_26994, n_26995, n_26996, n_26997, n_26998, n_26999, n_27000, n_27001, n_27002, n_27003, n_27004, n_27005, n_27006, n_27007, n_27008, n_27009, n_27010, n_27011, n_27012, n_27013, n_27014, n_27015, n_27016, n_27017, n_27018, n_27019, n_27020, n_27021, n_27022, n_27023, n_27024, n_27025, n_27026, n_27027, n_27028, n_27029, n_27030, n_27031, n_27032, n_27033, n_27034, n_27035, n_27036, n_27037, n_27038, n_27039, n_27040, n_27041, n_27042, n_27043, n_27044, n_27045, n_27046, n_27047, n_27048, n_27049, n_27050, n_27051, n_27052, n_27053, n_27054, n_27055, n_27056, n_27057, n_27058, n_27059, n_27060, n_27061, n_27062, n_27063, n_27064, n_27065, n_27066, n_27067, n_27068, n_27069, n_27070, n_27071, n_27072, n_27073, n_27074, n_27075, n_27076, n_27077, n_27078, n_27079, n_27080, n_27081, n_27082, n_27083, n_27084, n_27085, n_27086, n_27087, n_27088, n_27089, n_27090, n_27091, n_27092, n_27093, n_27094, n_27095, n_27096, n_27097, n_27098, n_27099, n_27100, n_27101, n_27102, n_27103, n_27104, n_27105, n_27106, n_27107, n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114, n_27115, n_27116, n_27117, n_27118, n_27119, n_27120, n_27121, n_27122, n_27123, n_27124, n_27125, n_27126, n_27127, n_27128, n_27129, n_27130, n_27131, n_27132, n_27133, n_27134, n_27135, n_27136, n_27137, n_27138, n_27139, n_27140, n_27141, n_27142, n_27143, n_27144, n_27145, n_27146, n_27147, n_27148, n_27149, n_27150, n_27151, n_27152, n_27153, n_27154, n_27155, n_27156, n_27157, n_27158, n_27159, n_27160, n_27161, n_27162, n_27163, n_27164, n_27165, n_27166, n_27167, n_27168, n_27169, n_27170, n_27171, n_27172, n_27173, n_27174, n_27175, n_27176, n_27177, n_27178, n_27179, n_27180, n_27181, n_27182, n_27183, n_27184, n_27185, n_27186, n_27187, n_27188, n_27189, n_27190, n_27191, n_27192, n_27193, n_27194, n_27195, n_27196, n_27197, n_27198, n_27199, n_27200, n_27201, n_27202, n_27203, n_27204, n_27205, n_27206, n_27207, n_27208, n_27209, n_27210, n_27211, n_27212, n_27213, n_27214, n_27215, n_27216, n_27217, n_27218, n_27219, n_27220, n_27221, n_27222, n_27223, n_27224, n_27225, n_27226, n_27227, n_27228, n_27229, n_27230, n_27231, n_27232, n_27233, n_27234, n_27235, n_27236, n_27237, n_27238, n_27239, n_27240, n_27241, n_27242, n_27243, n_27244, n_27245, n_27246, n_27247, n_27248, n_27249, n_27250, n_27251, n_27252, n_27253, n_27254, n_27255, n_27256, n_27257, n_27258, n_27259, n_27260, n_27261, n_27262, n_27263, n_27264, n_27265, n_27266, n_27267, n_27268, n_27269, n_27270, n_27271, n_27272, n_27273, n_27274, n_27275, n_27276, n_27277, n_27278, n_27279, n_27280, n_27281, n_27282, n_27283, n_27284, n_27285, n_27286, n_27287, n_27288, n_27289, n_27290, n_27291, n_27292, n_27293, n_27294, n_27295, n_27296, n_27297, n_27298, n_27299, n_27300, n_27301, n_27302, n_27303, n_27304, n_27305, n_27306, n_27307, n_27308, n_27309, n_27310, n_27311, n_27312, n_27313, n_27314, n_27315, n_27316, n_27317, n_27318, n_27319, n_27320, n_27321, n_27322, n_27323, n_27324, n_27325, n_27326, n_27327, n_27328, n_27329, n_27330, n_27331, n_27332, n_27333, n_27334, n_27335, n_27336, n_27337, n_27338, n_27339, n_27340, n_27341, n_27342, n_27343, n_27344, n_27345, n_27346, n_27347, n_27348, n_27349, n_27350, n_27351, n_27352, n_27353, n_27354, n_27355, n_27356, n_27357, n_27358, n_27359, n_27360, n_27361, n_27362, n_27363, n_27364, n_27365, n_27366, n_27367, n_27368, n_27369, n_27370, n_27371, n_27372, n_27373, n_27374, n_27375, n_27376, n_27377, n_27378, n_27379, n_27380, n_27381, n_27382, n_27383, n_27384, n_27385, n_27386, n_27387, n_27388, n_27389, n_27390, n_27391, n_27392, n_27393, n_27394, n_27395, n_27396, n_27397, n_27398, n_27399, n_27400, n_27401, n_27402, n_27403, n_27404, n_27405, n_27406, n_27407, n_27408, n_27409, n_27410, n_27411, n_27412, n_27413, n_27414, n_27415, n_27416, n_27417, n_27418, n_27419, n_27420, n_27421, n_27422, n_27423, n_27424, n_27425, n_27426, n_27427, n_27428, n_27429, n_27430, n_27431, n_27432, n_27433, n_27434, n_27435, n_27436, n_27437, n_27438, n_27439, n_27440, n_27441, n_27442, n_27443, n_27444, n_27445, n_27446, n_27447, n_27448, n_27449, n_27450, n_27451, n_27452, n_27453, n_27454, n_27455, n_27456, n_27457, n_27458, n_27459, n_27460, n_27461, n_27462, n_27463, n_27464, n_27465, n_27466, n_27467, n_27468, n_27469, n_27470, n_27471, n_27472, n_27473, n_27474, n_27475, n_27476, n_27477, n_27478, n_27479, n_27480, n_27481, n_27482, n_27483, n_27484, n_27485, n_27486, n_27487, n_27488, n_27489, n_27490, n_27491, n_27492, n_27493, n_27494, n_27495, n_27496, n_27497, n_27498, n_27499, n_27500, n_27501, n_27502, n_27503, n_27504, n_27505, n_27506, n_27507, n_27508, n_27509, n_27510, n_27511, n_27512, n_27513, n_27514, n_27515, n_27516, n_27517, n_27518, n_27519, n_27520, n_27521, n_27522, n_27523, n_27524, n_27525, n_27526, n_27527, n_27528, n_27529, n_27530, n_27531, n_27532, n_27533, n_27534, n_27535, n_27536, n_27537, n_27538, n_27539, n_27540, n_27541, n_27542, n_27543, n_27544, n_27545, n_27546, n_27547, n_27548, n_27549, n_27550, n_27551, n_27552, n_27553, n_27554, n_27555, n_27556, n_27557, n_27558, n_27559, n_27560, n_27561, n_27562, n_27563, n_27564, n_27565, n_27566, n_27567, n_27568, n_27569, n_27570, n_27571, n_27572, n_27573, n_27574, n_27575, n_27576, n_27577, n_27578, n_27579, n_27580, n_27581, n_27582, n_27583, n_27584, n_27585, n_27586, n_27587, n_27588, n_27589, n_27590, n_27591, n_27592, n_27593, n_27594, n_27595, n_27596, n_27597, n_27598, n_27599, n_27600, n_27601, n_27602, n_27603, n_27604, n_27605, n_27606, n_27607, n_27608, n_27609, n_27610, n_27611, n_27612, n_27613, n_27614, n_27615, n_27616, n_27617, n_27618, n_27619, n_27620, n_27621, n_27622, n_27623, n_27624, n_27625, n_27626, n_27627, n_27628, n_27629, n_27630, n_27631, n_27632, n_27633, n_27634, n_27635, n_27636, n_27637, n_27638, n_27639, n_27640, n_27641, n_27642, n_27643, n_27644, n_27645, n_27646, n_27647, n_27648, n_27649, n_27650, n_27651, n_27652, n_27653, n_27654, n_27655, n_27656, n_27657, n_27658, n_27659, n_27660, n_27661, n_27662, n_27663, n_27664, n_27665, n_27666, n_27667, n_27668, n_27669, n_27670, n_27671, n_27672, n_27673, n_27674, n_27675, n_27676, n_27677, n_27678, n_27679, n_27680, n_27681, n_27682, n_27683, n_27684, n_27685, n_27686, n_27687, n_27688, n_27689, n_27690, n_27691, n_27692, n_27693, n_27694, n_27695, n_27696, n_27697, n_27698, n_27699, n_27700, n_27701, n_27702, n_27703, n_27704, n_27705, n_27706, n_27707, n_27708, n_27709, n_27710, n_27711, n_27712, n_27713, n_27714, n_27715, n_27716, n_27717, n_27718, n_27719, n_27720, n_27721, n_27722, n_27723, n_27724, n_27725, n_27726, n_27727, n_27728, n_27729, n_27730, n_27731, n_27732, n_27733, n_27734, n_27735, n_27736, n_27737, n_27738, n_27739, n_27740, n_27741, n_27742, n_27743, n_27744, n_27745, n_27746, n_27747, n_27748, n_27749, n_27750, n_27751, n_27752, n_27753, n_27754, n_27755, n_27756, n_27757, n_27758, n_27759, n_27760, n_27761, n_27762, n_27763, n_27764, n_27765, n_27766, n_27767, n_27768, n_27769, n_27770, n_27771, n_27772, n_27773, n_27774, n_27775, n_27776, n_27777, n_27778, n_27779, n_27780, n_27781, n_27782, n_27783, n_27784, n_27785, n_27786, n_27787, n_27788, n_27789, n_27790, n_27791, n_27792, n_27793, n_27794, n_27795, n_27796, n_27797, n_27798, n_27799, n_27800, n_27801, n_27802, n_27803, n_27804, n_27805, n_27806, n_27807, n_27808, n_27809, n_27810, n_27811, n_27812, n_27813, n_27814, n_27815, n_27816, n_27817, n_27818, n_27819, n_27820, n_27821, n_27822, n_27823, n_27824, n_27825, n_27826, n_27827, n_27828, n_27829, n_27830, n_27831, n_27832, n_27833, n_27834, n_27835, n_27836, n_27837, n_27838, n_27839, n_27840, n_27841, n_27842, n_27843, n_27844, n_27845, n_27846, n_27847, n_27848, n_27849, n_27850, n_27851, n_27852, n_27853, n_27854, n_27855, n_27856, n_27857, n_27858, n_27859, n_27860, n_27861, n_27862, n_27863, n_27864, n_27865, n_27866, n_27867, n_27868, n_27869, n_27870, n_27871, n_27872, n_27873, n_27874, n_27875, n_27876, n_27877, n_27878, n_27879, n_27880, n_27881, n_27882, n_27883, n_27884, n_27885, n_27886, n_27887, n_27888, n_27889, n_27890, n_27891, n_27892, n_27893, n_27894, n_27895, n_27896, n_27897, n_27898, n_27899, n_27900, n_27901, n_27902, n_27903, n_27904, n_27905, n_27906, n_27907, n_27908, n_27909, n_27910, n_27911, n_27912, n_27913, n_27914, n_27915, n_27916, n_27917, n_27918, n_27919, n_27920, n_27921, n_27922, n_27923, n_27924, n_27925, n_27926, n_27927, n_27928, n_27929, n_27930, n_27931, n_27932, n_27933, n_27934, n_27935, n_27936, n_27937, n_27938, n_27939, n_27940, n_27941, n_27942, n_27943, n_27944, n_27945, n_27946, n_27947, n_27948, n_27949, n_27950, n_27951, n_27952, n_27953, n_27954, n_27955, n_27956, n_27957, n_27958, n_27959, n_27960, n_27961, n_27962, n_27963, n_27964, n_27965, n_27966, n_27967, n_27968, n_27969, n_27970, n_27971, n_27972, n_27973, n_27974, n_27975, n_27976, n_27977, n_27978, n_27979, n_27980, n_27981, n_27982, n_27983, n_27984, n_27985, n_27986, n_27987, n_27988, n_27989, n_27990, n_27991, n_27992, n_27993, n_27994, n_27995, n_27996, n_27997, n_27998, n_27999, n_28000, n_28001, n_28002, n_28003, n_28004, n_28005, n_28006, n_28007, n_28008, n_28009, n_28010, n_28011, n_28012, n_28013, n_28014, n_28015, n_28016, n_28017, n_28018, n_28019, n_28020, n_28021, n_28022, n_28023, n_28024, n_28025, n_28026, n_28027, n_28028, n_28029, n_28030, n_28031, n_28032, n_28033, n_28034, n_28035, n_28036, n_28037, n_28038, n_28039, n_28040, n_28041, n_28042, n_28043, n_28044, n_28045, n_28046, n_28047, n_28048, n_28049, n_28050, n_28051, n_28052, n_28053, n_28054, n_28055, n_28056, n_28057, n_28058, n_28059, n_28060, n_28061, n_28062, n_28063, n_28064, n_28065, n_28066, n_28067, n_28068, n_28069, n_28070, n_28071, n_28072, n_28073, n_28074, n_28075, n_28076, n_28077, n_28078, n_28079, n_28080, n_28081, n_28082, n_28083, n_28084, n_28085, n_28086, n_28087, n_28088, n_28089, n_28090, n_28091, n_28092, n_28093, n_28094, n_28095, n_28096, n_28097, n_28098, n_28099, n_28100, n_28101, n_28102, n_28103, n_28104, n_28105, n_28106, n_28107, n_28108, n_28109, n_28110, n_28111, n_28112, n_28113, n_28114, n_28115, n_28116, n_28117, n_28118, n_28119, n_28120, n_28121, n_28122, n_28123, n_28124, n_28125, n_28126, n_28127, n_28128, n_28129, n_28130, n_28131, n_28132, n_28133, n_28134, n_28135, n_28136, n_28137, n_28138, n_28139, n_28140, n_28141, n_28142, n_28143, n_28144, n_28145, n_28146, n_28147, n_28148, n_28149, n_28150, n_28151, n_28152, n_28153, n_28154, n_28155, n_28156, n_28157, n_28158, n_28159, n_28160, n_28161, n_28162, n_28163, n_28164, n_28165, n_28166, n_28167, n_28168, n_28169, n_28170, n_28171, n_28172, n_28173, n_28174, n_28175, n_28176, n_28177, n_28178, n_28179, n_28180, n_28181, n_28182, n_28183, n_28184, n_28185, n_28186, n_28187, n_28188, n_28189, n_28190, n_28191, n_28192, n_28193, n_28194, n_28195, n_28196, n_28197, n_28198, n_28199, n_28200, n_28201, n_28202, n_28203, n_28204, n_28205, n_28206, n_28207, n_28208, n_28209, n_28210, n_28211, n_28212, n_28213, n_28214, n_28215, n_28216, n_28217, n_28218, n_28219, n_28220, n_28221, n_28222, n_28223, n_28224, n_28225, n_28226, n_28227, n_28228, n_28229, n_28230, n_28231, n_28232, n_28233, n_28234, n_28235, n_28236, n_28237, n_28238, n_28239, n_28240, n_28241, n_28242, n_28243, n_28244, n_28245, n_28246, n_28247, n_28248, n_28249, n_28250, n_28251, n_28252, n_28253, n_28254, n_28255, n_28256, n_28257, n_28258, n_28259, n_28260, n_28261, n_28262, n_28263, n_28264, n_28265, n_28266, n_28267, n_28268, n_28269, n_28270, n_28271, n_28272, n_28273, n_28274, n_28275, n_28276, n_28277, n_28278, n_28279, n_28280, n_28281, n_28282, n_28283, n_28284, n_28285, n_28286, n_28287, n_28288, n_28289, n_28290, n_28291, n_28292, n_28293, n_28294, n_28295, n_28296, n_28297, n_28298, n_28299, n_28300, n_28301, n_28302, n_28303, n_28304, n_28305, n_28306, n_28307, n_28308, n_28309, n_28310, n_28311, n_28312, n_28313, n_28314, n_28315, n_28316, n_28317, n_28318, n_28319, n_28320, n_28321, n_28322, n_28323, n_28324, n_28325, n_28326, n_28327, n_28328, n_28329, n_28330, n_28331, n_28332, n_28333, n_28334, n_28335, n_28336, n_28337, n_28338, n_28339, n_28340, n_28341, n_28342, n_28343, n_28344, n_28345, n_28346, n_28347, n_28348, n_28349, n_28350, n_28351, n_28352, n_28353, n_28354, n_28355, n_28356, n_28357, n_28358, n_28359, n_28360, n_28361, n_28362, n_28363, n_28364, n_28365, n_28366, n_28367, n_28368, n_28369, n_28370, n_28371, n_28372, n_28373, n_28374, n_28375, n_28376, n_28377, n_28378, n_28379, n_28380, n_28381, n_28382, n_28383, n_28384, n_28385, n_28386, n_28387, n_28388, n_28389, n_28390, n_28391, n_28392, n_28393, n_28394, n_28395, n_28396, n_28397, n_28398, n_28399, n_28400, n_28401, n_28402, n_28403, n_28404, n_28405, n_28406, n_28407, n_28408, n_28409, n_28410, n_28411, n_28412, n_28413, n_28414, n_28415, n_28416, n_28417, n_28418, n_28419, n_28420, n_28421, n_28422, n_28423, n_28424, n_28425, n_28426, n_28427, n_28428, n_28429, n_28430, n_28431, n_28432, n_28433, n_28434, n_28435, n_28436, n_28437, n_28438, n_28439, n_28440, n_28441, n_28442, n_28443, n_28444, n_28445, n_28446, n_28447, n_28448, n_28449, n_28450, n_28451, n_28452, n_28453, n_28454, n_28455, n_28456, n_28457, n_28458, n_28459, n_28460, n_28461, n_28462, n_28463, n_28464, n_28465, n_28466, n_28467, n_28468, n_28469, n_28470, n_28471, n_28472, n_28473, n_28474, n_28475, n_28476, n_28477, n_28478, n_28479, n_28480, n_28481, n_28482, n_28483, n_28484, n_28485, n_28486, n_28487, n_28488, n_28489, n_28490, n_28491, n_28492, n_28493, n_28494, n_28495, n_28496, n_28497, n_28498, n_28499, n_28500, n_28501, n_28502, n_28503, n_28504, n_28505, n_28506, n_28507, n_28508, n_28509, n_28510, n_28511, n_28512, n_28513, n_28514, n_28515, n_28516, n_28517, n_28518, n_28519, n_28520, n_28521, n_28522, n_28523, n_28524, n_28525, n_28526, n_28527, n_28528, n_28529, n_28530, n_28531, n_28532, n_28533, n_28534, n_28535, n_28536, n_28537, n_28538, n_28539, n_28540, n_28541, n_28542, n_28543, n_28544, n_28545, n_28546, n_28547, n_28548, n_28549, n_28550, n_28551, n_28552, n_28553, n_28554, n_28555, n_28556, n_28557, n_28558, n_28559, n_28560, n_28561, n_28562, n_28563, n_28564, n_28565, n_28566, n_28567, n_28568, n_28569, n_28570, n_28571, n_28572, n_28573, n_28574, n_28575, n_28576, n_28577, n_28578, n_28579, n_28580, n_28581, n_28582, n_28583, n_28584, n_28585, n_28586, n_28587, n_28588, n_28589, n_28590, n_28591, n_28592, n_28593, n_28594, n_28595, n_28596, n_28597, n_28598, n_28599, n_28600, n_28601, n_28602, n_28603, n_28604, n_28605, n_28606, n_28607, n_28608, n_28609, n_28610, n_28611, n_28612, n_28613, n_28614, n_28615, n_28616, n_28617, n_28618, n_28619, n_28620, n_28621, n_28622, n_28623, n_28624, n_28625, n_28626, n_28627, n_28628, n_28629, n_28630, n_28631, n_28632, n_28633, n_28634, n_28635, n_28636, n_28637, n_28638, n_28639, n_28640, n_28641, n_28642, n_28643, n_28644, n_28645, n_28646, n_28647, n_28648, n_28649, n_28650, n_28651, n_28652, n_28653, n_28654, n_28655, n_28656, n_28657, n_28658, n_28659, n_28660, n_28661, n_28662, n_28663, n_28664, n_28665, n_28666, n_28667, n_28668, n_28669, n_28670, n_28671, n_28672, n_28673, n_28674, n_28675, n_28676, n_28677, n_28678, n_28679, n_28680, n_28681, n_28682, n_28683, n_28684, n_28685, n_28686, n_28687, n_28688, n_28689, n_28690, n_28691, n_28692, n_28693, n_28694, n_28695, n_28696, n_28697, n_28698, n_28699, n_28700, n_28701, n_28702, n_28703, n_28704, n_28705, n_28706, n_28707, n_28708, n_28709, n_28710, n_28711, n_28712, n_28713, n_28714, n_28715, n_28716, n_28717, n_28718, n_28719, n_28720, n_28721, n_28722, n_28723, n_28724, n_28725, n_28726, n_28727, n_28728, n_28729, n_28730, n_28731, n_28732, n_28733, n_28734, n_28735, n_28736, n_28737, n_28738, n_28739, n_28740, n_28741, n_28742, n_28743, n_28744, n_28745, n_28746, n_28747, n_28748, n_28749, n_28750, n_28751, n_28752, n_28753, n_28754, n_28755, n_28756, n_28757, n_28758, n_28759, n_28760, n_28761, n_28762, n_28763, n_28764, n_28765, n_28766, n_28767, n_28768, n_28769, n_28770, n_28771, n_28772, n_28773, n_28774, n_28775, n_28776, n_28777, n_28778, n_28779, n_28780, n_28781, n_28782, n_28783, n_28784, n_28785, n_28786, n_28787, n_28788, n_28789, n_28790, n_28791, n_28792, n_28793, n_28794, n_28795, n_28796, n_28797, n_28798, n_28799, n_28800, n_28801, n_28802, n_28803, n_28804, n_28805, n_28806, n_28807, n_28808, n_28809, n_28810, n_28811, n_28812, n_28813, n_28814, n_28815, n_28816, n_28817, n_28818, n_28819, n_28820, n_28821, n_28822, n_28823, n_28824, n_28825, n_28826, n_28827, n_28828, n_28829, n_28830, n_28831, n_28832, n_28833, n_28834, n_28835, n_28836, n_28837, n_28838, n_28839, n_28840, n_28841, n_28842, n_28843, n_28844, n_28845, n_28846, n_28847, n_28848, n_28849, n_28850, n_28851, n_28852, n_28853, n_28854, n_28855, n_28856, n_28857, n_28858, n_28859, n_28860, n_28861, n_28862, n_28863, n_28864, n_28865, n_28866, n_28867, n_28868, n_28869, n_28870, n_28871, n_28872, n_28873, n_28874, n_28875, n_28876, n_28877, n_28878, n_28879, n_28880, n_28881, n_28882, n_28883, n_28884, n_28885, n_28886, n_28887, n_28888, n_28889, n_28890, n_28891, n_28892, n_28893, n_28894, n_28895, n_28896, n_28897, n_28898, n_28899, n_28900, n_28901, n_28902, n_28903, n_28904, n_28905, n_28906, n_28907, n_28908, n_28909, n_28910, n_28911, n_28912, n_28913, n_28914, n_28915, n_28916, n_28917, n_28918, n_28919, n_28920, n_28921, n_28922, n_28923, n_28924, n_28925, n_28926, n_28927, n_28928, n_28929, n_28930, n_28931, n_28932, n_28933, n_28934, n_28935, n_28936, n_28937, n_28938, n_28939, n_28940, n_28941, n_28942, n_28943, n_28944, n_28945, n_28946, n_28947, n_28948, n_28949, n_28950, n_28951, n_28952, n_28953, n_28954, n_28955, n_28956, n_28957, n_28958, n_28959, n_28960, n_28961, n_28962, n_28963, n_28964, n_28965, n_28966, n_28967, n_28968, n_28969, n_28970, n_28971, n_28972, n_28973, n_28974, n_28975, n_28976, n_28977, n_28978, n_28979, n_28980, n_28981, n_28982, n_28983, n_28984, n_28985, n_28986, n_28987, n_28988, n_28989, n_28990, n_28991, n_28992, n_28993, n_28994, n_28995, n_28996, n_28997, n_28998, n_28999, n_29000, n_29001, n_29002, n_29003, n_29004, n_29005, n_29006, n_29007, n_29008, n_29009, n_29010, n_29011, n_29012, n_29013, n_29014, n_29015, n_29016, n_29017, n_29018, n_29019, n_29020, n_29021, n_29022, n_29023, n_29024, n_29025, n_29026, n_29027, n_29028, n_29029, n_29030, n_29031, n_29032, n_29033, n_29034, n_29035, n_29036, n_29037, n_29038, n_29039, n_29040, n_29041, n_29042, n_29043, n_29044, n_29045, n_29046, n_29047, n_29048, n_29049, n_29050, n_29051, n_29052, n_29053, n_29054, n_29055, n_29056, n_29057, n_29058, n_29059, n_29060, n_29061, n_29062, n_29063, n_29064, n_29065, n_29066, n_29067, n_29068, n_29069, n_29070, n_29071, n_29072, n_29073, n_29074, n_29075, n_29076, n_29077, n_29078, n_29079, n_29080, n_29081, n_29082, n_29083, n_29084, n_29085, n_29086, n_29087, n_29088, n_29089, n_29090, n_29091, n_29092, n_29093, n_29094, n_29095, n_29096, n_29097, n_29098, n_29099, n_29100, n_29101, n_29102, n_29103, n_29104, n_29105, n_29106, n_29107, n_29108, n_29109, n_29110, n_29111, n_29112, n_29113, n_29114, n_29115, n_29116, n_29117, n_29118, n_29119, n_29120, n_29121, n_29122, n_29123, n_29124, n_29125, n_29126, n_29127, n_29128, n_29129, n_29130, n_29131, n_29132, n_29133, n_29134, n_29135, n_29136, n_29137, n_29138, n_29139, n_29140, n_29141, n_29142, n_29143, n_29144, n_29145, n_29146, n_29147, n_29148, n_29149, n_29150, n_29151, n_29152, n_29153, n_29154, n_29155, n_29156, n_29157, n_29158, n_29159, n_29160, n_29161, n_29162, n_29163, n_29164, n_29165, n_29166, n_29167, n_29168, n_29169, n_29170, n_29171, n_29172, n_29173, n_29174, n_29175, n_29176, n_29177, n_29178, n_29179, n_29180, n_29181, n_29182, n_29183, n_29184, n_29185, n_29186, n_29187, n_29188, n_29189, n_29190, n_29191, n_29192, n_29193, n_29194, n_29195, n_29196, n_29197, n_29198, n_29199, n_29200, n_29201, n_29202, n_29203, n_29204, n_29205, n_29206, n_29207, n_29208, n_29209, n_29210, n_29211, n_29212, n_29213, n_29214, n_29215, n_29216, n_29217, n_29218, n_29219, n_29220, n_29221, n_29222, n_29223, n_29224, n_29225, n_29226, n_29227, n_29228, n_29229, n_29230, n_29231, n_29232, n_29233, n_29234, n_29235, n_29236, n_29237, n_29238, n_29239, n_29240, n_29241, n_29242, n_29243, n_29244, n_29245, n_29246, n_29247, n_29248, n_29249, n_29250, n_29251, n_29252, n_29253, n_29254, n_29255, n_29256, n_29257, n_29258, n_29259, n_29260, n_29261, n_29262, n_29263, n_29264, n_29265, n_29266, n_29267, n_29268, n_29269, n_29270, n_29271, n_29272, n_29273, n_29274, n_29275, n_29276, n_29277, n_29278, n_29279, n_29280, n_29281, n_29282, n_29283, n_29284, n_29285, n_29286, n_29287, n_29288, n_29289, n_29290, n_29291, n_29292, n_29293, n_29294, n_29295, n_29296, n_29297, n_29298, n_29299, n_29300, n_29301, n_29302, n_29303, n_29304, n_29305, n_29306, n_29307, n_29308, n_29309, n_29310, n_29311, n_29312, n_29313, n_29314, n_29315, n_29316, n_29317, n_29318, n_29319, n_29320, n_29321, n_29322, n_29323, n_29324, n_29325, n_29326, n_29327, n_29328, n_29329, n_29330, n_29331, n_29332, n_29333, n_29334, n_29335, n_29336, n_29337, n_29338, n_29339, n_29340, n_29341, n_29342, n_29343, n_29344, n_29345, n_29346, n_29347, n_29348, n_29349, n_29350, n_29351, n_29352, n_29353, n_29354, n_29355, n_29356, n_29357, n_29358, n_29359, n_29360, n_29361, n_29362, n_29363, n_29364, n_29365, n_29366, n_29367, n_29368, n_29369, n_29370, n_29371, n_29372, n_29373, n_29374, n_29375, n_29376, n_29377, n_29378, n_29379, n_29380, n_29381, n_29382, n_29383, n_29384, n_29385, n_29386, n_29387, n_29388, n_29389, n_29390, n_29391, n_29392, n_29393, n_29394, n_29395, n_29396, n_29397, n_29398, n_29399, n_29400, n_29401, n_29402, n_29403, n_29404, n_29405, n_29406, n_29407, n_29408, n_29409, n_29410, n_29411, n_29412, n_29413, n_29414, n_29415, n_29416, n_29417, n_29418, n_29419, n_29420, n_29421, n_29422, n_29423, n_29424, n_29425, n_29426, n_29427, n_29428, n_29429, n_29430, n_29431, n_29432, n_29433, n_29434, n_29435, n_29436, n_29437, n_29438, n_29439, n_29440, n_29441, n_29442, n_29443, n_29444, n_29445, n_29446, n_29447, n_29448, n_29449, n_29450, n_29451, n_29452, n_29453, n_29454, n_29455, n_29456, n_29457, n_29458, n_29459, n_29460, n_29461, n_29462, n_29463, n_29464, n_29465, n_29466, n_29467, n_29468, n_29469, n_29470, n_29471, n_29472, n_29473, n_29474, n_29475, n_29476, n_29477, n_29478, n_29479, n_29480, n_29481, n_29482, n_29483, n_29484, n_29485, n_29486, n_29487, n_29488, n_29489, n_29490, n_29491, n_29492, n_29493, n_29494, n_29495, n_29496, n_29497, n_29498, n_29499, n_29500, n_29501, n_29502, n_29503, n_29504, n_29505, n_29506, n_29507, n_29508, n_29509, n_29510, n_29511, n_29512, n_29513, n_29514, n_29515, n_29516, n_29517, n_29518, n_29519, n_29520, n_29521, n_29522, n_29523, n_29524, n_29525, n_29526, n_29527, n_29528, n_29529, n_29530, n_29531, n_29532, n_29533, n_29534, n_29535, n_29536, n_29537, n_29538, n_29539, n_29540, n_29541, n_29542, n_29543, n_29544, n_29545, n_29546, n_29547, n_29548, n_29549, n_29550, n_29551, n_29552, n_29553, n_29554, n_29555, n_29556, n_29557, n_29558, n_29559, n_29560, n_29561, n_29562, n_29563, n_29564, n_29565, n_29566, n_29567, n_29568, n_29569, n_29570, n_29571, n_29572, n_29573, n_29574, n_29575, n_29576, n_29577, n_29578, n_29579, n_29580, n_29581, n_29582, n_29583, n_29584, n_29585, n_29586, n_29587, n_29588, n_29589, n_29590, n_29591, n_29592, n_29593, n_29594, n_29595, n_29596, n_29597, n_29598, n_29599, n_29600, n_29601, n_29602, n_29603, n_29604, n_29605, n_29606, n_29607, n_29608, n_29609, n_29610, n_29611, n_29612, n_29613, n_29614, n_29615, n_29616, n_29617, n_29618, n_29619, n_29620, n_29621, n_29622, n_29623, n_29624, n_29625, n_29626, n_29627, n_29628, n_29629, n_29630, n_29631, n_29632, n_29633, n_29634, n_29635, n_29636, n_29637, n_29638, n_29639, n_29640, n_29641, n_29642, n_29643, n_29644, n_29645, n_29646, n_29647, n_29648, n_29649, n_29650, n_29651, n_29652, n_29653, n_29654, n_29655, n_29656, n_29657, n_29658, n_29659, n_29660, n_29661, n_29662, n_29663, n_29664, n_29665, n_29666, n_29667, n_29668, n_29669, n_29670, n_29671, n_29672, n_29673, n_29674, n_29675, n_29676, n_29677, n_29678, n_29679, n_29680, n_29681, n_29682, n_29683, n_29684, n_29685, n_29686, n_29687, n_29688, n_29689, n_29690, n_29691, n_29692, n_29693, n_29694, n_29695, n_29696, n_29697, n_29698, n_29699, n_29700, n_29701, n_29702, n_29703, n_29704, n_29705, n_29706, n_29707, n_29708, n_29709, n_29710, n_29711, n_29712, n_29713, n_29714, n_29715, n_29716, n_29717, n_29718, n_29719, n_29720, n_29721, n_29722, n_29723, n_29724, n_29725, n_29726, n_29727, n_29728, n_29729, n_29730, n_29731, n_29732, n_29733, n_29734, n_29735, n_29736, n_29737, n_29738, n_29739, n_29740, n_29741, n_29742, n_29743, n_29744, n_29745, n_29746, n_29747, n_29748, n_29749, n_29750, n_29751, n_29752, n_29753, n_29754, n_29755, n_29756, n_29757, n_29758, n_29759, n_29760, n_29761, n_29762, n_29763, n_29764, n_29765, n_29766, n_29767, n_29768, n_29769, n_29770, n_29771, n_29772, n_29773, n_29774, n_29775, n_29776, n_29777, n_29778, n_29779, n_29780, n_29781, n_29782, n_29783, n_29784, n_29785, n_29786, n_29787, n_29788, n_29789, n_29790, n_29791, n_29792, n_29793, n_29794, n_29795, n_29796, n_29797, n_29798, n_29799, n_29800, n_29801, n_29802, n_29803, n_29804, n_29805, n_29806, n_29807, n_29808, n_29809, n_29810, n_29811, n_29812, n_29813, n_29814, n_29815, n_29816, n_29817, n_29818, n_29819, n_29820, n_29821, n_29822, n_29823, n_29824, n_29825, n_29826, n_29827, n_29828, n_29829, n_29830, n_29831, n_29832, n_29833, n_29834, n_29835, n_29836, n_29837, n_29838, n_29839, n_29840, n_29841, n_29842, n_29843, n_29844, n_29845, n_29846, n_29847, n_29848, n_29849, n_29850, n_29851, n_29852, n_29853, n_29854, n_29855, n_29856, n_29857, n_29858, n_29859, n_29860, n_29861, n_29862, n_29863, n_29864, n_29865, n_29866, n_29867, n_29868, n_29869, n_29870, n_29871, n_29872, n_29873, n_29874, n_29875, n_29876, n_29877, n_29878, n_29879, n_29880, n_29881, n_29882, n_29883, n_29884, n_29885, n_29886, n_29887, n_29888, n_29889, n_29890, n_29891, n_29892, n_29893, n_29894, n_29895, n_29896, n_29897, n_29898, n_29899, n_29900, n_29901, n_29902, n_29903, n_29904, n_29905, n_29906, n_29907, n_29908, n_29909, n_29910, n_29911, n_29912, n_29913, n_29914, n_29915, n_29916, n_29917, n_29918, n_29919, n_29920, n_29921, n_29922, n_29923, n_29924, n_29925, n_29926, n_29927, n_29928, n_29929, n_29930, n_29931, n_29932, n_29933, n_29934, n_29935, n_29936, n_29937, n_29938, n_29939, n_29940, n_29941, n_29942, n_29943, n_29944, n_29945, n_29946, n_29947, n_29948, n_29949, n_29950, n_29951, n_29952, n_29953, n_29954, n_29955, n_29956, n_29957, n_29958, n_29959, n_29960, n_29961, n_29962, n_29963, n_29964, n_29965, n_29966, n_29967, n_29968, n_29969, n_29970, n_29971, n_29972, n_29973, n_29974, n_29975, n_29976, n_29977, n_29978, n_29979, n_29980, n_29981, n_29982, n_29983, n_29984, n_29985, n_29986, n_29987, n_29988, n_29989, n_29990, n_29991, n_29992, n_29993, n_29994, n_29995, n_29996, n_29997, n_29998, n_29999, n_30000, n_30001, n_30002, n_30003, n_30004, n_30005, n_30006, n_30007, n_30008, n_30009, n_30010, n_30011, n_30012, n_30013, n_30014, n_30015, n_30016, n_30017, n_30018, n_30019, n_30020, n_30021, n_30022, n_30023, n_30024, n_30025, n_30026, n_30027, n_30028, n_30029, n_30030, n_30031, n_30032, n_30033, n_30034, n_30035, n_30036, n_30037, n_30038, n_30039, n_30040, n_30041, n_30042, n_30043, n_30044, n_30045, n_30046, n_30047, n_30048, n_30049, n_30050, n_30051, n_30052, n_30053, n_30054, n_30055, n_30056, n_30057, n_30058, n_30059, n_30060, n_30061, n_30062, n_30063, n_30064, n_30065, n_30066, n_30067, n_30068, n_30069, n_30070, n_30071, n_30072, n_30073, n_30074, n_30075, n_30076, n_30077, n_30078, n_30079, n_30080, n_30081, n_30082, n_30083, n_30084, n_30085, n_30086, n_30087, n_30088, n_30089, n_30090, n_30091, n_30092, n_30093, n_30094, n_30095, n_30096, n_30097, n_30098, n_30099, n_30100, n_30101, n_30102, n_30103, n_30104, n_30105, n_30106, n_30107, n_30108, n_30109, n_30110, n_30111, n_30112, n_30113, n_30114, n_30115, n_30116, n_30117, n_30118, n_30119, n_30120, n_30121, n_30122, n_30123, n_30124, n_30125, n_30126, n_30127, n_30128, n_30129, n_30130, n_30131, n_30132, n_30133, n_30134, n_30135, n_30136, n_30137, n_30138, n_30139, n_30140, n_30141, n_30142, n_30143, n_30144, n_30145, n_30146, n_30147, n_30148, n_30149, n_30150, n_30151, n_30152, n_30153, n_30154, n_30155, n_30156, n_30157, n_30158, n_30159, n_30160, n_30161, n_30162, n_30163, n_30164, n_30165, n_30166, n_30167, n_30168, n_30169, n_30170, n_30171, n_30172, n_30173, n_30174, n_30175, n_30176, n_30177, n_30178, n_30179, n_30180, n_30181, n_30182, n_30183, n_30184, n_30185, n_30186, n_30187, n_30188, n_30189, n_30190, n_30191, n_30192, n_30193, n_30194, n_30195, n_30196, n_30197, n_30198, n_30199, n_30200, n_30201, n_30202, n_30203, n_30204, n_30205, n_30206, n_30207, n_30208, n_30209, n_30210, n_30211, n_30212, n_30213, n_30214, n_30215, n_30216, n_30217, n_30218, n_30219, n_30220, n_30221, n_30222, n_30223, n_30224, n_30225, n_30226, n_30227, n_30228, n_30229, n_30230, n_30231, n_30232, n_30233, n_30234, n_30235, n_30236, n_30237, n_30238, n_30239, n_30240, n_30241, n_30242, n_30243, n_30244, n_30245, n_30246, n_30247, n_30248, n_30249, n_30250, n_30251, n_30252, n_30253, n_30254, n_30255, n_30256, n_30257, n_30258, n_30259, n_30260, n_30261, n_30262, n_30263, n_30264, n_30265, n_30266, n_30267, n_30268, n_30269, n_30270, n_30271, n_30272, n_30273, n_30274, n_30275, n_30276, n_30277, n_30278, n_30279, n_30280, n_30281, n_30282, n_30283, n_30284, n_30285, n_30286, n_30287, n_30288, n_30289, n_30290, n_30291, n_30292, n_30293, n_30294, n_30295, n_30296, n_30297, n_30298, n_30299, n_30300, n_30301, n_30302, n_30303, n_30304, n_30305, n_30306, n_30307, n_30308, n_30309, n_30310, n_30311, n_30312, n_30313, n_30314, n_30315, n_30316, n_30317, n_30318, n_30319, n_30320, n_30321, n_30322, n_30323, n_30324, n_30325, n_30326, n_30327, n_30328, n_30329, n_30330, n_30331, n_30332, n_30333, n_30334, n_30335, n_30336, n_30337, n_30338, n_30339, n_30340, n_30341, n_30342, n_30343, n_30344, n_30345, n_30346, n_30347, n_30348, n_30349, n_30350, n_30351, n_30352, n_30353, n_30354, n_30355, n_30356, n_30357, n_30358, n_30359, n_30360, n_30361, n_30362, n_30363, n_30364, n_30365, n_30366, n_30367, n_30368, n_30369, n_30370, n_30371, n_30372, n_30373, n_30374, n_30375, n_30376, n_30377, n_30378, n_30379, n_30380, n_30381, n_30382, n_30383, n_30384, n_30385, n_30386, n_30387, n_30388, n_30389, n_30390, n_30391, n_30392, n_30393, n_30394, n_30395, n_30396, n_30397, n_30398, n_30399, n_30400, n_30401, n_30402, n_30403, n_30404, n_30405, n_30406, n_30407, n_30408, n_30409, n_30410, n_30411, n_30412, n_30413, n_30414, n_30415, n_30416, n_30417, n_30418, n_30419, n_30420, n_30421, n_30422, n_30423, n_30424, n_30425, n_30426, n_30427, n_30428, n_30429, n_30430, n_30431, n_30432, n_30433, n_30434, n_30435, n_30436, n_30437, n_30438, n_30439, n_30440, n_30441, n_30442, n_30443, n_30444, n_30445, n_30446, n_30447, n_30448, n_30449, n_30450, n_30451, n_30452, n_30453, n_30454, n_30455, n_30456, n_30457, n_30458, n_30459, n_30460, n_30461, n_30462, n_30463, n_30464, n_30465, n_30466, n_30467, n_30468, n_30469, n_30470, n_30471, n_30472, n_30473, n_30474, n_30475, n_30476, n_30477, n_30478, n_30479, n_30480, n_30481, n_30482, n_30483, n_30484, n_30485, n_30486, n_30487, n_30488, n_30489, n_30490, n_30491, n_30492, n_30493, n_30494, n_30495, n_30496, n_30497, n_30498, n_30499, n_30500, n_30501, n_30502, n_30503, n_30504, n_30505, n_30506, n_30507, n_30508, n_30509, n_30510, n_30511, n_30512, n_30513, n_30514, n_30515, n_30516, n_30517, n_30518, n_30519, n_30520, n_30521, n_30522, n_30523, n_30524, n_30525, n_30526, n_30527, n_30528, n_30529, n_30530, n_30531, n_30532, n_30533, n_30534, n_30535, n_30536, n_30537, n_30538, n_30539, n_30540, n_30541, n_30542, n_30543, n_30544, n_30545, n_30546, n_30547, n_30548, n_30549, n_30550, n_30551, n_30552, n_30553, n_30554, n_30555, n_30556, n_30557, n_30558, n_30559, n_30560, n_30561, n_30562, n_30563, n_30564, n_30565, n_30566, n_30567, n_30568, n_30569, n_30570, n_30571, n_30572, n_30573, n_30574, n_30575, n_30576, n_30577, n_30578, n_30579, n_30580, n_30581, n_30582, n_30583, n_30584, n_30585, n_30586, n_30587, n_30588, n_30589, n_30590, n_30591, n_30592, n_30593, n_30594, n_30595, n_30596, n_30597, n_30598, n_30599, n_30600, n_30601, n_30602, n_30603, n_30604, n_30605, n_30606, n_30607, n_30608, n_30609, n_30610, n_30611, n_30612, n_30613, n_30614, n_30615, n_30616, n_30617, n_30618, n_30619, n_30620, n_30621, n_30622, n_30623, n_30624, n_30625, n_30626, n_30627, n_30628, n_30629, n_30630, n_30631, n_30632, n_30633, n_30634, n_30635, n_30636, n_30637, n_30638, n_30639, n_30640, n_30641, n_30642, n_30643, n_30644, n_30645, n_30646, n_30647, n_30648, n_30649, n_30650, n_30651, n_30652, n_30653, n_30654, n_30655, n_30656, n_30657, n_30658, n_30659, n_30660, n_30661, n_30662, n_30663, n_30664, n_30665, n_30666, n_30667, n_30668, n_30669, n_30670, n_30671, n_30672, n_30673, n_30674, n_30675, n_30676, n_30677, n_30678, n_30679, n_30680, n_30681, n_30682, n_30683, n_30684, n_30685, n_30686, n_30687, n_30688, n_30689, n_30690, n_30691, n_30692, n_30693, n_30694, n_30695, n_30696, n_30697, n_30698, n_30699, n_30700, n_30701, n_30702, n_30703, n_30704, n_30705, n_30706, n_30707, n_30708, n_30709, n_30710, n_30711, n_30712, n_30713, n_30714, n_30715, n_30716, n_30717, n_30718, n_30719, n_30720, n_30721, n_30722, n_30723, n_30724, n_30725, n_30726, n_30727, n_30728, n_30729, n_30730, n_30731, n_30732, n_30733, n_30734, n_30735, n_30736, n_30737, n_30738, n_30739, n_30740, n_30741, n_30742, n_30743, n_30744, n_30745, n_30746, n_30747, n_30748, n_30749, n_30750, n_30751, n_30752, n_30753, n_30754, n_30755, n_30756, n_30757, n_30758, n_30759, n_30760, n_30761, n_30762, n_30763, n_30764, n_30765, n_30766, n_30767, n_30768, n_30769, n_30770, n_30771, n_30772, n_30773, n_30774, n_30775, n_30776, n_30777, n_30778, n_30779, n_30780, n_30781, n_30782, n_30783, n_30784, n_30785, n_30786, n_30787, n_30788, n_30789, n_30790, n_30791, n_30792, n_30793, n_30794, n_30795, n_30796, n_30797, n_30798, n_30799, n_30800, n_30801, n_30802, n_30803, n_30804, n_30805, n_30806, n_30807, n_30808, n_30809, n_30810, n_30811, n_30812, n_30813, n_30814, n_30815, n_30816, n_30817, n_30818, n_30819, n_30820, n_30821, n_30822, n_30823, n_30824, n_30825, n_30826, n_30827, n_30828, n_30829, n_30830, n_30831, n_30832, n_30833, n_30834, n_30835, n_30836, n_30837, n_30838, n_30839, n_30840, n_30841, n_30842, n_30843, n_30844, n_30845, n_30846, n_30847, n_30848, n_30849, n_30850, n_30851, n_30852, n_30853, n_30854, n_30855, n_30856, n_30857, n_30858, n_30859, n_30860, n_30861, n_30862, n_30863, n_30864, n_30865, n_30866, n_30867, n_30868, n_30869, n_30870, n_30871, n_30872, n_30873, n_30874, n_30875, n_30876, n_30877, n_30878, n_30879, n_30880, n_30881, n_30882, n_30883, n_30884, n_30885, n_30886, n_30887, n_30888, n_30889, n_30890, n_30891, n_30892, n_30893, n_30894, n_30895, n_30896, n_30897, n_30898, n_30899, n_30900, n_30901, n_30902, n_30903, n_30904, n_30905, n_30906, n_30907, n_30908, n_30909, n_30910, n_30911, n_30912, n_30913, n_30914, n_30915, n_30916, n_30917, n_30918, n_30919, n_30920, n_30921, n_30922, n_30923, n_30924, n_30925, n_30926, n_30927, n_30928, n_30929, n_30930, n_30931, n_30932, n_30933, n_30934, n_30935, n_30936, n_30937, n_30938, n_30939, n_30940, n_30941, n_30942, n_30943, n_30944, n_30945, n_30946, n_30947, n_30948, n_30949, n_30950, n_30951, n_30952, n_30953, n_30954, n_30955, n_30956, n_30957, n_30958, n_30959, n_30960, n_30961, n_30962, n_30963, n_30964, n_30965, n_30966, n_30967, n_30968, n_30969, n_30970, n_30971, n_30972, n_30973, n_30974, n_30975, n_30976, n_30977, n_30978, n_30979, n_30980, n_30981, n_30982, n_30983, n_30984, n_30985, n_30986, n_30987, n_30988, n_30989, n_30990, n_30991, n_30992, n_30993, n_30994, n_30995, n_30996, n_30997, n_30998, n_30999, n_31000, n_31001, n_31002, n_31003, n_31004, n_31005, n_31006, n_31007, n_31008, n_31009, n_31010, n_31011, n_31012, n_31013, n_31014, n_31015, n_31016, n_31017, n_31018, n_31019, n_31020, n_31021, n_31022, n_31023, n_31024, n_31025, n_31026, n_31027, n_31028, n_31029, n_31030, n_31031, n_31032, n_31033, n_31034, n_31035, n_31036, n_31037, n_31038, n_31039, n_31040, n_31041, n_31042, n_31043, n_31044, n_31045, n_31046, n_31047, n_31048, n_31049, n_31050, n_31051, n_31052, n_31053, n_31054, n_31055, n_31056, n_31057, n_31058, n_31059, n_31060, n_31061, n_31062, n_31063, n_31064, n_31065, n_31066, n_31067, n_31068, n_31069, n_31070, n_31071, n_31072, n_31073, n_31074, n_31075, n_31076, n_31077, n_31078, n_31079, n_31080, n_31081, n_31082, n_31083, n_31084, n_31085, n_31086, n_31087, n_31088, n_31089, n_31090, n_31091, n_31092, n_31093, n_31094, n_31095, n_31096, n_31097, n_31098, n_31099, n_31100, n_31101, n_31102, n_31103, n_31104, n_31105, n_31106, n_31107, n_31108, n_31109, n_31110, n_31111, n_31112, n_31113, n_31114, n_31115, n_31116, n_31117, n_31118, n_31119, n_31120, n_31121, n_31122, n_31123, n_31124, n_31125, n_31126, n_31127, n_31128, n_31129, n_31130, n_31131, n_31132, n_31133, n_31134, n_31135, n_31136, n_31137, n_31138, n_31139, n_31140, n_31141, n_31142, n_31143, n_31144, n_31145, n_31146, n_31147, n_31148, n_31149, n_31150, n_31151, n_31152, n_31153, n_31154, n_31155, n_31156, n_31157, n_31158, n_31159, n_31160, n_31161, n_31162, n_31163, n_31164, n_31165, n_31166, n_31167, n_31168, n_31169, n_31170, n_31171, n_31172, n_31173, n_31174, n_31175, n_31176, n_31177, n_31178, n_31179, n_31180, n_31181, n_31182, n_31183, n_31184, n_31185, n_31186, n_31187, n_31188, n_31189, n_31190, n_31191, n_31192, n_31193, n_31194, n_31195, n_31196, n_31197, n_31198, n_31199, n_31200, n_31201, n_31202, n_31203, n_31204, n_31205, n_31206, n_31207, n_31208, n_31209, n_31210, n_31211, n_31212, n_31213, n_31214, n_31215, n_31216, n_31217, n_31218, n_31219, n_31220, n_31221, n_31222, n_31223, n_31224, n_31225, n_31226, n_31227, n_31228, n_31229, n_31230, n_31231, n_31232, n_31233, n_31234, n_31235, n_31236, n_31237, n_31238, n_31239, n_31240, n_31241, n_31242, n_31243, n_31244, n_31245, n_31246, n_31247, n_31248, n_31249, n_31250, n_31251, n_31252, n_31253, n_31254, n_31255, n_31256, n_31257, n_31258, n_31259, n_31260, n_31261, n_31262, n_31263, n_31264, n_31265, n_31266, n_31267, n_31268, n_31269, n_31270, n_31271, n_31272, n_31273, n_31274, n_31275, n_31276, n_31277, n_31278, n_31279, n_31280, n_31281, n_31282, n_31283, n_31284, n_31285, n_31286, n_31287, n_31288, n_31289, n_31290, n_31291, n_31292, n_31293, n_31294, n_31295, n_31296, n_31297, n_31298, n_31299, n_31300, n_31301, n_31302, n_31303, n_31304, n_31305, n_31306, n_31307, n_31308, n_31309, n_31310, n_31311, n_31312, n_31313, n_31314, n_31315, n_31316, n_31317, n_31318, n_31319, n_31320, n_31321, n_31322, n_31323, n_31324, n_31325, n_31326, n_31327, n_31328, n_31329, n_31330, n_31331, n_31332, n_31333, n_31334, n_31335, n_31336, n_31337, n_31338, n_31339, n_31340, n_31341, n_31342, n_31343, n_31344, n_31345, n_31346, n_31347, n_31348, n_31349, n_31350, n_31351, n_31352, n_31353, n_31354, n_31355, n_31356, n_31357, n_31358, n_31359, n_31360, n_31361, n_31362, n_31363, n_31364, n_31365, n_31366, n_31367, n_31368, n_31369, n_31370, n_31371, n_31372, n_31373, n_31374, n_31375, n_31376, n_31377, n_31378, n_31379, n_31380, n_31381, n_31382, n_31383, n_31384, n_31385, n_31386, n_31387, n_31388, n_31389, n_31390, n_31391, n_31392, n_31393, n_31394, n_31395, n_31396, n_31397, n_31398, n_31399, n_31400, n_31401, n_31402, n_31403, n_31404, n_31405, n_31406, n_31407, n_31408, n_31409, n_31410, n_31411, n_31412, n_31413, n_31414, n_31415, n_31416, n_31417, n_31418, n_31419, n_31420, n_31421, n_31422, n_31423, n_31424, n_31425, n_31426, n_31427, n_31428, n_31429, n_31430, n_31431, n_31432, n_31433, n_31434, n_31435, n_31436, n_31437, n_31438, n_31439, n_31440, n_31441, n_31442, n_31443, n_31444, n_31445, n_31446, n_31447, n_31448, n_31449, n_31450, n_31451, n_31452, n_31453, n_31454, n_31455, n_31456, n_31457, n_31458, n_31459, n_31460, n_31461, n_31462, n_31463, n_31464, n_31465, n_31466, n_31467, n_31468, n_31469, n_31470, n_31471, n_31472, n_31473, n_31474, n_31475, n_31476, n_31477, n_31478, n_31479, n_31480, n_31481, n_31482, n_31483, n_31484, n_31485, n_31486, n_31487, n_31488, n_31489, n_31490, n_31491, n_31492, n_31493, n_31494, n_31495, n_31496, n_31497, n_31498, n_31499, n_31500, n_31501, n_31502, n_31503, n_31504, n_31505, n_31506, n_31507, n_31508, n_31509, n_31510, n_31511, n_31512, n_31513, n_31514, n_31515, n_31516, n_31517, n_31518, n_31519, n_31520, n_31521, n_31522, n_31523, n_31524, n_31525, n_31526, n_31527, n_31528, n_31529, n_31530, n_31531, n_31532, n_31533, n_31534, n_31535, n_31536, n_31537, n_31538, n_31539, n_31540, n_31541, n_31542, n_31543, n_31544, n_31545, n_31546, n_31547, n_31548, n_31549, n_31550, n_31551, n_31552, n_31553, n_31554, n_31555, n_31556, n_31557, n_31558, n_31559, n_31560, n_31561, n_31562, n_31563, n_31564, n_31565, n_31566, n_31567, n_31568, n_31569, n_31570, n_31571, n_31572, n_31573, n_31574, n_31575, n_31576, n_31577, n_31578, n_31579, n_31580, n_31581, n_31582, n_31583, n_31584, n_31585, n_31586, n_31587, n_31588, n_31589, n_31590, n_31591, n_31592, n_31593, n_31594, n_31595, n_31596, n_31597, n_31598, n_31599, n_31600, n_31601, n_31602, n_31603, n_31604, n_31605, n_31606, n_31607, n_31608, n_31609, n_31610, n_31611, n_31612, n_31613, n_31614, n_31615, n_31616, n_31617, n_31618, n_31619, n_31620, n_31621, n_31622, n_31623, n_31624, n_31625, n_31626, n_31627, n_31628, n_31629, n_31630, n_31631, n_31632, n_31633, n_31634, n_31635, n_31636, n_31637, n_31638, n_31639, n_31640, n_31641, n_31642, n_31643, n_31644, n_31645, n_31646, n_31647, n_31648, n_31649, n_31650, n_31651, n_31652, n_31653, n_31654, n_31655, n_31656, n_31657, n_31658, n_31659, n_31660, n_31661, n_31662, n_31663, n_31664, n_31665, n_31666, n_31667, n_31668, n_31669, n_31670, n_31671, n_31672, n_31673, n_31674, n_31675, n_31676, n_31677, n_31678, n_31679, n_31680, n_31681, n_31682, n_31683, n_31684, n_31685, n_31686, n_31687, n_31688, n_31689, n_31690, n_31691, n_31692, n_31693, n_31694, n_31695, n_31696, n_31697, n_31698, n_31699, n_31700, n_31701, n_31702, n_31703, n_31704, n_31705, n_31706, n_31707, n_31708, n_31709, n_31710, n_31711, n_31712, n_31713, n_31714, n_31715, n_31716, n_31717, n_31718, n_31719, n_31720, n_31721, n_31722, n_31723, n_31724, n_31725, n_31726, n_31727, n_31728, n_31729, n_31730, n_31731, n_31732, n_31733, n_31734, n_31735, n_31736, n_31737, n_31738, n_31739, n_31740, n_31741, n_31742, n_31743, n_31744, n_31745, n_31746, n_31747, n_31748, n_31749, n_31750, n_31751, n_31752, n_31753, n_31754, n_31755, n_31756, n_31757, n_31758, n_31759, n_31760, n_31761, n_31762, n_31763, n_31764, n_31765, n_31766, n_31767, n_31768, n_31769, n_31770, n_31771, n_31772, n_31773, n_31774, n_31775, n_31776, n_31777, n_31778, n_31779, n_31780, n_31781, n_31782, n_31783, n_31784, n_31785, n_31786, n_31787, n_31788, n_31789, n_31790, n_31791, n_31792, n_31793, n_31794, n_31795, n_31796, n_31797, n_31798, n_31799, n_31800, n_31801, n_31802, n_31803, n_31804, n_31805, n_31806, n_31807, n_31808, n_31809, n_31810, n_31811, n_31812, n_31813, n_31814, n_31815, n_31816, n_31817, n_31818, n_31819, n_31820, n_31821, n_31822, n_31823, n_31824, n_31825, n_31826, n_31827, n_31828, n_31829, n_31830, n_31831, n_31832, n_31833, n_31834, n_31835, n_31836, n_31837, n_31838, n_31839, n_31840, n_31841, n_31842, n_31843, n_31844, n_31845, n_31846, n_31847, n_31848, n_31849, n_31850, n_31851, n_31852, n_31853, n_31854, n_31855, n_31856, n_31857, n_31858, n_31859, n_31860, n_31861, n_31862, n_31863, n_31864, n_31865, n_31866, n_31867, n_31868, n_31869, n_31870, n_31871, n_31872, n_31873, n_31874, n_31875, n_31876, n_31877, n_31878, n_31879, n_31880, n_31881, n_31882, n_31883, n_31884, n_31885, n_31886, n_31887, n_31888, n_31889, n_31890, n_31891, n_31892, n_31893, n_31894, n_31895, n_31896, n_31897, n_31898, n_31899, n_31900, n_31901, n_31902, n_31903, n_31904, n_31905, n_31906, n_31907, n_31908, n_31909, n_31910, n_31911, n_31912, n_31913, n_31914, n_31915, n_31916, n_31917, n_31918, n_31919, n_31920, n_31921, n_31922, n_31923, n_31924, n_31925, n_31926, n_31927, n_31928, n_31929, n_31930, n_31931, n_31932, n_31933, n_31934, n_31935, n_31936, n_31937, n_31938, n_31939, n_31940, n_31941, n_31942, n_31943, n_31944, n_31945, n_31946, n_31947, n_31948, n_31949, n_31950, n_31951, n_31952, n_31953, n_31954, n_31955, n_31956, n_31957, n_31958, n_31959, n_31960, n_31961, n_31962, n_31963, n_31964, n_31965, n_31966, n_31967, n_31968, n_31969, n_31970, n_31971, n_31972, n_31973, n_31974, n_31975, n_31976, n_31977, n_31978, n_31979, n_31980, n_31981, n_31982, n_31983, n_31984, n_31985, n_31986, n_31987, n_31988, n_31989, n_31990, n_31991, n_31992, n_31993, n_31994, n_31995, n_31996, n_31997, n_31998, n_31999, n_32000, n_32001, n_32002, n_32003, n_32004, n_32005, n_32006, n_32007, n_32008, n_32009, n_32010, n_32011, n_32012, n_32013, n_32014, n_32015, n_32016, n_32017, n_32018, n_32019, n_32020, n_32021, n_32022, n_32023, n_32024, n_32025, n_32026, n_32027, n_32028, n_32029, n_32030, n_32031, n_32032, n_32033, n_32034, n_32035, n_32036, n_32037, n_32038, n_32039, n_32040, n_32041, n_32042, n_32043, n_32044, n_32045, n_32046, n_32047, n_32048, n_32049, n_32050, n_32051, n_32052, n_32053, n_32054, n_32055, n_32056, n_32057, n_32058, n_32059, n_32060, n_32061, n_32062, n_32063, n_32064, n_32065, n_32066, n_32067, n_32068, n_32069, n_32070, n_32071, n_32072, n_32073, n_32074, n_32075, n_32076, n_32077, n_32078, n_32079, n_32080, n_32081, n_32082, n_32083, n_32084, n_32085, n_32086, n_32087, n_32088, n_32089, n_32090, n_32091, n_32092, n_32093, n_32094, n_32095, n_32096, n_32097, n_32098, n_32099, n_32100, n_32101, n_32102, n_32103, n_32104, n_32105, n_32106, n_32107, n_32108, n_32109, n_32110, n_32111, n_32112, n_32113, n_32114, n_32115, n_32116, n_32117, n_32118, n_32119, n_32120, n_32121, n_32122, n_32123, n_32124, n_32125, n_32126, n_32127, n_32128, n_32129, n_32130, n_32131, n_32132, n_32133, n_32134, n_32135, n_32136, n_32137, n_32138, n_32139, n_32140, n_32141, n_32142, n_32143, n_32144, n_32145, n_32146, n_32147, n_32148, n_32149, n_32150, n_32151, n_32152, n_32153, n_32154, n_32155, n_32156, n_32157, n_32158, n_32159, n_32160, n_32161, n_32162, n_32163, n_32164, n_32165, n_32166, n_32167, n_32168, n_32169, n_32170, n_32171, n_32172, n_32173, n_32174, n_32175, n_32176, n_32177, n_32178, n_32179, n_32180, n_32181, n_32182, n_32183, n_32184, n_32185, n_32186, n_32187, n_32188, n_32189, n_32190, n_32191, n_32192, n_32193, n_32194, n_32195, n_32196, n_32197, n_32198, n_32199, n_32200, n_32201, n_32202, n_32203, n_32204, n_32205, n_32206, n_32207, n_32208, n_32209, n_32210, n_32211, n_32212, n_32213, n_32214, n_32215, n_32216, n_32217, n_32218, n_32219, n_32220, n_32221, n_32222, n_32223, n_32224, n_32225, n_32226, n_32227, n_32228, n_32229, n_32230, n_32231, n_32232, n_32233, n_32234, n_32235, n_32236, n_32237, n_32238, n_32239, n_32240, n_32241, n_32242, n_32243, n_32244, n_32245, n_32246, n_32247, n_32248, n_32249, n_32250, n_32251, n_32252, n_32253, n_32254, n_32255, n_32256, n_32257, n_32258, n_32259, n_32260, n_32261, n_32262, n_32263, n_32264, n_32265, n_32266, n_32267, n_32268, n_32269, n_32270, n_32271, n_32272, n_32273, n_32274, n_32275, n_32276, n_32277, n_32278, n_32279, n_32280, n_32281, n_32282, n_32283, n_32284, n_32285, n_32286, n_32287, n_32288, n_32289, n_32290, n_32291, n_32292, n_32293, n_32294, n_32295, n_32296, n_32297, n_32298, n_32299, n_32300, n_32301, n_32302, n_32303, n_32304, n_32305, n_32306, n_32307, n_32308, n_32309, n_32310, n_32311, n_32312, n_32313, n_32314, n_32315, n_32316, n_32317, n_32318, n_32319, n_32320, n_32321, n_32322, n_32323, n_32324, n_32325, n_32326, n_32327, n_32328, n_32329, n_32330, n_32331, n_32332, n_32333, n_32334, n_32335, n_32336, n_32337, n_32338, n_32339, n_32340, n_32341, n_32342, n_32343, n_32344, n_32345, n_32346, n_32347, n_32348, n_32349, n_32350, n_32351, n_32352, n_32353, n_32354, n_32355, n_32356, n_32357, n_32358, n_32359, n_32360, n_32361, n_32362, n_32363, n_32364, n_32365, n_32366, n_32367, n_32368, n_32369, n_32370, n_32371, n_32372, n_32373, n_32374, n_32375, n_32376, n_32377, n_32378, n_32379, n_32380, n_32381, n_32382, n_32383, n_32384, n_32385, n_32386, n_32387, n_32388, n_32389, n_32390, n_32391, n_32392, n_32393, n_32394, n_32395, n_32396, n_32397, n_32398, n_32399, n_32400, n_32401, n_32402, n_32403, n_32404, n_32405, n_32406, n_32407, n_32408, n_32409, n_32410, n_32411, n_32412, n_32413, n_32414, n_32415, n_32416, n_32417, n_32418, n_32419, n_32420, n_32421, n_32422, n_32423, n_32424, n_32425, n_32426, n_32427, n_32428, n_32429, n_32430, n_32431, n_32432, n_32433, n_32434, n_32435, n_32436, n_32437, n_32438, n_32439, n_32440, n_32441, n_32442, n_32443, n_32444, n_32445, n_32446, n_32447, n_32448, n_32449, n_32450, n_32451, n_32452, n_32453, n_32454, n_32455, n_32456, n_32457, n_32458, n_32459, n_32460, n_32461, n_32462, n_32463, n_32464, n_32465, n_32466, n_32467, n_32468, n_32469, n_32470, n_32471, n_32472, n_32473, n_32474, n_32475, n_32476, n_32477, n_32478, n_32479, n_32480, n_32481, n_32482, n_32483, n_32484, n_32485, n_32486, n_32487, n_32488, n_32489, n_32490, n_32491, n_32492, n_32493, n_32494, n_32495, n_32496, n_32497, n_32498, n_32499, n_32500, n_32501, n_32502, n_32503, n_32504, n_32505, n_32506, n_32507, n_32508, n_32509, n_32510, n_32511, n_32512, n_32513, n_32514, n_32515, n_32516, n_32517, n_32518, n_32519, n_32520, n_32521, n_32522, n_32523, n_32524, n_32525, n_32526, n_32527, n_32528, n_32529, n_32530, n_32531, n_32532, n_32533, n_32534, n_32535, n_32536, n_32537, n_32538, n_32539, n_32540, n_32541, n_32542, n_32543, n_32544, n_32545, n_32546, n_32547, n_32548, n_32549, n_32550, n_32551, n_32552, n_32553, n_32554, n_32555, n_32556, n_32557, n_32558, n_32559, n_32560, n_32561, n_32562, n_32563, n_32564, n_32565, n_32566, n_32567, n_32568, n_32569, n_32570, n_32571, n_32572, n_32573, n_32574, n_32575, n_32576, n_32577, n_32578, n_32579, n_32580, n_32581, n_32582, n_32583, n_32584, n_32585, n_32586, n_32587, n_32588, n_32589, n_32590, n_32591, n_32592, n_32593, n_32594, n_32595, n_32596, n_32597, n_32598, n_32599, n_32600, n_32601, n_32602, n_32603, n_32604, n_32605, n_32606, n_32607, n_32608, n_32609, n_32610, n_32611, n_32612, n_32613, n_32614, n_32615, n_32616, n_32617, n_32618, n_32619, n_32620, n_32621, n_32622, n_32623, n_32624, n_32625, n_32626, n_32627, n_32628, n_32629, n_32630, n_32631, n_32632, n_32633, n_32634, n_32635, n_32636, n_32637, n_32638, n_32639, n_32640, n_32641, n_32642, n_32643, n_32644, n_32645, n_32646, n_32647, n_32648, n_32649, n_32650, n_32651, n_32652, n_32653, n_32654, n_32655, n_32656, n_32657, n_32658, n_32659, n_32660, n_32661, n_32662, n_32663, n_32664, n_32665, n_32666, n_32667, n_32668, n_32669, n_32670, n_32671, n_32672, n_32673, n_32674, n_32675, n_32676, n_32677, n_32678, n_32679, n_32680, n_32681, n_32682, n_32683, n_32684, n_32685, n_32686, n_32687, n_32688, n_32689, n_32690, n_32691, n_32692, n_32693, n_32694, n_32695, n_32696, n_32697, n_32698, n_32699, n_32700, n_32701, n_32702, n_32703, n_32704, n_32705, n_32706, n_32707, n_32708, n_32709, n_32710, n_32711, n_32712, n_32713, n_32714, n_32715, n_32716, n_32717, n_32718, n_32719, n_32720, n_32721, n_32722, n_32723, n_32724, n_32725, n_32726, n_32727, n_32728, n_32729, n_32730, n_32731, n_32732, n_32733, n_32734, n_32735, n_32736, n_32737, n_32738, n_32739, n_32740, n_32741, n_32742, n_32743, n_32744, n_32745, n_32746, n_32747, n_32748, n_32749, n_32750, n_32751, n_32752, n_32753, n_32754, n_32755, n_32756, n_32757, n_32758, n_32759, n_32760, n_32761, n_32762, n_32763, n_32764, n_32765, n_32766, n_32767, n_32768, n_32769, n_32770, n_32771, n_32772, n_32773, n_32774, n_32775, n_32776, n_32777, n_32778, n_32779, n_32780, n_32781, n_32782, n_32783, n_32784, n_32785, n_32786, n_32787, n_32788, n_32789, n_32790, n_32791, n_32792, n_32793, n_32794, n_32795, n_32796, n_32797, n_32798, n_32799, n_32800, n_32801, n_32802, n_32803, n_32804, n_32805, n_32806, n_32807, n_32808, n_32809, n_32810, n_32811, n_32812, n_32813, n_32814, n_32815, n_32816, n_32817, n_32818, n_32819, n_32820, n_32821, n_32822, n_32823, n_32824, n_32825, n_32826, n_32827, n_32828, n_32829, n_32830, n_32831, n_32832, n_32833, n_32834, n_32835, n_32836, n_32837, n_32838, n_32839, n_32840, n_32841, n_32842, n_32843, n_32844, n_32845, n_32846, n_32847, n_32848, n_32849, n_32850, n_32851, n_32852, n_32853, n_32854, n_32855, n_32856, n_32857, n_32858, n_32859, n_32860, n_32861, n_32862, n_32863, n_32864, n_32865, n_32866, n_32867, n_32868, n_32869, n_32870, n_32871, n_32872, n_32873, n_32874, n_32875, n_32876, n_32877, n_32878, n_32879, n_32880, n_32881, n_32882, n_32883, n_32884, n_32885, n_32886, n_32887, n_32888, n_32889, n_32890, n_32891, n_32892, n_32893, n_32894, n_32895, n_32896, n_32897, n_32898, n_32899, n_32900, n_32901, n_32902, n_32903, n_32904, n_32905, n_32906, n_32907, n_32908, n_32909, n_32910, n_32911, n_32912, n_32913, n_32914, n_32915, n_32916, n_32917, n_32918, n_32919, n_32920, n_32921, n_32922, n_32923, n_32924, n_32925, n_32926, n_32927, n_32928, n_32929, n_32930, n_32931, n_32932, n_32933, n_32934, n_32935, n_32936, n_32937, n_32938, n_32939, n_32940, n_32941, n_32942, n_32943, n_32944, n_32945, n_32946, n_32947, n_32948, n_32949, n_32950, n_32951, n_32952, n_32953, n_32954, n_32955, n_32956, n_32957, n_32958, n_32959, n_32960, n_32961, n_32962, n_32963, n_32964, n_32965, n_32966, n_32967, n_32968, n_32969, n_32970, n_32971, n_32972, n_32973, n_32974, n_32975, n_32976, n_32977, n_32978, n_32979, n_32980, n_32981, n_32982, n_32983, n_32984, n_32985, n_32986, n_32987, n_32988, n_32989, n_32990, n_32991, n_32992, n_32993, n_32994, n_32995, n_32996, n_32997, n_32998, n_32999, n_33000, n_33001, n_33002, n_33003, n_33004, n_33005, n_33006, n_33007, n_33008, n_33009, n_33010, n_33011, n_33012, n_33013, n_33014, n_33015, n_33016, n_33017, n_33018, n_33019, n_33020, n_33021, n_33022, n_33023, n_33024, n_33025, n_33026, n_33027, n_33028, n_33029, n_33030, n_33031, n_33032, n_33033, n_33034, n_33035, n_33036, n_33037, n_33038, n_33039, n_33040, n_33041, n_33042, n_33043, n_33044, n_33045, n_33046, n_33047, n_33048, n_33049, n_33050, n_33051, n_33052, n_33053, n_33054, n_33055, n_33056, n_33057, n_33058, n_33059, n_33060, n_33061, n_33062, n_33063, n_33064, n_33065, n_33066, n_33067, n_33068, n_33069, n_33070, n_33071, n_33072, n_33073, n_33074, n_33075, n_33076, n_33077, n_33078, n_33079, n_33080, n_33081, n_33082, n_33083, n_33084, n_33085, n_33086, n_33087, n_33088, n_33089, n_33090, n_33091, n_33092, n_33093, n_33094, n_33095, n_33096, n_33097, n_33098, n_33099, n_33100, n_33101, n_33102, n_33103, n_33104, n_33105, n_33106, n_33107, n_33108, n_33109, n_33110, n_33111, n_33112, n_33113, n_33114, n_33115, n_33116, n_33117, n_33118, n_33119, n_33120, n_33121, n_33122, n_33123, n_33124, n_33125, n_33126, n_33127, n_33128, n_33129, n_33130, n_33131, n_33132, n_33133, n_33134, n_33135, n_33136, n_33137, n_33138, n_33139, n_33140, n_33141, n_33142, n_33143, n_33144, n_33145, n_33146, n_33147, n_33148, n_33149, n_33150, n_33151, n_33152, n_33153, n_33154, n_33155, n_33156, n_33157, n_33158, n_33159, n_33160, n_33161, n_33162, n_33163, n_33164, n_33165, n_33166, n_33167, n_33168, n_33169, n_33170, n_33171, n_33172, n_33173, n_33174, n_33175, n_33176, n_33177, n_33178, n_33179, n_33180, n_33181, n_33182, n_33183, n_33184, n_33185, n_33186, n_33187, n_33188, n_33189, n_33190, n_33191, n_33192, n_33193, n_33194, n_33195, n_33196, n_33197, n_33198, n_33199, n_33200, n_33201, n_33202, n_33203, n_33204, n_33205, n_33206, n_33207, n_33208, n_33209, n_33210, n_33211, n_33212, n_33213, n_33214, n_33215, n_33216, n_33217, n_33218, n_33219, n_33220, n_33221, n_33222, n_33223, n_33224, n_33225, n_33226, n_33227, n_33228, n_33229, n_33230, n_33231, n_33232, n_33233, n_33234, n_33235, n_33236, n_33237, n_33238, n_33239, n_33240, n_33241, n_33242, n_33243, n_33244, n_33245, n_33246, n_33247, n_33248, n_33249, n_33250, n_33251, n_33252, n_33253, n_33254, n_33255, n_33256, n_33257, n_33258, n_33259, n_33260, n_33261, n_33262, n_33263, n_33264, n_33265, n_33266, n_33267, n_33268, n_33269, n_33270, n_33271, n_33272, n_33273, n_33274, n_33275, n_33276, n_33277, n_33278, n_33279, n_33280, n_33281, n_33282, n_33283, n_33284, n_33285, n_33286, n_33287, n_33288, n_33289, n_33290, n_33291, n_33292, n_33293, n_33294, n_33295, n_33296, n_33297, n_33298, n_33299, n_33300, n_33301, n_33302, n_33303, n_33304, n_33305, n_33306, n_33307, n_33308, n_33309, n_33310, n_33311, n_33312, n_33313, n_33314, n_33315, n_33316, n_33317, n_33318, n_33319, n_33320, n_33321, n_33322, n_33323, n_33324, n_33325, n_33326, n_33327, n_33328, n_33329, n_33330, n_33331, n_33332, n_33333, n_33334, n_33335, n_33336, n_33337, n_33338, n_33339, n_33340, n_33341, n_33342, n_33343, n_33344, n_33345, n_33346, n_33347, n_33348, n_33349, n_33350, n_33351, n_33352, n_33353, n_33354, n_33355, n_33356, n_33357, n_33358, n_33359, n_33360, n_33361, n_33362, n_33363, n_33364, n_33365, n_33366, n_33367, n_33368, n_33369, n_33370, n_33371, n_33372, n_33373, n_33374, n_33375, n_33376, n_33377, n_33378, n_33379, n_33380, n_33381, n_33382, n_33383, n_33384, n_33385, n_33386, n_33387, n_33388, n_33389, n_33390, n_33391, n_33392, n_33393, n_33394, n_33395, n_33396, n_33397, n_33398, n_33399, n_33400, n_33401, n_33402, n_33403, n_33404, n_33405, n_33406, n_33407, n_33408, n_33409, n_33410, n_33411, n_33412, n_33413, n_33414, n_33415, n_33416, n_33417, n_33418, n_33419, n_33420, n_33421, n_33422, n_33423, n_33424, n_33425, n_33426, n_33427, n_33428, n_33429, n_33430, n_33431, n_33432, n_33433, n_33434, n_33435, n_33436, n_33437, n_33438, n_33439, n_33440, n_33441, n_33442, n_33443, n_33444, n_33445, n_33446, n_33447, n_33448, n_33449, n_33450, n_33451, n_33452, n_33453, n_33454, n_33455, n_33456, n_33457, n_33458, n_33459, n_33460, n_33461, n_33462, n_33463, n_33464, n_33465, n_33466, n_33467, n_33468, n_33469, n_33470, n_33471, n_33472, n_33473, n_33474, n_33475, n_33476, n_33477, n_33478, n_33479, n_33480, n_33481, n_33482, n_33483, n_33484, n_33485, n_33486, n_33487, n_33488, n_33489, n_33490, n_33491, n_33492, n_33493, n_33494, n_33495, n_33496, n_33497, n_33498, n_33499, n_33500, n_33501, n_33502, n_33503, n_33504, n_33505, n_33506, n_33507, n_33508, n_33509, n_33510, n_33511, n_33512, n_33513, n_33514, n_33515, n_33516, n_33517, n_33518, n_33519, n_33520, n_33521, n_33522, n_33523, n_33524, n_33525, n_33526, n_33527, n_33528, n_33529, n_33530, n_33531, n_33532, n_33533, n_33534, n_33535, n_33536, n_33537, n_33538, n_33539, n_33540, n_33541, n_33542, n_33543, n_33544, n_33545, n_33546, n_33547, n_33548, n_33549, n_33550, n_33551, n_33552, n_33553, n_33554, n_33555, n_33556, n_33557, n_33558, n_33559, n_33560, n_33561, n_33562, n_33563, n_33564, n_33565, n_33566, n_33567, n_33568, n_33569, n_33570, n_33571, n_33572, n_33573, n_33574, n_33575, n_33576, n_33577, n_33578, n_33579, n_33580, n_33581, n_33582, n_33583, n_33584, n_33585, n_33586, n_33587, n_33588, n_33589, n_33590, n_33591, n_33592, n_33593, n_33594, n_33595, n_33596, n_33597, n_33598, n_33599, n_33600, n_33601, n_33602, n_33603, n_33604, n_33605, n_33606, n_33607, n_33608, n_33609, n_33610, n_33611, n_33612, n_33613, n_33614, n_33615, n_33616, n_33617, n_33618, n_33619, n_33620, n_33621, n_33622, n_33623, n_33624, n_33625, n_33626, n_33627, n_33628, n_33629, n_33630, n_33631, n_33632, n_33633, n_33634, n_33635, n_33636, n_33637, n_33638, n_33639, n_33640, n_33641, n_33642, n_33643, n_33644, n_33645, n_33646, n_33647, n_33648, n_33649, n_33650, n_33651, n_33652, n_33653, n_33654, n_33655, n_33656, n_33657, n_33658, n_33659, n_33660, n_33661, n_33662, n_33663, n_33664, n_33665, n_33666, n_33667, n_33668, n_33669, n_33670, n_33671, n_33672, n_33673, n_33674, n_33675, n_33676, n_33677, n_33678, n_33679, n_33680, n_33681, n_33682, n_33683, n_33684, n_33685, n_33686, n_33687, n_33688, n_33689, n_33690, n_33691, n_33692, n_33693, n_33694, n_33695, n_33696, n_33697, n_33698, n_33699, n_33700, n_33701, n_33702, n_33703, n_33704, n_33705, n_33706, n_33707, n_33708, n_33709, n_33710, n_33711, n_33712, n_33713, n_33714, n_33715, n_33716, n_33717, n_33718, n_33719, n_33720, n_33721, n_33722, n_33723, n_33724, n_33725, n_33726, n_33727, n_33728, n_33729, n_33730, n_33731, n_33732, n_33733, n_33734, n_33735, n_33736, n_33737, n_33738, n_33739, n_33740, n_33741, n_33742, n_33743, n_33744, n_33745, n_33746, n_33747, n_33748, n_33749, n_33750, n_33751, n_33752, n_33753, n_33754, n_33755, n_33756, n_33757, n_33758, n_33759, n_33760, n_33761, n_33762, n_33763, n_33764, n_33765, n_33766, n_33767, n_33768, n_33769, n_33770, n_33771, n_33772, n_33773, n_33774, n_33775, n_33776, n_33777, n_33778, n_33779, n_33780, n_33781, n_33782, n_33783, n_33784, n_33785, n_33786, n_33787, n_33788, n_33789, n_33790, n_33791, n_33792, n_33793, n_33794, n_33795, n_33796, n_33797, n_33798, n_33799, n_33800, n_33801, n_33802, n_33803, n_33804, n_33805, n_33806, n_33807, n_33808, n_33809, n_33810, n_33811, n_33812, n_33813, n_33814, n_33815, n_33816, n_33817, n_33818, n_33819, n_33820, n_33821, n_33822, n_33823, n_33824, n_33825, n_33826, n_33827, n_33828, n_33829, n_33830, n_33831, n_33832, n_33833, n_33834, n_33835, n_33836, n_33837, n_33838, n_33839, n_33840, n_33841, n_33842, n_33843, n_33844, n_33845, n_33846, n_33847, n_33848, n_33849, n_33850, n_33851, n_33852, n_33853, n_33854, n_33855, n_33856, n_33857, n_33858, n_33859, n_33860, n_33861, n_33862, n_33863, n_33864, n_33865, n_33866, n_33867, n_33868, n_33869, n_33870, n_33871, n_33872, n_33873, n_33874, n_33875, n_33876, n_33877, n_33878, n_33879, n_33880, n_33881, n_33882, n_33883, n_33884, n_33885, n_33886, n_33887, n_33888, n_33889, n_33890, n_33891, n_33892, n_33893, n_33894, n_33895, n_33896, n_33897, n_33898, n_33899, n_33900, n_33901, n_33902, n_33903, n_33904, n_33905, n_33906, n_33907, n_33908, n_33909, n_33910, n_33911, n_33912, n_33913, n_33914, n_33915, n_33916, n_33917, n_33918, n_33919, n_33920, n_33921, n_33922, n_33923, n_33924, n_33925, n_33926, n_33927, n_33928, n_33929, n_33930, n_33931, n_33932, n_33933, n_33934, n_33935, n_33936, n_33937, n_33938, n_33939, n_33940, n_33941, n_33942, n_33943, n_33944, n_33945, n_33946, n_33947, n_33948, n_33949, n_33950, n_33951, n_33952, n_33953, n_33954, n_33955, n_33956, n_33957, n_33958, n_33959, n_33960, n_33961, n_33962, n_33963, n_33964, n_33965, n_33966, n_33967, n_33968, n_33969, n_33970, n_33971, n_33972, n_33973, n_33974, n_33975, n_33976, n_33977, n_33978, n_33979, n_33980, n_33981, n_33982, n_33983, n_33984, n_33985, n_33986, n_33987, n_33988, n_33989, n_33990, n_33991, n_33992, n_33993, n_33994, n_33995, n_33996, n_33997, n_33998, n_33999, n_34000, n_34001, n_34002, n_34003, n_34004, n_34005, n_34006, n_34007, n_34008, n_34009, n_34010, n_34011, n_34012, n_34013, n_34014, n_34015, n_34016, n_34017, n_34018, n_34019, n_34020, n_34021, n_34022, n_34023, n_34024, n_34025, n_34026, n_34027, n_34028, n_34029, n_34030, n_34031, n_34032, n_34033, n_34034, n_34035, n_34036, n_34037, n_34038, n_34039, n_34040, n_34041, n_34042, n_34043, n_34044, n_34045, n_34046, n_34047, n_34048, n_34049, n_34050, n_34051, n_34052, n_34053, n_34054, n_34055, n_34056, n_34057, n_34058, n_34059, n_34060, n_34061, n_34062, n_34063, n_34064, n_34065, n_34066, n_34067, n_34068, n_34069, n_34070, n_34071, n_34072, n_34073, n_34074, n_34075, n_34076, n_34077, n_34078, n_34079, n_34080, n_34081, n_34082, n_34083, n_34084, n_34085, n_34086, n_34087, n_34088, n_34089, n_34090, n_34091, n_34092, n_34093, n_34094, n_34095, n_34096, n_34097, n_34098, n_34099, n_34100, n_34101, n_34102, n_34103, n_34104, n_34105, n_34106, n_34107, n_34108, n_34109, n_34110, n_34111, n_34112, n_34113, n_34114, n_34115, n_34116, n_34117, n_34118, n_34119, n_34120, n_34121, n_34122, n_34123, n_34124, n_34125, n_34126, n_34127, n_34128, n_34129, n_34130, n_34131, n_34132, n_34133, n_34134, n_34135, n_34136, n_34137, n_34138, n_34139, n_34140, n_34141, n_34142, n_34143, n_34144, n_34145, n_34146, n_34147, n_34148, n_34149, n_34150, n_34151, n_34152, n_34153, n_34154, n_34155, n_34156, n_34157, n_34158, n_34159, n_34160, n_34161, n_34162, n_34163, n_34164, n_34165, n_34166, n_34167, n_34168, n_34169, n_34170, n_34171, n_34172, n_34173, n_34174, n_34175, n_34176, n_34177, n_34178, n_34179, n_34180, n_34181, n_34182, n_34183, n_34184, n_34185, n_34186, n_34187, n_34188, n_34189, n_34190, n_34191, n_34192, n_34193, n_34194, n_34195, n_34196, n_34197, n_34198, n_34199, n_34200, n_34201, n_34202, n_34203, n_34204, n_34205, n_34206, n_34207, n_34208, n_34209, n_34210, n_34211, n_34212, n_34213, n_34214, n_34215, n_34216, n_34217, n_34218, n_34219, n_34220, n_34221, n_34222, n_34223, n_34224, n_34225, n_34226, n_34227, n_34228, n_34229, n_34230, n_34231, n_34232, n_34233, n_34234, n_34235, n_34236, n_34237, n_34238, n_34239, n_34240, n_34241, n_34242, n_34243, n_34244, n_34245, n_34246, n_34247, n_34248, n_34249, n_34250, n_34251, n_34252, n_34253, n_34254, n_34255, n_34256, n_34257, n_34258, n_34259, n_34260, n_34261, n_34262, n_34263, n_34264, n_34265, n_34266, n_34267, n_34268, n_34269, n_34270, n_34271, n_34272, n_34273, n_34274, n_34275, n_34276, n_34277, n_34278, n_34279, n_34280, n_34281, n_34282, n_34283, n_34284, n_34285, n_34286, n_34287, n_34288, n_34289, n_34290, n_34291, n_34292, n_34293, n_34294, n_34295, n_34296, n_34297, n_34298, n_34299, n_34300, n_34301, n_34302, n_34303, n_34304, n_34305, n_34306, n_34307, n_34308, n_34309, n_34310, n_34311, n_34312, n_34313, n_34314, n_34315, n_34316, n_34317, n_34318, n_34319, n_34320, n_34321, n_34322, n_34323, n_34324, n_34325, n_34326, n_34327, n_34328, n_34329, n_34330, n_34331, n_34332, n_34333, n_34334, n_34335, n_34336, n_34337, n_34338, n_34339, n_34340, n_34341, n_34342, n_34343, n_34344, n_34345, n_34346, n_34347, n_34348, n_34349, n_34350, n_34351, n_34352, n_34353, n_34354, n_34355, n_34356, n_34357, n_34358, n_34359, n_34360, n_34361, n_34362, n_34363, n_34364, n_34365, n_34366, n_34367, n_34368, n_34369, n_34370, n_34371, n_34372, n_34373, n_34374, n_34375, n_34376, n_34377, n_34378, n_34379, n_34380, n_34381, n_34382, n_34383, n_34384, n_34385, n_34386, n_34387, n_34388, n_34389, n_34390, n_34391, n_34392, n_34393, n_34394, n_34395, n_34396, n_34397, n_34398, n_34399, n_34400, n_34401, n_34402, n_34403, n_34404, n_34405, n_34406, n_34407, n_34408, n_34409, n_34410, n_34411, n_34412, n_34413, n_34414, n_34415, n_34416, n_34417, n_34418, n_34419, n_34420, n_34421, n_34422, n_34423, n_34424, n_34425, n_34426, n_34427, n_34428, n_34429, n_34430, n_34431, n_34432, n_34433, n_34434, n_34435, n_34436, n_34437, n_34438, n_34439, n_34440, n_34441, n_34442, n_34443, n_34444, n_34445, n_34446, n_34447, n_34448, n_34449, n_34450, n_34451, n_34452, n_34453, n_34454, n_34455, n_34456, n_34457, n_34458, n_34459, n_34460, n_34461, n_34462, n_34463, n_34464, n_34465, n_34466, n_34467, n_34468, n_34469, n_34470, n_34471, n_34472, n_34473, n_34474, n_34475, n_34476, n_34477, n_34478, n_34479, n_34480, n_34481, n_34482, n_34483, n_34484, n_34485, n_34486, n_34487, n_34488, n_34489, n_34490, n_34491, n_34492, n_34493, n_34494, n_34495, n_34496, n_34497, n_34498, n_34499, n_34500, n_34501, n_34502, n_34503, n_34504, n_34505, n_34506, n_34507, n_34508, n_34509, n_34510, n_34511, n_34512, n_34513, n_34514, n_34515, n_34516, n_34517, n_34518, n_34519, n_34520, n_34521, n_34522, n_34523, n_34524, n_34525, n_34526, n_34527, n_34528, n_34529, n_34530, n_34531, n_34532, n_34533, n_34534, n_34535, n_34536, n_34537, n_34538, n_34539, n_34540, n_34541, n_34542, n_34543, n_34544, n_34545, n_34546, n_34547, n_34548, n_34549, n_34550, n_34551, n_34552, n_34553, n_34554, n_34555, n_34556, n_34557, n_34558, n_34559, n_34560, n_34561, n_34562, n_34563, n_34564, n_34565, n_34566, n_34567, n_34568, n_34569, n_34570, n_34571, n_34572, n_34573, n_34574, n_34575, n_34576, n_34577, n_34578, n_34579, n_34580, n_34581, n_34582, n_34583, n_34584, n_34585, n_34586, n_34587, n_34588, n_34589, n_34590, n_34591, n_34592, n_34593, n_34594, n_34595, n_34596, n_34597, n_34598, n_34599, n_34600, n_34601, n_34602, n_34603, n_34604, n_34605, n_34606, n_34607, n_34608, n_34609, n_34610, n_34611, n_34612, n_34613, n_34614, n_34615, n_34616, n_34617, n_34618, n_34619, n_34620, n_34621, n_34622, n_34623, n_34624, n_34625, n_34626, n_34627, n_34628, n_34629, n_34630, n_34631, n_34632, n_34633, n_34634, n_34635, n_34636, n_34637, n_34638, n_34639, n_34640, n_34641, n_34642, n_34643, n_34644, n_34645, n_34646, n_34647, n_34648, n_34649, n_34650, n_34651, n_34652, n_34653, n_34654, n_34655, n_34656, n_34657, n_34658, n_34659, n_34660, n_34661, n_34662, n_34663, n_34664, n_34665, n_34666, n_34667, n_34668, n_34669, n_34670, n_34671, n_34672, n_34673, n_34674, n_34675, n_34676, n_34677, n_34678, n_34679, n_34680, n_34681, n_34682, n_34683, n_34684, n_34685, n_34686, n_34687, n_34688, n_34689, n_34690, n_34691, n_34692, n_34693, n_34694, n_34695, n_34696, n_34697, n_34698, n_34699, n_34700, n_34701, n_34702, n_34703, n_34704, n_34705, n_34706, n_34707, n_34708, n_34709, n_34710, n_34711, n_34712, n_34713, n_34714, n_34715, n_34716, n_34717, n_34718, n_34719, n_34720, n_34721, n_34722, n_34723, n_34724, n_34725, n_34726, n_34727, n_34728, n_34729, n_34730, n_34731, n_34732, n_34733, n_34734, n_34735, n_34736, n_34737, n_34738, n_34739, n_34740, n_34741, n_34742, n_34743, n_34744, n_34745, n_34746, n_34747, n_34748, n_34749, n_34750, n_34751, n_34752, n_34753, n_34754, n_34755, n_34756, n_34757, n_34758, n_34759, n_34760, n_34761, n_34762, n_34763, n_34764, n_34765, n_34766, n_34767, n_34768, n_34769, n_34770, n_34771, n_34772, n_34773, n_34774, n_34775, n_34776, n_34777, n_34778, n_34779, n_34780, n_34781, n_34782, n_34783, n_34784, n_34785, n_34786, n_34787, n_34788, n_34789, n_34790, n_34791, n_34792, n_34793, n_34794, n_34795, n_34796, n_34797, n_34798, n_34799, n_34800, n_34801, n_34802, n_34803, n_34804, n_34805, n_34806, n_34807, n_34808, n_34809, n_34810, n_34811, n_34812, n_34813, n_34814, n_34815, n_34816, n_34817, n_34818, n_34819, n_34820, n_34821, n_34822, n_34823, n_34824, n_34825, n_34826, n_34827, n_34828, n_34829, n_34830, n_34831, n_34832, n_34833, n_34834, n_34835, n_34836, n_34837, n_34838, n_34839, n_34840, n_34841, n_34842, n_34843, n_34844, n_34845, n_34846, n_34847, n_34848, n_34849, n_34850, n_34851, n_34852, n_34853, n_34854, n_34855, n_34856, n_34857, n_34858, n_34859, n_34860, n_34861, n_34862, n_34863, n_34864, n_34865, n_34866, n_34867, n_34868, n_34869, n_34870, n_34871, n_34872, n_34873, n_34874, n_34875, n_34876, n_34877, n_34878, n_34879, n_34880, n_34881, n_34882, n_34883, n_34884, n_34885, n_34886, n_34887, n_34888, n_34889, n_34890, n_34891, n_34892, n_34893, n_34894, n_34895, n_34896, n_34897, n_34898, n_34899, n_34900, n_34901, n_34902, n_34903, n_34904, n_34905, n_34906, n_34907, n_34908, n_34909, n_34910, n_34911, n_34912, n_34913, n_34914, n_34915, n_34916, n_34917, n_34918, n_34919, n_34920, n_34921, n_34922, n_34923, n_34924, n_34925, n_34926, n_34927, n_34928, n_34929, n_34930, n_34931, n_34932, n_34933, n_34934, n_34935, n_34936, n_34937, n_34938, n_34939, n_34940, n_34941, n_34942, n_34943, n_34944, n_34945, n_34946, n_34947, n_34948, n_34949, n_34950, n_34951, n_34952, n_34953, n_34954, n_34955, n_34956, n_34957, n_34958, n_34959, n_34960, n_34961, n_34962, n_34963, n_34964, n_34965, n_34966, n_34967, n_34968, n_34969, n_34970, n_34971, n_34972, n_34973, n_34974, n_34975, n_34976, n_34977, n_34978, n_34979, n_34980, n_34981, n_34982, n_34983, n_34984, n_34985, n_34986, n_34987, n_34988, n_34989, n_34990, n_34991, n_34992, n_34993, n_34994, n_34995, n_34996, n_34997, n_34998, n_34999, n_35000, n_35001, n_35002, n_35003, n_35004, n_35005, n_35006, n_35007, n_35008, n_35009, n_35010, n_35011, n_35012, n_35013, n_35014, n_35015, n_35016, n_35017, n_35018, n_35019, n_35020, n_35021, n_35022, n_35023, n_35024, n_35025, n_35026, n_35027, n_35028, n_35029, n_35030, n_35031, n_35032, n_35033, n_35034, n_35035, n_35036, n_35037, n_35038, n_35039, n_35040, n_35041, n_35042, n_35043, n_35044, n_35045, n_35046, n_35047, n_35048, n_35049, n_35050, n_35051, n_35052, n_35053, n_35054, n_35055, n_35056, n_35057, n_35058, n_35059, n_35060, n_35061, n_35062, n_35063, n_35064, n_35065, n_35066, n_35067, n_35068, n_35069, n_35070, n_35071, n_35072, n_35073, n_35074, n_35075, n_35076, n_35077, n_35078, n_35079, n_35080, n_35081, n_35082, n_35083, n_35084, n_35085, n_35086, n_35087, n_35088, n_35089, n_35090, n_35091, n_35092, n_35093, n_35094, n_35095, n_35096, n_35097, n_35098, n_35099, n_35100, n_35101, n_35102, n_35103, n_35104, n_35105, n_35106, n_35107, n_35108, n_35109, n_35110, n_35111, n_35112, n_35113, n_35114, n_35115, n_35116, n_35117, n_35118, n_35119, n_35120, n_35121, n_35122, n_35123, n_35124, n_35125, n_35126, n_35127, n_35128, n_35129, n_35130, n_35131, n_35132, n_35133, n_35134, n_35135, n_35136, n_35137, n_35138, n_35139, n_35140, n_35141, n_35142, n_35143, n_35144, n_35145, n_35146, n_35147, n_35148, n_35149, n_35150, n_35151, n_35152, n_35153, n_35154, n_35155, n_35156, n_35157, n_35158, n_35159, n_35160, n_35161, n_35162, n_35163, n_35164, n_35165, n_35166, n_35167, n_35168, n_35169, n_35170, n_35171, n_35172, n_35173, n_35174, n_35175, n_35176, n_35177, n_35178, n_35179, n_35180, n_35181, n_35182, n_35183, n_35184, n_35185, n_35186, n_35187, n_35188, n_35189, n_35190, n_35191, n_35192, n_35193, n_35194, n_35195, n_35196, n_35197, n_35198, n_35199, n_35200, n_35201, n_35202, n_35203, n_35204, n_35205, n_35206, n_35207, n_35208, n_35209, n_35210, n_35211, n_35212, n_35213, n_35214, n_35215, n_35216, n_35217, n_35218, n_35219, n_35220, n_35221, n_35222, n_35223, n_35224, n_35225, n_35226, n_35227, n_35228, n_35229, n_35230, n_35231, n_35232, n_35233, n_35234, n_35235, n_35236, n_35237, n_35238, n_35239, n_35240, n_35241, n_35242, n_35243, n_35244, n_35245, n_35246, n_35247, n_35248, n_35249, n_35250, n_35251, n_35252, n_35253, n_35254, n_35255, n_35256, n_35257, n_35258, n_35259, n_35260, n_35261, n_35262, n_35263, n_35264, n_35265, n_35266, n_35267, n_35268, n_35269, n_35270, n_35271, n_35272, n_35273, n_35274, n_35275, n_35276, n_35277, n_35278, n_35279, n_35280, n_35281, n_35282, n_35283, n_35284, n_35285, n_35286, n_35287, n_35288, n_35289, n_35290, n_35291, n_35292, n_35293, n_35294, n_35295, n_35296, n_35297, n_35298, n_35299, n_35300, n_35301, n_35302, n_35303, n_35304, n_35305, n_35306, n_35307, n_35308, n_35309, n_35310, n_35311, n_35312, n_35313, n_35314, n_35315, n_35316, n_35317, n_35318, n_35319, n_35320, n_35321, n_35322, n_35323, n_35324, n_35325, n_35326, n_35327, n_35328, n_35329, n_35330, n_35331, n_35332, n_35333, n_35334, n_35335, n_35336, n_35337, n_35338, n_35339, n_35340, n_35341, n_35342, n_35343, n_35344, n_35345, n_35346, n_35347, n_35348, n_35349, n_35350, n_35351, n_35352, n_35353, n_35354, n_35355, n_35356, n_35357, n_35358, n_35359, n_35360, n_35361, n_35362, n_35363, n_35364, n_35365, n_35366, n_35367, n_35368, n_35369, n_35370, n_35371, n_35372, n_35373, n_35374, n_35375, n_35376, n_35377, n_35378, n_35379, n_35380, n_35381, n_35382, n_35383, n_35384, n_35385, n_35386, n_35387, n_35388, n_35389, n_35390, n_35391, n_35392, n_35393, n_35394, n_35395, n_35396, n_35397, n_35398, n_35399, n_35400, n_35401, n_35402, n_35403, n_35404, n_35405, n_35406, n_35407, n_35408, n_35409, n_35410, n_35411, n_35412, n_35413, n_35414, n_35415, n_35416, n_35417, n_35418, n_35419, n_35420, n_35421, n_35422, n_35423, n_35424, n_35425, n_35426, n_35427, n_35428, n_35429, n_35430, n_35431, n_35432, n_35433, n_35434, n_35435, n_35436, n_35437, n_35438, n_35439, n_35440, n_35441, n_35442, n_35443, n_35444, n_35445, n_35446, n_35447, n_35448, n_35449, n_35450, n_35451, n_35452, n_35453, n_35454, n_35455, n_35456, n_35457, n_35458, n_35459, n_35460, n_35461, n_35462, n_35463, n_35464, n_35465, n_35466, n_35467, n_35468, n_35469, n_35470, n_35471, n_35472, n_35473, n_35474, n_35475, n_35476, n_35477, n_35478, n_35479, n_35480, n_35481, n_35482, n_35483, n_35484, n_35485, n_35486, n_35487, n_35488, n_35489, n_35490, n_35491, n_35492, n_35493, n_35494, n_35495, n_35496, n_35497, n_35498, n_35499, n_35500, n_35501, n_35502, n_35503, n_35504, n_35505, n_35506, n_35507, n_35508, n_35509, n_35510, n_35511, n_35512, n_35513, n_35514, n_35515, n_35516, n_35517, n_35518, n_35519, n_35520, n_35521, n_35522, n_35523, n_35524, n_35525, n_35526, n_35527, n_35528, n_35529, n_35530, n_35531, n_35532, n_35533, n_35534, n_35535, n_35536, n_35537, n_35538, n_35539, n_35540, n_35541, n_35542, n_35543, n_35544, n_35545, n_35546, n_35547, n_35548, n_35549, n_35550, n_35551, n_35552, n_35553, n_35554, n_35555, n_35556, n_35557, n_35558, n_35559, n_35560, n_35561, n_35562, n_35563, n_35564, n_35565, n_35566, n_35567, n_35568, n_35569, n_35570, n_35571, n_35572, n_35573, n_35574, n_35575, n_35576, n_35577, n_35578, n_35579, n_35580, n_35581, n_35582, n_35583, n_35584, n_35585, n_35586, n_35587, n_35588, n_35589, n_35590, n_35591, n_35592, n_35593, n_35594, n_35595, n_35596, n_35597, n_35598, n_35599, n_35600, n_35601, n_35602, n_35603, n_35604, n_35605, n_35606, n_35607, n_35608, n_35609, n_35610, n_35611, n_35612, n_35613, n_35614, n_35615, n_35616, n_35617, n_35618, n_35619, n_35620, n_35621, n_35622, n_35623, n_35624, n_35625, n_35626, n_35627, n_35628, n_35629, n_35630, n_35631, n_35632, n_35633, n_35634, n_35635, n_35636, n_35637, n_35638, n_35639, n_35640, n_35641, n_35642, n_35643, n_35644, n_35645, n_35646, n_35647, n_35648, n_35649, n_35650, n_35651, n_35652, n_35653, n_35654, n_35655, n_35656, n_35657, n_35658, n_35659, n_35660, n_35661, n_35662, n_35663, n_35664, n_35665, n_35666, n_35667, n_35668, n_35669, n_35670, n_35671, n_35672, n_35673, n_35674, n_35675, n_35676, n_35677, n_35678, n_35679, n_35680, n_35681, n_35682, n_35683, n_35684, n_35685, n_35686, n_35687, n_35688, n_35689, n_35690, n_35691, n_35692, n_35693, n_35694, n_35695, n_35696, n_35697, n_35698, n_35699, n_35700, n_35701, n_35702, n_35703, n_35704, n_35705, n_35706, n_35707, n_35708, n_35709, n_35710, n_35711, n_35712, n_35713, n_35714, n_35715, n_35716, n_35717, n_35718, n_35719, n_35720, n_35721, n_35722, n_35723, n_35724, n_35725, n_35726, n_35727, n_35728, n_35729, n_35730, n_35731, n_35732, n_35733, n_35734, n_35735, n_35736, n_35737, n_35738, n_35739, n_35740, n_35741, n_35742, n_35743, n_35744, n_35745, n_35746, n_35747, n_35748, n_35749, n_35750, n_35751, n_35752, n_35753, n_35754, n_35755, n_35756, n_35757, n_35758, n_35759, n_35760, n_35761, n_35762, n_35763, n_35764, n_35765, n_35766, n_35767, n_35768, n_35769, n_35770, n_35771, n_35772, n_35773, n_35774, n_35775, n_35776, n_35777, n_35778, n_35779, n_35780, n_35781, n_35782, n_35783, n_35784, n_35785, n_35786, n_35787, n_35788, n_35789, n_35790, n_35791, n_35792, n_35793, n_35794, n_35795, n_35796, n_35797, n_35798, n_35799, n_35800, n_35801, n_35802, n_35803, n_35804, n_35805, n_35806, n_35807, n_35808, n_35809, n_35810, n_35811, n_35812, n_35813, n_35814, n_35815, n_35816, n_35817, n_35818, n_35819, n_35820, n_35821, n_35822, n_35823, n_35824, n_35825, n_35826, n_35827, n_35828, n_35829, n_35830, n_35831, n_35832, n_35833, n_35834, n_35835, n_35836, n_35837, n_35838, n_35839, n_35840, n_35841, n_35842, n_35843, n_35844, n_35845, n_35846, n_35847, n_35848, n_35849, n_35850, n_35851, n_35852, n_35853, n_35854, n_35855, n_35856, n_35857, n_35858, n_35859, n_35860, n_35861, n_35862, n_35863, n_35864, n_35865, n_35866, n_35867, n_35868, n_35869, n_35870, n_35871, n_35872, n_35873, n_35874, n_35875, n_35876, n_35877, n_35878, n_35879, n_35880, n_35881, n_35882, n_35883, n_35884, n_35885, n_35886, n_35887, n_35888, n_35889, n_35890, n_35891, n_35892, n_35893, n_35894, n_35895, n_35896, n_35897, n_35898, n_35899, n_35900, n_35901, n_35902, n_35903, n_35904, n_35905, n_35906, n_35907, n_35908, n_35909, n_35910, n_35911, n_35912, n_35913, n_35914, n_35915, n_35916, n_35917, n_35918, n_35919, n_35920, n_35921, n_35922, n_35923, n_35924, n_35925, n_35926, n_35927, n_35928, n_35929, n_35930, n_35931, n_35932, n_35933, n_35934, n_35935, n_35936, n_35937, n_35938, n_35939, n_35940, n_35941, n_35942, n_35943, n_35944, n_35945, n_35946, n_35947, n_35948, n_35949, n_35950, n_35951, n_35952, n_35953, n_35954, n_35955, n_35956, n_35957, n_35958, n_35959, n_35960, n_35961, n_35962, n_35963, n_35964, n_35965, n_35966, n_35967, n_35968, n_35969, n_35970, n_35971, n_35972, n_35973, n_35974, n_35975, n_35976, n_35977, n_35978, n_35979, n_35980, n_35981, n_35982, n_35983, n_35984, n_35985, n_35986, n_35987, n_35988, n_35989, n_35990, n_35991, n_35992, n_35993, n_35994, n_35995, n_35996, n_35997, n_35998, n_35999, n_36000, n_36001, n_36002, n_36003, n_36004, n_36005, n_36006, n_36007, n_36008, n_36009, n_36010, n_36011, n_36012, n_36013, n_36014, n_36015, n_36016, n_36017, n_36018, n_36019, n_36020, n_36021, n_36022, n_36023, n_36024, n_36025, n_36026, n_36027, n_36028, n_36029, n_36030, n_36031, n_36032, n_36033, n_36034, n_36035, n_36036, n_36037, n_36038, n_36039, n_36040, n_36041, n_36042, n_36043, n_36044, n_36045, n_36046, n_36047, n_36048, n_36049, n_36050, n_36051, n_36052, n_36053, n_36054, n_36055, n_36056, n_36057, n_36058, n_36059, n_36060, n_36061, n_36062, n_36063, n_36064, n_36065, n_36066, n_36067, n_36068, n_36069, n_36070, n_36071, n_36072, n_36073, n_36074, n_36075, n_36076, n_36077, n_36078, n_36079, n_36080, n_36081, n_36082, n_36083, n_36084, n_36085, n_36086, n_36087, n_36088, n_36089, n_36090, n_36091, n_36092, n_36093, n_36094, n_36095, n_36096, n_36097, n_36098, n_36099, n_36100, n_36101, n_36102, n_36103, n_36104, n_36105, n_36106, n_36107, n_36108, n_36109, n_36110, n_36111, n_36112, n_36113, n_36114, n_36115, n_36116, n_36117, n_36118, n_36119, n_36120, n_36121, n_36122, n_36123, n_36124, n_36125, n_36126, n_36127, n_36128, n_36129, n_36130, n_36131, n_36132, n_36133, n_36134, n_36135, n_36136, n_36137, n_36138, n_36139, n_36140, n_36141, n_36142, n_36143, n_36144, n_36145, n_36146, n_36147, n_36148, n_36149, n_36150, n_36151, n_36152, n_36153, n_36154, n_36155, n_36156, n_36157, n_36158, n_36159, n_36160, n_36161, n_36162, n_36163, n_36164, n_36165, n_36166, n_36167, n_36168, n_36169, n_36170, n_36171, n_36172, n_36173, n_36174, n_36175, n_36176, n_36177, n_36178, n_36179, n_36180, n_36181, n_36182, n_36183, n_36184, n_36185, n_36186, n_36187, n_36188, n_36189, n_36190, n_36191, n_36192, n_36193, n_36194, n_36195, n_36196, n_36197, n_36198, n_36199, n_36200, n_36201, n_36202, n_36203, n_36204, n_36205, n_36206, n_36207, n_36208, n_36209, n_36210, n_36211, n_36212, n_36213, n_36214, n_36215, n_36216, n_36217, n_36218, n_36219, n_36220, n_36221, n_36222, n_36223, n_36224, n_36225, n_36226, n_36227, n_36228, n_36229, n_36230, n_36231, n_36232, n_36233, n_36234, n_36235, n_36236, n_36237, n_36238, n_36239, n_36240, n_36241, n_36242, n_36243, n_36244, n_36245, n_36246, n_36247, n_36248, n_36249, n_36250, n_36251, n_36252, n_36253, n_36254, n_36255, n_36256, n_36257, n_36258, n_36259, n_36260, n_36261, n_36262, n_36263, n_36264, n_36265, n_36266, n_36267, n_36268, n_36269, n_36270, n_36271, n_36272, n_36273, n_36274, n_36275, n_36276, n_36277, n_36278, n_36279, n_36280, n_36281, n_36282, n_36283, n_36284, n_36285, n_36286, n_36287, n_36288, n_36289, n_36290, n_36291, n_36292, n_36293, n_36294, n_36295, n_36296, n_36297, n_36298, n_36299, n_36300, n_36301, n_36302, n_36303, n_36304, n_36305, n_36306, n_36307, n_36308, n_36309, n_36310, n_36311, n_36312, n_36313, n_36314, n_36315, n_36316, n_36317, n_36318, n_36319, n_36320, n_36321, n_36322, n_36323, n_36324, n_36325, n_36326, n_36327, n_36328, n_36329, n_36330, n_36331, n_36332, n_36333, n_36334, n_36335, n_36336, n_36337, n_36338, n_36339, n_36340, n_36341, n_36342, n_36343, n_36344, n_36345, n_36346, n_36347, n_36348, n_36349, n_36350, n_36351, n_36352, n_36353, n_36354, n_36355, n_36356, n_36357, n_36358, n_36359, n_36360, n_36361, n_36362, n_36363, n_36364, n_36365, n_36366, n_36367, n_36368, n_36369, n_36370, n_36371, n_36372, n_36373, n_36374, n_36375, n_36376, n_36377, n_36378, n_36379, n_36380, n_36381, n_36382, n_36383, n_36384, n_36385, n_36386, n_36387, n_36388, n_36389, n_36390, n_36391, n_36392, n_36393, n_36394, n_36395, n_36396, n_36397, n_36398, n_36399, n_36400, n_36401, n_36402, n_36403, n_36404, n_36405, n_36406, n_36407, n_36408, n_36409, n_36410, n_36411, n_36412, n_36413, n_36414, n_36415, n_36416, n_36417, n_36418, n_36419, n_36420, n_36421, n_36422, n_36423, n_36424, n_36425, n_36426, n_36427, n_36428, n_36429, n_36430, n_36431, n_36432, n_36433, n_36434, n_36435, n_36436, n_36437, n_36438, n_36439, n_36440, n_36441, n_36442, n_36443, n_36444, n_36445, n_36446, n_36447, n_36448, n_36449, n_36450, n_36451, n_36452, n_36453, n_36454, n_36455, n_36456, n_36457, n_36458, n_36459, n_36460, n_36461, n_36462, n_36463, n_36464, n_36465, n_36466, n_36467, n_36468, n_36469, n_36470, n_36471, n_36472, n_36473, n_36474, n_36475, n_36476, n_36477, n_36478, n_36479, n_36480, n_36481, n_36482, n_36483, n_36484, n_36485, n_36486, n_36487, n_36488, n_36489, n_36490, n_36491, n_36492, n_36493, n_36494, n_36495, n_36496, n_36497, n_36498, n_36499, n_36500, n_36501, n_36502, n_36503, n_36504, n_36505, n_36506, n_36507, n_36508, n_36509, n_36510, n_36511, n_36512, n_36513, n_36514, n_36515, n_36516, n_36517, n_36518, n_36519, n_36520, n_36521, n_36522, n_36523, n_36524, n_36525, n_36526, n_36527, n_36528, n_36529, n_36530, n_36531, n_36532, n_36533, n_36534, n_36535, n_36536, n_36537, n_36538, n_36539, n_36540, n_36541, n_36542, n_36543, n_36544, n_36545, n_36546, n_36547, n_36548, n_36549, n_36550, n_36551, n_36552, n_36553, n_36554, n_36555, n_36556, n_36557, n_36558, n_36559, n_36560, n_36561, n_36562, n_36563, n_36564, n_36565, n_36566, n_36567, n_36568, n_36569, n_36570, n_36571, n_36572, n_36573, n_36574, n_36575, n_36576, n_36577, n_36578, n_36579, n_36580, n_36581, n_36582, n_36583, n_36584, n_36585, n_36586, n_36587, n_36588, n_36589, n_36590, n_36591, n_36592, n_36593, n_36594, n_36595, n_36596, n_36597, n_36598, n_36599, n_36600, n_36601, n_36602, n_36603, n_36604, n_36605, n_36606, n_36607, n_36608, n_36609, n_36610, n_36611, n_36612, n_36613, n_36614, n_36615, n_36616, n_36617, n_36618, n_36619, n_36620, n_36621, n_36622, n_36623, n_36624, n_36625, n_36626, n_36627, n_36628, n_36629, n_36630, n_36631, n_36632, n_36633, n_36634, n_36635, n_36636, n_36637, n_36638, n_36639, n_36640, n_36641, n_36642, n_36643, n_36644, n_36645, n_36646, n_36647, n_36648, n_36649, n_36650, n_36651, n_36652, n_36653, n_36654, n_36655, n_36656, n_36657, n_36658, n_36659, n_36660, n_36661, n_36662, n_36663, n_36664, n_36665, n_36666, n_36667, n_36668, n_36669, n_36670, n_36671, n_36672, n_36673, n_36674, n_36675, n_36676, n_36677, n_36678, n_36679, n_36680, n_36681, n_36682, n_36683, n_36684, n_36685, n_36686, n_36687, n_36688, n_36689, n_36690, n_36691, n_36692, n_36693, n_36694, n_36695, n_36696, n_36697, n_36698, n_36699, n_36700, n_36701, n_36702, n_36703, n_36704, n_36705, n_36706, n_36707, n_36708, n_36709, n_36710, n_36711, n_36712, n_36713, n_36714, n_36715, n_36716, n_36717, n_36718, n_36719, n_36720, n_36721, n_36722, n_36723, n_36724, n_36725, n_36726, n_36727, n_36728, n_36729, n_36730, n_36731, n_36732, n_36733, n_36734, n_36735, n_36736, n_36737, n_36738, n_36739, n_36740, n_36741, n_36742, n_36743, n_36744, n_36745, n_36746, n_36747, n_36748, n_36749, n_36750, n_36751, n_36752, n_36753, n_36754, n_36755, n_36756, n_36757, n_36758, n_36759, n_36760, n_36761, n_36762, n_36763, n_36764, n_36765, n_36766, n_36767, n_36768, n_36769, n_36770, n_36771, n_36772, n_36773, n_36774, n_36775, n_36776, n_36777, n_36778, n_36779, n_36780, n_36781, n_36782, n_36783, n_36784, n_36785, n_36786, n_36787, n_36788, n_36789, n_36790, n_36791, n_36792, n_36793, n_36794, n_36795, n_36796, n_36797, n_36798, n_36799, n_36800, n_36801, n_36802, n_36803, n_36804, y7, n_36805, n_36806, n_36807, n_36808, n_36809, n_36810, n_36811, n_36812, n_36813, n_36814, n_36815, n_36816, n_36817, n_36818, n_36819, n_36820, n_36821, n_36822, n_36823, n_36824, n_36825, n_36826, n_36827, n_36828, n_36829, n_36830, n_36831, n_36832, n_36833, n_36834, n_36835, n_36836, n_36837, n_36838, n_36839, n_36840, n_36841, n_36842, n_36843, n_36844, n_36845, n_36846, n_36847, n_36848, n_36849, n_36850, n_36851, n_36852, n_36853, n_36854, y6, n_36855, n_36856, n_36857, n_36858, n_36859, n_36860, n_36861, n_36862, n_36863, n_36864, n_36865, n_36866, n_36867, n_36868, n_36869, n_36870, n_36871, n_36872, n_36873, n_36874, n_36875, n_36876, n_36877, n_36878, n_36879, n_36880, y5, n_36881, n_36882, n_36883, n_36884, n_36885, n_36886, n_36887, n_36888, n_36889, n_36890, n_36891, n_36892, n_36893, n_36894, n_36895, n_36896, n_36897, n_36898, n_36899, n_36900, n_36901, n_36902, n_36903, n_36904, n_36905, n_36906, n_36907, n_36908, n_36909, n_36910, n_36911, n_36912, y4, n_36913, n_36914, n_36915, n_36916, n_36917, n_36918, n_36919, n_36920, n_36921, n_36922, n_36923, n_36924, n_36925, n_36926, n_36927, n_36928, n_36929, n_36930, n_36931, n_36932, n_36933, n_36934, n_36935, y3, n_36936, n_36937, n_36938, n_36939, n_36940, n_36941, n_36942, n_36943, n_36944, n_36945, n_36946, n_36947, n_36948, n_36949, n_36950, n_36951, n_36952, n_36953, n_36954, n_36955, n_36956, y2, n_36957, n_36958, n_36959, n_36960, n_36961, n_36962, n_36963, n_36964, n_36965, n_36966, n_36967, n_36968, n_36969, n_36970, n_36971, n_36972, n_36973, n_36974, n_36975, n_36976, n_36977, y1, n_36978, n_36979, n_36980, n_36981, n_36982, n_36983, n_36984, n_36985, n_36986, n_36987, n_36988, n_36989, n_36990, y0, n_36991, n_36992, n_36993, n_36994, n_36995, n_36996, n_36997, n_36998, n_36999, n_37000, n_37001, n_37002, n_37003, n_37004, n_37005, n_37006, n_37007, n_37008, n_37009, n_37010, n_37011, n_37012, n_37013, n_37014, n_37015, n_37016, n_37017, y15, n_37018, n_37019, n_37020, n_37021, n_37022, n_37023, n_37024, n_37025, n_37026, n_37027, n_37028, n_37029, n_37030, n_37031, n_37032, n_37033, n_37034, n_37035, n_37036, n_37037, n_37038, n_37039, y14, n_37040, n_37041, n_37042, n_37043, n_37044, n_37045, n_37046, n_37047, n_37048, n_37049, n_37050, n_37051, n_37052, n_37053, n_37054, n_37055, n_37056, n_37057, n_37058, n_37059, n_37060, n_37061, y13, n_37062, n_37063, n_37064, n_37065, n_37066, n_37067, n_37068, n_37069, n_37070, n_37071, n_37072, n_37073, n_37074, n_37075, n_37076, n_37077, n_37078, n_37079, n_37080, n_37081, n_37082, n_37083, n_37084, y12, n_37085, n_37086, n_37087, n_37088, n_37089, n_37090, n_37091, n_37092, n_37093, n_37094, n_37095, n_37096, n_37097, n_37098, n_37099, n_37100, n_37101, n_37102, n_37103, n_37104, n_37105, n_37106, y11, n_37107, n_37108, n_37109, n_37110, n_37111, n_37112, n_37113, n_37114, n_37115, n_37116, n_37117, n_37118, n_37119, n_37120, n_37121, n_37122, n_37123, n_37124, n_37125, n_37126, n_37127, n_37128, y10, n_37129, n_37130, n_37131, n_37132, n_37133, n_37134, n_37135, n_37136, n_37137, n_37138, n_37139, n_37140, n_37141, n_37142, n_37143, n_37144, n_37145, n_37146, n_37147, n_37148, n_37149, n_37150, y9, n_37151, n_37152, n_37153, n_37154, n_37155, n_37156, n_37157, n_37158, n_37159, n_37160, n_37161, n_37162, n_37163, n_37164, n_37165, n_37166, n_37167, n_37168, n_37169, n_37170, n_37171, y8, n_37172, n_37173, n_37174, n_37175, n_37176, n_37177, n_37178, n_37179, n_37180, n_37181, n_37182, n_37183, n_37184, n_37185, n_37186, n_37187, n_37188, y23, n_37189, n_37190, n_37191, n_37192, n_37193, n_37194, n_37195, n_37196, n_37197, n_37198, n_37199, n_37200, n_37201, n_37202, n_37203, n_37204, n_37205, n_37206, n_37207, n_37208, n_37209, n_37210, n_37211, n_37212, n_37213, n_37214, n_37215, n_37216, n_37217, y22, n_37218, n_37219, n_37220, n_37221, n_37222, n_37223, n_37224, n_37225, n_37226, n_37227, n_37228, n_37229, n_37230, n_37231, n_37232, n_37233, n_37234, n_37235, n_37236, n_37237, n_37238, n_37239, y21, n_37240, n_37241, n_37242, n_37243, n_37244, n_37245, n_37246, n_37247, n_37248, n_37249, n_37250, n_37251, n_37252, n_37253, n_37254, n_37255, n_37256, n_37257, n_37258, n_37259, n_37260, n_37261, y20, n_37262, n_37263, n_37264, n_37265, n_37266, n_37267, n_37268, n_37269, n_37270, n_37271, n_37272, n_37273, n_37274, n_37275, n_37276, n_37277, n_37278, n_37279, n_37280, n_37281, n_37282, n_37283, y19, n_37284, n_37285, n_37286, n_37287, n_37288, n_37289, n_37290, n_37291, n_37292, n_37293, n_37294, n_37295, n_37296, n_37297, n_37298, n_37299, n_37300, n_37301, n_37302, n_37303, n_37304, n_37305, n_37306, y18, n_37307, n_37308, n_37309, n_37310, n_37311, n_37312, n_37313, n_37314, n_37315, n_37316, n_37317, n_37318, n_37319, n_37320, n_37321, y17, n_37322, n_37323, n_37324, n_37325, n_37326, n_37327, n_37328, n_37329, n_37330, n_37331, n_37332, n_37333, n_37334, n_37335, n_37336, n_37337, n_37338, n_37339, n_37340, n_37341, n_37342, y16, n_37343, n_37344, n_37345, n_37346, n_37347, n_37348, n_37349, n_37350, n_37351, n_37352, n_37353, n_37354, n_37355, n_37356, n_37357, n_37358, n_37359, n_37360, n_37361, n_37362, n_37363, n_37364, n_37365, y31, n_37366, n_37367, n_37368, n_37369, n_37370, n_37371, n_37372, n_37373, n_37374, n_37375, n_37376, n_37377, n_37378, n_37379, n_37380, n_37381, n_37382, n_37383, n_37384, n_37385, n_37386, n_37387, n_37388, n_37389, n_37390, n_37391, n_37392, n_37393, n_37394, n_37395, n_37396, y103, n_37397, y30, n_37398, n_37399, n_37400, n_37401, n_37402, n_37403, n_37404, n_37405, n_37406, n_37407, n_37408, n_37409, n_37410, n_37411, n_37412, n_37413, y102, n_37414, n_37415, n_37416, n_37417, n_37418, n_37419, n_37420, n_37421, n_37422, n_37423, n_37424, n_37425, n_37426, n_37427, n_37428, n_37429, n_37430, y29, n_37431, n_37432, n_37433, n_37434, n_37435, n_37436, n_37437, n_37438, n_37439, n_37440, n_37441, n_37442, n_37443, n_37444, n_37445, n_37446, n_37447, n_37448, n_37449, n_37450, n_37451, n_37452, n_37453, n_37454, n_37455, n_37456, n_37457, n_37458, n_37459, n_37460, n_37461, n_37462, n_37463, n_37464, n_37465, n_37466, y28, n_37467, n_37468, n_37469, n_37470, n_37471, n_37472, y101, n_37473, n_37474, n_37475, n_37476, n_37477, n_37478, n_37479, n_37480, n_37481, n_37482, n_37483, n_37484, n_37485, n_37486, n_37487, n_37488, n_37489, n_37490, n_37491, n_37492, n_37493, n_37494, n_37495, n_37496, n_37497, n_37498, n_37499, n_37500, n_37501, n_37502, n_37503, n_37504, n_37505, n_37506, n_37507, n_37508, n_37509, y27, n_37510, n_37511, n_37512, n_37513, y100, n_37514, n_37515, n_37516, n_37517, n_37518, n_37519, n_37520, n_37521, n_37522, n_37523, n_37524, n_37525, n_37526, n_37527, n_37528, n_37529, n_37530, n_37531, n_37532, n_37533, n_37534, n_37535, n_37536, n_37537, y26, n_37538, n_37539, n_37540, n_37541, n_37542, n_37543, n_37544, n_37545, n_37546, n_37547, n_37548, n_37549, n_37550, n_37551, n_37552, n_37553, n_37554, n_37555, n_37556, n_37557, n_37558, n_37559, n_37560, y99, n_37561, n_37562, n_37563, n_37564, n_37565, n_37566, n_37567, n_37568, n_37569, n_37570, n_37571, n_37572, n_37573, n_37574, n_37575, n_37576, n_37577, n_37578, y25, n_37579, n_37580, n_37581, n_37582, n_37583, n_37584, n_37585, n_37586, n_37587, n_37588, n_37589, n_37590, n_37591, n_37592, n_37593, n_37594, n_37595, n_37596, n_37597, n_37598, n_37599, n_37600, n_37601, n_37602, n_37603, n_37604, y98, n_37605, n_37606, n_37607, n_37608, n_37609, n_37610, n_37611, n_37612, n_37613, n_37614, n_37615, n_37616, n_37617, n_37618, n_37619, n_37620, n_37621, n_37622, n_37623, n_37624, n_37625, n_37626, n_37627, n_37628, n_37629, n_37630, n_37631, n_37632, n_37633, y24, n_37634, n_37635, n_37636, n_37637, n_37638, n_37639, n_37640, y97, n_37641, n_37642, n_37643, n_37644, n_37645, n_37646, n_37647, n_37648, n_37649, n_37650, n_37651, n_37652, n_37653, n_37654, n_37655, n_37656, n_37657, n_37658, n_37659, n_37660, n_37661, n_37662, n_37663, n_37664, n_37665, n_37666, n_37667, n_37668, y96, n_37669, n_37670, n_37671, n_37672, n_37673, n_37674, n_37675, n_37676, n_37677, n_37678, n_37679, n_37680, n_37681, n_37682, n_37683, n_37684, n_37685, n_37686, n_37687, n_37688, n_37689, n_37690, n_37691, n_37692, n_37693, n_37694, n_37695, n_37696, n_37697, y111, n_37698, n_37699, n_37700, n_37701, n_37702, n_37703, n_37704, n_37705, n_37706, n_37707, n_37708, n_37709, n_37710, n_37711, n_37712, n_37713, n_37714, n_37715, n_37716, n_37717, n_37718, n_37719, y110, n_37720, n_37721, n_37722, n_37723, n_37724, n_37725, n_37726, n_37727, n_37728, n_37729, n_37730, n_37731, n_37732, n_37733, n_37734, n_37735, n_37736, n_37737, n_37738, n_37739, y109, n_37740, n_37741, n_37742, n_37743, n_37744, n_37745, n_37746, n_37747, n_37748, n_37749, n_37750, n_37751, n_37752, n_37753, n_37754, n_37755, n_37756, n_37757, n_37758, n_37759, n_37760, n_37761, n_37762, y108, n_37763, n_37764, n_37765, n_37766, n_37767, n_37768, n_37769, n_37770, n_37771, n_37772, n_37773, n_37774, n_37775, n_37776, y107, n_37777, n_37778, n_37779, n_37780, n_37781, n_37782, n_37783, n_37784, n_37785, n_37786, n_37787, n_37788, n_37789, n_37790, n_37791, n_37792, n_37793, n_37794, n_37795, n_37796, n_37797, n_37798, n_37799, n_37800, n_37801, n_37802, n_37803, n_37804, y106, n_37805, n_37806, n_37807, n_37808, n_37809, n_37810, n_37811, n_37812, n_37813, n_37814, n_37815, n_37816, n_37817, n_37818, n_37819, n_37820, n_37821, n_37822, n_37823, n_37824, n_37825, n_37826, y105, n_37827, n_37828, n_37829, n_37830, n_37831, n_37832, n_37833, n_37834, n_37835, n_37836, n_37837, n_37838, n_37839, n_37840, y104, n_37841, n_37842, n_37843, n_37844, n_37845, n_37846, n_37847, n_37848, n_37849, n_37850, n_37851, n_37852, n_37853, n_37854, n_37855, n_37856, n_37857, n_37858, n_37859, n_37860, n_37861, n_37862, n_37863, n_37864, n_37865, n_37866, n_37867, n_37868, n_37869, n_37870, y119, n_37871, n_37872, n_37873, n_37874, n_37875, n_37876, n_37877, n_37878, n_37879, n_37880, n_37881, n_37882, n_37883, n_37884, y118, n_37885, n_37886, n_37887, n_37888, n_37889, n_37890, n_37891, n_37892, n_37893, n_37894, n_37895, n_37896, n_37897, n_37898, n_37899, n_37900, n_37901, n_37902, n_37903, n_37904, n_37905, n_37906, n_37907, n_37908, n_37909, n_37910, n_37911, n_37912, y117, n_37913, n_37914, n_37915, n_37916, n_37917, n_37918, n_37919, n_37920, n_37921, n_37922, n_37923, n_37924, n_37925, n_37926, n_37927, n_37928, n_37929, n_37930, n_37931, n_37932, n_37933, n_37934, n_37935, n_37936, y116, n_37937, n_37938, n_37939, n_37940, n_37941, y71, n_37942, n_37943, n_37944, n_37945, n_37946, n_37947, n_37948, n_37949, n_37950, n_37951, n_37952, n_37953, n_37954, n_37955, n_37956, n_37957, n_37958, n_37959, n_37960, n_37961, n_37962, n_37963, n_37964, n_37965, y115, n_37966, n_37967, n_37968, n_37969, n_37970, n_37971, n_37972, n_37973, n_37974, n_37975, n_37976, n_37977, n_37978, y70, n_37979, n_37980, n_37981, n_37982, n_37983, n_37984, n_37985, n_37986, n_37987, n_37988, n_37989, n_37990, n_37991, n_37992, n_37993, n_37994, n_37995, y114, n_37996, n_37997, n_37998, n_37999, n_38000, n_38001, n_38002, n_38003, n_38004, n_38005, n_38006, n_38007, n_38008, n_38009, n_38010, n_38011, n_38012, n_38013, n_38014, n_38015, n_38016, n_38017, n_38018, n_38019, y113, n_38020, n_38021, n_38022, n_38023, n_38024, n_38025, n_38026, n_38027, n_38028, n_38029, n_38030, n_38031, n_38032, n_38033, n_38034, n_38035, n_38036, n_38037, n_38038, n_38039, n_38040, n_38041, y69, n_38042, n_38043, n_38044, n_38045, n_38046, n_38047, n_38048, n_38049, n_38050, n_38051, n_38052, n_38053, n_38054, n_38055, n_38056, n_38057, n_38058, y112, n_38059, n_38060, n_38061, n_38062, n_38063, n_38064, n_38065, n_38066, n_38067, n_38068, n_38069, n_38070, n_38071, n_38072, n_38073, n_38074, n_38075, n_38076, n_38077, n_38078, n_38079, n_38080, n_38081, y68, n_38082, n_38083, n_38084, n_38085, n_38086, n_38087, n_38088, n_38089, n_38090, n_38091, n_38092, n_38093, n_38094, n_38095, n_38096, n_38097, n_38098, n_38099, y127, n_38100, n_38101, n_38102, n_38103, n_38104, n_38105, n_38106, n_38107, n_38108, n_38109, n_38110, n_38111, n_38112, n_38113, n_38114, n_38115, n_38116, n_38117, n_38118, n_38119, y67, n_38120, n_38121, n_38122, n_38123, n_38124, n_38125, n_38126, n_38127, n_38128, n_38129, n_38130, n_38131, n_38132, n_38133, n_38134, n_38135, n_38136, n_38137, n_38138, n_38139, n_38140, n_38141, n_38142, n_38143, y126, n_38144, n_38145, n_38146, n_38147, n_38148, n_38149, n_38150, n_38151, n_38152, n_38153, n_38154, n_38155, n_38156, n_38157, n_38158, n_38159, n_38160, n_38161, n_38162, n_38163, n_38164, n_38165, n_38166, y66, n_38167, n_38168, n_38169, n_38170, n_38171, n_38172, n_38173, n_38174, n_38175, n_38176, n_38177, n_38178, n_38179, n_38180, n_38181, n_38182, n_38183, n_38184, n_38185, n_38186, n_38187, n_38188, n_38189, n_38190, n_38191, n_38192, n_38193, n_38194, n_38195, n_38196, n_38197, n_38198, n_38199, n_38200, n_38201, n_38202, n_38203, n_38204, y125, n_38205, n_38206, n_38207, n_38208, n_38209, n_38210, y65, n_38211, n_38212, n_38213, n_38214, n_38215, n_38216, n_38217, n_38218, n_38219, n_38220, n_38221, n_38222, n_38223, n_38224, n_38225, n_38226, n_38227, n_38228, n_38229, n_38230, n_38231, n_38232, n_38233, n_38234, n_38235, n_38236, n_38237, n_38238, n_38239, n_38240, n_38241, n_38242, n_38243, n_38244, n_38245, n_38246, n_38247, n_38248, n_38249, n_38250, y124, n_38251, n_38252, n_38253, n_38254, n_38255, y64, n_38256, n_38257, n_38258, n_38259, n_38260, n_38261, n_38262, n_38263, n_38264, n_38265, n_38266, n_38267, n_38268, n_38269, n_38270, n_38271, n_38272, n_38273, n_38274, n_38275, n_38276, n_38277, n_38278, y123, n_38279, n_38280, n_38281, n_38282, n_38283, n_38284, n_38285, n_38286, n_38287, n_38288, n_38289, n_38290, n_38291, n_38292, n_38293, n_38294, n_38295, n_38296, n_38297, n_38298, n_38299, n_38300, n_38301, n_38302, y79, n_38303, n_38304, n_38305, n_38306, n_38307, n_38308, n_38309, n_38310, n_38311, n_38312, n_38313, n_38314, n_38315, n_38316, n_38317, n_38318, n_38319, n_38320, n_38321, n_38322, n_38323, n_38324, n_38325, n_38326, n_38327, n_38328, n_38329, n_38330, n_38331, n_38332, n_38333, n_38334, n_38335, n_38336, n_38337, n_38338, y122, n_38339, n_38340, n_38341, y78, n_38342, n_38343, n_38344, n_38345, n_38346, n_38347, n_38348, n_38349, n_38350, n_38351, n_38352, n_38353, n_38354, n_38355, n_38356, n_38357, n_38358, n_38359, n_38360, n_38361, n_38362, n_38363, n_38364, n_38365, n_38366, n_38367, n_38368, n_38369, n_38370, n_38371, n_38372, n_38373, n_38374, n_38375, n_38376, n_38377, n_38378, n_38379, n_38380, y121, n_38381, n_38382, n_38383, n_38384, n_38385, n_38386, n_38387, n_38388, n_38389, n_38390, y77, n_38391, n_38392, n_38393, n_38394, n_38395, n_38396, n_38397, y120, n_38398, n_38399, n_38400, n_38401, n_38402, n_38403, n_38404, n_38405, n_38406, n_38407, n_38408, n_38409, n_38410, n_38411, n_38412, n_38413, n_38414, n_38415, n_38416, n_38417, n_38418, n_38419, n_38420, n_38421, n_38422, n_38423, n_38424, n_38425, n_38426, n_38427, y76, n_38428, n_38429, n_38430, n_38431, n_38432, n_38433, n_38434, n_38435, n_38436, n_38437, n_38438, n_38439, n_38440, n_38441, n_38442, n_38443, n_38444, n_38445, n_38446, n_38447, n_38448, n_38449, n_38450, n_38451, n_38452, n_38453, n_38454, n_38455, n_38456, n_38457, y75, n_38458, n_38459, n_38460, n_38461, n_38462, n_38463, n_38464, n_38465, n_38466, n_38467, n_38468, n_38469, n_38470, n_38471, n_38472, n_38473, n_38474, n_38475, n_38476, n_38477, n_38478, n_38479, n_38480, n_38481, y74, n_38482, n_38483, n_38484, n_38485, n_38486, n_38487, n_38488, n_38489, n_38490, n_38491, n_38492, y39, n_38493, n_38494, n_38495, n_38496, n_38497, n_38498, n_38499, n_38500, n_38501, n_38502, n_38503, n_38504, n_38505, n_38506, y73, n_38507, n_38508, n_38509, n_38510, n_38511, n_38512, n_38513, n_38514, n_38515, n_38516, n_38517, n_38518, n_38519, n_38520, n_38521, n_38522, n_38523, n_38524, y72, n_38525, n_38526, n_38527, n_38528, n_38529, n_38530, n_38531, y38, n_38532, n_38533, n_38534, n_38535, n_38536, n_38537, n_38538, n_38539, n_38540, n_38541, n_38542, n_38543, n_38544, n_38545, n_38546, n_38547, n_38548, n_38549, n_38550, n_38551, n_38552, y87, n_38553, n_38554, n_38555, n_38556, n_38557, n_38558, n_38559, n_38560, n_38561, n_38562, n_38563, n_38564, n_38565, n_38566, n_38567, n_38568, n_38569, y37, n_38570, n_38571, n_38572, n_38573, n_38574, n_38575, n_38576, n_38577, n_38578, n_38579, n_38580, n_38581, n_38582, n_38583, n_38584, n_38585, n_38586, n_38587, n_38588, n_38589, y86, n_38590, n_38591, n_38592, n_38593, n_38594, n_38595, y36, n_38596, n_38597, n_38598, n_38599, n_38600, n_38601, n_38602, n_38603, n_38604, n_38605, n_38606, n_38607, n_38608, n_38609, n_38610, n_38611, n_38612, n_38613, n_38614, n_38615, n_38616, y85, n_38617, n_38618, n_38619, n_38620, n_38621, n_38622, n_38623, n_38624, y35, n_38625, n_38626, n_38627, n_38628, n_38629, n_38630, n_38631, n_38632, n_38633, n_38634, n_38635, n_38636, n_38637, y84, n_38638, n_38639, n_38640, n_38641, n_38642, n_38643, n_38644, n_38645, n_38646, n_38647, n_38648, n_38649, n_38650, n_38651, n_38652, n_38653, y34, n_38654, n_38655, n_38656, n_38657, n_38658, n_38659, n_38660, n_38661, n_38662, n_38663, n_38664, n_38665, y83, n_38666, n_38667, n_38668, n_38669, n_38670, n_38671, n_38672, n_38673, n_38674, n_38675, n_38676, y33, n_38677, n_38678, n_38679, n_38680, n_38681, n_38682, n_38683, n_38684, n_38685, n_38686, n_38687, n_38688, n_38689, n_38690, n_38691, n_38692, n_38693, n_38694, n_38695, n_38696, n_38697, n_38698, n_38699, n_38700, n_38701, n_38702, n_38703, n_38704, y82, n_38705, n_38706, n_38707, n_38708, y32, n_38709, n_38710, n_38711, n_38712, n_38713, n_38714, n_38715, n_38716, n_38717, n_38718, n_38719, n_38720, n_38721, n_38722, n_38723, y81, n_38724, n_38725, n_38726, n_38727, n_38728, n_38729, n_38730, n_38731, n_38732, n_38733, n_38734, n_38735, n_38736, y47, n_38737, n_38738, n_38739, n_38740, n_38741, n_38742, n_38743, n_38744, n_38745, n_38746, n_38747, n_38748, n_38749, n_38750, n_38751, n_38752, n_38753, n_38754, n_38755, n_38756, n_38757, n_38758, n_38759, y80, n_38760, n_38761, n_38762, n_38763, n_38764, n_38765, n_38766, n_38767, n_38768, n_38769, y46, n_38770, n_38771, n_38772, n_38773, n_38774, n_38775, n_38776, n_38777, n_38778, n_38779, n_38780, n_38781, n_38782, y95, n_38783, n_38784, n_38785, n_38786, n_38787, n_38788, n_38789, n_38790, n_38791, n_38792, n_38793, n_38794, n_38795, n_38796, n_38797, n_38798, n_38799, y45, n_38800, n_38801, n_38802, n_38803, n_38804, n_38805, n_38806, n_38807, n_38808, n_38809, n_38810, n_38811, n_38812, n_38813, n_38814, n_38815, n_38816, n_38817, n_38818, n_38819, n_38820, n_38821, n_38822, y94, n_38823, n_38824, n_38825, n_38826, n_38827, n_38828, n_38829, y44, n_38830, n_38831, n_38832, n_38833, n_38834, n_38835, n_38836, n_38837, n_38838, n_38839, n_38840, n_38841, n_38842, n_38843, n_38844, n_38845, n_38846, n_38847, n_38848, n_38849, n_38850, n_38851, n_38852, y93, n_38853, n_38854, n_38855, n_38856, n_38857, n_38858, y43, n_38859, n_38860, n_38861, n_38862, n_38863, n_38864, n_38865, n_38866, n_38867, n_38868, n_38869, n_38870, n_38871, n_38872, n_38873, n_38874, n_38875, n_38876, n_38877, n_38878, n_38879, n_38880, n_38881, y92, n_38882, n_38883, n_38884, n_38885, n_38886, n_38887, n_38888, n_38889, y42, n_38890, n_38891, n_38892, n_38893, n_38894, n_38895, n_38896, n_38897, n_38898, n_38899, n_38900, n_38901, n_38902, n_38903, n_38904, n_38905, n_38906, n_38907, n_38908, n_38909, n_38910, n_38911, n_38912, y91, n_38913, n_38914, n_38915, n_38916, n_38917, n_38918, n_38919, n_38920, n_38921, y41, n_38922, n_38923, n_38924, n_38925, n_38926, n_38927, n_38928, n_38929, n_38930, n_38931, n_38932, n_38933, n_38934, y90, n_38935, n_38936, n_38937, n_38938, n_38939, n_38940, n_38941, n_38942, n_38943, n_38944, n_38945, n_38946, n_38947, n_38948, n_38949, n_38950, y40, n_38951, n_38952, n_38953, n_38954, n_38955, n_38956, n_38957, n_38958, n_38959, n_38960, n_38961, n_38962, n_38963, n_38964, n_38965, n_38966, n_38967, n_38968, n_38969, n_38970, n_38971, n_38972, n_38973, y89, n_38974, n_38975, n_38976, n_38977, n_38978, n_38979, n_38980, y55, n_38981, n_38982, n_38983, y88, n_38984, n_38985, n_38986, n_38987, n_38988, n_38989, n_38990, n_38991, n_38992, n_38993, n_38994, n_38995, n_38996, n_38997, n_38998, n_38999, n_39000, n_39001, y54, n_39002, n_39003, n_39004, n_39005, n_39006, n_39007, n_39008, n_39009, n_39010, n_39011, n_39012, n_39013, n_39014, n_39015, n_39016, n_39017, y53, n_39018, n_39019, n_39020, n_39021, n_39022, n_39023, n_39024, n_39025, y52, n_39026, n_39027, n_39028, n_39029, n_39030, n_39031, n_39032, n_39033, y51, n_39034, n_39035, n_39036, n_39037, y50, n_39038, n_39039, n_39040, n_39041, n_39042, n_39043, n_39044, y49, n_39045, n_39046, n_39047, n_39048, n_39049, y48, n_39050, n_39051, n_39052, n_39053, n_39054, n_39055, n_39056, n_39057, y63, n_39058, n_39059, n_39060, n_39061, n_39062, n_39063, n_39064, y62, n_39065, n_39066, n_39067, n_39068, n_39069, n_39070, y61, n_39071, n_39072, n_39073, n_39074, n_39075, n_39076, y60, n_39077, n_39078, n_39079, n_39080, n_39081, n_39082, n_39083, y59, n_39084, n_39085, n_39086, n_39087, y58, n_39088, n_39089, n_39090, n_39091, n_39092, n_39093, n_39094, y57, n_39095, y56;
assign n_0 = ~x6 & ~x7;
assign n_1 = x25 ^ x24;
assign n_2 = ~x5 & n_0;
assign n_3 = n_0 ^ x5;
assign n_4 = ~x4 & n_2;
assign n_5 = n_2 ^ x4;
assign n_6 = ~x3 & n_4;
assign n_7 = n_4 ^ x3;
assign n_8 = ~x2 & n_6;
assign n_9 = n_6 ^ x2;
assign n_10 = ~n_5 & ~n_7;
assign n_11 = ~x1 & n_8;
assign n_12 = n_8 ^ x1;
assign n_13 = ~n_9 & n_10;
assign n_14 = n_10 ^ n_9;
assign n_15 = ~x0 & n_11;
assign n_16 = n_11 ^ x0;
assign n_17 = n_13 & ~n_12;
assign n_18 = n_12 ^ n_13;
assign n_19 = ~x15 & n_15;
assign n_20 = n_15 ^ x15;
assign n_21 = n_16 & ~n_17;
assign n_22 = n_17 ^ n_16;
assign n_23 = ~x14 & n_19;
assign n_24 = n_19 ^ x14;
assign n_25 = n_20 & n_21;
assign n_26 = n_21 ^ n_20;
assign n_27 = ~x13 & n_23;
assign n_28 = n_23 ^ x13;
assign n_29 = n_24 & n_25;
assign n_30 = n_25 ^ n_24;
assign n_31 = ~x12 & n_27;
assign n_32 = n_27 ^ x12;
assign n_33 = ~n_29 & ~n_28;
assign n_34 = n_28 ^ n_29;
assign n_35 = ~x11 & n_31;
assign n_36 = n_31 ^ x11;
assign n_37 = ~n_33 & n_32;
assign n_38 = n_32 ^ n_33;
assign n_39 = n_35 ^ x10;
assign n_40 = ~x10 & n_35;
assign n_41 = n_36 & n_37;
assign n_42 = n_37 ^ n_36;
assign n_43 = ~x9 & n_40;
assign n_44 = n_40 ^ x9;
assign n_45 = n_39 ^ n_41;
assign n_46 = ~n_41 & ~n_39;
assign n_47 = ~x8 & n_43;
assign n_48 = n_43 ^ x8;
assign n_49 = n_44 & ~n_46;
assign n_50 = ~x23 & n_47;
assign n_51 = n_47 ^ x23;
assign n_52 = ~n_48 & ~n_49;
assign n_53 = n_49 ^ n_48;
assign n_54 = ~x22 & n_50;
assign n_55 = n_50 ^ x22;
assign n_56 = n_51 & ~n_52;
assign n_57 = n_52 ^ n_51;
assign n_58 = ~x21 & n_54;
assign n_59 = n_54 ^ x21;
assign n_60 = ~n_56 & ~n_55;
assign n_61 = n_55 ^ n_56;
assign n_62 = ~x20 & n_58;
assign n_63 = n_58 ^ x20;
assign n_64 = ~n_60 & n_59;
assign n_65 = n_59 ^ n_60;
assign n_66 = ~x19 & n_62;
assign n_67 = n_62 ^ x19;
assign n_68 = ~n_63 & ~n_64;
assign n_69 = n_64 ^ n_63;
assign n_70 = ~x18 & n_66;
assign n_71 = n_66 ^ x18;
assign n_72 = n_67 & ~n_68;
assign n_73 = n_68 ^ n_67;
assign n_74 = ~x17 & n_70;
assign n_75 = n_70 ^ x17;
assign n_76 = ~n_71 & ~n_72;
assign n_77 = n_72 ^ n_71;
assign n_78 = ~x16 & n_74;
assign n_79 = n_74 ^ x16;
assign n_80 = ~n_75 & n_76;
assign n_81 = n_76 ^ n_75;
assign n_82 = ~x31 & n_78;
assign n_83 = n_78 ^ x31;
assign n_84 = n_79 & ~n_80;
assign n_85 = n_80 ^ n_79;
assign n_86 = ~x30 & n_82;
assign n_87 = n_82 ^ x30;
assign n_88 = ~n_83 & ~n_84;
assign n_89 = n_84 ^ n_83;
assign n_90 = n_86 ^ x29;
assign n_91 = ~x29 & n_86;
assign n_92 = ~n_87 & n_88;
assign n_93 = n_88 ^ n_87;
assign n_94 = n_91 ^ x28;
assign n_95 = ~x28 & n_91;
assign n_96 = ~n_90 & n_92;
assign n_97 = n_92 ^ n_90;
assign n_98 = x39 & ~n_93;
assign n_99 = n_93 ^ x39;
assign n_100 = n_95 ^ x27;
assign n_101 = ~x27 & n_95;
assign n_102 = n_96 ^ n_94;
assign n_103 = n_94 & ~n_96;
assign n_104 = n_93 & n_97;
assign n_105 = n_97 ^ n_93;
assign n_106 = n_101 ^ x26;
assign n_107 = ~x26 & n_101;
assign n_108 = n_103 ^ n_100;
assign n_109 = ~n_100 & ~n_103;
assign n_110 = ~n_102 & n_104;
assign n_111 = n_104 ^ n_102;
assign n_112 = n_105 ^ x38;
assign n_113 = n_98 ^ n_105;
assign n_114 = n_107 ^ x25;
assign n_115 = n_109 ^ n_106;
assign n_116 = n_106 & ~n_109;
assign n_117 = ~n_110 & n_108;
assign n_118 = n_108 ^ n_110;
assign n_119 = n_111 ^ n_105;
assign n_120 = n_105 & ~n_111;
assign n_121 = n_98 ^ n_112;
assign n_122 = n_112 & ~n_113;
assign n_123 = n_114 ^ n_116;
assign n_124 = n_107 ^ n_116;
assign n_125 = ~n_117 & ~n_115;
assign n_126 = n_115 ^ n_117;
assign n_127 = n_119 ^ x37;
assign n_128 = n_120 ^ x36;
assign n_129 = n_122 ^ x38;
assign n_130 = ~n_114 & n_124;
assign n_131 = n_125 & ~n_123;
assign n_132 = n_123 ^ n_125;
assign n_133 = n_126 ^ n_120;
assign n_134 = n_120 & n_126;
assign n_135 = n_129 ^ n_119;
assign n_136 = n_130 ^ n_1;
assign n_137 = n_133 ^ x35;
assign n_138 = n_132 ^ n_134;
assign n_139 = n_134 & ~n_132;
assign n_140 = ~n_135 & n_127;
assign n_141 = n_135 ^ x37;
assign n_142 = n_131 & ~n_136;
assign n_143 = n_136 ^ n_131;
assign n_144 = n_138 ^ x34;
assign n_145 = n_140 ^ x37;
assign n_146 = ~n_141 & ~n_121;
assign n_147 = n_121 ^ n_141;
assign n_148 = x7 & ~n_142;
assign n_149 = n_142 ^ x7;
assign n_150 = n_143 ^ n_139;
assign n_151 = n_139 & ~n_143;
assign n_152 = n_145 ^ n_120;
assign n_153 = ~x6 & n_148;
assign n_154 = n_148 ^ x7;
assign n_155 = n_150 ^ x33;
assign n_156 = n_151 ^ x32;
assign n_157 = ~n_152 & n_128;
assign n_158 = n_152 ^ x36;
assign n_159 = ~n_3 & n_153;
assign n_160 = n_153 ^ n_3;
assign n_161 = n_154 ^ x6;
assign n_162 = n_157 ^ x36;
assign n_163 = ~n_146 & n_158;
assign n_164 = n_158 ^ n_146;
assign n_165 = n_159 ^ n_7;
assign n_166 = n_159 ^ n_5;
assign n_167 = n_161 ^ n_151;
assign n_168 = ~n_151 & ~n_161;
assign n_169 = n_162 ^ n_133;
assign n_170 = ~n_5 & ~n_165;
assign n_171 = n_167 ^ x47;
assign n_172 = n_168 ^ n_160;
assign n_173 = n_160 & n_168;
assign n_174 = n_169 & ~n_137;
assign n_175 = n_169 ^ x35;
assign n_176 = n_170 ^ n_7;
assign n_177 = n_172 ^ x46;
assign n_178 = ~n_173 & n_166;
assign n_179 = n_166 ^ n_173;
assign n_180 = n_174 ^ x35;
assign n_181 = ~n_163 & n_175;
assign n_182 = n_175 ^ n_163;
assign n_183 = ~n_10 & ~n_176;
assign n_184 = n_176 ^ n_10;
assign n_185 = n_178 ^ x44;
assign n_186 = n_179 ^ x45;
assign n_187 = n_180 ^ n_138;
assign n_188 = n_14 & ~n_183;
assign n_189 = n_183 ^ n_14;
assign n_190 = n_184 ^ n_159;
assign n_191 = ~n_187 & n_144;
assign n_192 = n_187 ^ x34;
assign n_193 = ~n_188 & ~n_18;
assign n_194 = n_18 ^ n_188;
assign n_195 = n_99 ^ n_189;
assign n_196 = ~n_189 & n_178;
assign n_197 = n_178 ^ n_189;
assign n_198 = n_190 ^ n_159;
assign n_199 = n_191 ^ x34;
assign n_200 = ~n_181 & n_192;
assign n_201 = n_192 ^ n_181;
assign n_202 = ~n_193 & ~n_22;
assign n_203 = n_22 ^ n_193;
assign n_204 = n_121 ^ n_194;
assign n_205 = ~n_194 & ~n_196;
assign n_206 = n_196 ^ n_194;
assign n_207 = n_197 ^ x43;
assign n_208 = n_199 ^ n_150;
assign n_209 = ~n_26 & ~n_202;
assign n_210 = n_202 ^ n_26;
assign n_211 = n_147 ^ n_203;
assign n_212 = ~n_205 & n_203;
assign n_213 = n_203 ^ n_205;
assign n_214 = n_206 ^ x42;
assign n_215 = n_208 ^ x33;
assign n_216 = ~n_208 & n_155;
assign n_217 = ~n_30 & n_209;
assign n_218 = n_209 ^ n_30;
assign n_219 = n_164 ^ n_210;
assign n_220 = n_212 ^ x40;
assign n_221 = n_213 ^ x41;
assign n_222 = ~n_215 & ~n_200;
assign n_223 = n_200 ^ n_215;
assign n_224 = n_216 ^ x33;
assign n_225 = ~n_217 & ~n_34;
assign n_226 = n_34 ^ n_217;
assign n_227 = n_182 ^ n_218;
assign n_228 = ~n_212 & n_218;
assign n_229 = n_218 ^ n_212;
assign n_230 = n_224 ^ n_151;
assign n_231 = ~n_225 & n_38;
assign n_232 = n_38 ^ n_225;
assign n_233 = n_201 ^ n_226;
assign n_234 = n_226 & ~n_228;
assign n_235 = n_228 ^ n_226;
assign n_236 = n_229 ^ x55;
assign n_237 = n_230 ^ x32;
assign n_238 = ~n_230 & n_156;
assign n_239 = ~n_42 & n_231;
assign n_240 = n_231 ^ n_42;
assign n_241 = n_232 ^ n_223;
assign n_242 = n_232 & ~n_234;
assign n_243 = n_234 ^ n_232;
assign n_244 = n_235 ^ x54;
assign n_245 = ~n_222 & n_237;
assign n_246 = n_237 ^ n_222;
assign n_247 = n_238 ^ x32;
assign n_248 = ~n_45 & ~n_239;
assign n_249 = n_239 ^ n_45;
assign n_250 = n_242 ^ x52;
assign n_251 = ~x53 & n_243;
assign n_252 = n_243 ^ x53;
assign n_253 = n_246 ^ n_240;
assign n_254 = n_247 ^ n_167;
assign n_255 = n_248 ^ n_44;
assign n_256 = n_44 & n_248;
assign n_257 = ~n_242 & n_249;
assign n_258 = n_249 ^ n_242;
assign n_259 = n_251 ^ n_252;
assign n_260 = n_254 ^ x47;
assign n_261 = ~n_254 & n_171;
assign n_262 = n_255 ^ n_46;
assign n_263 = n_53 & ~n_256;
assign n_264 = n_256 ^ n_53;
assign n_265 = n_258 ^ x51;
assign n_266 = ~n_245 & ~n_260;
assign n_267 = n_260 ^ n_245;
assign n_268 = n_261 ^ x47;
assign n_269 = ~n_262 & n_257;
assign n_270 = n_257 ^ n_262;
assign n_271 = n_57 & n_263;
assign n_272 = n_263 ^ n_57;
assign n_273 = n_267 ^ n_249;
assign n_274 = n_268 ^ n_172;
assign n_275 = ~n_269 & n_264;
assign n_276 = n_264 ^ n_269;
assign n_277 = n_270 ^ x50;
assign n_278 = n_61 & n_271;
assign n_279 = n_271 ^ n_61;
assign n_280 = n_274 ^ x46;
assign n_281 = ~n_274 & n_177;
assign n_282 = n_275 ^ x48;
assign n_283 = n_276 ^ x49;
assign n_284 = ~x49 & n_276;
assign n_285 = n_278 ^ n_65;
assign n_286 = n_65 & n_278;
assign n_287 = ~n_279 & n_275;
assign n_288 = n_275 ^ n_279;
assign n_289 = n_266 ^ n_280;
assign n_290 = ~n_280 & n_266;
assign n_291 = n_281 ^ x46;
assign n_292 = n_283 ^ n_284;
assign n_293 = n_286 ^ n_69;
assign n_294 = n_69 & n_286;
assign n_295 = ~n_285 & n_287;
assign n_296 = n_287 ^ n_285;
assign n_297 = ~x63 & n_288;
assign n_298 = n_288 ^ x63;
assign n_299 = n_262 ^ n_289;
assign n_300 = n_291 ^ n_179;
assign n_301 = n_73 & n_294;
assign n_302 = n_294 ^ n_73;
assign n_303 = n_295 ^ n_293;
assign n_304 = ~n_293 & n_295;
assign n_305 = n_296 ^ x62;
assign n_306 = n_298 ^ n_297;
assign n_307 = ~n_300 & n_186;
assign n_308 = n_300 ^ x45;
assign n_309 = n_301 ^ n_77;
assign n_310 = ~n_77 & ~n_301;
assign n_311 = n_303 ^ x61;
assign n_312 = n_304 ^ x60;
assign n_313 = ~x60 & n_304;
assign n_314 = n_307 ^ x45;
assign n_315 = n_290 & ~n_308;
assign n_316 = n_308 ^ n_290;
assign n_317 = n_304 ^ n_309;
assign n_318 = n_309 & ~n_304;
assign n_319 = n_81 ^ n_310;
assign n_320 = ~n_310 & ~n_81;
assign n_321 = n_312 ^ n_313;
assign n_322 = n_314 ^ n_178;
assign n_323 = n_314 ^ n_185;
assign n_324 = n_264 ^ n_316;
assign n_325 = n_317 ^ x59;
assign n_326 = n_318 ^ n_319;
assign n_327 = ~n_319 & ~n_318;
assign n_328 = n_320 ^ n_85;
assign n_329 = n_85 & n_320;
assign n_330 = n_185 & ~n_322;
assign n_331 = ~n_315 & n_323;
assign n_332 = n_323 ^ n_315;
assign n_333 = n_326 ^ x58;
assign n_334 = n_327 ^ n_328;
assign n_335 = ~n_328 & n_327;
assign n_336 = n_329 ^ n_89;
assign n_337 = n_330 ^ x44;
assign n_338 = n_272 ^ n_332;
assign n_339 = n_334 ^ x57;
assign n_340 = n_335 ^ x56;
assign n_341 = n_337 ^ n_197;
assign n_342 = ~n_341 & n_207;
assign n_343 = n_341 ^ x43;
assign n_344 = n_342 ^ x43;
assign n_345 = ~n_331 & ~n_343;
assign n_346 = n_343 ^ n_331;
assign n_347 = n_344 ^ n_206;
assign n_348 = n_279 ^ n_346;
assign n_349 = ~n_347 & n_214;
assign n_350 = n_347 ^ x42;
assign n_351 = n_349 ^ x42;
assign n_352 = n_345 & ~n_350;
assign n_353 = n_350 ^ n_345;
assign n_354 = n_351 ^ n_213;
assign n_355 = n_285 ^ n_353;
assign n_356 = ~n_354 & n_221;
assign n_357 = n_354 ^ x41;
assign n_358 = n_356 ^ x41;
assign n_359 = ~n_352 & n_357;
assign n_360 = n_357 ^ n_352;
assign n_361 = n_358 ^ n_212;
assign n_362 = n_293 ^ n_360;
assign n_363 = ~n_361 & n_220;
assign n_364 = n_361 ^ x40;
assign n_365 = n_363 ^ x40;
assign n_366 = ~n_359 & ~n_364;
assign n_367 = n_364 ^ n_359;
assign n_368 = n_365 ^ n_229;
assign n_369 = n_302 ^ n_367;
assign n_370 = n_368 & ~n_236;
assign n_371 = n_368 ^ x55;
assign n_372 = n_370 ^ x55;
assign n_373 = n_371 & n_366;
assign n_374 = n_366 ^ n_371;
assign n_375 = n_372 ^ n_235;
assign n_376 = n_374 ^ n_309;
assign n_377 = ~n_375 & n_244;
assign n_378 = n_375 ^ x54;
assign n_379 = n_377 ^ x54;
assign n_380 = n_373 & ~n_378;
assign n_381 = n_378 ^ n_373;
assign n_382 = ~n_251 & n_379;
assign n_383 = n_379 ^ n_252;
assign n_384 = n_381 ^ n_319;
assign n_385 = n_382 ^ n_242;
assign n_386 = ~n_259 & ~n_382;
assign n_387 = n_380 & n_383;
assign n_388 = n_383 ^ n_380;
assign n_389 = ~n_250 & n_385;
assign n_390 = n_386 ^ n_250;
assign n_391 = n_336 ^ n_387;
assign n_392 = n_388 ^ n_328;
assign n_393 = n_389 ^ x52;
assign n_394 = ~n_387 & n_390;
assign n_395 = n_391 ^ n_390;
assign n_396 = ~n_259 & ~n_393;
assign n_397 = n_258 ^ n_396;
assign n_398 = n_397 & n_265;
assign n_399 = n_397 ^ x51;
assign n_400 = n_398 ^ x51;
assign n_401 = ~n_399 & n_394;
assign n_402 = n_394 ^ n_399;
assign n_403 = n_400 ^ n_270;
assign n_404 = ~n_93 & ~n_402;
assign n_405 = n_402 ^ n_93;
assign n_406 = ~n_403 & n_277;
assign n_407 = n_403 ^ x50;
assign n_408 = n_404 ^ n_105;
assign n_409 = n_404 ^ n_402;
assign n_410 = n_406 ^ x50;
assign n_411 = n_401 & n_407;
assign n_412 = n_407 ^ n_401;
assign n_413 = n_409 ^ x71;
assign n_414 = x71 & n_409;
assign n_415 = ~n_284 & n_410;
assign n_416 = n_410 ^ n_283;
assign n_417 = n_412 ^ n_404;
assign n_418 = n_412 ^ n_408;
assign n_419 = n_414 ^ x70;
assign n_420 = n_415 ^ n_275;
assign n_421 = ~n_292 & ~n_415;
assign n_422 = n_416 & ~n_411;
assign n_423 = n_411 ^ n_416;
assign n_424 = n_408 & ~n_417;
assign n_425 = n_105 & n_418;
assign n_426 = ~n_282 & n_420;
assign n_427 = n_421 ^ n_282;
assign n_428 = n_423 ^ n_111;
assign n_429 = n_424 ^ n_105;
assign n_430 = n_414 ^ n_425;
assign n_431 = n_426 ^ x48;
assign n_432 = ~n_427 & n_422;
assign n_433 = n_422 ^ n_427;
assign n_434 = n_429 ^ n_423;
assign n_435 = n_429 ^ n_111;
assign n_436 = n_430 ^ x70;
assign n_437 = n_430 & n_419;
assign n_438 = ~n_292 & ~n_431;
assign n_439 = n_118 ^ n_433;
assign n_440 = ~n_428 & ~n_434;
assign n_441 = n_435 ^ n_423;
assign n_442 = ~n_413 & n_436;
assign n_443 = n_436 ^ n_413;
assign n_444 = n_437 ^ x70;
assign n_445 = ~n_297 & ~n_438;
assign n_446 = n_298 ^ n_438;
assign n_447 = n_440 ^ n_111;
assign n_448 = ~n_111 & ~n_441;
assign n_449 = ~n_445 & ~n_306;
assign n_450 = n_445 & n_313;
assign n_451 = ~n_432 & n_446;
assign n_452 = n_446 ^ n_432;
assign n_453 = n_447 ^ n_433;
assign n_454 = n_447 ^ n_118;
assign n_455 = n_448 ^ n_425;
assign n_456 = ~n_425 & ~n_448;
assign n_457 = n_449 ^ n_296;
assign n_458 = n_449 ^ n_305;
assign n_459 = n_450 ^ n_449;
assign n_460 = n_452 ^ n_126;
assign n_461 = n_439 & n_453;
assign n_462 = n_454 ^ n_433;
assign n_463 = n_444 ^ n_455;
assign n_464 = n_455 ^ x69;
assign n_465 = ~n_305 & ~n_457;
assign n_466 = n_458 & n_451;
assign n_467 = n_451 ^ n_458;
assign n_468 = n_459 ^ n_296;
assign n_469 = n_461 ^ n_118;
assign n_470 = ~n_118 & ~n_462;
assign n_471 = n_463 ^ x69;
assign n_472 = n_463 & ~n_464;
assign n_473 = n_465 ^ x62;
assign n_474 = n_467 ^ n_132;
assign n_475 = ~n_305 & ~n_468;
assign n_476 = n_469 ^ n_452;
assign n_477 = n_456 ^ n_470;
assign n_478 = n_470 & n_456;
assign n_479 = ~n_442 & ~n_471;
assign n_480 = n_471 ^ n_442;
assign n_481 = n_472 ^ x69;
assign n_482 = n_473 ^ n_303;
assign n_483 = n_473 ^ n_311;
assign n_484 = x62 ^ n_475;
assign n_485 = n_476 & ~n_460;
assign n_486 = n_126 & n_476;
assign n_487 = n_476 ^ n_126;
assign n_488 = n_477 ^ x68;
assign n_489 = n_481 ^ n_477;
assign n_490 = ~n_311 & n_482;
assign n_491 = n_466 & ~n_483;
assign n_492 = n_483 ^ n_466;
assign n_493 = n_484 ^ n_303;
assign n_494 = n_485 ^ n_126;
assign n_495 = n_486 ^ n_478;
assign n_496 = n_478 & ~n_486;
assign n_497 = n_489 ^ x68;
assign n_498 = n_489 & ~n_488;
assign n_499 = n_490 ^ x61;
assign n_500 = n_492 ^ n_143;
assign n_501 = ~n_311 & ~n_493;
assign n_502 = n_494 ^ n_467;
assign n_503 = n_494 ^ n_132;
assign n_504 = n_495 ^ x67;
assign n_505 = ~n_479 & n_497;
assign n_506 = n_497 ^ n_479;
assign n_507 = n_498 ^ x68;
assign n_508 = n_499 ^ n_312;
assign n_509 = n_303 ^ n_501;
assign n_510 = ~n_474 & ~n_502;
assign n_511 = n_503 ^ n_467;
assign n_512 = n_507 ^ x67;
assign n_513 = n_507 ^ n_495;
assign n_514 = n_508 & ~n_491;
assign n_515 = n_491 ^ n_508;
assign n_516 = n_509 & ~n_321;
assign n_517 = n_510 ^ n_132;
assign n_518 = ~n_132 & ~n_511;
assign n_519 = n_512 ^ n_495;
assign n_520 = n_504 & ~n_513;
assign n_521 = n_149 ^ n_515;
assign n_522 = n_317 ^ n_516;
assign n_523 = n_517 ^ n_492;
assign n_524 = n_517 ^ n_143;
assign n_525 = n_518 ^ n_496;
assign n_526 = n_496 & ~n_518;
assign n_527 = n_505 & ~n_519;
assign n_528 = n_519 ^ n_505;
assign n_529 = n_520 ^ x67;
assign n_530 = n_522 ^ x59;
assign n_531 = n_522 & n_325;
assign n_532 = n_500 & ~n_523;
assign n_533 = n_524 ^ n_492;
assign n_534 = n_525 ^ x66;
assign n_535 = n_529 ^ n_525;
assign n_536 = ~n_514 & ~n_530;
assign n_537 = n_530 ^ n_514;
assign n_538 = n_531 ^ x59;
assign n_539 = n_532 ^ n_143;
assign n_540 = ~n_143 & ~n_533;
assign n_541 = n_535 ^ x66;
assign n_542 = ~n_535 & n_534;
assign n_543 = n_537 ^ n_161;
assign n_544 = n_538 ^ n_326;
assign n_545 = n_539 ^ n_515;
assign n_546 = ~n_540 & n_526;
assign n_547 = n_526 ^ n_540;
assign n_548 = n_527 ^ n_541;
assign n_549 = n_541 & ~n_527;
assign n_550 = n_542 ^ x66;
assign n_551 = n_544 ^ x58;
assign n_552 = ~n_544 & n_333;
assign n_553 = n_545 & n_521;
assign n_554 = ~n_545 & ~n_149;
assign n_555 = n_149 ^ n_545;
assign n_556 = n_547 ^ x65;
assign n_557 = n_550 ^ n_547;
assign n_558 = ~n_536 & ~n_551;
assign n_559 = n_551 ^ n_536;
assign n_560 = n_552 ^ x58;
assign n_561 = n_553 ^ n_149;
assign n_562 = n_554 & n_546;
assign n_563 = n_546 ^ n_554;
assign n_564 = ~n_557 & n_556;
assign n_565 = n_557 ^ x65;
assign n_566 = n_559 ^ n_160;
assign n_567 = n_560 ^ n_334;
assign n_568 = n_561 ^ n_537;
assign n_569 = n_563 ^ x64;
assign n_570 = n_564 ^ x65;
assign n_571 = ~n_549 & ~n_565;
assign n_572 = n_565 ^ n_549;
assign n_573 = n_567 ^ x57;
assign n_574 = n_567 & ~n_339;
assign n_575 = ~n_568 & ~n_543;
assign n_576 = n_161 & n_568;
assign n_577 = n_568 ^ n_161;
assign n_578 = n_570 ^ n_563;
assign n_579 = n_558 ^ n_573;
assign n_580 = n_573 & n_558;
assign n_581 = n_574 ^ x57;
assign n_582 = n_575 ^ n_161;
assign n_583 = ~n_562 & ~n_576;
assign n_584 = n_576 ^ n_562;
assign n_585 = n_578 & ~n_569;
assign n_586 = n_578 ^ x64;
assign n_587 = n_579 ^ n_166;
assign n_588 = n_581 ^ n_340;
assign n_589 = n_582 ^ n_559;
assign n_590 = n_582 ^ n_160;
assign n_591 = n_584 ^ x79;
assign n_592 = n_585 ^ x64;
assign n_593 = n_571 & n_586;
assign n_594 = n_586 ^ n_571;
assign n_595 = n_588 ^ n_580;
assign n_596 = ~n_566 & ~n_589;
assign n_597 = n_590 ^ n_559;
assign n_598 = n_592 ^ n_584;
assign n_599 = n_592 ^ x79;
assign n_600 = n_198 ^ n_595;
assign n_601 = n_596 ^ n_160;
assign n_602 = ~n_160 & n_597;
assign n_603 = n_591 & ~n_598;
assign n_604 = n_599 ^ n_584;
assign n_605 = n_601 ^ n_579;
assign n_606 = n_601 ^ n_166;
assign n_607 = ~n_602 & n_583;
assign n_608 = n_583 ^ n_602;
assign n_609 = n_603 ^ x79;
assign n_610 = ~n_593 & n_604;
assign n_611 = n_604 ^ n_593;
assign n_612 = ~n_587 & n_605;
assign n_613 = n_606 ^ n_579;
assign n_614 = n_608 ^ x78;
assign n_615 = n_609 ^ n_608;
assign n_616 = n_612 ^ n_166;
assign n_617 = n_166 & ~n_613;
assign n_618 = n_615 & ~n_614;
assign n_619 = n_615 ^ x78;
assign n_620 = n_616 ^ n_595;
assign n_621 = ~n_607 & ~n_617;
assign n_622 = n_617 ^ n_607;
assign n_623 = n_618 ^ x78;
assign n_624 = ~n_619 & n_610;
assign n_625 = n_610 ^ n_619;
assign n_626 = n_620 & n_600;
assign n_627 = ~n_620 & n_198;
assign n_628 = n_198 ^ n_620;
assign n_629 = n_622 ^ x77;
assign n_630 = n_623 ^ n_622;
assign n_631 = n_626 ^ n_198;
assign n_632 = n_621 & n_627;
assign n_633 = n_627 ^ n_621;
assign n_634 = n_630 & ~n_629;
assign n_635 = n_630 ^ x77;
assign n_636 = n_631 ^ n_189;
assign n_637 = n_631 ^ n_99;
assign n_638 = n_633 ^ x76;
assign n_639 = n_634 ^ x77;
assign n_640 = n_624 & ~n_635;
assign n_641 = n_635 ^ n_624;
assign n_642 = n_195 & ~n_636;
assign n_643 = ~n_189 & ~n_637;
assign n_644 = n_637 ^ n_189;
assign n_645 = n_639 ^ n_633;
assign n_646 = n_642 ^ n_99;
assign n_647 = n_632 & ~n_643;
assign n_648 = n_643 ^ n_632;
assign n_649 = n_645 & ~n_638;
assign n_650 = n_645 ^ x76;
assign n_651 = n_646 ^ n_194;
assign n_652 = n_646 ^ n_121;
assign n_653 = n_648 ^ x75;
assign n_654 = n_649 ^ x76;
assign n_655 = n_640 & ~n_650;
assign n_656 = n_650 ^ n_640;
assign n_657 = n_204 & ~n_651;
assign n_658 = n_194 & n_652;
assign n_659 = n_652 ^ n_194;
assign n_660 = n_654 ^ n_648;
assign n_661 = n_657 ^ n_121;
assign n_662 = ~n_658 & ~n_647;
assign n_663 = n_647 ^ n_658;
assign n_664 = ~n_660 & n_653;
assign n_665 = n_660 ^ x75;
assign n_666 = n_661 ^ n_203;
assign n_667 = n_663 ^ x74;
assign n_668 = n_664 ^ x75;
assign n_669 = ~n_665 & ~n_655;
assign n_670 = n_655 ^ n_665;
assign n_671 = n_666 & ~n_211;
assign n_672 = n_147 ^ n_666;
assign n_673 = n_668 ^ n_663;
assign n_674 = n_671 ^ n_147;
assign n_675 = n_203 & n_672;
assign n_676 = n_672 ^ n_203;
assign n_677 = ~n_673 & n_667;
assign n_678 = n_673 ^ x74;
assign n_679 = n_674 ^ n_210;
assign n_680 = n_674 ^ n_164;
assign n_681 = ~n_675 & ~n_662;
assign n_682 = n_662 ^ n_675;
assign n_683 = n_677 ^ x74;
assign n_684 = n_669 & ~n_678;
assign n_685 = n_678 ^ n_669;
assign n_686 = n_219 & ~n_679;
assign n_687 = n_210 & n_680;
assign n_688 = n_680 ^ n_210;
assign n_689 = n_682 ^ x73;
assign n_690 = n_683 ^ n_682;
assign n_691 = n_686 ^ n_164;
assign n_692 = n_681 & n_687;
assign n_693 = n_687 ^ n_681;
assign n_694 = n_690 & ~n_689;
assign n_695 = n_690 ^ x73;
assign n_696 = n_691 ^ n_218;
assign n_697 = n_691 ^ n_227;
assign n_698 = n_693 ^ x72;
assign n_699 = n_694 ^ x73;
assign n_700 = n_684 & n_695;
assign n_701 = n_227 & n_696;
assign n_702 = ~n_218 & ~n_697;
assign n_703 = n_697 ^ n_218;
assign n_704 = n_699 ^ n_693;
assign n_705 = n_701 ^ n_182;
assign n_706 = ~n_692 & ~n_702;
assign n_707 = n_702 ^ n_692;
assign n_708 = n_704 & ~n_698;
assign n_709 = n_704 ^ x72;
assign n_710 = n_705 ^ n_226;
assign n_711 = n_707 ^ x87;
assign n_712 = n_708 ^ x72;
assign n_713 = ~n_700 & ~n_709;
assign n_714 = n_709 ^ n_700;
assign n_715 = ~n_710 & ~n_233;
assign n_716 = n_201 ^ n_710;
assign n_717 = n_712 ^ n_707;
assign n_718 = n_712 ^ n_711;
assign n_719 = n_714 & n_405;
assign n_720 = n_714 ^ n_93;
assign n_721 = n_405 ^ n_714;
assign n_722 = n_715 ^ n_201;
assign n_723 = n_413 ^ n_716;
assign n_724 = n_226 & ~n_716;
assign n_725 = n_716 ^ n_226;
assign n_726 = n_711 & ~n_717;
assign n_727 = n_718 & n_713;
assign n_728 = n_713 ^ n_718;
assign n_729 = n_719 ^ n_418;
assign n_730 = ~n_402 & n_720;
assign n_731 = n_722 ^ n_232;
assign n_732 = n_722 ^ n_223;
assign n_733 = ~n_706 & ~n_724;
assign n_734 = n_724 ^ n_706;
assign n_735 = n_726 ^ x87;
assign n_736 = n_728 ^ n_719;
assign n_737 = n_728 ^ n_729;
assign n_738 = n_730 ^ n_93;
assign n_739 = ~n_241 & n_731;
assign n_740 = ~n_232 & n_732;
assign n_741 = n_732 ^ n_232;
assign n_742 = n_734 ^ x86;
assign n_743 = n_735 ^ n_734;
assign n_744 = n_729 & ~n_736;
assign n_745 = n_417 & n_737;
assign n_746 = x103 & n_738;
assign n_747 = n_738 ^ x103;
assign n_748 = n_739 ^ n_223;
assign n_749 = ~n_740 & ~n_733;
assign n_750 = n_733 ^ n_740;
assign n_751 = n_443 ^ n_741;
assign n_752 = n_743 & ~n_742;
assign n_753 = n_743 ^ x86;
assign n_754 = n_744 ^ n_418;
assign n_755 = n_745 ^ n_105;
assign n_756 = n_746 ^ x102;
assign n_757 = n_240 ^ n_748;
assign n_758 = n_750 ^ x85;
assign n_759 = n_752 ^ x86;
assign n_760 = n_727 & ~n_753;
assign n_761 = n_753 ^ n_727;
assign n_762 = n_754 ^ n_441;
assign n_763 = ~n_738 & n_755;
assign n_764 = n_755 ^ n_738;
assign n_765 = n_757 & ~n_253;
assign n_766 = n_246 ^ n_757;
assign n_767 = n_759 ^ n_750;
assign n_768 = n_761 ^ n_441;
assign n_769 = n_754 ^ n_761;
assign n_770 = n_762 ^ n_761;
assign n_771 = n_764 ^ n_746;
assign n_772 = n_764 ^ n_756;
assign n_773 = n_765 ^ n_246;
assign n_774 = ~n_240 & n_766;
assign n_775 = n_480 ^ n_766;
assign n_776 = n_766 ^ n_240;
assign n_777 = ~n_767 & n_758;
assign n_778 = n_767 ^ x85;
assign n_779 = n_768 & n_769;
assign n_780 = n_434 & n_770;
assign n_781 = n_756 & n_771;
assign n_782 = n_773 ^ n_249;
assign n_783 = n_774 & ~n_749;
assign n_784 = n_749 ^ n_774;
assign n_785 = n_777 ^ x85;
assign n_786 = n_760 & n_778;
assign n_787 = n_778 ^ n_760;
assign n_788 = n_779 ^ n_441;
assign n_789 = n_780 ^ n_111;
assign n_790 = n_781 ^ x102;
assign n_791 = n_782 & ~n_273;
assign n_792 = n_267 ^ n_782;
assign n_793 = n_784 ^ x84;
assign n_794 = n_785 ^ n_784;
assign n_795 = n_787 ^ n_462;
assign n_796 = n_788 ^ n_787;
assign n_797 = n_763 & ~n_789;
assign n_798 = n_789 ^ n_763;
assign n_799 = n_791 ^ n_267;
assign n_800 = n_249 & n_792;
assign n_801 = n_506 ^ n_792;
assign n_802 = n_792 ^ n_249;
assign n_803 = ~n_794 & n_793;
assign n_804 = n_794 ^ x84;
assign n_805 = n_796 & ~n_795;
assign n_806 = n_796 ^ n_462;
assign n_807 = n_790 ^ n_798;
assign n_808 = n_798 ^ x101;
assign n_809 = n_799 ^ n_289;
assign n_810 = n_799 ^ n_262;
assign n_811 = ~n_800 & n_783;
assign n_812 = n_783 ^ n_800;
assign n_813 = n_803 ^ x84;
assign n_814 = n_804 & n_786;
assign n_815 = n_786 ^ n_804;
assign n_816 = n_805 ^ n_462;
assign n_817 = ~n_453 & n_806;
assign n_818 = n_807 ^ x101;
assign n_819 = n_807 & ~n_808;
assign n_820 = ~n_299 & n_809;
assign n_821 = n_810 ^ n_289;
assign n_822 = n_812 ^ x83;
assign n_823 = n_813 ^ n_812;
assign n_824 = n_487 ^ n_815;
assign n_825 = n_816 ^ n_815;
assign n_826 = n_816 ^ n_487;
assign n_827 = n_817 ^ n_118;
assign n_828 = n_818 & n_772;
assign n_829 = n_772 ^ n_818;
assign n_830 = n_819 ^ x101;
assign n_831 = n_820 ^ n_262;
assign n_832 = ~n_262 & n_821;
assign n_833 = n_528 ^ n_821;
assign n_834 = ~n_823 & n_822;
assign n_835 = n_823 ^ x83;
assign n_836 = ~n_824 & n_825;
assign n_837 = n_826 ^ n_815;
assign n_838 = ~n_827 & ~n_797;
assign n_839 = n_797 ^ n_827;
assign n_840 = n_830 ^ x100;
assign n_841 = n_831 ^ n_316;
assign n_842 = n_811 & ~n_832;
assign n_843 = n_832 ^ n_811;
assign n_844 = n_834 ^ x83;
assign n_845 = n_835 & n_814;
assign n_846 = n_814 ^ n_835;
assign n_847 = n_836 ^ n_487;
assign n_848 = ~n_476 & n_837;
assign n_849 = n_839 ^ x100;
assign n_850 = n_830 ^ n_839;
assign n_851 = n_840 ^ n_839;
assign n_852 = n_841 & n_324;
assign n_853 = ~n_264 & ~n_841;
assign n_854 = n_841 ^ n_264;
assign n_855 = n_843 ^ x82;
assign n_856 = n_844 ^ n_843;
assign n_857 = n_846 ^ n_511;
assign n_858 = n_847 ^ n_846;
assign n_859 = n_848 ^ n_126;
assign n_860 = ~n_849 & n_850;
assign n_861 = n_851 & n_828;
assign n_862 = n_828 ^ n_851;
assign n_863 = n_852 ^ n_264;
assign n_864 = ~n_842 & ~n_853;
assign n_865 = n_853 ^ n_842;
assign n_866 = n_548 ^ n_854;
assign n_867 = ~n_856 & n_855;
assign n_868 = n_856 ^ x82;
assign n_869 = n_858 & ~n_857;
assign n_870 = n_858 ^ n_511;
assign n_871 = ~n_838 & n_859;
assign n_872 = n_859 ^ n_838;
assign n_873 = n_860 ^ x100;
assign n_874 = n_863 ^ n_332;
assign n_875 = n_865 ^ x81;
assign n_876 = n_867 ^ x82;
assign n_877 = ~n_845 & ~n_868;
assign n_878 = n_868 ^ n_845;
assign n_879 = n_869 ^ n_511;
assign n_880 = n_502 & n_870;
assign n_881 = n_872 ^ x99;
assign n_882 = n_873 ^ n_872;
assign n_883 = ~n_874 & n_272;
assign n_884 = n_874 & n_338;
assign n_885 = n_272 ^ n_874;
assign n_886 = n_876 ^ n_865;
assign n_887 = n_878 ^ n_533;
assign n_888 = n_879 ^ n_878;
assign n_889 = n_879 ^ n_533;
assign n_890 = n_880 ^ n_132;
assign n_891 = n_882 & ~n_881;
assign n_892 = n_882 ^ x99;
assign n_893 = n_883 ^ n_864;
assign n_894 = ~n_864 & n_883;
assign n_895 = n_884 ^ n_272;
assign n_896 = n_572 ^ n_885;
assign n_897 = ~n_886 & n_875;
assign n_898 = n_886 ^ x81;
assign n_899 = n_887 & ~n_888;
assign n_900 = n_889 ^ n_878;
assign n_901 = ~n_890 & n_871;
assign n_902 = n_871 ^ n_890;
assign n_903 = n_891 ^ x99;
assign n_904 = ~n_861 & ~n_892;
assign n_905 = n_892 ^ n_861;
assign n_906 = n_893 ^ x80;
assign n_907 = n_895 ^ n_279;
assign n_908 = n_895 ^ n_346;
assign n_909 = n_897 ^ x81;
assign n_910 = ~n_877 & n_898;
assign n_911 = n_898 ^ n_877;
assign n_912 = n_899 ^ n_533;
assign n_913 = n_523 & ~n_900;
assign n_914 = n_902 ^ x98;
assign n_915 = n_903 ^ n_902;
assign n_916 = n_907 ^ n_346;
assign n_917 = n_348 & ~n_908;
assign n_918 = n_909 ^ n_893;
assign n_919 = n_909 ^ x80;
assign n_920 = n_555 ^ n_911;
assign n_921 = n_912 ^ n_911;
assign n_922 = n_912 ^ n_555;
assign n_923 = n_913 ^ n_143;
assign n_924 = n_915 & ~n_914;
assign n_925 = n_915 ^ x98;
assign n_926 = n_279 & ~n_916;
assign n_927 = n_594 ^ n_916;
assign n_928 = n_917 ^ n_279;
assign n_929 = n_906 & ~n_918;
assign n_930 = n_919 ^ n_893;
assign n_931 = n_920 & ~n_921;
assign n_932 = n_922 ^ n_911;
assign n_933 = n_901 & ~n_923;
assign n_934 = n_923 ^ n_901;
assign n_935 = n_924 ^ x98;
assign n_936 = n_925 & ~n_904;
assign n_937 = n_904 ^ n_925;
assign n_938 = n_926 ^ n_894;
assign n_939 = ~n_894 & ~n_926;
assign n_940 = n_928 ^ n_353;
assign n_941 = n_929 ^ x80;
assign n_942 = n_910 & n_930;
assign n_943 = n_930 ^ n_910;
assign n_944 = n_931 ^ n_555;
assign n_945 = ~n_545 & ~n_932;
assign n_946 = n_934 ^ x97;
assign n_947 = n_935 ^ n_934;
assign n_948 = n_938 ^ x95;
assign n_949 = n_285 & ~n_940;
assign n_950 = n_940 & ~n_355;
assign n_951 = n_940 ^ n_285;
assign n_952 = n_941 ^ n_938;
assign n_953 = n_577 ^ n_943;
assign n_954 = n_944 ^ n_943;
assign n_955 = n_944 ^ n_577;
assign n_956 = n_945 ^ n_149;
assign n_957 = n_947 & ~n_946;
assign n_958 = n_947 ^ x97;
assign n_959 = n_939 ^ n_949;
assign n_960 = ~n_949 & n_939;
assign n_961 = n_950 ^ n_285;
assign n_962 = n_611 ^ n_951;
assign n_963 = ~n_952 & n_948;
assign n_964 = n_952 ^ x95;
assign n_965 = ~n_953 & n_954;
assign n_966 = n_955 ^ n_943;
assign n_967 = ~n_933 & ~n_956;
assign n_968 = n_956 ^ n_933;
assign n_969 = n_957 ^ x97;
assign n_970 = n_936 & n_958;
assign n_971 = n_958 ^ n_936;
assign n_972 = n_959 ^ x94;
assign n_973 = n_961 ^ n_360;
assign n_974 = n_963 ^ x95;
assign n_975 = n_942 & n_964;
assign n_976 = n_964 ^ n_942;
assign n_977 = n_965 ^ n_577;
assign n_978 = n_568 & n_966;
assign n_979 = n_968 ^ x96;
assign n_980 = n_969 ^ n_968;
assign n_981 = n_293 & n_973;
assign n_982 = ~n_973 & n_362;
assign n_983 = n_973 ^ n_293;
assign n_984 = n_974 ^ n_959;
assign n_985 = n_976 ^ n_597;
assign n_986 = n_977 ^ n_976;
assign n_987 = n_977 ^ n_597;
assign n_988 = n_978 ^ n_161;
assign n_989 = n_980 & ~n_979;
assign n_990 = n_980 ^ x96;
assign n_991 = n_981 ^ n_960;
assign n_992 = n_960 & ~n_981;
assign n_993 = n_982 ^ n_293;
assign n_994 = n_983 ^ n_625;
assign n_995 = n_984 & ~n_972;
assign n_996 = n_984 ^ x94;
assign n_997 = n_985 & n_986;
assign n_998 = n_987 ^ n_976;
assign n_999 = n_967 & n_988;
assign n_1000 = n_988 ^ n_967;
assign n_1001 = n_989 ^ x96;
assign n_1002 = n_970 & n_990;
assign n_1003 = n_990 ^ n_970;
assign n_1004 = n_991 ^ x93;
assign n_1005 = n_993 ^ n_367;
assign n_1006 = n_995 ^ x94;
assign n_1007 = ~n_996 & n_975;
assign n_1008 = n_975 ^ n_996;
assign n_1009 = n_997 ^ n_597;
assign n_1010 = n_589 & ~n_998;
assign n_1011 = n_1000 ^ x111;
assign n_1012 = n_1001 ^ n_1000;
assign n_1013 = n_1005 & n_302;
assign n_1014 = ~n_1005 & n_369;
assign n_1015 = n_302 ^ n_1005;
assign n_1016 = n_1006 ^ n_991;
assign n_1017 = n_1008 ^ n_613;
assign n_1018 = n_1009 ^ n_1008;
assign n_1019 = n_1009 ^ n_613;
assign n_1020 = n_1010 ^ n_160;
assign n_1021 = n_1012 & ~n_1011;
assign n_1022 = n_1012 ^ x111;
assign n_1023 = n_992 ^ n_1013;
assign n_1024 = n_1013 & ~n_992;
assign n_1025 = n_1014 ^ n_302;
assign n_1026 = n_641 ^ n_1015;
assign n_1027 = n_1016 & ~n_1004;
assign n_1028 = n_1016 ^ x93;
assign n_1029 = n_1017 & n_1018;
assign n_1030 = n_1019 ^ n_1008;
assign n_1031 = n_999 & ~n_1020;
assign n_1032 = n_1020 ^ n_999;
assign n_1033 = n_1021 ^ x111;
assign n_1034 = ~n_1002 & ~n_1022;
assign n_1035 = n_1022 ^ n_1002;
assign n_1036 = n_1023 ^ x92;
assign n_1037 = n_1025 ^ n_309;
assign n_1038 = n_1025 ^ n_374;
assign n_1039 = n_1027 ^ x93;
assign n_1040 = n_1028 & ~n_1007;
assign n_1041 = n_1007 ^ n_1028;
assign n_1042 = n_1029 ^ n_613;
assign n_1043 = ~n_605 & n_1030;
assign n_1044 = n_1032 ^ x110;
assign n_1045 = n_1033 ^ n_1032;
assign n_1046 = n_1037 ^ n_374;
assign n_1047 = ~n_1038 & ~n_376;
assign n_1048 = n_1039 ^ n_1023;
assign n_1049 = n_628 ^ n_1041;
assign n_1050 = n_1042 ^ n_1041;
assign n_1051 = n_1042 ^ n_628;
assign n_1052 = n_1043 ^ n_166;
assign n_1053 = ~n_1045 & n_1044;
assign n_1054 = n_1045 ^ x110;
assign n_1055 = n_309 & n_1046;
assign n_1056 = n_656 ^ n_1046;
assign n_1057 = n_1047 ^ n_309;
assign n_1058 = ~n_1048 & n_1036;
assign n_1059 = n_1048 ^ x92;
assign n_1060 = n_1049 & n_1050;
assign n_1061 = n_1051 ^ n_1041;
assign n_1062 = n_1052 & ~n_1031;
assign n_1063 = n_1031 ^ n_1052;
assign n_1064 = n_1053 ^ x110;
assign n_1065 = ~n_1034 & ~n_1054;
assign n_1066 = n_1054 ^ n_1034;
assign n_1067 = n_1024 ^ n_1055;
assign n_1068 = ~n_1055 & n_1024;
assign n_1069 = n_1057 ^ n_381;
assign n_1070 = n_1058 ^ x92;
assign n_1071 = n_1059 & ~n_1040;
assign n_1072 = n_1040 ^ n_1059;
assign n_1073 = n_1060 ^ n_628;
assign n_1074 = ~n_620 & ~n_1061;
assign n_1075 = n_1063 ^ x109;
assign n_1076 = n_1064 ^ n_1063;
assign n_1077 = n_1067 ^ x91;
assign n_1078 = n_319 & n_1069;
assign n_1079 = ~n_1069 & ~n_384;
assign n_1080 = n_1069 ^ n_319;
assign n_1081 = n_1070 ^ n_1067;
assign n_1082 = n_644 ^ n_1072;
assign n_1083 = n_1073 ^ n_1072;
assign n_1084 = n_1073 ^ n_644;
assign n_1085 = n_1074 ^ n_198;
assign n_1086 = n_1076 & ~n_1075;
assign n_1087 = n_1076 ^ x109;
assign n_1088 = n_1078 ^ n_1068;
assign n_1089 = ~n_1068 & ~n_1078;
assign n_1090 = n_1079 ^ n_319;
assign n_1091 = n_1080 ^ n_670;
assign n_1092 = ~n_1081 & n_1077;
assign n_1093 = n_1081 ^ x91;
assign n_1094 = n_1082 & n_1083;
assign n_1095 = n_1084 ^ n_1072;
assign n_1096 = n_1085 & ~n_1062;
assign n_1097 = n_1062 ^ n_1085;
assign n_1098 = n_1086 ^ x109;
assign n_1099 = n_1087 & n_1065;
assign n_1100 = n_1065 ^ n_1087;
assign n_1101 = n_1088 ^ x90;
assign n_1102 = n_1090 ^ n_388;
assign n_1103 = n_1092 ^ x91;
assign n_1104 = n_1071 & n_1093;
assign n_1105 = n_1093 ^ n_1071;
assign n_1106 = n_1094 ^ n_644;
assign n_1107 = n_637 & n_1095;
assign n_1108 = n_1097 ^ x108;
assign n_1109 = n_1098 ^ n_1097;
assign n_1110 = n_721 & ~n_1100;
assign n_1111 = n_1100 ^ n_721;
assign n_1112 = n_328 & n_1102;
assign n_1113 = ~n_1102 & n_392;
assign n_1114 = n_1102 ^ n_328;
assign n_1115 = n_1103 ^ n_1088;
assign n_1116 = n_659 ^ n_1105;
assign n_1117 = n_1106 ^ n_1105;
assign n_1118 = n_1106 ^ n_659;
assign n_1119 = n_1107 ^ n_189;
assign n_1120 = ~n_1109 & n_1108;
assign n_1121 = n_1109 ^ x108;
assign n_1122 = n_1110 ^ n_737;
assign n_1123 = n_714 & ~n_1111;
assign n_1124 = n_1112 ^ n_1089;
assign n_1125 = n_1089 & ~n_1112;
assign n_1126 = n_1113 ^ n_328;
assign n_1127 = n_1114 ^ n_685;
assign n_1128 = ~n_1115 & n_1101;
assign n_1129 = n_1115 ^ x90;
assign n_1130 = ~n_1116 & n_1117;
assign n_1131 = n_1118 ^ n_1105;
assign n_1132 = ~n_1119 & ~n_1096;
assign n_1133 = n_1096 ^ n_1119;
assign n_1134 = n_1120 ^ x108;
assign n_1135 = ~n_1121 & n_1099;
assign n_1136 = n_1099 ^ n_1121;
assign n_1137 = n_1123 ^ n_405;
assign n_1138 = n_1124 ^ x89;
assign n_1139 = n_1126 ^ n_395;
assign n_1140 = n_1128 ^ x90;
assign n_1141 = ~n_1129 & ~n_1104;
assign n_1142 = n_1104 ^ n_1129;
assign n_1143 = n_1130 ^ n_659;
assign n_1144 = n_652 & n_1131;
assign n_1145 = n_1133 ^ x107;
assign n_1146 = n_1134 ^ n_1133;
assign n_1147 = n_1136 ^ n_1110;
assign n_1148 = n_1136 ^ n_1122;
assign n_1149 = ~n_93 & n_1137;
assign n_1150 = n_1137 ^ n_93;
assign n_1151 = n_336 & ~n_1139;
assign n_1152 = n_1139 ^ n_684;
assign n_1153 = n_1139 ^ n_336;
assign n_1154 = n_1140 ^ n_1124;
assign n_1155 = n_1142 ^ n_672;
assign n_1156 = n_1143 ^ n_1142;
assign n_1157 = n_1143 ^ n_672;
assign n_1158 = n_1144 ^ n_194;
assign n_1159 = ~n_1146 & n_1145;
assign n_1160 = n_1146 ^ x107;
assign n_1161 = n_1122 & ~n_1147;
assign n_1162 = n_736 & n_1148;
assign n_1163 = n_1149 ^ n_105;
assign n_1164 = x135 & ~n_1150;
assign n_1165 = n_1150 ^ x135;
assign n_1166 = n_1151 ^ n_1125;
assign n_1167 = n_1152 ^ n_695;
assign n_1168 = n_1154 & ~n_1138;
assign n_1169 = n_1154 ^ x89;
assign n_1170 = ~n_1155 & ~n_1156;
assign n_1171 = n_1157 ^ n_1142;
assign n_1172 = n_1158 & ~n_1132;
assign n_1173 = n_1132 ^ n_1158;
assign n_1174 = n_1159 ^ x107;
assign n_1175 = n_1160 & ~n_1135;
assign n_1176 = n_1135 ^ n_1160;
assign n_1177 = n_1161 ^ n_737;
assign n_1178 = n_1162 ^ n_418;
assign n_1179 = n_1164 ^ x134;
assign n_1180 = n_1168 ^ x89;
assign n_1181 = ~n_1141 & ~n_1169;
assign n_1182 = n_1169 ^ n_1141;
assign n_1183 = n_1170 ^ n_672;
assign n_1184 = n_1171 & n_676;
assign n_1185 = n_1173 ^ x106;
assign n_1186 = n_1174 ^ n_1173;
assign n_1187 = n_1177 ^ n_1176;
assign n_1188 = n_1177 ^ n_770;
assign n_1189 = n_1178 ^ n_1149;
assign n_1190 = n_1178 ^ n_1163;
assign n_1191 = n_1180 ^ n_1166;
assign n_1192 = n_688 ^ n_1182;
assign n_1193 = n_1182 ^ n_1183;
assign n_1194 = n_688 ^ n_1183;
assign n_1195 = n_1184 ^ n_203;
assign n_1196 = ~n_1186 & n_1185;
assign n_1197 = n_1186 ^ x106;
assign n_1198 = n_1187 ^ n_770;
assign n_1199 = n_1187 & n_1188;
assign n_1200 = n_1163 & ~n_1189;
assign n_1201 = n_1190 ^ n_1164;
assign n_1202 = n_1190 ^ n_1179;
assign n_1203 = n_1191 ^ x88;
assign n_1204 = ~n_1193 & ~n_1192;
assign n_1205 = n_1194 ^ n_1182;
assign n_1206 = n_1195 & ~n_1172;
assign n_1207 = n_1172 ^ n_1195;
assign n_1208 = n_1196 ^ x106;
assign n_1209 = n_1197 & n_1175;
assign n_1210 = n_1175 ^ n_1197;
assign n_1211 = ~n_769 & ~n_1198;
assign n_1212 = n_1199 ^ n_770;
assign n_1213 = n_1200 ^ n_105;
assign n_1214 = n_1179 & ~n_1201;
assign n_1215 = ~n_1202 & n_1165;
assign n_1216 = n_1165 ^ n_1202;
assign n_1217 = n_1203 ^ n_1181;
assign n_1218 = n_1204 ^ n_688;
assign n_1219 = n_680 & ~n_1205;
assign n_1220 = n_1207 ^ x105;
assign n_1221 = n_1208 ^ n_1207;
assign n_1222 = n_1210 ^ n_806;
assign n_1223 = n_1211 ^ n_441;
assign n_1224 = n_1212 ^ n_1210;
assign n_1225 = n_1212 ^ n_806;
assign n_1226 = n_1214 ^ x134;
assign n_1227 = n_1217 ^ n_697;
assign n_1228 = n_1218 ^ n_1217;
assign n_1229 = n_1218 ^ n_697;
assign n_1230 = n_1219 ^ n_210;
assign n_1231 = n_1208 ^ n_1220;
assign n_1232 = ~n_1220 & n_1221;
assign n_1233 = n_1213 ^ n_1223;
assign n_1234 = n_1223 ^ n_111;
assign n_1235 = n_1222 & ~n_1224;
assign n_1236 = n_1225 ^ n_1210;
assign n_1237 = ~n_1227 & n_1228;
assign n_1238 = n_1229 ^ n_1217;
assign n_1239 = ~n_1206 & n_1230;
assign n_1240 = n_1230 ^ n_1206;
assign n_1241 = n_1231 & ~n_1209;
assign n_1242 = n_1209 ^ n_1231;
assign n_1243 = n_1232 ^ x105;
assign n_1244 = n_1233 ^ n_111;
assign n_1245 = n_1233 & n_1234;
assign n_1246 = n_1235 ^ n_806;
assign n_1247 = ~n_796 & n_1236;
assign n_1248 = n_1237 ^ n_697;
assign n_1249 = n_1238 & ~n_703;
assign n_1250 = n_1240 ^ x104;
assign n_1251 = n_1242 ^ n_837;
assign n_1252 = n_1243 ^ n_1240;
assign n_1253 = n_1226 ^ n_1244;
assign n_1254 = n_1244 ^ x133;
assign n_1255 = n_1245 ^ n_111;
assign n_1256 = n_1246 ^ n_1242;
assign n_1257 = n_1246 ^ n_837;
assign n_1258 = n_1247 ^ n_462;
assign n_1259 = n_1248 ^ n_716;
assign n_1260 = n_1248 ^ n_413;
assign n_1261 = n_1249 ^ n_218;
assign n_1262 = ~n_1252 & n_1250;
assign n_1263 = n_1252 ^ x104;
assign n_1264 = n_1253 ^ x133;
assign n_1265 = ~n_1253 & n_1254;
assign n_1266 = n_1251 & ~n_1256;
assign n_1267 = n_1257 ^ n_1242;
assign n_1268 = n_1255 ^ n_1258;
assign n_1269 = n_1258 ^ n_118;
assign n_1270 = n_723 & ~n_1259;
assign n_1271 = n_1260 ^ n_716;
assign n_1272 = n_1239 & ~n_1261;
assign n_1273 = n_1261 ^ n_1239;
assign n_1274 = n_1262 ^ x104;
assign n_1275 = ~n_1263 & n_1241;
assign n_1276 = n_1241 ^ n_1263;
assign n_1277 = ~n_1264 & n_1215;
assign n_1278 = n_1215 ^ n_1264;
assign n_1279 = n_1265 ^ x133;
assign n_1280 = n_1266 ^ n_837;
assign n_1281 = ~n_825 & n_1267;
assign n_1282 = n_1268 ^ n_118;
assign n_1283 = ~n_1268 & ~n_1269;
assign n_1284 = n_1270 ^ n_413;
assign n_1285 = ~n_1271 & ~n_725;
assign n_1286 = n_1273 ^ x119;
assign n_1287 = n_1274 ^ n_1273;
assign n_1288 = n_1276 ^ n_870;
assign n_1289 = n_1280 ^ n_1276;
assign n_1290 = n_1280 ^ n_870;
assign n_1291 = n_1281 ^ n_487;
assign n_1292 = n_1279 ^ n_1282;
assign n_1293 = n_1282 ^ x132;
assign n_1294 = n_1283 ^ n_118;
assign n_1295 = n_1284 ^ n_741;
assign n_1296 = n_1285 ^ n_226;
assign n_1297 = n_1274 ^ n_1286;
assign n_1298 = n_1286 & ~n_1287;
assign n_1299 = n_1288 & ~n_1289;
assign n_1300 = n_1290 ^ n_1276;
assign n_1301 = n_1291 ^ n_126;
assign n_1302 = n_1292 ^ x132;
assign n_1303 = ~n_1292 & n_1293;
assign n_1304 = n_1294 ^ n_1291;
assign n_1305 = n_1295 & n_751;
assign n_1306 = n_443 ^ n_1295;
assign n_1307 = n_1296 & ~n_1272;
assign n_1308 = n_1272 ^ n_1296;
assign n_1309 = ~n_1297 & n_1275;
assign n_1310 = n_1275 ^ n_1297;
assign n_1311 = n_1298 ^ x119;
assign n_1312 = n_1299 ^ n_870;
assign n_1313 = ~n_858 & n_1300;
assign n_1314 = n_1277 & ~n_1302;
assign n_1315 = n_1302 ^ n_1277;
assign n_1316 = n_1303 ^ x132;
assign n_1317 = n_1304 & ~n_1301;
assign n_1318 = n_1304 ^ n_126;
assign n_1319 = n_1305 ^ n_443;
assign n_1320 = n_732 & ~n_1306;
assign n_1321 = n_1306 ^ n_741;
assign n_1322 = n_1308 ^ x118;
assign n_1323 = n_1310 ^ n_900;
assign n_1324 = n_1311 ^ n_1308;
assign n_1325 = n_1312 ^ n_1310;
assign n_1326 = n_1312 ^ n_900;
assign n_1327 = n_1313 ^ n_511;
assign n_1328 = n_1317 ^ n_126;
assign n_1329 = n_1316 ^ n_1318;
assign n_1330 = n_1318 ^ x131;
assign n_1331 = n_1319 ^ n_766;
assign n_1332 = n_1320 ^ n_232;
assign n_1333 = n_1324 & ~n_1322;
assign n_1334 = n_1324 ^ x118;
assign n_1335 = ~n_1323 & ~n_1325;
assign n_1336 = n_1326 ^ n_1310;
assign n_1337 = n_1327 ^ n_132;
assign n_1338 = n_1328 ^ n_1327;
assign n_1339 = n_1328 ^ n_132;
assign n_1340 = n_1329 ^ x131;
assign n_1341 = n_1329 & ~n_1330;
assign n_1342 = ~n_1331 & n_775;
assign n_1343 = n_480 ^ n_1331;
assign n_1344 = ~n_1307 & ~n_1332;
assign n_1345 = n_1332 ^ n_1307;
assign n_1346 = n_1333 ^ x118;
assign n_1347 = ~n_1334 & ~n_1309;
assign n_1348 = n_1309 ^ n_1334;
assign n_1349 = n_1335 ^ n_900;
assign n_1350 = n_888 & ~n_1336;
assign n_1351 = n_1337 & n_1338;
assign n_1352 = n_1339 ^ n_1327;
assign n_1353 = ~n_1340 & ~n_1314;
assign n_1354 = n_1314 ^ n_1340;
assign n_1355 = n_1341 ^ x131;
assign n_1356 = n_1342 ^ n_480;
assign n_1357 = n_1343 & n_776;
assign n_1358 = n_1343 ^ n_766;
assign n_1359 = n_1345 ^ x117;
assign n_1360 = n_1346 ^ n_1345;
assign n_1361 = n_1348 ^ n_932;
assign n_1362 = n_1349 ^ n_1348;
assign n_1363 = n_1350 ^ n_533;
assign n_1364 = n_1351 ^ n_132;
assign n_1365 = n_1352 ^ x130;
assign n_1366 = n_1355 ^ n_1352;
assign n_1367 = n_1356 ^ n_792;
assign n_1368 = n_1357 ^ n_240;
assign n_1369 = n_1360 & ~n_1359;
assign n_1370 = n_1360 ^ x117;
assign n_1371 = n_1362 & ~n_1361;
assign n_1372 = n_1362 ^ n_932;
assign n_1373 = n_1363 ^ n_1364;
assign n_1374 = n_1364 ^ n_143;
assign n_1375 = ~n_1366 & n_1365;
assign n_1376 = n_1366 ^ x130;
assign n_1377 = ~n_1367 & n_801;
assign n_1378 = n_506 ^ n_1367;
assign n_1379 = ~n_1368 & n_1344;
assign n_1380 = n_1344 ^ n_1368;
assign n_1381 = n_1369 ^ x117;
assign n_1382 = ~n_1347 & n_1370;
assign n_1383 = n_1370 ^ n_1347;
assign n_1384 = n_1371 ^ n_932;
assign n_1385 = n_921 & n_1372;
assign n_1386 = n_1165 ^ n_1372;
assign n_1387 = n_1373 ^ n_143;
assign n_1388 = ~n_1373 & n_1374;
assign n_1389 = n_1375 ^ x130;
assign n_1390 = ~n_1353 & ~n_1376;
assign n_1391 = n_1376 ^ n_1353;
assign n_1392 = n_1377 ^ n_506;
assign n_1393 = n_1378 & n_802;
assign n_1394 = n_1378 ^ n_792;
assign n_1395 = n_1380 ^ x116;
assign n_1396 = n_1381 ^ n_1380;
assign n_1397 = n_1383 ^ n_966;
assign n_1398 = n_1384 ^ n_1383;
assign n_1399 = n_1384 ^ n_966;
assign n_1400 = n_1385 ^ n_555;
assign n_1401 = n_1387 ^ x129;
assign n_1402 = n_1388 ^ n_143;
assign n_1403 = n_1389 ^ n_1387;
assign n_1404 = n_1392 ^ n_821;
assign n_1405 = n_1393 ^ n_249;
assign n_1406 = ~n_1396 & n_1395;
assign n_1407 = n_1396 ^ x116;
assign n_1408 = n_1397 & n_1398;
assign n_1409 = n_1399 ^ n_1383;
assign n_1410 = n_1400 ^ n_149;
assign n_1411 = n_1402 ^ n_1400;
assign n_1412 = n_1403 & ~n_1401;
assign n_1413 = n_1403 ^ x129;
assign n_1414 = ~n_1404 & n_833;
assign n_1415 = n_528 ^ n_1404;
assign n_1416 = n_1405 & ~n_1379;
assign n_1417 = n_1379 ^ n_1405;
assign n_1418 = n_1406 ^ x116;
assign n_1419 = ~n_1407 & n_1382;
assign n_1420 = n_1382 ^ n_1407;
assign n_1421 = n_1408 ^ n_966;
assign n_1422 = ~n_954 & ~n_1409;
assign n_1423 = n_1216 ^ n_1409;
assign n_1424 = ~n_1411 & ~n_1410;
assign n_1425 = n_1411 ^ n_149;
assign n_1426 = n_1412 ^ x129;
assign n_1427 = ~n_1390 & ~n_1413;
assign n_1428 = n_1413 ^ n_1390;
assign n_1429 = n_1414 ^ n_528;
assign n_1430 = ~n_809 & n_1415;
assign n_1431 = n_1415 ^ n_821;
assign n_1432 = n_1417 ^ x115;
assign n_1433 = n_1418 ^ n_1417;
assign n_1434 = n_1420 ^ n_998;
assign n_1435 = n_1421 ^ n_1420;
assign n_1436 = n_1421 ^ n_998;
assign n_1437 = n_1422 ^ n_577;
assign n_1438 = n_1424 ^ n_149;
assign n_1439 = n_1425 ^ x128;
assign n_1440 = n_1426 ^ n_1425;
assign n_1441 = n_1429 ^ n_854;
assign n_1442 = n_1430 ^ n_262;
assign n_1443 = n_1433 & ~n_1432;
assign n_1444 = n_1433 ^ x115;
assign n_1445 = ~n_1434 & ~n_1435;
assign n_1446 = n_1436 ^ n_1420;
assign n_1447 = n_1437 ^ n_161;
assign n_1448 = n_1438 ^ n_1437;
assign n_1449 = ~n_1440 & n_1439;
assign n_1450 = n_1440 ^ x128;
assign n_1451 = n_548 ^ n_1441;
assign n_1452 = n_1441 & n_866;
assign n_1453 = n_1416 & ~n_1442;
assign n_1454 = n_1442 ^ n_1416;
assign n_1455 = n_1443 ^ x115;
assign n_1456 = n_1419 & n_1444;
assign n_1457 = n_1444 ^ n_1419;
assign n_1458 = n_1445 ^ n_998;
assign n_1459 = ~n_986 & ~n_1446;
assign n_1460 = n_1278 ^ n_1446;
assign n_1461 = n_1448 & n_1447;
assign n_1462 = n_1448 ^ n_161;
assign n_1463 = n_1449 ^ x128;
assign n_1464 = ~n_1450 & ~n_1427;
assign n_1465 = n_1427 ^ n_1450;
assign n_1466 = ~n_841 & n_1451;
assign n_1467 = n_1451 ^ n_854;
assign n_1468 = n_747 ^ n_1451;
assign n_1469 = n_1452 ^ n_548;
assign n_1470 = n_1454 ^ x114;
assign n_1471 = n_1455 ^ n_1454;
assign n_1472 = n_1455 ^ x114;
assign n_1473 = n_1457 ^ n_1030;
assign n_1474 = n_1458 ^ n_1457;
assign n_1475 = n_1458 ^ n_1030;
assign n_1476 = n_1459 ^ n_597;
assign n_1477 = n_1461 ^ n_161;
assign n_1478 = n_1462 ^ x143;
assign n_1479 = n_1463 ^ n_1462;
assign n_1480 = n_1466 ^ n_264;
assign n_1481 = n_1469 ^ n_885;
assign n_1482 = ~n_1470 & n_1471;
assign n_1483 = n_1472 ^ n_1454;
assign n_1484 = ~n_1473 & ~n_1474;
assign n_1485 = n_1475 ^ n_1457;
assign n_1486 = n_1476 ^ n_160;
assign n_1487 = n_1477 ^ n_1476;
assign n_1488 = ~n_1479 & n_1478;
assign n_1489 = n_1479 ^ x143;
assign n_1490 = n_1480 ^ n_1453;
assign n_1491 = ~n_1453 & ~n_1480;
assign n_1492 = n_572 ^ n_1481;
assign n_1493 = n_1481 & ~n_896;
assign n_1494 = n_1482 ^ x114;
assign n_1495 = n_1456 & n_1483;
assign n_1496 = n_1483 ^ n_1456;
assign n_1497 = n_1484 ^ n_1030;
assign n_1498 = ~n_1018 & n_1485;
assign n_1499 = n_1315 ^ n_1485;
assign n_1500 = n_1487 & n_1486;
assign n_1501 = n_1487 ^ n_160;
assign n_1502 = n_1488 ^ x143;
assign n_1503 = ~n_1489 & n_1464;
assign n_1504 = n_1464 ^ n_1489;
assign n_1505 = n_1490 ^ x113;
assign n_1506 = ~n_874 & n_1492;
assign n_1507 = n_1492 ^ n_885;
assign n_1508 = n_772 ^ n_1492;
assign n_1509 = n_1493 ^ n_572;
assign n_1510 = n_1494 ^ n_1490;
assign n_1511 = n_1494 ^ x113;
assign n_1512 = n_1496 ^ n_1061;
assign n_1513 = n_1497 ^ n_1496;
assign n_1514 = n_1497 ^ n_1061;
assign n_1515 = n_1498 ^ n_613;
assign n_1516 = n_1500 ^ n_160;
assign n_1517 = n_1501 ^ x142;
assign n_1518 = n_1502 ^ n_1501;
assign n_1519 = n_1506 ^ n_272;
assign n_1520 = n_1509 ^ n_927;
assign n_1521 = n_1509 ^ n_916;
assign n_1522 = ~n_1505 & n_1510;
assign n_1523 = n_1511 ^ n_1490;
assign n_1524 = n_1513 & n_1512;
assign n_1525 = n_1514 ^ n_1496;
assign n_1526 = n_1515 ^ n_166;
assign n_1527 = n_1516 ^ n_1515;
assign n_1528 = n_1518 & ~n_1517;
assign n_1529 = n_1518 ^ x142;
assign n_1530 = n_1519 ^ n_1491;
assign n_1531 = n_1491 & n_1519;
assign n_1532 = n_908 & ~n_1520;
assign n_1533 = n_829 ^ n_1520;
assign n_1534 = n_1520 ^ n_916;
assign n_1535 = n_927 & ~n_1521;
assign n_1536 = n_1522 ^ x113;
assign n_1537 = ~n_1523 & ~n_1495;
assign n_1538 = n_1495 ^ n_1523;
assign n_1539 = n_1524 ^ n_1061;
assign n_1540 = ~n_1050 & n_1525;
assign n_1541 = n_1354 ^ n_1525;
assign n_1542 = n_1527 & ~n_1526;
assign n_1543 = n_1527 ^ n_166;
assign n_1544 = n_1528 ^ x142;
assign n_1545 = n_1503 & n_1529;
assign n_1546 = n_1529 ^ n_1503;
assign n_1547 = n_1530 ^ x112;
assign n_1548 = n_1532 ^ n_279;
assign n_1549 = n_1535 ^ n_594;
assign n_1550 = n_1536 ^ n_1530;
assign n_1551 = n_1538 ^ n_1095;
assign n_1552 = n_1539 ^ n_1538;
assign n_1553 = n_1539 ^ n_1095;
assign n_1554 = n_1540 ^ n_628;
assign n_1555 = n_1542 ^ n_166;
assign n_1556 = n_1543 ^ x141;
assign n_1557 = n_1544 ^ n_1543;
assign n_1558 = n_1548 ^ n_1531;
assign n_1559 = n_1531 & n_1548;
assign n_1560 = n_1549 ^ n_611;
assign n_1561 = n_1549 ^ n_951;
assign n_1562 = n_1550 & ~n_1547;
assign n_1563 = n_1550 ^ x112;
assign n_1564 = n_1551 & n_1552;
assign n_1565 = n_1553 ^ n_1538;
assign n_1566 = n_1554 ^ n_198;
assign n_1567 = n_1555 ^ n_1554;
assign n_1568 = n_1557 & ~n_1556;
assign n_1569 = n_1557 ^ x141;
assign n_1570 = n_1558 ^ x127;
assign n_1571 = n_1560 ^ n_951;
assign n_1572 = ~n_962 & n_1561;
assign n_1573 = n_1562 ^ x112;
assign n_1574 = n_1563 & ~n_1537;
assign n_1575 = n_1537 ^ n_1563;
assign n_1576 = n_1564 ^ n_1095;
assign n_1577 = ~n_1083 & ~n_1565;
assign n_1578 = n_1391 ^ n_1565;
assign n_1579 = ~n_1567 & ~n_1566;
assign n_1580 = n_1567 ^ n_198;
assign n_1581 = n_1568 ^ x141;
assign n_1582 = n_1569 & n_1545;
assign n_1583 = n_1545 ^ n_1569;
assign n_1584 = ~n_940 & n_1571;
assign n_1585 = n_862 ^ n_1571;
assign n_1586 = n_1572 ^ n_611;
assign n_1587 = n_1573 ^ n_1558;
assign n_1588 = n_1575 ^ n_1131;
assign n_1589 = n_1576 ^ n_1575;
assign n_1590 = n_1576 ^ n_1131;
assign n_1591 = n_1577 ^ n_644;
assign n_1592 = n_1579 ^ n_198;
assign n_1593 = n_1580 ^ x140;
assign n_1594 = n_1581 ^ n_1580;
assign n_1595 = n_1584 ^ n_285;
assign n_1596 = n_1586 ^ n_625;
assign n_1597 = n_983 ^ n_1586;
assign n_1598 = n_1587 & ~n_1570;
assign n_1599 = n_1587 ^ x127;
assign n_1600 = n_1588 & ~n_1589;
assign n_1601 = n_1590 ^ n_1575;
assign n_1602 = n_1591 ^ n_189;
assign n_1603 = n_1592 ^ n_1591;
assign n_1604 = n_1594 & ~n_1593;
assign n_1605 = n_1594 ^ x140;
assign n_1606 = n_1559 ^ n_1595;
assign n_1607 = n_1595 & n_1559;
assign n_1608 = n_983 ^ n_1596;
assign n_1609 = n_994 & ~n_1597;
assign n_1610 = n_1598 ^ x127;
assign n_1611 = n_1599 & n_1574;
assign n_1612 = n_1574 ^ n_1599;
assign n_1613 = n_1600 ^ n_1131;
assign n_1614 = ~n_1117 & n_1601;
assign n_1615 = n_1428 ^ n_1601;
assign n_1616 = ~n_1603 & n_1602;
assign n_1617 = n_1603 ^ n_189;
assign n_1618 = n_1604 ^ x140;
assign n_1619 = n_1582 & n_1605;
assign n_1620 = n_1605 ^ n_1582;
assign n_1621 = n_1606 ^ x126;
assign n_1622 = n_973 & ~n_1608;
assign n_1623 = n_905 ^ n_1608;
assign n_1624 = n_1609 ^ n_625;
assign n_1625 = n_1610 ^ n_1606;
assign n_1626 = n_1612 ^ n_1171;
assign n_1627 = n_1613 ^ n_1612;
assign n_1628 = n_1613 ^ n_1171;
assign n_1629 = n_1614 ^ n_659;
assign n_1630 = n_1616 ^ n_189;
assign n_1631 = n_1617 ^ x139;
assign n_1632 = n_1618 ^ n_1617;
assign n_1633 = n_1622 ^ n_293;
assign n_1634 = n_1624 ^ n_1015;
assign n_1635 = n_1625 & ~n_1621;
assign n_1636 = n_1625 ^ x126;
assign n_1637 = ~n_1626 & n_1627;
assign n_1638 = n_1628 ^ n_1612;
assign n_1639 = n_1629 ^ n_194;
assign n_1640 = n_1630 ^ n_1629;
assign n_1641 = n_1632 & ~n_1631;
assign n_1642 = n_1632 ^ x139;
assign n_1643 = n_1633 ^ n_1607;
assign n_1644 = n_1607 & n_1633;
assign n_1645 = n_641 ^ n_1634;
assign n_1646 = ~n_1634 & n_1026;
assign n_1647 = n_1635 ^ x126;
assign n_1648 = ~n_1636 & ~n_1611;
assign n_1649 = n_1611 ^ n_1636;
assign n_1650 = n_1637 ^ n_1171;
assign n_1651 = n_1156 & ~n_1638;
assign n_1652 = n_1465 ^ n_1638;
assign n_1653 = ~n_1640 & n_1639;
assign n_1654 = n_1640 ^ n_194;
assign n_1655 = n_1641 ^ x139;
assign n_1656 = ~n_1619 & ~n_1642;
assign n_1657 = n_1642 ^ n_1619;
assign n_1658 = n_1643 ^ x125;
assign n_1659 = n_1005 & ~n_1645;
assign n_1660 = n_1645 ^ n_1015;
assign n_1661 = n_937 ^ n_1645;
assign n_1662 = n_1646 ^ n_641;
assign n_1663 = n_1647 ^ n_1643;
assign n_1664 = n_1649 ^ n_1205;
assign n_1665 = n_1649 ^ n_1650;
assign n_1666 = n_1650 ^ n_1205;
assign n_1667 = n_1651 ^ n_672;
assign n_1668 = n_1653 ^ n_194;
assign n_1669 = n_1654 ^ x138;
assign n_1670 = n_1655 ^ n_1654;
assign n_1671 = n_1659 ^ n_302;
assign n_1672 = n_1662 ^ n_656;
assign n_1673 = n_1662 ^ n_1046;
assign n_1674 = n_1663 & ~n_1658;
assign n_1675 = n_1663 ^ x125;
assign n_1676 = ~n_1665 & ~n_1664;
assign n_1677 = n_1649 ^ n_1666;
assign n_1678 = n_1667 ^ n_203;
assign n_1679 = n_1668 ^ n_1667;
assign n_1680 = n_1668 ^ n_203;
assign n_1681 = n_1670 & ~n_1669;
assign n_1682 = n_1670 ^ x138;
assign n_1683 = n_1644 ^ n_1671;
assign n_1684 = n_1671 & n_1644;
assign n_1685 = n_1672 ^ n_1046;
assign n_1686 = ~n_1056 & n_1673;
assign n_1687 = n_1674 ^ x125;
assign n_1688 = n_1648 & ~n_1675;
assign n_1689 = n_1675 ^ n_1648;
assign n_1690 = n_1676 ^ n_1205;
assign n_1691 = n_1193 & ~n_1677;
assign n_1692 = n_1504 ^ n_1677;
assign n_1693 = n_1678 & n_1679;
assign n_1694 = n_1680 ^ n_1667;
assign n_1695 = n_1681 ^ x138;
assign n_1696 = n_1656 & ~n_1682;
assign n_1697 = n_1682 ^ n_1656;
assign n_1698 = n_1683 ^ x124;
assign n_1699 = n_1038 & n_1685;
assign n_1700 = n_971 ^ n_1685;
assign n_1701 = n_1686 ^ n_656;
assign n_1702 = n_1687 ^ n_1683;
assign n_1703 = n_1689 ^ n_1238;
assign n_1704 = n_1689 ^ n_1690;
assign n_1705 = n_1690 ^ n_1238;
assign n_1706 = n_1691 ^ n_688;
assign n_1707 = n_1693 ^ n_203;
assign n_1708 = n_1694 ^ x137;
assign n_1709 = n_1695 ^ n_1694;
assign n_1710 = n_1699 ^ n_309;
assign n_1711 = n_1701 ^ n_1080;
assign n_1712 = n_1702 & ~n_1698;
assign n_1713 = n_1702 ^ x124;
assign n_1714 = ~n_1703 & ~n_1704;
assign n_1715 = n_1689 ^ n_1705;
assign n_1716 = n_1706 ^ n_210;
assign n_1717 = n_1707 ^ n_1706;
assign n_1718 = n_1709 & ~n_1708;
assign n_1719 = n_1709 ^ x137;
assign n_1720 = n_1684 ^ n_1710;
assign n_1721 = n_1710 & ~n_1684;
assign n_1722 = n_1711 ^ n_670;
assign n_1723 = ~n_1711 & n_1091;
assign n_1724 = n_1712 ^ x124;
assign n_1725 = ~n_1713 & n_1688;
assign n_1726 = n_1688 ^ n_1713;
assign n_1727 = n_1714 ^ n_1238;
assign n_1728 = ~n_1228 & n_1715;
assign n_1729 = n_1546 ^ n_1715;
assign n_1730 = n_1717 & n_1716;
assign n_1731 = n_1717 ^ n_210;
assign n_1732 = n_1718 ^ x137;
assign n_1733 = n_1696 & ~n_1719;
assign n_1734 = n_1719 ^ n_1696;
assign n_1735 = n_1720 ^ x123;
assign n_1736 = n_1069 & ~n_1722;
assign n_1737 = n_1722 ^ n_1080;
assign n_1738 = n_1003 ^ n_1722;
assign n_1739 = n_1723 ^ n_670;
assign n_1740 = n_1724 ^ n_1720;
assign n_1741 = n_1726 ^ n_1271;
assign n_1742 = n_1727 ^ n_1726;
assign n_1743 = n_1728 ^ n_697;
assign n_1744 = n_1730 ^ n_210;
assign n_1745 = n_1731 ^ x136;
assign n_1746 = n_1732 ^ n_1731;
assign n_1747 = n_1736 ^ n_319;
assign n_1748 = n_1739 ^ n_1114;
assign n_1749 = n_1740 & ~n_1735;
assign n_1750 = n_1740 ^ x123;
assign n_1751 = n_1742 & n_1741;
assign n_1752 = n_1742 ^ n_1271;
assign n_1753 = n_1743 ^ n_218;
assign n_1754 = n_1743 ^ n_1744;
assign n_1755 = ~n_1746 & n_1745;
assign n_1756 = n_1746 ^ x136;
assign n_1757 = n_1721 ^ n_1747;
assign n_1758 = n_1747 & ~n_1721;
assign n_1759 = n_1748 ^ n_685;
assign n_1760 = ~n_1748 & ~n_1127;
assign n_1761 = n_1749 ^ x123;
assign n_1762 = ~n_1750 & n_1725;
assign n_1763 = n_1725 ^ n_1750;
assign n_1764 = n_1751 ^ n_1271;
assign n_1765 = n_1260 & n_1752;
assign n_1766 = n_1752 ^ n_1583;
assign n_1767 = ~n_1754 & ~n_1753;
assign n_1768 = n_1754 ^ n_218;
assign n_1769 = n_1755 ^ x136;
assign n_1770 = n_1733 & n_1756;
assign n_1771 = n_1756 ^ n_1733;
assign n_1772 = n_1757 ^ x122;
assign n_1773 = n_1102 & n_1759;
assign n_1774 = n_1759 ^ n_1114;
assign n_1775 = n_1035 ^ n_1759;
assign n_1776 = n_1760 ^ n_685;
assign n_1777 = n_1761 ^ n_1757;
assign n_1778 = n_1763 ^ n_1306;
assign n_1779 = n_1764 ^ n_1763;
assign n_1780 = n_1764 ^ n_1306;
assign n_1781 = n_1765 ^ n_716;
assign n_1782 = n_1767 ^ n_218;
assign n_1783 = n_1768 ^ x151;
assign n_1784 = n_1769 ^ n_1768;
assign n_1785 = n_1773 ^ n_328;
assign n_1786 = n_1776 ^ n_1167;
assign n_1787 = n_1777 ^ x122;
assign n_1788 = ~n_1777 & n_1772;
assign n_1789 = n_1778 & ~n_1779;
assign n_1790 = n_1780 ^ n_1763;
assign n_1791 = n_1781 ^ n_226;
assign n_1792 = n_1782 ^ n_1781;
assign n_1793 = n_1782 ^ n_226;
assign n_1794 = ~n_1784 & n_1783;
assign n_1795 = n_1784 ^ x151;
assign n_1796 = n_1785 ^ n_1758;
assign n_1797 = n_1758 & n_1785;
assign n_1798 = n_1786 & n_1153;
assign n_1799 = n_1066 ^ n_1786;
assign n_1800 = n_1786 ^ n_1139;
assign n_1801 = n_1787 ^ n_1762;
assign n_1802 = n_1762 & n_1787;
assign n_1803 = n_1788 ^ x122;
assign n_1804 = n_1789 ^ n_1306;
assign n_1805 = ~n_1790 & ~n_1321;
assign n_1806 = n_1620 ^ n_1790;
assign n_1807 = ~n_1791 & n_1792;
assign n_1808 = n_1793 ^ n_1781;
assign n_1809 = n_1794 ^ x151;
assign n_1810 = n_1795 & n_1770;
assign n_1811 = n_1770 ^ n_1795;
assign n_1812 = n_1796 ^ x121;
assign n_1813 = n_1798 ^ n_336;
assign n_1814 = n_1801 ^ n_1343;
assign n_1815 = n_1803 ^ n_1796;
assign n_1816 = n_1804 ^ n_1801;
assign n_1817 = n_1804 ^ n_1343;
assign n_1818 = n_1805 ^ n_741;
assign n_1819 = n_1807 ^ n_226;
assign n_1820 = n_1808 ^ x150;
assign n_1821 = n_1809 ^ n_1808;
assign n_1822 = n_1813 ^ n_1797;
assign n_1823 = n_1815 ^ x121;
assign n_1824 = n_1815 & ~n_1812;
assign n_1825 = n_1814 & n_1816;
assign n_1826 = n_1817 ^ n_1801;
assign n_1827 = n_1818 ^ n_232;
assign n_1828 = n_1819 ^ n_1818;
assign n_1829 = n_1821 & ~n_1820;
assign n_1830 = n_1821 ^ x150;
assign n_1831 = n_1802 ^ n_1823;
assign n_1832 = n_1823 & ~n_1802;
assign n_1833 = n_1824 ^ x121;
assign n_1834 = n_1825 ^ n_1343;
assign n_1835 = ~n_1826 & n_1358;
assign n_1836 = n_1657 ^ n_1826;
assign n_1837 = ~n_1828 & n_1827;
assign n_1838 = n_1828 ^ n_232;
assign n_1839 = n_1829 ^ x150;
assign n_1840 = ~n_1830 & n_1810;
assign n_1841 = n_1810 ^ n_1830;
assign n_1842 = n_1831 ^ n_1378;
assign n_1843 = n_1833 ^ n_1822;
assign n_1844 = n_1834 ^ n_1378;
assign n_1845 = n_1834 ^ n_1831;
assign n_1846 = n_1835 ^ n_766;
assign n_1847 = n_1837 ^ n_232;
assign n_1848 = n_1838 ^ x149;
assign n_1849 = n_1839 ^ n_1838;
assign n_1850 = n_1843 ^ x120;
assign n_1851 = n_1844 ^ n_1831;
assign n_1852 = ~n_1845 & n_1842;
assign n_1853 = n_1846 ^ n_240;
assign n_1854 = n_1847 ^ n_1846;
assign n_1855 = ~n_1849 & n_1848;
assign n_1856 = n_1849 ^ x149;
assign n_1857 = n_1850 ^ n_1832;
assign n_1858 = n_1851 & n_1394;
assign n_1859 = n_1697 ^ n_1851;
assign n_1860 = n_1852 ^ n_1378;
assign n_1861 = ~n_1854 & n_1853;
assign n_1862 = n_1854 ^ n_240;
assign n_1863 = n_1855 ^ x149;
assign n_1864 = ~n_1840 & ~n_1856;
assign n_1865 = n_1856 ^ n_1840;
assign n_1866 = n_1857 ^ n_1415;
assign n_1867 = n_1858 ^ n_792;
assign n_1868 = n_1860 ^ n_1415;
assign n_1869 = n_1860 ^ n_1857;
assign n_1870 = n_1861 ^ n_240;
assign n_1871 = n_1862 ^ x148;
assign n_1872 = n_1863 ^ n_1862;
assign n_1873 = n_1867 ^ n_249;
assign n_1874 = n_1868 ^ n_1857;
assign n_1875 = ~n_1866 & n_1869;
assign n_1876 = n_1870 ^ n_1867;
assign n_1877 = n_1870 ^ n_249;
assign n_1878 = ~n_1872 & n_1871;
assign n_1879 = n_1872 ^ x148;
assign n_1880 = ~n_1874 & n_1431;
assign n_1881 = n_1734 ^ n_1874;
assign n_1882 = n_1875 ^ n_1415;
assign n_1883 = n_1873 & ~n_1876;
assign n_1884 = n_1877 ^ n_1867;
assign n_1885 = n_1878 ^ x148;
assign n_1886 = n_1864 & ~n_1879;
assign n_1887 = n_1879 ^ n_1864;
assign n_1888 = n_1880 ^ n_821;
assign n_1889 = n_1882 ^ n_747;
assign n_1890 = n_1882 ^ n_1451;
assign n_1891 = n_1883 ^ n_249;
assign n_1892 = n_1884 ^ x147;
assign n_1893 = n_1885 ^ n_1884;
assign n_1894 = n_1888 ^ n_262;
assign n_1895 = n_1889 ^ n_1451;
assign n_1896 = n_1468 & ~n_1890;
assign n_1897 = n_1891 ^ n_1888;
assign n_1898 = ~n_1893 & n_1892;
assign n_1899 = n_1893 ^ x147;
assign n_1900 = n_1895 & ~n_1467;
assign n_1901 = n_1771 ^ n_1895;
assign n_1902 = n_1896 ^ n_747;
assign n_1903 = n_1897 ^ n_262;
assign n_1904 = ~n_1897 & ~n_1894;
assign n_1905 = n_1898 ^ x147;
assign n_1906 = n_1886 & ~n_1899;
assign n_1907 = n_1899 ^ n_1886;
assign n_1908 = n_1900 ^ n_854;
assign n_1909 = n_1902 ^ n_1492;
assign n_1910 = n_1903 ^ x146;
assign n_1911 = n_1904 ^ n_262;
assign n_1912 = n_1905 ^ n_1903;
assign n_1913 = n_1905 ^ x146;
assign n_1914 = n_1908 ^ n_264;
assign n_1915 = n_1909 ^ n_772;
assign n_1916 = ~n_1909 & n_1508;
assign n_1917 = n_1911 ^ n_1908;
assign n_1918 = ~n_1910 & n_1912;
assign n_1919 = n_1913 ^ n_1903;
assign n_1920 = n_1915 & n_1507;
assign n_1921 = n_1915 ^ n_1492;
assign n_1922 = n_1915 ^ n_1811;
assign n_1923 = n_1916 ^ n_772;
assign n_1924 = n_1917 ^ n_264;
assign n_1925 = ~n_1917 & ~n_1914;
assign n_1926 = n_1918 ^ x146;
assign n_1927 = n_1906 & n_1919;
assign n_1928 = n_1919 ^ n_1906;
assign n_1929 = n_1920 ^ n_885;
assign n_1930 = n_1923 ^ n_1533;
assign n_1931 = n_1923 ^ n_1520;
assign n_1932 = n_1924 ^ x145;
assign n_1933 = n_1925 ^ n_264;
assign n_1934 = n_1926 ^ n_1924;
assign n_1935 = n_1930 & n_1534;
assign n_1936 = n_1930 ^ n_1520;
assign n_1937 = n_1841 ^ n_1930;
assign n_1938 = n_1533 & n_1931;
assign n_1939 = n_1929 ^ n_1933;
assign n_1940 = n_1933 ^ n_272;
assign n_1941 = ~n_1934 & n_1932;
assign n_1942 = n_1934 ^ x145;
assign n_1943 = n_1935 ^ n_916;
assign n_1944 = n_1938 ^ n_829;
assign n_1945 = n_1939 ^ n_272;
assign n_1946 = ~n_1939 & ~n_1940;
assign n_1947 = n_1941 ^ x145;
assign n_1948 = n_1927 & ~n_1942;
assign n_1949 = n_1942 ^ n_1927;
assign n_1950 = n_1943 ^ n_279;
assign n_1951 = n_1944 ^ n_862;
assign n_1952 = n_1944 ^ n_1571;
assign n_1953 = n_1945 ^ x144;
assign n_1954 = n_1946 ^ n_272;
assign n_1955 = n_1947 ^ n_1945;
assign n_1956 = n_1951 ^ n_1571;
assign n_1957 = ~n_1585 & n_1952;
assign n_1958 = n_1943 ^ n_1954;
assign n_1959 = n_1955 & ~n_1953;
assign n_1960 = n_1955 ^ x144;
assign n_1961 = n_1560 & n_1956;
assign n_1962 = n_1865 ^ n_1956;
assign n_1963 = n_1957 ^ n_862;
assign n_1964 = n_1958 ^ n_279;
assign n_1965 = ~n_1958 & n_1950;
assign n_1966 = n_1959 ^ x144;
assign n_1967 = ~n_1948 & ~n_1960;
assign n_1968 = n_1960 ^ n_1948;
assign n_1969 = n_1961 ^ n_951;
assign n_1970 = n_1963 ^ n_1608;
assign n_1971 = n_1964 ^ x159;
assign n_1972 = n_1965 ^ n_279;
assign n_1973 = n_1966 ^ n_1964;
assign n_1974 = n_1969 ^ n_285;
assign n_1975 = n_905 ^ n_1970;
assign n_1976 = ~n_1970 & ~n_1623;
assign n_1977 = n_1972 ^ n_1969;
assign n_1978 = n_1973 & ~n_1971;
assign n_1979 = n_1973 ^ x159;
assign n_1980 = n_1596 & n_1975;
assign n_1981 = n_1975 ^ n_1608;
assign n_1982 = n_1887 ^ n_1975;
assign n_1983 = n_1976 ^ n_905;
assign n_1984 = n_1977 ^ n_285;
assign n_1985 = n_1977 & ~n_1974;
assign n_1986 = n_1978 ^ x159;
assign n_1987 = n_1979 & ~n_1967;
assign n_1988 = n_1967 ^ n_1979;
assign n_1989 = n_1980 ^ n_983;
assign n_1990 = n_1983 ^ n_1645;
assign n_1991 = n_1984 ^ x158;
assign n_1992 = n_1985 ^ n_285;
assign n_1993 = n_1986 ^ n_1984;
assign n_1994 = n_1989 ^ n_293;
assign n_1995 = n_937 ^ n_1990;
assign n_1996 = n_1990 & ~n_1661;
assign n_1997 = n_1992 ^ n_1989;
assign n_1998 = n_1993 ^ x158;
assign n_1999 = ~n_1993 & n_1991;
assign n_2000 = ~n_1995 & n_1660;
assign n_2001 = n_1995 ^ n_1645;
assign n_2002 = n_1907 ^ n_1995;
assign n_2003 = n_1996 ^ n_937;
assign n_2004 = n_1997 ^ n_293;
assign n_2005 = ~n_1997 & n_1994;
assign n_2006 = n_1998 ^ n_1987;
assign n_2007 = ~n_1987 & n_1998;
assign n_2008 = n_1999 ^ x158;
assign n_2009 = n_2000 ^ n_1015;
assign n_2010 = n_2003 ^ n_1685;
assign n_2011 = n_2004 ^ x157;
assign n_2012 = n_2005 ^ n_293;
assign n_2013 = ~n_1111 & ~n_2006;
assign n_2014 = n_2006 ^ n_1111;
assign n_2015 = n_2008 ^ n_2004;
assign n_2016 = n_2009 ^ n_302;
assign n_2017 = n_971 ^ n_2010;
assign n_2018 = ~n_2010 & ~n_1700;
assign n_2019 = n_2012 ^ n_2009;
assign n_2020 = n_2013 ^ n_1148;
assign n_2021 = ~n_1100 & n_2014;
assign n_2022 = n_2015 & ~n_2011;
assign n_2023 = n_2015 ^ x157;
assign n_2024 = n_1672 & ~n_2017;
assign n_2025 = n_2017 ^ n_1685;
assign n_2026 = n_1928 ^ n_2017;
assign n_2027 = n_2018 ^ n_971;
assign n_2028 = n_2019 ^ n_302;
assign n_2029 = ~n_2019 & n_2016;
assign n_2030 = n_2021 ^ n_721;
assign n_2031 = n_2022 ^ x157;
assign n_2032 = n_2023 & ~n_2007;
assign n_2033 = n_2007 ^ n_2023;
assign n_2034 = n_2024 ^ n_1046;
assign n_2035 = n_2027 ^ n_1722;
assign n_2036 = n_2028 ^ x156;
assign n_2037 = n_2029 ^ n_302;
assign n_2038 = n_405 & n_2030;
assign n_2039 = n_2030 ^ n_405;
assign n_2040 = n_2031 ^ n_2028;
assign n_2041 = n_2033 ^ n_2013;
assign n_2042 = n_2033 ^ n_2020;
assign n_2043 = n_2034 ^ n_309;
assign n_2044 = n_1003 ^ n_2035;
assign n_2045 = ~n_2035 & n_1738;
assign n_2046 = n_2037 ^ n_2034;
assign n_2047 = n_2038 ^ n_418;
assign n_2048 = x167 & n_2039;
assign n_2049 = n_2039 ^ x167;
assign n_2050 = n_2040 & ~n_2036;
assign n_2051 = n_2040 ^ x156;
assign n_2052 = n_2020 & ~n_2041;
assign n_2053 = n_1147 & n_2042;
assign n_2054 = ~n_2044 & n_1737;
assign n_2055 = n_2044 ^ n_1722;
assign n_2056 = n_1949 ^ n_2044;
assign n_2057 = n_2045 ^ n_1003;
assign n_2058 = n_2046 ^ n_309;
assign n_2059 = n_2046 & n_2043;
assign n_2060 = n_2048 ^ x166;
assign n_2061 = n_2050 ^ x156;
assign n_2062 = ~n_2032 & ~n_2051;
assign n_2063 = n_2051 ^ n_2032;
assign n_2064 = n_2052 ^ n_1148;
assign n_2065 = n_2053 ^ n_737;
assign n_2066 = n_2054 ^ n_1080;
assign n_2067 = n_2057 ^ n_1759;
assign n_2068 = n_2058 ^ x155;
assign n_2069 = n_2059 ^ n_309;
assign n_2070 = n_2061 ^ n_2058;
assign n_2071 = n_2063 ^ n_1198;
assign n_2072 = n_2064 ^ n_2063;
assign n_2073 = n_2064 ^ n_1198;
assign n_2074 = n_2065 ^ n_2038;
assign n_2075 = n_2065 ^ n_2047;
assign n_2076 = n_2066 ^ n_319;
assign n_2077 = n_1035 ^ n_2067;
assign n_2078 = n_2067 & n_1775;
assign n_2079 = n_2069 ^ n_2066;
assign n_2080 = n_2070 & ~n_2068;
assign n_2081 = n_2070 ^ x155;
assign n_2082 = ~n_2071 & ~n_2072;
assign n_2083 = n_2073 ^ n_2063;
assign n_2084 = n_2047 & ~n_2074;
assign n_2085 = n_2075 ^ n_2048;
assign n_2086 = n_2075 ^ n_2060;
assign n_2087 = ~n_2077 & ~n_1774;
assign n_2088 = n_2077 ^ n_1759;
assign n_2089 = n_1968 ^ n_2077;
assign n_2090 = n_2078 ^ n_1035;
assign n_2091 = n_2079 ^ n_319;
assign n_2092 = n_2079 & n_2076;
assign n_2093 = n_2080 ^ x155;
assign n_2094 = ~n_2062 & n_2081;
assign n_2095 = n_2081 ^ n_2062;
assign n_2096 = n_2082 ^ n_1198;
assign n_2097 = ~n_1187 & ~n_2083;
assign n_2098 = n_2084 ^ n_418;
assign n_2099 = n_2060 & ~n_2085;
assign n_2100 = n_2087 ^ n_1114;
assign n_2101 = n_2090 ^ n_1799;
assign n_2102 = n_2091 ^ x154;
assign n_2103 = n_2092 ^ n_319;
assign n_2104 = n_2093 ^ n_2091;
assign n_2105 = n_2095 ^ n_1236;
assign n_2106 = n_2095 ^ n_2096;
assign n_2107 = n_2096 ^ n_1236;
assign n_2108 = n_2097 ^ n_770;
assign n_2109 = n_2098 ^ n_441;
assign n_2110 = n_2099 ^ x166;
assign n_2111 = n_2100 ^ n_328;
assign n_2112 = ~n_2101 & ~n_1800;
assign n_2113 = n_1988 ^ n_2101;
assign n_2114 = n_2101 ^ n_1786;
assign n_2115 = n_2103 ^ n_2100;
assign n_2116 = ~n_2104 & n_2102;
assign n_2117 = n_2104 ^ x154;
assign n_2118 = n_2106 & n_2105;
assign n_2119 = n_2107 ^ n_2095;
assign n_2120 = n_2108 ^ n_441;
assign n_2121 = n_2098 ^ n_2108;
assign n_2122 = n_2109 ^ n_2108;
assign n_2123 = n_2112 ^ n_1139;
assign n_2124 = n_2115 ^ n_328;
assign n_2125 = ~n_2115 & n_2111;
assign n_2126 = n_2116 ^ x154;
assign n_2127 = n_2094 & ~n_2117;
assign n_2128 = n_2117 ^ n_2094;
assign n_2129 = n_2118 ^ n_1236;
assign n_2130 = n_1224 & ~n_2119;
assign n_2131 = ~n_2120 & ~n_2121;
assign n_2132 = n_2110 ^ n_2122;
assign n_2133 = n_2122 ^ x165;
assign n_2134 = n_2123 ^ n_336;
assign n_2135 = n_2124 ^ x153;
assign n_2136 = n_2125 ^ n_328;
assign n_2137 = n_2126 ^ n_2124;
assign n_2138 = n_2128 ^ n_1267;
assign n_2139 = n_2129 ^ n_2128;
assign n_2140 = n_2129 ^ n_1267;
assign n_2141 = n_2130 ^ n_806;
assign n_2142 = n_2131 ^ n_441;
assign n_2143 = n_2132 ^ x165;
assign n_2144 = n_2132 & ~n_2133;
assign n_2145 = n_2136 ^ x152;
assign n_2146 = n_2137 & ~n_2135;
assign n_2147 = n_2137 ^ x153;
assign n_2148 = n_2138 & ~n_2139;
assign n_2149 = n_2140 ^ n_2128;
assign n_2150 = n_2141 ^ n_462;
assign n_2151 = n_2142 ^ n_2141;
assign n_2152 = n_2142 ^ n_462;
assign n_2153 = ~n_2143 & n_2086;
assign n_2154 = n_2086 ^ n_2143;
assign n_2155 = n_2144 ^ x165;
assign n_2156 = n_2145 ^ n_2134;
assign n_2157 = n_2146 ^ x153;
assign n_2158 = n_2127 & n_2147;
assign n_2159 = n_2147 ^ n_2127;
assign n_2160 = n_2148 ^ n_1267;
assign n_2161 = n_1256 & n_2149;
assign n_2162 = ~n_2150 & n_2151;
assign n_2163 = n_2152 ^ n_2141;
assign n_2164 = n_2157 ^ n_2156;
assign n_2165 = n_2159 ^ n_1300;
assign n_2166 = n_2160 ^ n_2159;
assign n_2167 = n_2160 ^ n_1300;
assign n_2168 = n_2161 ^ n_837;
assign n_2169 = n_2162 ^ n_462;
assign n_2170 = n_2155 ^ n_2163;
assign n_2171 = n_2163 ^ x164;
assign n_2172 = n_2164 ^ n_2158;
assign n_2173 = ~n_2165 & n_2166;
assign n_2174 = n_2167 ^ n_2159;
assign n_2175 = n_2168 ^ n_487;
assign n_2176 = n_2169 ^ n_2168;
assign n_2177 = n_2169 ^ n_487;
assign n_2178 = n_2170 ^ x164;
assign n_2179 = ~n_2170 & n_2171;
assign n_2180 = n_2172 ^ n_1336;
assign n_2181 = n_2173 ^ n_1300;
assign n_2182 = n_1289 & ~n_2174;
assign n_2183 = ~n_2175 & n_2176;
assign n_2184 = n_2177 ^ n_2168;
assign n_2185 = ~n_2153 & ~n_2178;
assign n_2186 = n_2178 ^ n_2153;
assign n_2187 = n_2179 ^ x164;
assign n_2188 = n_2181 ^ n_2172;
assign n_2189 = n_2181 ^ n_1336;
assign n_2190 = n_2182 ^ n_870;
assign n_2191 = n_2183 ^ n_487;
assign n_2192 = n_2184 ^ x163;
assign n_2193 = n_2187 ^ n_2184;
assign n_2194 = n_2180 & n_2188;
assign n_2195 = n_2189 ^ n_2172;
assign n_2196 = n_2190 ^ n_511;
assign n_2197 = n_2191 ^ n_2190;
assign n_2198 = n_2191 ^ n_511;
assign n_2199 = ~n_2193 & n_2192;
assign n_2200 = n_2193 ^ x163;
assign n_2201 = n_2194 ^ n_1336;
assign n_2202 = n_1325 & n_2195;
assign n_2203 = ~n_2196 & n_2197;
assign n_2204 = n_2198 ^ n_2190;
assign n_2205 = n_2199 ^ x163;
assign n_2206 = ~n_2185 & n_2200;
assign n_2207 = n_2200 ^ n_2185;
assign n_2208 = n_2201 ^ n_1165;
assign n_2209 = n_2201 ^ n_1386;
assign n_2210 = n_2202 ^ n_900;
assign n_2211 = n_2203 ^ n_511;
assign n_2212 = n_2204 ^ x162;
assign n_2213 = n_2205 ^ n_2204;
assign n_2214 = n_1386 & n_2208;
assign n_2215 = ~n_1362 & ~n_2209;
assign n_2216 = n_2210 ^ n_533;
assign n_2217 = n_2211 ^ n_2210;
assign n_2218 = n_2211 ^ n_533;
assign n_2219 = ~n_2213 & n_2212;
assign n_2220 = n_2213 ^ x162;
assign n_2221 = n_2214 ^ n_1372;
assign n_2222 = n_2215 ^ n_932;
assign n_2223 = n_2216 & ~n_2217;
assign n_2224 = n_2218 ^ n_2210;
assign n_2225 = n_2219 ^ x162;
assign n_2226 = ~n_2206 & ~n_2220;
assign n_2227 = n_2220 ^ n_2206;
assign n_2228 = n_2221 ^ n_1409;
assign n_2229 = n_2223 ^ n_533;
assign n_2230 = n_2224 ^ x161;
assign n_2231 = n_2225 ^ n_2224;
assign n_2232 = n_2228 & ~n_1423;
assign n_2233 = n_1216 ^ n_2228;
assign n_2234 = n_2229 ^ n_555;
assign n_2235 = n_2222 ^ n_2229;
assign n_2236 = n_2231 & ~n_2230;
assign n_2237 = n_2231 ^ x161;
assign n_2238 = n_2232 ^ n_1216;
assign n_2239 = ~n_1398 & ~n_2233;
assign n_2240 = n_2233 ^ n_1409;
assign n_2241 = n_2222 ^ n_2234;
assign n_2242 = n_2234 & ~n_2235;
assign n_2243 = n_2236 ^ x161;
assign n_2244 = ~n_2226 & ~n_2237;
assign n_2245 = n_2237 ^ n_2226;
assign n_2246 = n_2238 ^ n_1446;
assign n_2247 = n_2239 ^ n_966;
assign n_2248 = n_2241 ^ x160;
assign n_2249 = n_2242 ^ n_555;
assign n_2250 = n_2243 ^ n_2241;
assign n_2251 = n_2246 & ~n_1460;
assign n_2252 = n_1278 ^ n_2246;
assign n_2253 = n_2247 ^ n_577;
assign n_2254 = n_2249 ^ n_2247;
assign n_2255 = n_2249 ^ n_577;
assign n_2256 = n_2250 & ~n_2248;
assign n_2257 = n_2250 ^ x160;
assign n_2258 = n_2251 ^ n_1278;
assign n_2259 = n_1435 & ~n_2252;
assign n_2260 = n_2252 ^ n_1446;
assign n_2261 = ~n_2253 & n_2254;
assign n_2262 = n_2255 ^ n_2247;
assign n_2263 = n_2256 ^ x160;
assign n_2264 = n_2244 & ~n_2257;
assign n_2265 = n_2257 ^ n_2244;
assign n_2266 = n_2258 ^ n_1485;
assign n_2267 = n_2259 ^ n_998;
assign n_2268 = n_2261 ^ n_577;
assign n_2269 = n_2262 ^ x175;
assign n_2270 = n_2263 ^ n_2262;
assign n_2271 = ~n_2266 & n_1499;
assign n_2272 = n_1315 ^ n_2266;
assign n_2273 = n_2267 ^ n_597;
assign n_2274 = n_2268 ^ n_2267;
assign n_2275 = n_2268 ^ n_597;
assign n_2276 = ~n_2270 & n_2269;
assign n_2277 = n_2270 ^ x175;
assign n_2278 = n_2271 ^ n_1315;
assign n_2279 = n_1474 & n_2272;
assign n_2280 = n_2272 ^ n_1485;
assign n_2281 = ~n_2273 & ~n_2274;
assign n_2282 = n_2275 ^ n_2267;
assign n_2283 = n_2276 ^ x175;
assign n_2284 = n_2264 & n_2277;
assign n_2285 = n_2277 ^ n_2264;
assign n_2286 = n_2278 ^ n_1525;
assign n_2287 = n_2279 ^ n_1030;
assign n_2288 = n_2281 ^ n_597;
assign n_2289 = n_2282 ^ x174;
assign n_2290 = n_2283 ^ n_2282;
assign n_2291 = n_1354 ^ n_2286;
assign n_2292 = ~n_2286 & n_1541;
assign n_2293 = n_2287 ^ n_613;
assign n_2294 = n_2288 ^ n_2287;
assign n_2295 = n_2288 ^ n_613;
assign n_2296 = ~n_2290 & n_2289;
assign n_2297 = n_2290 ^ x174;
assign n_2298 = ~n_1513 & n_2291;
assign n_2299 = n_2291 ^ n_1525;
assign n_2300 = n_2292 ^ n_1354;
assign n_2301 = ~n_2293 & ~n_2294;
assign n_2302 = n_2295 ^ n_2287;
assign n_2303 = n_2296 ^ x174;
assign n_2304 = ~n_2297 & ~n_2284;
assign n_2305 = n_2284 ^ n_2297;
assign n_2306 = n_2298 ^ n_1061;
assign n_2307 = n_2300 ^ n_1565;
assign n_2308 = n_2301 ^ n_613;
assign n_2309 = n_2302 ^ x173;
assign n_2310 = n_2303 ^ n_2302;
assign n_2311 = n_2306 ^ n_628;
assign n_2312 = n_1391 ^ n_2307;
assign n_2313 = n_2307 & n_1578;
assign n_2314 = n_2308 ^ n_2306;
assign n_2315 = n_2308 ^ n_628;
assign n_2316 = n_2310 & ~n_2309;
assign n_2317 = n_2310 ^ x173;
assign n_2318 = ~n_1552 & n_2312;
assign n_2319 = n_2312 ^ n_1565;
assign n_2320 = n_2049 ^ n_2312;
assign n_2321 = n_2313 ^ n_1391;
assign n_2322 = ~n_2311 & ~n_2314;
assign n_2323 = n_2315 ^ n_2306;
assign n_2324 = n_2316 ^ x173;
assign n_2325 = n_2304 & n_2317;
assign n_2326 = n_2317 ^ n_2304;
assign n_2327 = n_2318 ^ n_1095;
assign n_2328 = n_2321 ^ n_1601;
assign n_2329 = n_2322 ^ n_628;
assign n_2330 = n_2323 ^ x172;
assign n_2331 = n_2324 ^ n_2323;
assign n_2332 = n_2327 ^ n_644;
assign n_2333 = n_1428 ^ n_2328;
assign n_2334 = n_2328 & n_1615;
assign n_2335 = n_2329 ^ n_644;
assign n_2336 = n_2329 ^ n_2327;
assign n_2337 = ~n_2331 & n_2330;
assign n_2338 = n_2331 ^ x172;
assign n_2339 = n_1589 & ~n_2333;
assign n_2340 = n_2333 ^ n_1601;
assign n_2341 = n_2086 ^ n_2333;
assign n_2342 = n_2334 ^ n_1428;
assign n_2343 = n_2335 ^ n_2327;
assign n_2344 = ~n_2332 & ~n_2336;
assign n_2345 = n_2337 ^ x172;
assign n_2346 = ~n_2325 & n_2338;
assign n_2347 = n_2338 ^ n_2325;
assign n_2348 = n_2339 ^ n_1131;
assign n_2349 = n_2342 ^ n_1638;
assign n_2350 = n_2343 ^ x171;
assign n_2351 = n_2344 ^ n_644;
assign n_2352 = n_2345 ^ n_2343;
assign n_2353 = n_2345 ^ x171;
assign n_2354 = n_2348 ^ n_659;
assign n_2355 = n_1465 ^ n_2349;
assign n_2356 = n_2349 & n_1652;
assign n_2357 = n_2351 ^ n_659;
assign n_2358 = n_2351 ^ n_2348;
assign n_2359 = ~n_2350 & n_2352;
assign n_2360 = n_2353 ^ n_2343;
assign n_2361 = ~n_1627 & n_2355;
assign n_2362 = n_2355 ^ n_1638;
assign n_2363 = n_2154 ^ n_2355;
assign n_2364 = n_2356 ^ n_1465;
assign n_2365 = n_2357 ^ n_2348;
assign n_2366 = ~n_2354 & n_2358;
assign n_2367 = n_2359 ^ x171;
assign n_2368 = n_2346 & ~n_2360;
assign n_2369 = n_2360 ^ n_2346;
assign n_2370 = n_2361 ^ n_1171;
assign n_2371 = n_2364 ^ n_1677;
assign n_2372 = n_2365 ^ x170;
assign n_2373 = n_2366 ^ n_659;
assign n_2374 = n_2367 ^ n_2365;
assign n_2375 = n_2370 ^ n_672;
assign n_2376 = n_1504 ^ n_2371;
assign n_2377 = ~n_2371 & ~n_1692;
assign n_2378 = n_2373 ^ n_672;
assign n_2379 = n_2373 ^ n_2370;
assign n_2380 = ~n_2374 & n_2372;
assign n_2381 = n_2374 ^ x170;
assign n_2382 = n_1665 & n_2376;
assign n_2383 = n_2376 ^ n_1677;
assign n_2384 = n_2186 ^ n_2376;
assign n_2385 = n_2377 ^ n_1504;
assign n_2386 = n_2378 ^ n_2370;
assign n_2387 = n_2375 & n_2379;
assign n_2388 = n_2380 ^ x170;
assign n_2389 = n_2368 & n_2381;
assign n_2390 = n_2381 ^ n_2368;
assign n_2391 = n_2382 ^ n_1205;
assign n_2392 = n_2385 ^ n_1729;
assign n_2393 = n_2385 ^ n_1715;
assign n_2394 = n_2386 ^ x169;
assign n_2395 = n_2387 ^ n_672;
assign n_2396 = n_2388 ^ n_2386;
assign n_2397 = n_2391 ^ n_688;
assign n_2398 = n_1704 & ~n_2392;
assign n_2399 = n_2207 ^ n_2392;
assign n_2400 = n_2392 ^ n_1715;
assign n_2401 = ~n_1729 & ~n_2393;
assign n_2402 = n_2395 ^ n_688;
assign n_2403 = n_2395 ^ n_2391;
assign n_2404 = n_2396 & ~n_2394;
assign n_2405 = n_2396 ^ x169;
assign n_2406 = n_2398 ^ n_1238;
assign n_2407 = n_2401 ^ n_1546;
assign n_2408 = n_2402 ^ n_2391;
assign n_2409 = n_2397 & n_2403;
assign n_2410 = n_2404 ^ x169;
assign n_2411 = ~n_2389 & n_2405;
assign n_2412 = n_2405 ^ n_2389;
assign n_2413 = n_2406 ^ n_697;
assign n_2414 = n_2407 ^ n_1583;
assign n_2415 = n_2407 ^ n_1752;
assign n_2416 = n_2408 ^ x168;
assign n_2417 = n_2409 ^ n_688;
assign n_2418 = n_2410 ^ n_2408;
assign n_2419 = n_2414 ^ n_1752;
assign n_2420 = ~n_1766 & n_2415;
assign n_2421 = n_2417 ^ n_2406;
assign n_2422 = n_2418 ^ x168;
assign n_2423 = ~n_2418 & n_2416;
assign n_2424 = ~n_1742 & n_2419;
assign n_2425 = n_2227 ^ n_2419;
assign n_2426 = n_2420 ^ n_1583;
assign n_2427 = n_2421 ^ n_697;
assign n_2428 = n_2421 & ~n_2413;
assign n_2429 = ~n_2422 & n_2411;
assign n_2430 = n_2411 ^ n_2422;
assign n_2431 = n_2423 ^ x168;
assign n_2432 = n_2424 ^ n_1271;
assign n_2433 = n_2426 ^ n_1790;
assign n_2434 = n_2427 ^ x183;
assign n_2435 = n_2428 ^ n_697;
assign n_2436 = n_2431 ^ n_2427;
assign n_2437 = n_2432 ^ n_716;
assign n_2438 = n_1620 ^ n_2433;
assign n_2439 = ~n_2433 & n_1806;
assign n_2440 = n_2435 ^ n_2432;
assign n_2441 = n_2436 ^ x183;
assign n_2442 = ~n_2436 & n_2434;
assign n_2443 = n_1779 & ~n_2438;
assign n_2444 = n_2438 ^ n_1790;
assign n_2445 = n_2245 ^ n_2438;
assign n_2446 = n_2439 ^ n_1620;
assign n_2447 = n_2440 ^ n_716;
assign n_2448 = ~n_2440 & n_2437;
assign n_2449 = n_2429 & ~n_2441;
assign n_2450 = n_2441 ^ n_2429;
assign n_2451 = n_2442 ^ x183;
assign n_2452 = n_2443 ^ n_1306;
assign n_2453 = n_2446 ^ n_1826;
assign n_2454 = n_2447 ^ x182;
assign n_2455 = n_2448 ^ n_716;
assign n_2456 = n_2451 ^ x182;
assign n_2457 = n_2451 ^ n_2447;
assign n_2458 = n_2452 ^ n_741;
assign n_2459 = n_1657 ^ n_2453;
assign n_2460 = ~n_2453 & ~n_1836;
assign n_2461 = n_2455 ^ n_2452;
assign n_2462 = n_2456 ^ n_2447;
assign n_2463 = ~n_2454 & n_2457;
assign n_2464 = ~n_1816 & n_2459;
assign n_2465 = n_2459 ^ n_1826;
assign n_2466 = n_2265 ^ n_2459;
assign n_2467 = n_2460 ^ n_1657;
assign n_2468 = n_2461 ^ n_741;
assign n_2469 = ~n_2461 & ~n_2458;
assign n_2470 = n_2449 & n_2462;
assign n_2471 = n_2462 ^ n_2449;
assign n_2472 = n_2463 ^ x182;
assign n_2473 = n_2464 ^ n_1343;
assign n_2474 = n_2467 ^ n_1851;
assign n_2475 = n_2468 ^ x181;
assign n_2476 = n_2469 ^ n_741;
assign n_2477 = n_2472 ^ n_2468;
assign n_2478 = n_2473 ^ n_766;
assign n_2479 = n_1697 ^ n_2474;
assign n_2480 = ~n_2474 & ~n_1859;
assign n_2481 = n_2476 ^ n_766;
assign n_2482 = n_2476 ^ n_2473;
assign n_2483 = n_2477 ^ x181;
assign n_2484 = ~n_2477 & n_2475;
assign n_2485 = n_1845 & ~n_2479;
assign n_2486 = n_2479 ^ n_1851;
assign n_2487 = n_2285 ^ n_2479;
assign n_2488 = n_2480 ^ n_1697;
assign n_2489 = n_2481 ^ n_2473;
assign n_2490 = n_2478 & ~n_2482;
assign n_2491 = n_2470 & ~n_2483;
assign n_2492 = n_2483 ^ n_2470;
assign n_2493 = n_2484 ^ x181;
assign n_2494 = n_2485 ^ n_1378;
assign n_2495 = n_2488 ^ n_1874;
assign n_2496 = n_2489 ^ x180;
assign n_2497 = n_2490 ^ n_766;
assign n_2498 = n_2493 ^ n_2489;
assign n_2499 = n_2494 ^ n_792;
assign n_2500 = n_1734 ^ n_2495;
assign n_2501 = ~n_2495 & n_1881;
assign n_2502 = n_2497 ^ n_792;
assign n_2503 = n_2497 ^ n_2494;
assign n_2504 = n_2498 ^ x180;
assign n_2505 = ~n_2498 & n_2496;
assign n_2506 = ~n_1869 & ~n_2500;
assign n_2507 = n_2500 ^ n_1874;
assign n_2508 = n_2305 ^ n_2500;
assign n_2509 = n_2501 ^ n_1734;
assign n_2510 = n_2502 ^ n_2494;
assign n_2511 = n_2499 & ~n_2503;
assign n_2512 = ~n_2491 & n_2504;
assign n_2513 = n_2505 ^ x180;
assign n_2514 = n_2506 ^ n_1415;
assign n_2515 = n_2509 ^ n_1895;
assign n_2516 = n_2510 ^ x179;
assign n_2517 = n_2511 ^ n_792;
assign n_2518 = n_2513 ^ n_2510;
assign n_2519 = n_2514 ^ n_821;
assign n_2520 = n_1771 ^ n_2515;
assign n_2521 = n_2515 & n_1901;
assign n_2522 = n_2517 ^ n_2514;
assign n_2523 = n_2518 ^ x179;
assign n_2524 = ~n_2518 & n_2516;
assign n_2525 = n_1889 & ~n_2520;
assign n_2526 = n_2520 ^ n_1895;
assign n_2527 = n_2326 ^ n_2520;
assign n_2528 = n_2521 ^ n_1771;
assign n_2529 = n_2522 ^ n_821;
assign n_2530 = ~n_2522 & n_2519;
assign n_2531 = n_2512 ^ n_2523;
assign n_2532 = n_2523 & n_2512;
assign n_2533 = n_2524 ^ x179;
assign n_2534 = n_2525 ^ n_1451;
assign n_2535 = n_2528 ^ n_1811;
assign n_2536 = n_2528 ^ n_1915;
assign n_2537 = n_2530 ^ n_821;
assign n_2538 = n_2531 ^ n_2014;
assign n_2539 = n_2014 & n_2531;
assign n_2540 = n_2533 ^ n_2529;
assign n_2541 = n_2533 ^ x178;
assign n_2542 = n_2534 ^ n_854;
assign n_2543 = n_2535 ^ n_1915;
assign n_2544 = n_1922 & ~n_2536;
assign n_2545 = n_2537 ^ n_854;
assign n_2546 = n_2537 ^ n_2534;
assign n_2547 = ~n_2006 & n_2538;
assign n_2548 = n_2539 ^ n_2042;
assign n_2549 = n_2540 ^ x178;
assign n_2550 = ~n_2540 & n_2541;
assign n_2551 = n_2543 & n_1921;
assign n_2552 = n_2347 ^ n_2543;
assign n_2553 = n_2544 ^ n_1811;
assign n_2554 = n_2545 ^ n_2534;
assign n_2555 = ~n_2542 & ~n_2546;
assign n_2556 = n_2547 ^ n_1111;
assign n_2557 = n_2532 ^ n_2549;
assign n_2558 = n_2549 & n_2532;
assign n_2559 = n_2550 ^ x178;
assign n_2560 = n_2551 ^ n_1492;
assign n_2561 = n_2553 ^ n_1841;
assign n_2562 = n_2553 ^ n_1930;
assign n_2563 = n_2554 ^ x177;
assign n_2564 = n_2555 ^ n_854;
assign n_2565 = n_2556 ^ n_721;
assign n_2566 = n_721 & ~n_2556;
assign n_2567 = n_2548 ^ n_2557;
assign n_2568 = n_2557 ^ n_2539;
assign n_2569 = n_2559 ^ n_2554;
assign n_2570 = n_2560 ^ n_885;
assign n_2571 = n_2561 ^ n_1930;
assign n_2572 = ~n_1937 & ~n_2562;
assign n_2573 = n_2564 ^ n_885;
assign n_2574 = n_2564 ^ n_2560;
assign n_2575 = x199 & ~n_2565;
assign n_2576 = n_2565 ^ x199;
assign n_2577 = n_2566 ^ n_737;
assign n_2578 = n_2041 & n_2567;
assign n_2579 = ~n_2568 & n_2548;
assign n_2580 = n_2569 ^ x177;
assign n_2581 = n_2569 & ~n_2563;
assign n_2582 = ~n_1936 & ~n_2571;
assign n_2583 = n_2369 ^ n_2571;
assign n_2584 = n_2572 ^ n_1841;
assign n_2585 = n_2573 ^ n_2560;
assign n_2586 = n_2570 & n_2574;
assign n_2587 = n_2575 ^ x198;
assign n_2588 = n_2578 ^ n_1148;
assign n_2589 = n_2579 ^ n_2042;
assign n_2590 = n_2558 ^ n_2580;
assign n_2591 = ~n_2580 & n_2558;
assign n_2592 = n_2581 ^ x177;
assign n_2593 = n_2582 ^ n_1520;
assign n_2594 = n_2584 ^ n_1956;
assign n_2595 = n_2585 ^ x176;
assign n_2596 = n_2586 ^ n_885;
assign n_2597 = n_2588 ^ n_2577;
assign n_2598 = n_2588 ^ n_2566;
assign n_2599 = n_2589 ^ n_2083;
assign n_2600 = n_2589 ^ n_2590;
assign n_2601 = n_2590 ^ n_2083;
assign n_2602 = n_2592 ^ n_2585;
assign n_2603 = n_2593 ^ n_916;
assign n_2604 = n_1865 ^ n_2594;
assign n_2605 = n_2594 & ~n_1962;
assign n_2606 = n_2593 ^ n_2596;
assign n_2607 = n_2597 ^ n_2575;
assign n_2608 = n_2597 ^ n_2587;
assign n_2609 = n_2577 & ~n_2598;
assign n_2610 = n_2599 ^ n_2590;
assign n_2611 = n_2600 & n_2601;
assign n_2612 = n_2602 ^ x176;
assign n_2613 = n_2602 & ~n_2595;
assign n_2614 = n_1951 & n_2604;
assign n_2615 = n_2604 ^ n_1956;
assign n_2616 = n_2390 ^ n_2604;
assign n_2617 = n_2605 ^ n_1865;
assign n_2618 = n_2606 ^ n_916;
assign n_2619 = n_2606 & n_2603;
assign n_2620 = n_2587 & ~n_2607;
assign n_2621 = ~n_2608 & n_2576;
assign n_2622 = n_2576 ^ n_2608;
assign n_2623 = n_2609 ^ n_737;
assign n_2624 = n_2072 & n_2610;
assign n_2625 = n_2611 ^ n_2083;
assign n_2626 = n_2591 ^ n_2612;
assign n_2627 = n_2612 & ~n_2591;
assign n_2628 = n_2613 ^ x176;
assign n_2629 = n_2614 ^ n_1571;
assign n_2630 = n_2617 ^ n_1975;
assign n_2631 = n_2618 ^ x191;
assign n_2632 = n_2619 ^ n_916;
assign n_2633 = n_2620 ^ x198;
assign n_2634 = n_2623 ^ n_770;
assign n_2635 = n_2624 ^ n_1198;
assign n_2636 = n_2625 ^ n_2119;
assign n_2637 = n_2625 ^ n_2626;
assign n_2638 = n_2626 ^ n_2119;
assign n_2639 = n_2628 ^ n_2618;
assign n_2640 = n_2629 ^ n_951;
assign n_2641 = n_1887 ^ n_2630;
assign n_2642 = n_2630 & n_1982;
assign n_2643 = n_2632 ^ n_2629;
assign n_2644 = n_2634 ^ n_2635;
assign n_2645 = n_2635 ^ n_770;
assign n_2646 = n_2623 ^ n_2635;
assign n_2647 = n_2636 ^ n_2626;
assign n_2648 = n_2637 & ~n_2638;
assign n_2649 = n_2639 ^ x191;
assign n_2650 = ~n_2639 & n_2631;
assign n_2651 = ~n_2641 & ~n_1981;
assign n_2652 = n_2641 ^ n_1975;
assign n_2653 = n_2412 ^ n_2641;
assign n_2654 = n_2642 ^ n_1887;
assign n_2655 = n_2643 ^ n_951;
assign n_2656 = n_2643 & n_2640;
assign n_2657 = n_2633 ^ n_2644;
assign n_2658 = n_2644 ^ x197;
assign n_2659 = ~n_2645 & n_2646;
assign n_2660 = ~n_2106 & n_2647;
assign n_2661 = n_2648 ^ n_2119;
assign n_2662 = n_2627 ^ n_2649;
assign n_2663 = ~n_2649 & n_2627;
assign n_2664 = n_2650 ^ x191;
assign n_2665 = n_2651 ^ n_1608;
assign n_2666 = n_2654 ^ n_1995;
assign n_2667 = n_2655 ^ x190;
assign n_2668 = n_2656 ^ n_951;
assign n_2669 = n_2657 ^ x197;
assign n_2670 = n_2657 & ~n_2658;
assign n_2671 = n_2659 ^ n_770;
assign n_2672 = n_2660 ^ n_1236;
assign n_2673 = n_2661 ^ n_2149;
assign n_2674 = n_2662 ^ n_2149;
assign n_2675 = n_2661 ^ n_2662;
assign n_2676 = n_2664 ^ n_2655;
assign n_2677 = n_2665 ^ n_983;
assign n_2678 = n_1907 ^ n_2666;
assign n_2679 = n_2666 & ~n_2002;
assign n_2680 = n_2668 ^ n_983;
assign n_2681 = n_2668 ^ n_2665;
assign n_2682 = ~n_2669 & ~n_2621;
assign n_2683 = n_2621 ^ n_2669;
assign n_2684 = n_2670 ^ x197;
assign n_2685 = n_2671 ^ n_806;
assign n_2686 = n_2672 ^ n_806;
assign n_2687 = n_2671 ^ n_2672;
assign n_2688 = n_2673 ^ n_2662;
assign n_2689 = n_2674 & n_2675;
assign n_2690 = n_2676 ^ x190;
assign n_2691 = n_2676 & ~n_2667;
assign n_2692 = ~n_2678 & n_2001;
assign n_2693 = n_2678 ^ n_1995;
assign n_2694 = n_2430 ^ n_2678;
assign n_2695 = n_2679 ^ n_1907;
assign n_2696 = n_2680 ^ n_2665;
assign n_2697 = n_2677 & n_2681;
assign n_2698 = n_2685 ^ n_2672;
assign n_2699 = n_2686 & ~n_2687;
assign n_2700 = n_2139 & ~n_2688;
assign n_2701 = n_2689 ^ n_2149;
assign n_2702 = n_2663 ^ n_2690;
assign n_2703 = n_2690 & n_2663;
assign n_2704 = n_2691 ^ x190;
assign n_2705 = n_2692 ^ n_1645;
assign n_2706 = n_2695 ^ n_2017;
assign n_2707 = n_2696 ^ x189;
assign n_2708 = n_2697 ^ n_983;
assign n_2709 = n_2684 ^ n_2698;
assign n_2710 = n_2698 ^ x196;
assign n_2711 = n_2699 ^ n_806;
assign n_2712 = n_2700 ^ n_1267;
assign n_2713 = n_2701 ^ n_2174;
assign n_2714 = n_2702 ^ n_2174;
assign n_2715 = n_2701 ^ n_2702;
assign n_2716 = n_2704 ^ n_2696;
assign n_2717 = n_2705 ^ n_1015;
assign n_2718 = n_1928 ^ n_2706;
assign n_2719 = n_2706 & n_2026;
assign n_2720 = n_2708 ^ n_1015;
assign n_2721 = n_2708 ^ n_2705;
assign n_2722 = n_2709 ^ x196;
assign n_2723 = ~n_2709 & n_2710;
assign n_2724 = n_2711 ^ n_837;
assign n_2725 = n_2712 ^ n_837;
assign n_2726 = n_2711 ^ n_2712;
assign n_2727 = n_2713 ^ n_2702;
assign n_2728 = n_2714 & n_2715;
assign n_2729 = n_2716 ^ x189;
assign n_2730 = ~n_2716 & n_2707;
assign n_2731 = n_2718 & ~n_2025;
assign n_2732 = n_2718 ^ n_2017;
assign n_2733 = n_2450 ^ n_2718;
assign n_2734 = n_2719 ^ n_1928;
assign n_2735 = n_2720 ^ n_2705;
assign n_2736 = n_2717 & ~n_2721;
assign n_2737 = n_2722 & n_2682;
assign n_2738 = n_2682 ^ n_2722;
assign n_2739 = n_2723 ^ x196;
assign n_2740 = n_2724 ^ n_2712;
assign n_2741 = n_2725 & ~n_2726;
assign n_2742 = ~n_2166 & n_2727;
assign n_2743 = n_2728 ^ n_2174;
assign n_2744 = n_2703 ^ n_2729;
assign n_2745 = ~n_2729 & n_2703;
assign n_2746 = n_2730 ^ x189;
assign n_2747 = n_2731 ^ n_1685;
assign n_2748 = n_2734 ^ n_2044;
assign n_2749 = n_2735 ^ x188;
assign n_2750 = n_2736 ^ n_1015;
assign n_2751 = n_2739 ^ n_2740;
assign n_2752 = n_2740 ^ x195;
assign n_2753 = n_2741 ^ n_837;
assign n_2754 = n_2742 ^ n_1300;
assign n_2755 = n_2743 ^ n_2195;
assign n_2756 = n_2744 ^ n_2195;
assign n_2757 = n_2743 ^ n_2744;
assign n_2758 = n_2746 ^ x188;
assign n_2759 = n_2746 ^ n_2735;
assign n_2760 = n_2747 ^ n_1046;
assign n_2761 = n_1949 ^ n_2748;
assign n_2762 = ~n_2748 & ~n_2056;
assign n_2763 = n_2750 ^ n_1046;
assign n_2764 = n_2750 ^ n_2747;
assign n_2765 = n_2751 ^ x195;
assign n_2766 = ~n_2751 & n_2752;
assign n_2767 = n_2753 ^ n_870;
assign n_2768 = n_2754 ^ n_870;
assign n_2769 = n_2753 ^ n_2754;
assign n_2770 = n_2755 ^ n_2744;
assign n_2771 = n_2756 & n_2757;
assign n_2772 = n_2758 ^ n_2735;
assign n_2773 = ~n_2749 & n_2759;
assign n_2774 = n_2761 & n_2055;
assign n_2775 = n_2761 ^ n_2044;
assign n_2776 = n_2471 ^ n_2761;
assign n_2777 = n_2762 ^ n_1949;
assign n_2778 = n_2763 ^ n_2747;
assign n_2779 = n_2760 & n_2764;
assign n_2780 = ~n_2737 & ~n_2765;
assign n_2781 = n_2765 ^ n_2737;
assign n_2782 = n_2766 ^ x195;
assign n_2783 = n_2767 ^ n_2754;
assign n_2784 = n_2768 & ~n_2769;
assign n_2785 = ~n_2188 & ~n_2770;
assign n_2786 = n_2771 ^ n_2195;
assign n_2787 = n_2772 ^ n_2745;
assign n_2788 = ~n_2745 & ~n_2772;
assign n_2789 = n_2773 ^ x188;
assign n_2790 = n_2774 ^ n_1722;
assign n_2791 = n_2777 ^ n_2077;
assign n_2792 = n_2778 ^ x187;
assign n_2793 = n_2779 ^ n_1046;
assign n_2794 = n_2782 ^ n_2783;
assign n_2795 = n_2783 ^ x194;
assign n_2796 = n_2784 ^ n_870;
assign n_2797 = n_2785 ^ n_1336;
assign n_2798 = n_2786 ^ n_2209;
assign n_2799 = n_2786 ^ n_2787;
assign n_2800 = n_2787 ^ n_2209;
assign n_2801 = n_2789 ^ n_2778;
assign n_2802 = n_2790 ^ n_1080;
assign n_2803 = n_1968 ^ n_2791;
assign n_2804 = n_2791 & ~n_2089;
assign n_2805 = n_2793 ^ n_1080;
assign n_2806 = n_2793 ^ n_2790;
assign n_2807 = n_2794 ^ x194;
assign n_2808 = ~n_2794 & n_2795;
assign n_2809 = n_2796 ^ n_900;
assign n_2810 = n_2797 ^ n_900;
assign n_2811 = n_2796 ^ n_2797;
assign n_2812 = n_2798 ^ n_2787;
assign n_2813 = ~n_2799 & ~n_2800;
assign n_2814 = n_2801 ^ x187;
assign n_2815 = n_2801 & ~n_2792;
assign n_2816 = ~n_2803 & ~n_2088;
assign n_2817 = n_2803 ^ n_2077;
assign n_2818 = n_2492 ^ n_2803;
assign n_2819 = n_2804 ^ n_1968;
assign n_2820 = n_2805 ^ n_2790;
assign n_2821 = n_2802 & n_2806;
assign n_2822 = ~n_2780 & n_2807;
assign n_2823 = n_2807 ^ n_2780;
assign n_2824 = n_2808 ^ x194;
assign n_2825 = n_2809 ^ n_2797;
assign n_2826 = n_2810 & n_2811;
assign n_2827 = ~n_2208 & ~n_2812;
assign n_2828 = n_2813 ^ n_2209;
assign n_2829 = n_2788 ^ n_2814;
assign n_2830 = ~n_2814 & n_2788;
assign n_2831 = n_2815 ^ x187;
assign n_2832 = n_2816 ^ n_1759;
assign n_2833 = n_2819 ^ n_2113;
assign n_2834 = n_2820 ^ x186;
assign n_2835 = n_2821 ^ n_1080;
assign n_2836 = n_2824 ^ n_2825;
assign n_2837 = n_2825 ^ x193;
assign n_2838 = n_2826 ^ n_900;
assign n_2839 = n_2827 ^ n_1372;
assign n_2840 = n_2828 ^ n_2233;
assign n_2841 = n_2829 ^ n_2233;
assign n_2842 = n_2828 ^ n_2829;
assign n_2843 = n_2831 ^ n_2820;
assign n_2844 = n_2832 ^ n_1114;
assign n_2845 = ~n_2833 & ~n_2114;
assign n_2846 = n_2833 ^ n_2491;
assign n_2847 = n_2833 ^ n_2101;
assign n_2848 = n_2835 ^ n_1114;
assign n_2849 = n_2835 ^ n_2832;
assign n_2850 = n_2836 ^ x193;
assign n_2851 = ~n_2836 & n_2837;
assign n_2852 = n_2838 ^ n_932;
assign n_2853 = n_2839 ^ n_932;
assign n_2854 = n_2838 ^ n_2839;
assign n_2855 = n_2840 ^ n_2829;
assign n_2856 = n_2841 & ~n_2842;
assign n_2857 = n_2843 ^ x186;
assign n_2858 = ~n_2843 & n_2834;
assign n_2859 = n_2845 ^ n_1786;
assign n_2860 = n_2846 ^ n_2504;
assign n_2861 = n_2848 ^ n_2832;
assign n_2862 = ~n_2844 & n_2849;
assign n_2863 = n_2822 & n_2850;
assign n_2864 = n_2850 ^ n_2822;
assign n_2865 = n_2851 ^ x193;
assign n_2866 = n_2852 ^ n_2839;
assign n_2867 = ~n_2853 & n_2854;
assign n_2868 = ~n_2855 & n_2240;
assign n_2869 = n_2856 ^ n_2233;
assign n_2870 = n_2830 ^ n_2857;
assign n_2871 = n_2857 & n_2830;
assign n_2872 = n_2858 ^ x186;
assign n_2873 = n_2859 ^ n_1139;
assign n_2874 = n_2861 ^ x185;
assign n_2875 = n_2862 ^ n_1114;
assign n_2876 = n_2865 ^ n_2866;
assign n_2877 = n_2866 ^ x192;
assign n_2878 = n_2867 ^ n_932;
assign n_2879 = n_2868 ^ n_1409;
assign n_2880 = n_2869 ^ n_2252;
assign n_2881 = n_2870 ^ n_2252;
assign n_2882 = n_2869 ^ n_2870;
assign n_2883 = n_2872 ^ n_2861;
assign n_2884 = n_2875 ^ x184;
assign n_2885 = n_2876 ^ x192;
assign n_2886 = ~n_2876 & n_2877;
assign n_2887 = n_2878 ^ n_966;
assign n_2888 = n_2879 ^ n_966;
assign n_2889 = n_2878 ^ n_2879;
assign n_2890 = n_2880 ^ n_2870;
assign n_2891 = ~n_2881 & n_2882;
assign n_2892 = n_2883 ^ x185;
assign n_2893 = ~n_2883 & n_2874;
assign n_2894 = n_2884 ^ n_2873;
assign n_2895 = n_2863 & n_2885;
assign n_2896 = n_2885 ^ n_2863;
assign n_2897 = n_2886 ^ x192;
assign n_2898 = n_2887 ^ n_2879;
assign n_2899 = ~n_2888 & ~n_2889;
assign n_2900 = n_2890 & n_2260;
assign n_2901 = n_2891 ^ n_2252;
assign n_2902 = n_2871 ^ n_2892;
assign n_2903 = ~n_2892 & ~n_2871;
assign n_2904 = n_2893 ^ x185;
assign n_2905 = n_2897 ^ n_2898;
assign n_2906 = n_2898 ^ x207;
assign n_2907 = n_2899 ^ n_966;
assign n_2908 = n_2900 ^ n_1446;
assign n_2909 = n_2901 ^ n_2272;
assign n_2910 = n_2902 ^ n_2272;
assign n_2911 = n_2901 ^ n_2902;
assign n_2912 = n_2904 ^ n_2903;
assign n_2913 = n_2905 ^ x207;
assign n_2914 = ~n_2905 & n_2906;
assign n_2915 = n_2907 ^ n_998;
assign n_2916 = n_2908 ^ n_998;
assign n_2917 = n_2907 ^ n_2908;
assign n_2918 = n_2909 ^ n_2902;
assign n_2919 = ~n_2910 & ~n_2911;
assign n_2920 = n_2912 ^ n_2894;
assign n_2921 = n_2895 & n_2913;
assign n_2922 = n_2913 ^ n_2895;
assign n_2923 = n_2914 ^ x207;
assign n_2924 = n_2915 ^ n_2908;
assign n_2925 = n_2916 & n_2917;
assign n_2926 = n_2918 & n_2280;
assign n_2927 = n_2919 ^ n_2272;
assign n_2928 = n_2920 ^ n_2291;
assign n_2929 = n_2923 ^ n_2924;
assign n_2930 = n_2924 ^ x206;
assign n_2931 = n_2925 ^ n_998;
assign n_2932 = n_2926 ^ n_1485;
assign n_2933 = n_2927 ^ n_2291;
assign n_2934 = n_2927 ^ n_2920;
assign n_2935 = n_2929 ^ x206;
assign n_2936 = ~n_2929 & n_2930;
assign n_2937 = n_2931 ^ n_1030;
assign n_2938 = n_2932 ^ n_1030;
assign n_2939 = n_2931 ^ n_2932;
assign n_2940 = n_2933 ^ n_2920;
assign n_2941 = ~n_2928 & n_2934;
assign n_2942 = ~n_2921 & ~n_2935;
assign n_2943 = n_2935 ^ n_2921;
assign n_2944 = n_2936 ^ x206;
assign n_2945 = n_2937 ^ n_2932;
assign n_2946 = n_2938 & n_2939;
assign n_2947 = ~n_2940 & n_2299;
assign n_2948 = n_2941 ^ n_2291;
assign n_2949 = n_2944 ^ n_2945;
assign n_2950 = n_2945 ^ x205;
assign n_2951 = n_2946 ^ n_1030;
assign n_2952 = n_2947 ^ n_1525;
assign n_2953 = n_2948 ^ n_2312;
assign n_2954 = n_2949 ^ x205;
assign n_2955 = n_2949 & ~n_2950;
assign n_2956 = n_2951 ^ n_1061;
assign n_2957 = n_2952 ^ n_1061;
assign n_2958 = n_2951 ^ n_2952;
assign n_2959 = n_2049 ^ n_2953;
assign n_2960 = ~n_2953 & n_2320;
assign n_2961 = n_2942 & n_2954;
assign n_2962 = n_2954 ^ n_2942;
assign n_2963 = n_2955 ^ x205;
assign n_2964 = n_2956 ^ n_2952;
assign n_2965 = ~n_2957 & ~n_2958;
assign n_2966 = n_2959 & ~n_2319;
assign n_2967 = n_2959 ^ n_2312;
assign n_2968 = n_2960 ^ n_2049;
assign n_2969 = n_2963 ^ n_2964;
assign n_2970 = n_2964 ^ x204;
assign n_2971 = n_2965 ^ n_1061;
assign n_2972 = n_2966 ^ n_1565;
assign n_2973 = n_2968 ^ n_2333;
assign n_2974 = n_2968 ^ n_2086;
assign n_2975 = n_2969 ^ x204;
assign n_2976 = n_2969 & ~n_2970;
assign n_2977 = n_2971 ^ n_1095;
assign n_2978 = n_2972 ^ n_1095;
assign n_2979 = n_2971 ^ n_2972;
assign n_2980 = n_2973 ^ n_2086;
assign n_2981 = n_2974 & n_2341;
assign n_2982 = ~n_2961 & ~n_2975;
assign n_2983 = n_2975 ^ n_2961;
assign n_2984 = n_2976 ^ x204;
assign n_2985 = n_2977 ^ n_2972;
assign n_2986 = ~n_2978 & ~n_2979;
assign n_2987 = n_2980 & ~n_2340;
assign n_2988 = n_2981 ^ n_2333;
assign n_2989 = n_2984 ^ n_2985;
assign n_2990 = n_2985 ^ x203;
assign n_2991 = n_2986 ^ n_1095;
assign n_2992 = n_2987 ^ n_1601;
assign n_2993 = n_2988 ^ n_2355;
assign n_2994 = n_2989 ^ x203;
assign n_2995 = ~n_2989 & n_2990;
assign n_2996 = n_2991 ^ n_1131;
assign n_2997 = n_2992 ^ n_1131;
assign n_2998 = n_2991 ^ n_2992;
assign n_2999 = n_2154 ^ n_2993;
assign n_3000 = n_2993 & ~n_2363;
assign n_3001 = n_2982 & n_2994;
assign n_3002 = n_2994 ^ n_2982;
assign n_3003 = n_2995 ^ x203;
assign n_3004 = n_2996 ^ n_2992;
assign n_3005 = n_2997 & ~n_2998;
assign n_3006 = n_2999 & ~n_2362;
assign n_3007 = n_2999 ^ n_2355;
assign n_3008 = n_3000 ^ n_2154;
assign n_3009 = n_3003 ^ n_3004;
assign n_3010 = n_3004 ^ x202;
assign n_3011 = n_3005 ^ n_1131;
assign n_3012 = n_3006 ^ n_1638;
assign n_3013 = n_3008 ^ n_2376;
assign n_3014 = n_3009 ^ x202;
assign n_3015 = ~n_3009 & n_3010;
assign n_3016 = n_3011 ^ n_1171;
assign n_3017 = n_3012 ^ n_1171;
assign n_3018 = n_3011 ^ n_3012;
assign n_3019 = n_2186 ^ n_3013;
assign n_3020 = n_3013 & ~n_2384;
assign n_3021 = n_3001 & n_3014;
assign n_3022 = n_3014 ^ n_3001;
assign n_3023 = n_3015 ^ x202;
assign n_3024 = n_3016 ^ n_3012;
assign n_3025 = ~n_3017 & n_3018;
assign n_3026 = n_3019 & ~n_2383;
assign n_3027 = n_3019 ^ n_2376;
assign n_3028 = n_3020 ^ n_2186;
assign n_3029 = n_3023 ^ n_3024;
assign n_3030 = n_3024 ^ x201;
assign n_3031 = n_3025 ^ n_1171;
assign n_3032 = n_3026 ^ n_1677;
assign n_3033 = n_3028 ^ n_2399;
assign n_3034 = n_3028 ^ n_2392;
assign n_3035 = n_3029 ^ x201;
assign n_3036 = n_3029 & ~n_3030;
assign n_3037 = n_3031 ^ n_1205;
assign n_3038 = n_3032 ^ n_1205;
assign n_3039 = n_3031 ^ n_3032;
assign n_3040 = ~n_3033 & ~n_2400;
assign n_3041 = n_3033 ^ n_2392;
assign n_3042 = n_2399 & ~n_3034;
assign n_3043 = ~n_3021 & n_3035;
assign n_3044 = n_3035 ^ n_3021;
assign n_3045 = n_3036 ^ x201;
assign n_3046 = n_3037 ^ n_3032;
assign n_3047 = n_3038 & n_3039;
assign n_3048 = n_3040 ^ n_1715;
assign n_3049 = n_3042 ^ n_2207;
assign n_3050 = n_3045 ^ n_3046;
assign n_3051 = n_3046 ^ x200;
assign n_3052 = n_3047 ^ n_1205;
assign n_3053 = n_3048 ^ n_1238;
assign n_3054 = n_3049 ^ n_2419;
assign n_3055 = n_3050 ^ x200;
assign n_3056 = ~n_3050 & n_3051;
assign n_3057 = n_3052 ^ n_3048;
assign n_3058 = n_3052 ^ n_3053;
assign n_3059 = n_2227 ^ n_3054;
assign n_3060 = n_3054 & ~n_2425;
assign n_3061 = n_3043 ^ n_3055;
assign n_3062 = n_3055 & ~n_3043;
assign n_3063 = n_3056 ^ x200;
assign n_3064 = n_3053 & n_3057;
assign n_3065 = n_2414 & n_3059;
assign n_3066 = n_2576 ^ n_3059;
assign n_3067 = n_3059 ^ n_2419;
assign n_3068 = n_3060 ^ n_2227;
assign n_3069 = n_2538 & ~n_3061;
assign n_3070 = n_3061 ^ n_2538;
assign n_3071 = n_3058 ^ n_3063;
assign n_3072 = n_3063 ^ x215;
assign n_3073 = n_3064 ^ n_1238;
assign n_3074 = n_3065 ^ n_1752;
assign n_3075 = n_3068 ^ n_2245;
assign n_3076 = n_3068 ^ n_2438;
assign n_3077 = n_3069 ^ n_2567;
assign n_3078 = n_2531 & ~n_3070;
assign n_3079 = n_3071 ^ x215;
assign n_3080 = n_3071 & n_3072;
assign n_3081 = n_3073 ^ n_3074;
assign n_3082 = n_3074 ^ n_1271;
assign n_3083 = n_3075 ^ n_2438;
assign n_3084 = ~n_2445 & ~n_3076;
assign n_3085 = n_3078 ^ n_2014;
assign n_3086 = n_3079 ^ n_3062;
assign n_3087 = n_3062 & ~n_3079;
assign n_3088 = n_3080 ^ x215;
assign n_3089 = n_3081 ^ n_1271;
assign n_3090 = ~n_3081 & ~n_3082;
assign n_3091 = n_3083 & n_2444;
assign n_3092 = n_2622 ^ n_3083;
assign n_3093 = n_3084 ^ n_2245;
assign n_3094 = ~n_1111 & n_3085;
assign n_3095 = n_3085 ^ n_1111;
assign n_3096 = n_3086 ^ n_3069;
assign n_3097 = n_3086 ^ n_3077;
assign n_3098 = n_3088 ^ n_3089;
assign n_3099 = n_3089 ^ x214;
assign n_3100 = n_3090 ^ n_1271;
assign n_3101 = n_3091 ^ n_1790;
assign n_3102 = n_3093 ^ n_2459;
assign n_3103 = n_3094 ^ n_1148;
assign n_3104 = x231 & ~n_3095;
assign n_3105 = n_3095 ^ x231;
assign n_3106 = n_3077 & n_3096;
assign n_3107 = n_2568 & ~n_3097;
assign n_3108 = n_3098 ^ x214;
assign n_3109 = n_3098 & ~n_3099;
assign n_3110 = n_3100 ^ n_1306;
assign n_3111 = n_3101 ^ n_1306;
assign n_3112 = n_3100 ^ n_3101;
assign n_3113 = n_2265 ^ n_3102;
assign n_3114 = ~n_3102 & ~n_2466;
assign n_3115 = n_3104 ^ x230;
assign n_3116 = n_3106 ^ n_2567;
assign n_3117 = n_3107 ^ n_2042;
assign n_3118 = n_3087 ^ n_3108;
assign n_3119 = ~n_3108 & n_3087;
assign n_3120 = n_3109 ^ x214;
assign n_3121 = n_3110 ^ n_3101;
assign n_3122 = n_3111 & ~n_3112;
assign n_3123 = ~n_3113 & ~n_2465;
assign n_3124 = n_3113 ^ n_2459;
assign n_3125 = n_2683 ^ n_3113;
assign n_3126 = n_3114 ^ n_2265;
assign n_3127 = n_3116 ^ n_2610;
assign n_3128 = n_3117 ^ n_3094;
assign n_3129 = n_3117 ^ n_3103;
assign n_3130 = n_3118 ^ n_2610;
assign n_3131 = n_3116 ^ n_3118;
assign n_3132 = n_3120 ^ n_3121;
assign n_3133 = n_3121 ^ x213;
assign n_3134 = n_3122 ^ n_1306;
assign n_3135 = n_3123 ^ n_1826;
assign n_3136 = n_3126 ^ n_2479;
assign n_3137 = n_3127 ^ n_3118;
assign n_3138 = n_3103 & ~n_3128;
assign n_3139 = n_3129 ^ n_3104;
assign n_3140 = n_3129 ^ n_3115;
assign n_3141 = ~n_3130 & n_3131;
assign n_3142 = n_3132 ^ x213;
assign n_3143 = n_3132 & ~n_3133;
assign n_3144 = n_3134 ^ n_1343;
assign n_3145 = n_3135 ^ n_1343;
assign n_3146 = n_3134 ^ n_3135;
assign n_3147 = n_2285 ^ n_3136;
assign n_3148 = ~n_3136 & ~n_2487;
assign n_3149 = ~n_2600 & ~n_3137;
assign n_3150 = n_3138 ^ n_1148;
assign n_3151 = n_3115 & ~n_3139;
assign n_3152 = n_3140 & ~n_3105;
assign n_3153 = n_3105 ^ n_3140;
assign n_3154 = n_3141 ^ n_2610;
assign n_3155 = n_3142 ^ n_3119;
assign n_3156 = n_3119 & ~n_3142;
assign n_3157 = n_3143 ^ x213;
assign n_3158 = n_3144 ^ n_3135;
assign n_3159 = ~n_3145 & ~n_3146;
assign n_3160 = n_3147 & ~n_2486;
assign n_3161 = n_3147 ^ n_2479;
assign n_3162 = n_3147 ^ n_2738;
assign n_3163 = n_3148 ^ n_2285;
assign n_3164 = n_3149 ^ n_2083;
assign n_3165 = n_3150 ^ n_1198;
assign n_3166 = n_3151 ^ x230;
assign n_3167 = n_3154 ^ n_3155;
assign n_3168 = n_3155 ^ n_2647;
assign n_3169 = n_3157 ^ n_3158;
assign n_3170 = n_3158 ^ x212;
assign n_3171 = n_3159 ^ n_1343;
assign n_3172 = n_3160 ^ n_1851;
assign n_3173 = n_3163 ^ n_2305;
assign n_3174 = n_3163 ^ n_2500;
assign n_3175 = n_3164 ^ n_1198;
assign n_3176 = n_3150 ^ n_3164;
assign n_3177 = n_3165 ^ n_3164;
assign n_3178 = n_3167 ^ n_2647;
assign n_3179 = n_3167 & ~n_3168;
assign n_3180 = n_3169 ^ x212;
assign n_3181 = ~n_3169 & n_3170;
assign n_3182 = n_3171 ^ n_1378;
assign n_3183 = n_3172 ^ n_1378;
assign n_3184 = n_3171 ^ n_3172;
assign n_3185 = n_3173 ^ n_2500;
assign n_3186 = n_2508 & n_3174;
assign n_3187 = n_3175 & n_3176;
assign n_3188 = n_3166 ^ n_3177;
assign n_3189 = n_3177 ^ x229;
assign n_3190 = ~n_2637 & ~n_3178;
assign n_3191 = n_3179 ^ n_2647;
assign n_3192 = n_3156 ^ n_3180;
assign n_3193 = n_3180 & n_3156;
assign n_3194 = n_3181 ^ x212;
assign n_3195 = n_3182 ^ n_3172;
assign n_3196 = n_3183 & ~n_3184;
assign n_3197 = n_3185 & n_2507;
assign n_3198 = n_2781 ^ n_3185;
assign n_3199 = n_3186 ^ n_2305;
assign n_3200 = n_3187 ^ n_1198;
assign n_3201 = n_3188 ^ x229;
assign n_3202 = ~n_3188 & n_3189;
assign n_3203 = n_3190 ^ n_2119;
assign n_3204 = n_3191 ^ n_2688;
assign n_3205 = n_3192 ^ n_2688;
assign n_3206 = n_3191 ^ n_3192;
assign n_3207 = n_3194 ^ n_3195;
assign n_3208 = n_3195 ^ x211;
assign n_3209 = n_3196 ^ n_1378;
assign n_3210 = n_3197 ^ n_1874;
assign n_3211 = n_3199 ^ n_2520;
assign n_3212 = n_3200 ^ n_1236;
assign n_3213 = n_3152 & n_3201;
assign n_3214 = n_3201 ^ n_3152;
assign n_3215 = n_3202 ^ x229;
assign n_3216 = n_3203 ^ n_1236;
assign n_3217 = n_3200 ^ n_3203;
assign n_3218 = n_3204 ^ n_3192;
assign n_3219 = ~n_3205 & ~n_3206;
assign n_3220 = n_3207 ^ x211;
assign n_3221 = ~n_3207 & n_3208;
assign n_3222 = n_3209 ^ n_1415;
assign n_3223 = n_3210 ^ n_1415;
assign n_3224 = n_3209 ^ n_3210;
assign n_3225 = n_2326 ^ n_3211;
assign n_3226 = ~n_3211 & n_2527;
assign n_3227 = n_3212 ^ n_3203;
assign n_3228 = n_3215 ^ x228;
assign n_3229 = ~n_3216 & ~n_3217;
assign n_3230 = ~n_2675 & ~n_3218;
assign n_3231 = n_3219 ^ n_2688;
assign n_3232 = n_3193 ^ n_3220;
assign n_3233 = ~n_3220 & ~n_3193;
assign n_3234 = n_3221 ^ x211;
assign n_3235 = n_3222 ^ n_3210;
assign n_3236 = ~n_3223 & n_3224;
assign n_3237 = ~n_3225 & ~n_2526;
assign n_3238 = n_3225 ^ n_2520;
assign n_3239 = n_2823 ^ n_3225;
assign n_3240 = n_3226 ^ n_2326;
assign n_3241 = n_3227 ^ x228;
assign n_3242 = n_3215 ^ n_3227;
assign n_3243 = n_3228 ^ n_3227;
assign n_3244 = n_3229 ^ n_1236;
assign n_3245 = n_3230 ^ n_2149;
assign n_3246 = n_3231 ^ n_2727;
assign n_3247 = n_3232 ^ n_2727;
assign n_3248 = n_3231 ^ n_3232;
assign n_3249 = n_3234 ^ n_3235;
assign n_3250 = n_3235 ^ x210;
assign n_3251 = n_3236 ^ n_1415;
assign n_3252 = n_3237 ^ n_1895;
assign n_3253 = n_3240 ^ n_2543;
assign n_3254 = n_3241 & ~n_3242;
assign n_3255 = n_3243 & n_3213;
assign n_3256 = n_3213 ^ n_3243;
assign n_3257 = n_3244 ^ n_1267;
assign n_3258 = n_3245 ^ n_1267;
assign n_3259 = n_3244 ^ n_3245;
assign n_3260 = n_3246 ^ n_3232;
assign n_3261 = ~n_3247 & ~n_3248;
assign n_3262 = n_3249 ^ x210;
assign n_3263 = n_3249 & ~n_3250;
assign n_3264 = n_3251 ^ n_1451;
assign n_3265 = n_3252 ^ n_1451;
assign n_3266 = n_3251 ^ n_3252;
assign n_3267 = n_2347 ^ n_3253;
assign n_3268 = n_3253 & ~n_2552;
assign n_3269 = n_3254 ^ x228;
assign n_3270 = n_3257 ^ n_3245;
assign n_3271 = n_3258 & ~n_3259;
assign n_3272 = ~n_2715 & n_3260;
assign n_3273 = n_3261 ^ n_2727;
assign n_3274 = n_3233 ^ n_3262;
assign n_3275 = n_3262 & n_3233;
assign n_3276 = n_3263 ^ x210;
assign n_3277 = n_3264 ^ n_3252;
assign n_3278 = n_3265 & ~n_3266;
assign n_3279 = n_2535 & n_3267;
assign n_3280 = n_3267 ^ n_2543;
assign n_3281 = n_2864 ^ n_3267;
assign n_3282 = n_3268 ^ n_2347;
assign n_3283 = n_3269 ^ n_3270;
assign n_3284 = n_3270 ^ x227;
assign n_3285 = n_3271 ^ n_1267;
assign n_3286 = n_3272 ^ n_2174;
assign n_3287 = n_3273 ^ n_3274;
assign n_3288 = n_3274 ^ n_2770;
assign n_3289 = n_3276 ^ n_3277;
assign n_3290 = n_3277 ^ x209;
assign n_3291 = n_3278 ^ n_1451;
assign n_3292 = n_3279 ^ n_1915;
assign n_3293 = n_3282 ^ n_2571;
assign n_3294 = n_3283 ^ x227;
assign n_3295 = ~n_3283 & n_3284;
assign n_3296 = n_3285 ^ n_1300;
assign n_3297 = n_3286 ^ n_1300;
assign n_3298 = n_3285 ^ n_3286;
assign n_3299 = n_3287 ^ n_2770;
assign n_3300 = n_3287 & n_3288;
assign n_3301 = n_3289 ^ x209;
assign n_3302 = ~n_3289 & n_3290;
assign n_3303 = n_3291 ^ n_1492;
assign n_3304 = n_3292 ^ n_1492;
assign n_3305 = n_3291 ^ n_3292;
assign n_3306 = n_2369 ^ n_3293;
assign n_3307 = ~n_3293 & n_2583;
assign n_3308 = n_3255 & n_3294;
assign n_3309 = n_3294 ^ n_3255;
assign n_3310 = n_3295 ^ x227;
assign n_3311 = n_3296 ^ n_3286;
assign n_3312 = ~n_3297 & n_3298;
assign n_3313 = ~n_2757 & n_3299;
assign n_3314 = n_3300 ^ n_2770;
assign n_3315 = n_3301 ^ n_3275;
assign n_3316 = ~n_3275 & n_3301;
assign n_3317 = n_3302 ^ x209;
assign n_3318 = n_3303 ^ n_3292;
assign n_3319 = n_3304 & ~n_3305;
assign n_3320 = ~n_2561 & ~n_3306;
assign n_3321 = n_2896 ^ n_3306;
assign n_3322 = n_3306 ^ n_2571;
assign n_3323 = n_3307 ^ n_2369;
assign n_3324 = n_3310 ^ n_3311;
assign n_3325 = n_3311 ^ x226;
assign n_3326 = n_3312 ^ n_1300;
assign n_3327 = n_3313 ^ n_2195;
assign n_3328 = n_3314 ^ n_2812;
assign n_3329 = n_3315 ^ n_2812;
assign n_3330 = n_3314 ^ n_3315;
assign n_3331 = n_3317 ^ n_3318;
assign n_3332 = n_3318 ^ x208;
assign n_3333 = n_3319 ^ n_1492;
assign n_3334 = n_3320 ^ n_1930;
assign n_3335 = n_3323 ^ n_2390;
assign n_3336 = n_3323 ^ n_2604;
assign n_3337 = n_3324 ^ x226;
assign n_3338 = n_3324 & ~n_3325;
assign n_3339 = n_3326 ^ n_1336;
assign n_3340 = n_3327 ^ n_1336;
assign n_3341 = n_3326 ^ n_3327;
assign n_3342 = n_3328 ^ n_3315;
assign n_3343 = n_3329 & ~n_3330;
assign n_3344 = n_3331 ^ x208;
assign n_3345 = ~n_3331 & n_3332;
assign n_3346 = n_3334 ^ n_3333;
assign n_3347 = n_3334 ^ n_1520;
assign n_3348 = n_3335 ^ n_2604;
assign n_3349 = n_2616 & n_3336;
assign n_3350 = n_3308 & ~n_3337;
assign n_3351 = n_3337 ^ n_3308;
assign n_3352 = n_3338 ^ x226;
assign n_3353 = n_3339 ^ n_3327;
assign n_3354 = ~n_3340 & ~n_3341;
assign n_3355 = n_2799 & ~n_3342;
assign n_3356 = n_3343 ^ n_2812;
assign n_3357 = n_3344 ^ n_3316;
assign n_3358 = n_3316 & n_3344;
assign n_3359 = n_3345 ^ x208;
assign n_3360 = n_3346 ^ n_1520;
assign n_3361 = ~n_3346 & ~n_3347;
assign n_3362 = ~n_3348 & n_2615;
assign n_3363 = n_2922 ^ n_3348;
assign n_3364 = n_3349 ^ n_2390;
assign n_3365 = n_3352 ^ n_3353;
assign n_3366 = n_3353 ^ x225;
assign n_3367 = n_3354 ^ n_1336;
assign n_3368 = n_3355 ^ n_2209;
assign n_3369 = n_3356 ^ n_2855;
assign n_3370 = n_3357 ^ n_2855;
assign n_3371 = n_3356 ^ n_3357;
assign n_3372 = n_3359 ^ n_3360;
assign n_3373 = n_3360 ^ x223;
assign n_3374 = n_3361 ^ n_1520;
assign n_3375 = n_3362 ^ n_1956;
assign n_3376 = n_3364 ^ n_2641;
assign n_3377 = n_3365 ^ x225;
assign n_3378 = n_3365 & ~n_3366;
assign n_3379 = n_3367 ^ n_1372;
assign n_3380 = n_3368 ^ n_1372;
assign n_3381 = n_3367 ^ n_3368;
assign n_3382 = n_3369 ^ n_3357;
assign n_3383 = ~n_3370 & n_3371;
assign n_3384 = n_3372 ^ x223;
assign n_3385 = n_3372 & ~n_3373;
assign n_3386 = n_3374 ^ n_1571;
assign n_3387 = n_3375 ^ n_1571;
assign n_3388 = n_3374 ^ n_3375;
assign n_3389 = n_2412 ^ n_3376;
assign n_3390 = n_3376 & ~n_2653;
assign n_3391 = n_3350 & ~n_3377;
assign n_3392 = n_3377 ^ n_3350;
assign n_3393 = n_3378 ^ x225;
assign n_3394 = n_3379 ^ n_3368;
assign n_3395 = ~n_3380 & ~n_3381;
assign n_3396 = n_2842 & n_3382;
assign n_3397 = n_3383 ^ n_2855;
assign n_3398 = n_3384 ^ n_3358;
assign n_3399 = n_3358 & ~n_3384;
assign n_3400 = n_3385 ^ x223;
assign n_3401 = n_3386 ^ n_3375;
assign n_3402 = n_3387 & n_3388;
assign n_3403 = ~n_3389 & ~n_2652;
assign n_3404 = n_3389 ^ n_2641;
assign n_3405 = n_2943 ^ n_3389;
assign n_3406 = n_3390 ^ n_2412;
assign n_3407 = n_3393 ^ n_3394;
assign n_3408 = n_3394 ^ x224;
assign n_3409 = n_3395 ^ n_1372;
assign n_3410 = n_3396 ^ n_2233;
assign n_3411 = n_3397 ^ n_2890;
assign n_3412 = n_3398 ^ n_2890;
assign n_3413 = n_3397 ^ n_3398;
assign n_3414 = n_3400 ^ n_3401;
assign n_3415 = n_3401 ^ x222;
assign n_3416 = n_3402 ^ n_1571;
assign n_3417 = n_3403 ^ n_1975;
assign n_3418 = n_3406 ^ n_2678;
assign n_3419 = n_3407 ^ x224;
assign n_3420 = ~n_3407 & n_3408;
assign n_3421 = n_3409 ^ n_1409;
assign n_3422 = n_3410 ^ n_1409;
assign n_3423 = n_3409 ^ n_3410;
assign n_3424 = n_3411 ^ n_3398;
assign n_3425 = ~n_3412 & ~n_3413;
assign n_3426 = n_3414 ^ x222;
assign n_3427 = n_3414 & ~n_3415;
assign n_3428 = n_3416 ^ n_1608;
assign n_3429 = n_3417 ^ n_1608;
assign n_3430 = n_3416 ^ n_3417;
assign n_3431 = n_2430 ^ n_3418;
assign n_3432 = n_3418 & ~n_2694;
assign n_3433 = n_3391 & n_3419;
assign n_3434 = n_3419 ^ n_3391;
assign n_3435 = n_3420 ^ x224;
assign n_3436 = n_3421 ^ n_3410;
assign n_3437 = n_3422 & n_3423;
assign n_3438 = ~n_2882 & n_3424;
assign n_3439 = n_3425 ^ n_2890;
assign n_3440 = n_3399 ^ n_3426;
assign n_3441 = ~n_3426 & n_3399;
assign n_3442 = n_3427 ^ x222;
assign n_3443 = n_3428 ^ n_3417;
assign n_3444 = ~n_3429 & ~n_3430;
assign n_3445 = ~n_3431 & n_2693;
assign n_3446 = n_3431 ^ n_2678;
assign n_3447 = n_2962 ^ n_3431;
assign n_3448 = n_3432 ^ n_2430;
assign n_3449 = n_3435 ^ n_3436;
assign n_3450 = n_3436 ^ x239;
assign n_3451 = n_3437 ^ n_1409;
assign n_3452 = n_3438 ^ n_2252;
assign n_3453 = n_3439 ^ n_2918;
assign n_3454 = n_3440 ^ n_2918;
assign n_3455 = n_3439 ^ n_3440;
assign n_3456 = n_3442 ^ n_3443;
assign n_3457 = n_3443 ^ x221;
assign n_3458 = n_3444 ^ n_1608;
assign n_3459 = n_3445 ^ n_1995;
assign n_3460 = n_3448 ^ n_2718;
assign n_3461 = n_3449 ^ x239;
assign n_3462 = ~n_3449 & n_3450;
assign n_3463 = n_3451 ^ n_1446;
assign n_3464 = n_3452 ^ n_1446;
assign n_3465 = n_3451 ^ n_3452;
assign n_3466 = n_3453 ^ n_3440;
assign n_3467 = ~n_3454 & n_3455;
assign n_3468 = n_3456 ^ x221;
assign n_3469 = n_3456 & ~n_3457;
assign n_3470 = n_3458 ^ n_1645;
assign n_3471 = n_3459 ^ n_1645;
assign n_3472 = n_3458 ^ n_3459;
assign n_3473 = n_2450 ^ n_3460;
assign n_3474 = ~n_3460 & n_2733;
assign n_3475 = ~n_3433 & ~n_3461;
assign n_3476 = n_3461 ^ n_3433;
assign n_3477 = n_3462 ^ x239;
assign n_3478 = n_3463 ^ n_3452;
assign n_3479 = n_3464 & ~n_3465;
assign n_3480 = n_2911 & ~n_3466;
assign n_3481 = n_3467 ^ n_2918;
assign n_3482 = n_3468 ^ n_3441;
assign n_3483 = n_3441 & ~n_3468;
assign n_3484 = n_3469 ^ x221;
assign n_3485 = n_3470 ^ n_3459;
assign n_3486 = n_3471 & ~n_3472;
assign n_3487 = n_3473 & ~n_2732;
assign n_3488 = n_3473 ^ n_2718;
assign n_3489 = n_2983 ^ n_3473;
assign n_3490 = n_3474 ^ n_2450;
assign n_3491 = n_3477 ^ n_3478;
assign n_3492 = n_3478 ^ x238;
assign n_3493 = n_3479 ^ n_1446;
assign n_3494 = n_3480 ^ n_2272;
assign n_3495 = n_3481 ^ n_2940;
assign n_3496 = n_3482 ^ n_2940;
assign n_3497 = n_3481 ^ n_3482;
assign n_3498 = n_3484 ^ n_3485;
assign n_3499 = n_3485 ^ x220;
assign n_3500 = n_3486 ^ n_1645;
assign n_3501 = n_3487 ^ n_2017;
assign n_3502 = n_3490 ^ n_2761;
assign n_3503 = n_3491 ^ x238;
assign n_3504 = n_3491 & ~n_3492;
assign n_3505 = n_3493 ^ n_1485;
assign n_3506 = n_3494 ^ n_1485;
assign n_3507 = n_3493 ^ n_3494;
assign n_3508 = n_3495 ^ n_3482;
assign n_3509 = n_3496 & n_3497;
assign n_3510 = n_3498 ^ x220;
assign n_3511 = n_3498 & ~n_3499;
assign n_3512 = n_3500 ^ n_1685;
assign n_3513 = n_3501 ^ n_1685;
assign n_3514 = n_3500 ^ n_3501;
assign n_3515 = n_2471 ^ n_3502;
assign n_3516 = ~n_3502 & ~n_2776;
assign n_3517 = ~n_3475 & ~n_3503;
assign n_3518 = n_3504 ^ x238;
assign n_3519 = n_3505 ^ n_3494;
assign n_3520 = n_3506 & n_3507;
assign n_3521 = ~n_2934 & n_3508;
assign n_3522 = n_3509 ^ n_2940;
assign n_3523 = n_3510 ^ n_3483;
assign n_3524 = ~n_3483 & n_3510;
assign n_3525 = n_3511 ^ x220;
assign n_3526 = n_3512 ^ n_3501;
assign n_3527 = ~n_3513 & ~n_3514;
assign n_3528 = ~n_3515 & ~n_2775;
assign n_3529 = n_3515 ^ n_2761;
assign n_3530 = n_3002 ^ n_3515;
assign n_3531 = n_3516 ^ n_2471;
assign n_3532 = n_3518 ^ n_3519;
assign n_3533 = n_3519 ^ x237;
assign n_3534 = n_3520 ^ n_1485;
assign n_3535 = n_3521 ^ n_2291;
assign n_3536 = n_3522 ^ n_2959;
assign n_3537 = n_3523 ^ n_2959;
assign n_3538 = n_3522 ^ n_3523;
assign n_3539 = n_3525 ^ x219;
assign n_3540 = n_3526 ^ x219;
assign n_3541 = n_3525 ^ n_3526;
assign n_3542 = n_3527 ^ n_1685;
assign n_3543 = n_3528 ^ n_2044;
assign n_3544 = n_3531 ^ n_2803;
assign n_3545 = n_3532 ^ x237;
assign n_3546 = n_3532 & ~n_3533;
assign n_3547 = n_3534 ^ n_1525;
assign n_3548 = n_3535 ^ n_1525;
assign n_3549 = n_3534 ^ n_3535;
assign n_3550 = n_3536 ^ n_3523;
assign n_3551 = n_3537 & n_3538;
assign n_3552 = n_3539 ^ n_3526;
assign n_3553 = n_3540 & ~n_3541;
assign n_3554 = n_3542 ^ n_3543;
assign n_3555 = n_3543 ^ n_1722;
assign n_3556 = n_3544 ^ n_2492;
assign n_3557 = ~n_3544 & ~n_2818;
assign n_3558 = n_3545 ^ n_3517;
assign n_3559 = ~n_3517 & n_3545;
assign n_3560 = n_3546 ^ x237;
assign n_3561 = n_3547 ^ n_3535;
assign n_3562 = n_3548 & ~n_3549;
assign n_3563 = ~n_3550 & n_2967;
assign n_3564 = n_3551 ^ n_2959;
assign n_3565 = n_3552 ^ n_3524;
assign n_3566 = ~n_3524 & n_3552;
assign n_3567 = n_3553 ^ x219;
assign n_3568 = n_3554 ^ n_1722;
assign n_3569 = n_3554 & n_3555;
assign n_3570 = n_3556 & n_2817;
assign n_3571 = n_3556 ^ n_2803;
assign n_3572 = n_3022 ^ n_3556;
assign n_3573 = n_3557 ^ n_2492;
assign n_3574 = n_3558 ^ n_3070;
assign n_3575 = ~n_3070 & n_3558;
assign n_3576 = n_3560 ^ n_3561;
assign n_3577 = n_3561 ^ x236;
assign n_3578 = n_3562 ^ n_1525;
assign n_3579 = n_3563 ^ n_2312;
assign n_3580 = n_3564 ^ n_2980;
assign n_3581 = n_3565 ^ n_2980;
assign n_3582 = n_3564 ^ n_3565;
assign n_3583 = n_3567 ^ n_3568;
assign n_3584 = n_3568 ^ x218;
assign n_3585 = n_3569 ^ n_1722;
assign n_3586 = n_3570 ^ n_2077;
assign n_3587 = n_3573 ^ n_2860;
assign n_3588 = ~n_3061 & ~n_3574;
assign n_3589 = n_3575 ^ n_3097;
assign n_3590 = n_3576 ^ x236;
assign n_3591 = ~n_3576 & n_3577;
assign n_3592 = n_3578 ^ n_1565;
assign n_3593 = n_3579 ^ n_1565;
assign n_3594 = n_3578 ^ n_3579;
assign n_3595 = n_3580 ^ n_3565;
assign n_3596 = ~n_3581 & n_3582;
assign n_3597 = n_3583 ^ x218;
assign n_3598 = ~n_3583 & n_3584;
assign n_3599 = n_3585 ^ n_3586;
assign n_3600 = n_3586 ^ n_1759;
assign n_3601 = n_3587 & n_2847;
assign n_3602 = n_3587 ^ n_2833;
assign n_3603 = n_3588 ^ n_2538;
assign n_3604 = n_3559 ^ n_3590;
assign n_3605 = n_3590 & ~n_3559;
assign n_3606 = n_3591 ^ x236;
assign n_3607 = n_3592 ^ n_3579;
assign n_3608 = ~n_3593 & ~n_3594;
assign n_3609 = ~n_2974 & ~n_3595;
assign n_3610 = n_3596 ^ n_2980;
assign n_3611 = n_3566 ^ n_3597;
assign n_3612 = ~n_3597 & ~n_3566;
assign n_3613 = n_3598 ^ x218;
assign n_3614 = n_3599 ^ n_1759;
assign n_3615 = ~n_3599 & ~n_3600;
assign n_3616 = n_3601 ^ n_2101;
assign n_3617 = n_3603 ^ n_2014;
assign n_3618 = n_2014 & n_3603;
assign n_3619 = n_3604 ^ n_3589;
assign n_3620 = n_3604 ^ n_3575;
assign n_3621 = n_3606 ^ n_3607;
assign n_3622 = n_3607 ^ x235;
assign n_3623 = n_3608 ^ n_1565;
assign n_3624 = n_3609 ^ n_2333;
assign n_3625 = n_3610 ^ n_2999;
assign n_3626 = n_3611 ^ n_2999;
assign n_3627 = n_3610 ^ n_3611;
assign n_3628 = n_3613 ^ x217;
assign n_3629 = n_3614 ^ x217;
assign n_3630 = n_3614 ^ n_3613;
assign n_3631 = n_3615 ^ n_1759;
assign n_3632 = n_3616 ^ n_1786;
assign n_3633 = x263 & n_3617;
assign n_3634 = n_3617 ^ x263;
assign n_3635 = n_3618 ^ n_2042;
assign n_3636 = ~n_3096 & n_3619;
assign n_3637 = ~n_3589 & n_3620;
assign n_3638 = n_3621 ^ x235;
assign n_3639 = n_3621 & ~n_3622;
assign n_3640 = n_3623 ^ n_1601;
assign n_3641 = n_3624 ^ n_1601;
assign n_3642 = n_3623 ^ n_3624;
assign n_3643 = n_3625 ^ n_3611;
assign n_3644 = ~n_3626 & n_3627;
assign n_3645 = n_3614 ^ n_3628;
assign n_3646 = n_3629 & ~n_3630;
assign n_3647 = n_3631 ^ x216;
assign n_3648 = n_3633 ^ x262;
assign n_3649 = n_3636 ^ n_2567;
assign n_3650 = n_3637 ^ n_3097;
assign n_3651 = n_3605 ^ n_3638;
assign n_3652 = n_3638 & ~n_3605;
assign n_3653 = n_3639 ^ x235;
assign n_3654 = n_3640 ^ n_3624;
assign n_3655 = ~n_3641 & ~n_3642;
assign n_3656 = ~n_3643 & n_3007;
assign n_3657 = n_3644 ^ n_2999;
assign n_3658 = n_3612 ^ n_3645;
assign n_3659 = n_3645 & ~n_3612;
assign n_3660 = n_3646 ^ x217;
assign n_3661 = n_3647 ^ n_3632;
assign n_3662 = n_3649 ^ n_3635;
assign n_3663 = n_3649 ^ n_3618;
assign n_3664 = n_3650 ^ n_3651;
assign n_3665 = n_3651 ^ n_3137;
assign n_3666 = n_3653 ^ n_3654;
assign n_3667 = n_3654 ^ x234;
assign n_3668 = n_3655 ^ n_1601;
assign n_3669 = n_3656 ^ n_2355;
assign n_3670 = n_3657 ^ n_3019;
assign n_3671 = n_3658 ^ n_3019;
assign n_3672 = n_3657 ^ n_3658;
assign n_3673 = n_3660 ^ n_3661;
assign n_3674 = n_3662 ^ n_3633;
assign n_3675 = n_3662 ^ n_3648;
assign n_3676 = n_3635 & ~n_3663;
assign n_3677 = n_3664 ^ n_3137;
assign n_3678 = n_3664 & ~n_3665;
assign n_3679 = n_3666 ^ x234;
assign n_3680 = ~n_3666 & n_3667;
assign n_3681 = n_3668 ^ n_1638;
assign n_3682 = n_3669 ^ n_1638;
assign n_3683 = n_3668 ^ n_3669;
assign n_3684 = n_3670 ^ n_3658;
assign n_3685 = ~n_3671 & n_3672;
assign n_3686 = n_3673 ^ n_3659;
assign n_3687 = n_3648 & ~n_3674;
assign n_3688 = n_3676 ^ n_2042;
assign n_3689 = ~n_3131 & n_3677;
assign n_3690 = n_3678 ^ n_3137;
assign n_3691 = n_3652 ^ n_3679;
assign n_3692 = n_3679 & ~n_3652;
assign n_3693 = n_3680 ^ x234;
assign n_3694 = n_3681 ^ n_3669;
assign n_3695 = ~n_3682 & ~n_3683;
assign n_3696 = ~n_3684 & n_3027;
assign n_3697 = n_3685 ^ n_3019;
assign n_3698 = n_3686 ^ n_3033;
assign n_3699 = n_3687 ^ x262;
assign n_3700 = n_3688 ^ n_2083;
assign n_3701 = n_3689 ^ n_2610;
assign n_3702 = n_3690 ^ n_3178;
assign n_3703 = n_3691 ^ n_3690;
assign n_3704 = n_3693 ^ n_3694;
assign n_3705 = n_3694 ^ x233;
assign n_3706 = n_3695 ^ n_1638;
assign n_3707 = n_3696 ^ n_2376;
assign n_3708 = n_3697 ^ n_3033;
assign n_3709 = n_3697 ^ n_3686;
assign n_3710 = n_3700 ^ n_3701;
assign n_3711 = n_3701 ^ n_2083;
assign n_3712 = n_3688 ^ n_3701;
assign n_3713 = n_3691 ^ n_3702;
assign n_3714 = n_3702 & ~n_3703;
assign n_3715 = n_3704 ^ x233;
assign n_3716 = n_3704 & ~n_3705;
assign n_3717 = n_3706 ^ n_1677;
assign n_3718 = n_3707 ^ n_1677;
assign n_3719 = n_3706 ^ n_3707;
assign n_3720 = n_3708 ^ n_3686;
assign n_3721 = ~n_3698 & ~n_3709;
assign n_3722 = n_3699 ^ n_3710;
assign n_3723 = n_3710 ^ x261;
assign n_3724 = ~n_3711 & ~n_3712;
assign n_3725 = ~n_3167 & ~n_3713;
assign n_3726 = n_3714 ^ n_3178;
assign n_3727 = n_3692 ^ n_3715;
assign n_3728 = ~n_3715 & n_3692;
assign n_3729 = n_3716 ^ x233;
assign n_3730 = n_3717 ^ n_3707;
assign n_3731 = ~n_3718 & n_3719;
assign n_3732 = ~n_3720 & n_3041;
assign n_3733 = n_3721 ^ n_3033;
assign n_3734 = n_3722 ^ x261;
assign n_3735 = n_3722 & ~n_3723;
assign n_3736 = n_3724 ^ n_2083;
assign n_3737 = n_3725 ^ n_2647;
assign n_3738 = n_3726 ^ n_3218;
assign n_3739 = n_3727 ^ n_3218;
assign n_3740 = n_3726 ^ n_3727;
assign n_3741 = n_3729 ^ n_3730;
assign n_3742 = n_3730 ^ x232;
assign n_3743 = n_3731 ^ n_1677;
assign n_3744 = n_3732 ^ n_2392;
assign n_3745 = n_3733 ^ n_3066;
assign n_3746 = n_3733 ^ n_2576;
assign n_3747 = n_3735 ^ x261;
assign n_3748 = n_3736 ^ n_2119;
assign n_3749 = n_3737 ^ n_2119;
assign n_3750 = n_3736 ^ n_3737;
assign n_3751 = n_3738 ^ n_3727;
assign n_3752 = n_3739 & ~n_3740;
assign n_3753 = n_3741 ^ x232;
assign n_3754 = ~n_3741 & n_3742;
assign n_3755 = n_3743 ^ n_3744;
assign n_3756 = n_3744 ^ n_1715;
assign n_3757 = ~n_3745 & n_3067;
assign n_3758 = n_3066 & n_3746;
assign n_3759 = n_3748 ^ n_3737;
assign n_3760 = ~n_3749 & n_3750;
assign n_3761 = n_3206 & ~n_3751;
assign n_3762 = n_3752 ^ n_3218;
assign n_3763 = n_3753 ^ n_3728;
assign n_3764 = ~n_3728 & ~n_3753;
assign n_3765 = n_3754 ^ x232;
assign n_3766 = n_3755 ^ n_1715;
assign n_3767 = ~n_3755 & ~n_3756;
assign n_3768 = n_3757 ^ n_2419;
assign n_3769 = n_3758 ^ n_3059;
assign n_3770 = n_3747 ^ n_3759;
assign n_3771 = n_3759 ^ x260;
assign n_3772 = n_3760 ^ n_2119;
assign n_3773 = n_3761 ^ n_2688;
assign n_3774 = n_3762 ^ n_3260;
assign n_3775 = n_3763 ^ n_3260;
assign n_3776 = n_3762 ^ n_3763;
assign n_3777 = n_3765 ^ x247;
assign n_3778 = n_3766 ^ x247;
assign n_3779 = n_3765 ^ n_3766;
assign n_3780 = n_3767 ^ n_1715;
assign n_3781 = n_3769 ^ n_3083;
assign n_3782 = n_3770 ^ x260;
assign n_3783 = ~n_3770 & n_3771;
assign n_3784 = n_3772 ^ n_2149;
assign n_3785 = n_3773 ^ n_2149;
assign n_3786 = n_3772 ^ n_3773;
assign n_3787 = n_3774 ^ n_3763;
assign n_3788 = ~n_3775 & ~n_3776;
assign n_3789 = n_3777 ^ n_3766;
assign n_3790 = n_3778 & ~n_3779;
assign n_3791 = n_3780 ^ n_1752;
assign n_3792 = n_3768 ^ n_3780;
assign n_3793 = n_2622 ^ n_3781;
assign n_3794 = ~n_3781 & n_3092;
assign n_3795 = n_3783 ^ x260;
assign n_3796 = n_3784 ^ n_3773;
assign n_3797 = ~n_3785 & ~n_3786;
assign n_3798 = n_3248 & n_3787;
assign n_3799 = n_3788 ^ n_3260;
assign n_3800 = n_3764 ^ n_3789;
assign n_3801 = n_3789 & ~n_3764;
assign n_3802 = n_3790 ^ x247;
assign n_3803 = n_3768 ^ n_3791;
assign n_3804 = n_3791 & ~n_3792;
assign n_3805 = ~n_3075 & n_3793;
assign n_3806 = n_3793 ^ n_3083;
assign n_3807 = n_3794 ^ n_2622;
assign n_3808 = n_3795 ^ n_3796;
assign n_3809 = n_3796 ^ x259;
assign n_3810 = n_3797 ^ n_2149;
assign n_3811 = n_3798 ^ n_2727;
assign n_3812 = n_3799 ^ n_3299;
assign n_3813 = n_3800 ^ n_3299;
assign n_3814 = n_3799 ^ n_3800;
assign n_3815 = n_3802 ^ n_3803;
assign n_3816 = n_3803 ^ x246;
assign n_3817 = n_3804 ^ n_1752;
assign n_3818 = n_3805 ^ n_2438;
assign n_3819 = n_3807 ^ n_3113;
assign n_3820 = n_3808 ^ x259;
assign n_3821 = ~n_3808 & n_3809;
assign n_3822 = n_3810 ^ n_2174;
assign n_3823 = n_3811 ^ n_3810;
assign n_3824 = n_3812 ^ n_3800;
assign n_3825 = ~n_3813 & n_3814;
assign n_3826 = n_3815 ^ x246;
assign n_3827 = ~n_3815 & n_3816;
assign n_3828 = n_3817 ^ n_1790;
assign n_3829 = n_3818 ^ n_1790;
assign n_3830 = n_3817 ^ n_3818;
assign n_3831 = n_2683 ^ n_3819;
assign n_3832 = n_3819 & ~n_3125;
assign n_3833 = ~n_3782 & ~n_3820;
assign n_3834 = n_3820 ^ n_3782;
assign n_3835 = n_3821 ^ x259;
assign n_3836 = n_3811 ^ n_3822;
assign n_3837 = ~n_3822 & ~n_3823;
assign n_3838 = ~n_3287 & ~n_3824;
assign n_3839 = n_3825 ^ n_3299;
assign n_3840 = n_3801 ^ n_3826;
assign n_3841 = ~n_3826 & ~n_3801;
assign n_3842 = n_3827 ^ x246;
assign n_3843 = n_3828 ^ n_3818;
assign n_3844 = n_3829 & n_3830;
assign n_3845 = ~n_3831 & ~n_3124;
assign n_3846 = n_3831 ^ n_3113;
assign n_3847 = n_3832 ^ n_2683;
assign n_3848 = n_3835 ^ n_3836;
assign n_3849 = n_3836 ^ x258;
assign n_3850 = n_3837 ^ n_2174;
assign n_3851 = n_3838 ^ n_2770;
assign n_3852 = n_3839 ^ n_3342;
assign n_3853 = n_3840 ^ n_3342;
assign n_3854 = n_3839 ^ n_3840;
assign n_3855 = n_3842 ^ n_3843;
assign n_3856 = n_3843 ^ x245;
assign n_3857 = n_3844 ^ n_1790;
assign n_3858 = n_3845 ^ n_2459;
assign n_3859 = n_3847 ^ n_2738;
assign n_3860 = n_3847 ^ n_3147;
assign n_3861 = n_3848 ^ x258;
assign n_3862 = n_3848 & ~n_3849;
assign n_3863 = n_3850 ^ n_2195;
assign n_3864 = n_3851 ^ n_2195;
assign n_3865 = n_3850 ^ n_3851;
assign n_3866 = n_3852 ^ n_3840;
assign n_3867 = n_3853 & n_3854;
assign n_3868 = n_3855 ^ x245;
assign n_3869 = ~n_3855 & n_3856;
assign n_3870 = n_3857 ^ n_1826;
assign n_3871 = n_3858 ^ n_1826;
assign n_3872 = n_3857 ^ n_3858;
assign n_3873 = n_3859 ^ n_3147;
assign n_3874 = n_3162 & ~n_3860;
assign n_3875 = ~n_3833 & ~n_3861;
assign n_3876 = n_3861 ^ n_3833;
assign n_3877 = n_3862 ^ x258;
assign n_3878 = n_3863 ^ n_3851;
assign n_3879 = ~n_3864 & ~n_3865;
assign n_3880 = n_3330 & n_3866;
assign n_3881 = n_3634 ^ n_3866;
assign n_3882 = n_3867 ^ n_3342;
assign n_3883 = n_3868 ^ n_3841;
assign n_3884 = n_3841 & ~n_3868;
assign n_3885 = n_3869 ^ x245;
assign n_3886 = n_3870 ^ n_3858;
assign n_3887 = ~n_3871 & n_3872;
assign n_3888 = n_3873 & ~n_3161;
assign n_3889 = n_3874 ^ n_2738;
assign n_3890 = n_3877 ^ n_3878;
assign n_3891 = n_3878 ^ x257;
assign n_3892 = n_3879 ^ n_2195;
assign n_3893 = n_3880 ^ n_2812;
assign n_3894 = n_3882 ^ n_3382;
assign n_3895 = n_3883 ^ n_3382;
assign n_3896 = n_3882 ^ n_3883;
assign n_3897 = n_3885 ^ n_3886;
assign n_3898 = n_3886 ^ x244;
assign n_3899 = n_3887 ^ n_1826;
assign n_3900 = n_3888 ^ n_2479;
assign n_3901 = n_3889 ^ n_3185;
assign n_3902 = n_3890 ^ x257;
assign n_3903 = ~n_3890 & n_3891;
assign n_3904 = n_3892 ^ n_2209;
assign n_3905 = n_3893 ^ n_2209;
assign n_3906 = n_3892 ^ n_3893;
assign n_3907 = n_3894 ^ n_3883;
assign n_3908 = n_3895 & n_3896;
assign n_3909 = n_3897 ^ x244;
assign n_3910 = ~n_3897 & n_3898;
assign n_3911 = n_3899 ^ n_1851;
assign n_3912 = n_3900 ^ n_1851;
assign n_3913 = n_3899 ^ n_3900;
assign n_3914 = n_2781 ^ n_3901;
assign n_3915 = ~n_3901 & ~n_3198;
assign n_3916 = ~n_3875 & ~n_3902;
assign n_3917 = n_3902 ^ n_3875;
assign n_3918 = n_3903 ^ x257;
assign n_3919 = n_3904 ^ n_3893;
assign n_3920 = n_3905 & n_3906;
assign n_3921 = ~n_3371 & ~n_3907;
assign n_3922 = n_3675 ^ n_3907;
assign n_3923 = n_3908 ^ n_3382;
assign n_3924 = n_3909 ^ n_3884;
assign n_3925 = ~n_3884 & n_3909;
assign n_3926 = n_3910 ^ x244;
assign n_3927 = n_3911 ^ n_3900;
assign n_3928 = ~n_3912 & ~n_3913;
assign n_3929 = ~n_3173 & ~n_3914;
assign n_3930 = n_3914 ^ n_3185;
assign n_3931 = n_3915 ^ n_2781;
assign n_3932 = n_3918 ^ n_3919;
assign n_3933 = n_3919 ^ x256;
assign n_3934 = n_3920 ^ n_2209;
assign n_3935 = n_3921 ^ n_2855;
assign n_3936 = n_3923 ^ n_3424;
assign n_3937 = n_3924 ^ n_3424;
assign n_3938 = n_3923 ^ n_3924;
assign n_3939 = n_3926 ^ n_3927;
assign n_3940 = n_3927 ^ x243;
assign n_3941 = n_3928 ^ n_1851;
assign n_3942 = n_3929 ^ n_2500;
assign n_3943 = n_3931 ^ n_3225;
assign n_3944 = n_3932 ^ x256;
assign n_3945 = ~n_3932 & n_3933;
assign n_3946 = n_3934 ^ n_2233;
assign n_3947 = n_3935 ^ n_2233;
assign n_3948 = n_3934 ^ n_3935;
assign n_3949 = n_3936 ^ n_3924;
assign n_3950 = ~n_3937 & n_3938;
assign n_3951 = n_3939 ^ x243;
assign n_3952 = ~n_3939 & n_3940;
assign n_3953 = n_3941 ^ n_1874;
assign n_3954 = n_3942 ^ n_1874;
assign n_3955 = n_3941 ^ n_3942;
assign n_3956 = n_2823 ^ n_3943;
assign n_3957 = ~n_3943 & n_3239;
assign n_3958 = ~n_3944 & n_3916;
assign n_3959 = n_3916 ^ n_3944;
assign n_3960 = n_3945 ^ x256;
assign n_3961 = n_3946 ^ n_3935;
assign n_3962 = n_3947 & ~n_3948;
assign n_3963 = n_3413 & ~n_3949;
assign n_3964 = n_3734 ^ n_3949;
assign n_3965 = n_3950 ^ n_3424;
assign n_3966 = n_3925 ^ n_3951;
assign n_3967 = n_3951 & n_3925;
assign n_3968 = n_3952 ^ x243;
assign n_3969 = n_3953 ^ n_3942;
assign n_3970 = n_3954 & n_3955;
assign n_3971 = ~n_3956 & n_3238;
assign n_3972 = n_3956 ^ n_3105;
assign n_3973 = n_3956 ^ n_3225;
assign n_3974 = n_3957 ^ n_2823;
assign n_3975 = n_3960 ^ n_3961;
assign n_3976 = n_3961 ^ x271;
assign n_3977 = n_3962 ^ n_2233;
assign n_3978 = n_3963 ^ n_2890;
assign n_3979 = n_3965 ^ n_3466;
assign n_3980 = n_3966 ^ n_3466;
assign n_3981 = n_3965 ^ n_3966;
assign n_3982 = n_3968 ^ n_3969;
assign n_3983 = n_3969 ^ x242;
assign n_3984 = n_3970 ^ n_1874;
assign n_3985 = n_3971 ^ n_2520;
assign n_3986 = n_3974 ^ n_3267;
assign n_3987 = n_3975 ^ x271;
assign n_3988 = n_3975 & ~n_3976;
assign n_3989 = n_3977 ^ n_2252;
assign n_3990 = n_3978 ^ n_2252;
assign n_3991 = n_3977 ^ n_3978;
assign n_3992 = n_3979 ^ n_3966;
assign n_3993 = ~n_3980 & ~n_3981;
assign n_3994 = n_3982 ^ x242;
assign n_3995 = ~n_3982 & n_3983;
assign n_3996 = n_3984 ^ n_1895;
assign n_3997 = n_3985 ^ n_1895;
assign n_3998 = n_3984 ^ n_3985;
assign n_3999 = n_2864 ^ n_3986;
assign n_4000 = n_3986 & n_3281;
assign n_4001 = ~n_3958 & ~n_3987;
assign n_4002 = n_3987 ^ n_3958;
assign n_4003 = n_3988 ^ x271;
assign n_4004 = n_3989 ^ n_3978;
assign n_4005 = ~n_3990 & n_3991;
assign n_4006 = ~n_3455 & ~n_3992;
assign n_4007 = n_3782 ^ n_3992;
assign n_4008 = n_3993 ^ n_3466;
assign n_4009 = n_3994 ^ n_3967;
assign n_4010 = n_3967 & n_3994;
assign n_4011 = n_3995 ^ x242;
assign n_4012 = n_3996 ^ n_3985;
assign n_4013 = ~n_3997 & ~n_3998;
assign n_4014 = ~n_3999 & n_3280;
assign n_4015 = n_3999 ^ n_3267;
assign n_4016 = n_3153 ^ n_3999;
assign n_4017 = n_4000 ^ n_2864;
assign n_4018 = n_4003 ^ n_4004;
assign n_4019 = n_4004 ^ x270;
assign n_4020 = n_4005 ^ n_2252;
assign n_4021 = n_4006 ^ n_2918;
assign n_4022 = n_4008 ^ n_3508;
assign n_4023 = n_4009 ^ n_3508;
assign n_4024 = n_4008 ^ n_4009;
assign n_4025 = n_4011 ^ n_4012;
assign n_4026 = n_4012 ^ x241;
assign n_4027 = n_4013 ^ n_1895;
assign n_4028 = n_4014 ^ n_2543;
assign n_4029 = n_4017 ^ n_3321;
assign n_4030 = n_4017 ^ n_3306;
assign n_4031 = n_4018 ^ x270;
assign n_4032 = ~n_4018 & n_4019;
assign n_4033 = n_4020 ^ n_2272;
assign n_4034 = n_4021 ^ n_4020;
assign n_4035 = n_4022 ^ n_4009;
assign n_4036 = n_4023 & n_4024;
assign n_4037 = n_4025 ^ x241;
assign n_4038 = ~n_4025 & n_4026;
assign n_4039 = n_4027 ^ n_1915;
assign n_4040 = n_4028 ^ n_1915;
assign n_4041 = n_4027 ^ n_4028;
assign n_4042 = ~n_4029 & n_3322;
assign n_4043 = n_4029 ^ n_3306;
assign n_4044 = n_3214 ^ n_4029;
assign n_4045 = ~n_3321 & n_4030;
assign n_4046 = n_4001 & n_4031;
assign n_4047 = n_4031 ^ n_4001;
assign n_4048 = n_4032 ^ x270;
assign n_4049 = n_4021 ^ n_4033;
assign n_4050 = ~n_4033 & n_4034;
assign n_4051 = ~n_3497 & ~n_4035;
assign n_4052 = n_3834 ^ n_4035;
assign n_4053 = n_4036 ^ n_3508;
assign n_4054 = n_4010 ^ n_4037;
assign n_4055 = ~n_4037 & ~n_4010;
assign n_4056 = n_4038 ^ x241;
assign n_4057 = n_4039 ^ n_4028;
assign n_4058 = n_4040 & ~n_4041;
assign n_4059 = n_4042 ^ n_2571;
assign n_4060 = n_4045 ^ n_2896;
assign n_4061 = n_4048 ^ n_4049;
assign n_4062 = n_4049 ^ x269;
assign n_4063 = n_4050 ^ n_2272;
assign n_4064 = n_4051 ^ n_2940;
assign n_4065 = n_4053 ^ n_3550;
assign n_4066 = n_4054 ^ n_3550;
assign n_4067 = n_4053 ^ n_4054;
assign n_4068 = n_4056 ^ n_4057;
assign n_4069 = n_4057 ^ x240;
assign n_4070 = n_4058 ^ n_1915;
assign n_4071 = n_4059 ^ n_1930;
assign n_4072 = n_4060 ^ n_2922;
assign n_4073 = n_4060 ^ n_3348;
assign n_4074 = n_4061 ^ x269;
assign n_4075 = n_4061 & ~n_4062;
assign n_4076 = n_4063 ^ n_2291;
assign n_4077 = n_4064 ^ n_2291;
assign n_4078 = n_4063 ^ n_4064;
assign n_4079 = n_4065 ^ n_4054;
assign n_4080 = n_4066 & n_4067;
assign n_4081 = n_4068 ^ x240;
assign n_4082 = ~n_4068 & n_4069;
assign n_4083 = n_4059 ^ n_4070;
assign n_4084 = n_4072 ^ n_3348;
assign n_4085 = ~n_3363 & n_4073;
assign n_4086 = n_4046 & ~n_4074;
assign n_4087 = n_4074 ^ n_4046;
assign n_4088 = n_4075 ^ x269;
assign n_4089 = n_4076 ^ n_4064;
assign n_4090 = ~n_4077 & n_4078;
assign n_4091 = ~n_3538 & n_4079;
assign n_4092 = n_3876 ^ n_4079;
assign n_4093 = n_4080 ^ n_3550;
assign n_4094 = n_4055 ^ n_4081;
assign n_4095 = n_4081 & ~n_4055;
assign n_4096 = n_4082 ^ x240;
assign n_4097 = n_4083 ^ n_1930;
assign n_4098 = n_4083 & ~n_4071;
assign n_4099 = ~n_3335 & ~n_4084;
assign n_4100 = n_4084 ^ n_3256;
assign n_4101 = n_4085 ^ n_2922;
assign n_4102 = n_4088 ^ n_4089;
assign n_4103 = n_4089 ^ x268;
assign n_4104 = n_4090 ^ n_2291;
assign n_4105 = n_4091 ^ n_2959;
assign n_4106 = n_4093 ^ n_3595;
assign n_4107 = n_4093 ^ n_4094;
assign n_4108 = n_4094 ^ n_3595;
assign n_4109 = n_4096 ^ n_4097;
assign n_4110 = n_4097 ^ x255;
assign n_4111 = n_4098 ^ n_1930;
assign n_4112 = n_4099 ^ n_2604;
assign n_4113 = n_4101 ^ n_2943;
assign n_4114 = n_4101 ^ n_3389;
assign n_4115 = n_4102 ^ x268;
assign n_4116 = n_4102 & ~n_4103;
assign n_4117 = n_4104 ^ n_2312;
assign n_4118 = n_4105 ^ n_2312;
assign n_4119 = n_4104 ^ n_4105;
assign n_4120 = n_4106 ^ n_4094;
assign n_4121 = ~n_4107 & n_4108;
assign n_4122 = n_4109 ^ x255;
assign n_4123 = n_4109 & ~n_4110;
assign n_4124 = n_4111 ^ n_1956;
assign n_4125 = n_4112 ^ n_1956;
assign n_4126 = n_4111 ^ n_4112;
assign n_4127 = n_4113 ^ n_3389;
assign n_4128 = n_3405 & n_4114;
assign n_4129 = ~n_4086 & n_4115;
assign n_4130 = n_4115 ^ n_4086;
assign n_4131 = n_4116 ^ x268;
assign n_4132 = n_4117 ^ n_4105;
assign n_4133 = n_4118 & ~n_4119;
assign n_4134 = ~n_3582 & ~n_4120;
assign n_4135 = n_3917 ^ n_4120;
assign n_4136 = n_4121 ^ n_3595;
assign n_4137 = n_4122 ^ n_4095;
assign n_4138 = ~n_4095 & n_4122;
assign n_4139 = n_4123 ^ x255;
assign n_4140 = n_4124 ^ n_4112;
assign n_4141 = n_4125 & ~n_4126;
assign n_4142 = n_4127 & n_3404;
assign n_4143 = n_3309 ^ n_4127;
assign n_4144 = n_4128 ^ n_2943;
assign n_4145 = n_4131 ^ n_4132;
assign n_4146 = n_4132 ^ x267;
assign n_4147 = n_4133 ^ n_2312;
assign n_4148 = n_4134 ^ n_2980;
assign n_4149 = n_4136 ^ n_3643;
assign n_4150 = n_4137 ^ n_3643;
assign n_4151 = n_4136 ^ n_4137;
assign n_4152 = n_4139 ^ n_4140;
assign n_4153 = n_4140 ^ x254;
assign n_4154 = n_4141 ^ n_1956;
assign n_4155 = n_4142 ^ n_2641;
assign n_4156 = n_4144 ^ n_3431;
assign n_4157 = n_4145 ^ x267;
assign n_4158 = ~n_4145 & n_4146;
assign n_4159 = n_4147 ^ n_2333;
assign n_4160 = n_4148 ^ n_2333;
assign n_4161 = n_4147 ^ n_4148;
assign n_4162 = n_4149 ^ n_4137;
assign n_4163 = ~n_4150 & n_4151;
assign n_4164 = n_4152 ^ x254;
assign n_4165 = ~n_4152 & n_4153;
assign n_4166 = n_4154 ^ n_4155;
assign n_4167 = n_4155 ^ n_1975;
assign n_4168 = n_2962 ^ n_4156;
assign n_4169 = ~n_4156 & n_3447;
assign n_4170 = n_4129 & ~n_4157;
assign n_4171 = n_4157 ^ n_4129;
assign n_4172 = n_4158 ^ x267;
assign n_4173 = n_4159 ^ n_4148;
assign n_4174 = ~n_4160 & ~n_4161;
assign n_4175 = ~n_3627 & n_4162;
assign n_4176 = n_3959 ^ n_4162;
assign n_4177 = n_4163 ^ n_3643;
assign n_4178 = n_4164 ^ n_4138;
assign n_4179 = ~n_4138 & n_4164;
assign n_4180 = n_4165 ^ x254;
assign n_4181 = n_4166 ^ n_1975;
assign n_4182 = n_4166 & ~n_4167;
assign n_4183 = ~n_4168 & n_3446;
assign n_4184 = n_4168 ^ n_3431;
assign n_4185 = n_3351 ^ n_4168;
assign n_4186 = n_4169 ^ n_2962;
assign n_4187 = n_4172 ^ n_4173;
assign n_4188 = n_4173 ^ x266;
assign n_4189 = n_4174 ^ n_2333;
assign n_4190 = n_4175 ^ n_2999;
assign n_4191 = n_4177 ^ n_3684;
assign n_4192 = n_4178 ^ n_3684;
assign n_4193 = n_4177 ^ n_4178;
assign n_4194 = n_4180 ^ n_4181;
assign n_4195 = n_4181 ^ x253;
assign n_4196 = n_4182 ^ n_1975;
assign n_4197 = n_4183 ^ n_2678;
assign n_4198 = n_4186 ^ n_3473;
assign n_4199 = n_4187 ^ x266;
assign n_4200 = n_4187 & ~n_4188;
assign n_4201 = n_4189 ^ n_2355;
assign n_4202 = n_4190 ^ n_2355;
assign n_4203 = n_4189 ^ n_4190;
assign n_4204 = n_4191 ^ n_4178;
assign n_4205 = n_4192 & ~n_4193;
assign n_4206 = n_4194 ^ x253;
assign n_4207 = n_4194 & ~n_4195;
assign n_4208 = n_4196 ^ n_1995;
assign n_4209 = n_4197 ^ n_1995;
assign n_4210 = n_4196 ^ n_4197;
assign n_4211 = n_2983 ^ n_4198;
assign n_4212 = n_4198 & n_3489;
assign n_4213 = ~n_4170 & ~n_4199;
assign n_4214 = n_4199 ^ n_4170;
assign n_4215 = n_4200 ^ x266;
assign n_4216 = n_4201 ^ n_4190;
assign n_4217 = n_4202 & n_4203;
assign n_4218 = ~n_3672 & ~n_4204;
assign n_4219 = n_4002 ^ n_4204;
assign n_4220 = n_4205 ^ n_3684;
assign n_4221 = n_4179 ^ n_4206;
assign n_4222 = n_4206 & ~n_4179;
assign n_4223 = n_4207 ^ x253;
assign n_4224 = n_4208 ^ n_4197;
assign n_4225 = n_4209 & n_4210;
assign n_4226 = ~n_4211 & n_3488;
assign n_4227 = n_4211 ^ n_3473;
assign n_4228 = n_3392 ^ n_4211;
assign n_4229 = n_4212 ^ n_2983;
assign n_4230 = n_4215 ^ n_4216;
assign n_4231 = n_4216 ^ x265;
assign n_4232 = n_4217 ^ n_2355;
assign n_4233 = n_4218 ^ n_3019;
assign n_4234 = n_4220 ^ n_3720;
assign n_4235 = n_4221 ^ n_3720;
assign n_4236 = n_4220 ^ n_4221;
assign n_4237 = n_4223 ^ n_4224;
assign n_4238 = n_4224 ^ x252;
assign n_4239 = n_4225 ^ n_1995;
assign n_4240 = n_4226 ^ n_2718;
assign n_4241 = n_4229 ^ n_3515;
assign n_4242 = n_4230 ^ x265;
assign n_4243 = n_4230 & ~n_4231;
assign n_4244 = n_4232 ^ n_2376;
assign n_4245 = n_4233 ^ n_2376;
assign n_4246 = n_4232 ^ n_4233;
assign n_4247 = n_4234 ^ n_4221;
assign n_4248 = ~n_4235 & n_4236;
assign n_4249 = n_4237 ^ x252;
assign n_4250 = ~n_4237 & n_4238;
assign n_4251 = n_4239 ^ n_2017;
assign n_4252 = n_4240 ^ n_2017;
assign n_4253 = n_4239 ^ n_4240;
assign n_4254 = n_4241 ^ n_3002;
assign n_4255 = n_4241 & ~n_3530;
assign n_4256 = n_4213 & ~n_4242;
assign n_4257 = n_4242 ^ n_4213;
assign n_4258 = n_4243 ^ x265;
assign n_4259 = n_4244 ^ n_4233;
assign n_4260 = n_4245 & ~n_4246;
assign n_4261 = n_3709 & n_4247;
assign n_4262 = n_4047 ^ n_4247;
assign n_4263 = n_4248 ^ n_3720;
assign n_4264 = n_4222 ^ n_4249;
assign n_4265 = ~n_4249 & n_4222;
assign n_4266 = n_4250 ^ x252;
assign n_4267 = n_4251 ^ n_4240;
assign n_4268 = ~n_4252 & n_4253;
assign n_4269 = ~n_4254 & ~n_3529;
assign n_4270 = n_4254 ^ n_3515;
assign n_4271 = n_3434 ^ n_4254;
assign n_4272 = n_4255 ^ n_3002;
assign n_4273 = n_4258 ^ n_4259;
assign n_4274 = n_4259 ^ x264;
assign n_4275 = n_4260 ^ n_2376;
assign n_4276 = n_4261 ^ n_3033;
assign n_4277 = n_4263 ^ n_3745;
assign n_4278 = n_4264 ^ n_3745;
assign n_4279 = n_4263 ^ n_4264;
assign n_4280 = n_4266 ^ n_4267;
assign n_4281 = n_4267 ^ x251;
assign n_4282 = n_4268 ^ n_2017;
assign n_4283 = n_4269 ^ n_2761;
assign n_4284 = n_4272 ^ n_3556;
assign n_4285 = n_4273 ^ x264;
assign n_4286 = ~n_4273 & n_4274;
assign n_4287 = n_4275 ^ n_4276;
assign n_4288 = n_4276 ^ n_2392;
assign n_4289 = n_4277 ^ n_4264;
assign n_4290 = ~n_4278 & n_4279;
assign n_4291 = n_4280 ^ x251;
assign n_4292 = ~n_4280 & n_4281;
assign n_4293 = n_4282 ^ n_2044;
assign n_4294 = n_4283 ^ n_2044;
assign n_4295 = n_4282 ^ n_4283;
assign n_4296 = n_4284 ^ n_3022;
assign n_4297 = ~n_4284 & n_3572;
assign n_4298 = ~n_4256 & ~n_4285;
assign n_4299 = n_4285 ^ n_4256;
assign n_4300 = n_4286 ^ x264;
assign n_4301 = n_4287 ^ n_2392;
assign n_4302 = n_4287 & n_4288;
assign n_4303 = ~n_3746 & n_4289;
assign n_4304 = n_4087 ^ n_4289;
assign n_4305 = n_4290 ^ n_3745;
assign n_4306 = n_4291 ^ n_4265;
assign n_4307 = n_4265 & ~n_4291;
assign n_4308 = n_4292 ^ x251;
assign n_4309 = n_4293 ^ n_4283;
assign n_4310 = ~n_4294 & n_4295;
assign n_4311 = n_4296 & ~n_3571;
assign n_4312 = n_4296 ^ n_3556;
assign n_4313 = n_3476 ^ n_4296;
assign n_4314 = n_4297 ^ n_3022;
assign n_4315 = n_4300 ^ n_4301;
assign n_4316 = n_4301 ^ x279;
assign n_4317 = n_4302 ^ n_2392;
assign n_4318 = n_4303 ^ n_3059;
assign n_4319 = n_4305 ^ n_3793;
assign n_4320 = n_4306 ^ n_3793;
assign n_4321 = n_4305 ^ n_4306;
assign n_4322 = n_4308 ^ n_4309;
assign n_4323 = n_4309 ^ x250;
assign n_4324 = n_4310 ^ n_2044;
assign n_4325 = n_4311 ^ n_2803;
assign n_4326 = n_4314 ^ n_3587;
assign n_4327 = n_4315 ^ x279;
assign n_4328 = ~n_4315 & n_4316;
assign n_4329 = n_4317 ^ n_2419;
assign n_4330 = n_4318 ^ n_2419;
assign n_4331 = n_4317 ^ n_4318;
assign n_4332 = n_4319 ^ n_4306;
assign n_4333 = n_4320 & n_4321;
assign n_4334 = n_4322 ^ x250;
assign n_4335 = ~n_4322 & n_4323;
assign n_4336 = n_4324 ^ n_2077;
assign n_4337 = n_4325 ^ n_2077;
assign n_4338 = n_4325 ^ n_4324;
assign n_4339 = n_4326 ^ n_3044;
assign n_4340 = ~n_4298 & n_4327;
assign n_4341 = n_4327 ^ n_4298;
assign n_4342 = n_4328 ^ x279;
assign n_4343 = n_4329 ^ n_4318;
assign n_4344 = n_4330 & n_4331;
assign n_4345 = ~n_4332 & n_3806;
assign n_4346 = n_4130 ^ n_4332;
assign n_4347 = n_4333 ^ n_3793;
assign n_4348 = n_4334 ^ n_4307;
assign n_4349 = n_4307 & ~n_4334;
assign n_4350 = n_4335 ^ x250;
assign n_4351 = n_4325 ^ n_4336;
assign n_4352 = n_4337 & ~n_4338;
assign n_4353 = n_4339 & ~n_3602;
assign n_4354 = n_4339 ^ n_3503;
assign n_4355 = n_4339 ^ n_3587;
assign n_4356 = n_4342 ^ n_4343;
assign n_4357 = n_4343 ^ x278;
assign n_4358 = n_4344 ^ n_2419;
assign n_4359 = n_4345 ^ n_3083;
assign n_4360 = n_4347 ^ n_3831;
assign n_4361 = n_4348 ^ n_3831;
assign n_4362 = n_4347 ^ n_4348;
assign n_4363 = n_4350 ^ n_4351;
assign n_4364 = n_4351 ^ x249;
assign n_4365 = n_4352 ^ n_2077;
assign n_4366 = n_4353 ^ n_2833;
assign n_4367 = n_4354 ^ n_3475;
assign n_4368 = n_4356 ^ x278;
assign n_4369 = n_4356 & ~n_4357;
assign n_4370 = n_4358 ^ n_2438;
assign n_4371 = n_4359 ^ n_2438;
assign n_4372 = n_4358 ^ n_4359;
assign n_4373 = n_4360 ^ n_4348;
assign n_4374 = ~n_4361 & ~n_4362;
assign n_4375 = n_4363 ^ x249;
assign n_4376 = n_4363 & ~n_4364;
assign n_4377 = n_4366 ^ n_2101;
assign n_4378 = n_4340 & ~n_4368;
assign n_4379 = n_4368 ^ n_4340;
assign n_4380 = n_4369 ^ x278;
assign n_4381 = n_4370 ^ n_4359;
assign n_4382 = ~n_4371 & ~n_4372;
assign n_4383 = ~n_4373 & n_3846;
assign n_4384 = n_4171 ^ n_4373;
assign n_4385 = n_4374 ^ n_3831;
assign n_4386 = n_4349 ^ n_4375;
assign n_4387 = n_4375 & n_4349;
assign n_4388 = n_4376 ^ x249;
assign n_4389 = n_4377 ^ x248;
assign n_4390 = n_4380 ^ n_4381;
assign n_4391 = n_4381 ^ x277;
assign n_4392 = n_4382 ^ n_2438;
assign n_4393 = n_4383 ^ n_3113;
assign n_4394 = n_4385 ^ n_3873;
assign n_4395 = n_4385 ^ n_4386;
assign n_4396 = n_4386 ^ n_3873;
assign n_4397 = n_4365 ^ n_4389;
assign n_4398 = n_4390 ^ x277;
assign n_4399 = n_4390 & ~n_4391;
assign n_4400 = n_4392 ^ n_2459;
assign n_4401 = n_4393 ^ n_2459;
assign n_4402 = n_4392 ^ n_4393;
assign n_4403 = n_4394 ^ n_4386;
assign n_4404 = ~n_4395 & ~n_4396;
assign n_4405 = n_4388 ^ n_4397;
assign n_4406 = ~n_4398 & n_4378;
assign n_4407 = n_4378 ^ n_4398;
assign n_4408 = n_4399 ^ x277;
assign n_4409 = n_4400 ^ n_4393;
assign n_4410 = ~n_4401 & ~n_4402;
assign n_4411 = n_3859 & n_4403;
assign n_4412 = n_4214 ^ n_4403;
assign n_4413 = n_4404 ^ n_3873;
assign n_4414 = n_4405 ^ n_4387;
assign n_4415 = n_4408 ^ n_4409;
assign n_4416 = n_4409 ^ x276;
assign n_4417 = n_4410 ^ n_2459;
assign n_4418 = n_4411 ^ n_3147;
assign n_4419 = n_4413 ^ n_3914;
assign n_4420 = n_4413 ^ n_4414;
assign n_4421 = n_4414 ^ n_3914;
assign n_4422 = n_4415 ^ x276;
assign n_4423 = ~n_4415 & n_4416;
assign n_4424 = n_4417 ^ n_2479;
assign n_4425 = n_4418 ^ n_4417;
assign n_4426 = n_4419 ^ n_4414;
assign n_4427 = n_4420 & n_4421;
assign n_4428 = n_4406 & n_4422;
assign n_4429 = n_4422 ^ n_4406;
assign n_4430 = n_4423 ^ x276;
assign n_4431 = n_4418 ^ n_4424;
assign n_4432 = ~n_4424 & ~n_4425;
assign n_4433 = n_4426 & ~n_3930;
assign n_4434 = n_4257 ^ n_4426;
assign n_4435 = n_4427 ^ n_3914;
assign n_4436 = n_4430 ^ n_4431;
assign n_4437 = n_4431 ^ x275;
assign n_4438 = n_4432 ^ n_2479;
assign n_4439 = n_4433 ^ n_3185;
assign n_4440 = n_4435 ^ n_3972;
assign n_4441 = n_4435 ^ n_3956;
assign n_4442 = n_4436 ^ x275;
assign n_4443 = n_4436 & ~n_4437;
assign n_4444 = n_4438 ^ n_2500;
assign n_4445 = n_4439 ^ n_2500;
assign n_4446 = n_4438 ^ n_4439;
assign n_4447 = n_4440 & n_3973;
assign n_4448 = n_4440 ^ n_3956;
assign n_4449 = n_4299 ^ n_4440;
assign n_4450 = ~n_3972 & ~n_4441;
assign n_4451 = n_4428 & ~n_4442;
assign n_4452 = n_4442 ^ n_4428;
assign n_4453 = n_4443 ^ x275;
assign n_4454 = n_4444 ^ n_4439;
assign n_4455 = ~n_4445 & n_4446;
assign n_4456 = n_4447 ^ n_3225;
assign n_4457 = n_4450 ^ n_3105;
assign n_4458 = n_4453 ^ n_4454;
assign n_4459 = n_4454 ^ x274;
assign n_4460 = n_4455 ^ n_2500;
assign n_4461 = n_4457 ^ n_3999;
assign n_4462 = n_4458 ^ x274;
assign n_4463 = ~n_4458 & n_4459;
assign n_4464 = n_4460 ^ n_2520;
assign n_4465 = n_4456 ^ n_4460;
assign n_4466 = n_3153 ^ n_4461;
assign n_4467 = n_4461 & n_4016;
assign n_4468 = n_4451 & n_4462;
assign n_4469 = n_4462 ^ n_4451;
assign n_4470 = n_4463 ^ x274;
assign n_4471 = n_4456 ^ n_4464;
assign n_4472 = n_4464 & ~n_4465;
assign n_4473 = n_4466 & ~n_4015;
assign n_4474 = n_4466 ^ n_3999;
assign n_4475 = n_4341 ^ n_4466;
assign n_4476 = n_4467 ^ n_3153;
assign n_4477 = n_4470 ^ x273;
assign n_4478 = n_4470 ^ n_4471;
assign n_4479 = n_4472 ^ n_2520;
assign n_4480 = n_4473 ^ n_3267;
assign n_4481 = n_4476 ^ n_4029;
assign n_4482 = n_4478 ^ x273;
assign n_4483 = n_4478 & n_4477;
assign n_4484 = n_4479 ^ n_2543;
assign n_4485 = n_4480 ^ n_2543;
assign n_4486 = n_4479 ^ n_4480;
assign n_4487 = n_3214 ^ n_4481;
assign n_4488 = ~n_4481 & ~n_4044;
assign n_4489 = n_4468 & ~n_4482;
assign n_4490 = n_4482 ^ n_4468;
assign n_4491 = n_4483 ^ x273;
assign n_4492 = n_4484 ^ n_4480;
assign n_4493 = n_4485 & n_4486;
assign n_4494 = n_4487 & n_4043;
assign n_4495 = n_4487 ^ n_4029;
assign n_4496 = n_4379 ^ n_4487;
assign n_4497 = n_4488 ^ n_3214;
assign n_4498 = n_4491 ^ x272;
assign n_4499 = n_4491 ^ n_4492;
assign n_4500 = n_4493 ^ n_2543;
assign n_4501 = n_4494 ^ n_3306;
assign n_4502 = n_4497 ^ n_3256;
assign n_4503 = n_4497 ^ n_4084;
assign n_4504 = n_4499 ^ x272;
assign n_4505 = n_4499 & n_4498;
assign n_4506 = n_4500 ^ n_4501;
assign n_4507 = n_4501 ^ n_2571;
assign n_4508 = n_4502 ^ n_4084;
assign n_4509 = ~n_4100 & n_4503;
assign n_4510 = ~n_4489 & n_4504;
assign n_4511 = n_4504 ^ n_4489;
assign n_4512 = n_4505 ^ x272;
assign n_4513 = n_4506 ^ n_2571;
assign n_4514 = n_4506 & n_4507;
assign n_4515 = n_4072 & ~n_4508;
assign n_4516 = n_4508 ^ n_4407;
assign n_4517 = n_4509 ^ n_3256;
assign n_4518 = n_4512 ^ n_4513;
assign n_4519 = n_4513 ^ x287;
assign n_4520 = n_4514 ^ n_2571;
assign n_4521 = n_4515 ^ n_3348;
assign n_4522 = n_4517 ^ n_4127;
assign n_4523 = n_4518 ^ x287;
assign n_4524 = ~n_4518 & n_4519;
assign n_4525 = n_4520 ^ n_2604;
assign n_4526 = n_4521 ^ n_2604;
assign n_4527 = n_4520 ^ n_4521;
assign n_4528 = n_3309 ^ n_4522;
assign n_4529 = ~n_4522 & n_4143;
assign n_4530 = n_4510 & ~n_4523;
assign n_4531 = n_4523 ^ n_4510;
assign n_4532 = n_4524 ^ x287;
assign n_4533 = n_4525 ^ n_4521;
assign n_4534 = ~n_4526 & ~n_4527;
assign n_4535 = ~n_4113 & n_4528;
assign n_4536 = n_4528 ^ n_4127;
assign n_4537 = n_4429 ^ n_4528;
assign n_4538 = n_4529 ^ n_3309;
assign n_4539 = n_4532 ^ x286;
assign n_4540 = n_4533 ^ x286;
assign n_4541 = n_4532 ^ n_4533;
assign n_4542 = n_4534 ^ n_2604;
assign n_4543 = n_4535 ^ n_3389;
assign n_4544 = n_4538 ^ n_3351;
assign n_4545 = n_4538 ^ n_4168;
assign n_4546 = n_4539 ^ n_4533;
assign n_4547 = n_4540 & ~n_4541;
assign n_4548 = n_4542 ^ n_2641;
assign n_4549 = n_4543 ^ n_2641;
assign n_4550 = n_4542 ^ n_4543;
assign n_4551 = n_4544 ^ n_4168;
assign n_4552 = n_4185 & n_4545;
assign n_4553 = ~n_4530 & n_4546;
assign n_4554 = n_4546 ^ n_4530;
assign n_4555 = n_4547 ^ x286;
assign n_4556 = n_4548 ^ n_4543;
assign n_4557 = n_4549 & n_4550;
assign n_4558 = n_4551 & n_4184;
assign n_4559 = n_4452 ^ n_4551;
assign n_4560 = n_4552 ^ n_3351;
assign n_4561 = ~n_3574 & ~n_4554;
assign n_4562 = n_4554 ^ n_3574;
assign n_4563 = n_4555 ^ x285;
assign n_4564 = n_4556 ^ x285;
assign n_4565 = n_4555 ^ n_4556;
assign n_4566 = n_4557 ^ n_2641;
assign n_4567 = n_4558 ^ n_3431;
assign n_4568 = n_4560 ^ n_4211;
assign n_4569 = n_4561 ^ n_3619;
assign n_4570 = n_3558 & n_4562;
assign n_4571 = n_4563 ^ n_4556;
assign n_4572 = n_4564 & ~n_4565;
assign n_4573 = n_4566 ^ n_2678;
assign n_4574 = n_4567 ^ n_2678;
assign n_4575 = n_4566 ^ n_4567;
assign n_4576 = n_3392 ^ n_4568;
assign n_4577 = ~n_4568 & n_4228;
assign n_4578 = n_4570 ^ n_3070;
assign n_4579 = n_4553 ^ n_4571;
assign n_4580 = n_4571 & n_4553;
assign n_4581 = n_4572 ^ x285;
assign n_4582 = n_4573 ^ n_4567;
assign n_4583 = n_4574 & ~n_4575;
assign n_4584 = ~n_4576 & ~n_4227;
assign n_4585 = n_4576 ^ n_4211;
assign n_4586 = n_4469 ^ n_4576;
assign n_4587 = n_4577 ^ n_3392;
assign n_4588 = n_2538 & ~n_4578;
assign n_4589 = n_4578 ^ n_2538;
assign n_4590 = n_4579 ^ n_4561;
assign n_4591 = n_4569 ^ n_4579;
assign n_4592 = n_4581 ^ n_4582;
assign n_4593 = n_4582 ^ x284;
assign n_4594 = n_4583 ^ n_2678;
assign n_4595 = n_4584 ^ n_3473;
assign n_4596 = n_4587 ^ n_3434;
assign n_4597 = n_4587 ^ n_4254;
assign n_4598 = n_4588 ^ n_2567;
assign n_4599 = x295 & ~n_4589;
assign n_4600 = n_4589 ^ x295;
assign n_4601 = ~n_4590 & n_4569;
assign n_4602 = ~n_3620 & n_4591;
assign n_4603 = n_4592 ^ x284;
assign n_4604 = n_4592 & ~n_4593;
assign n_4605 = n_4594 ^ n_2718;
assign n_4606 = n_4595 ^ n_2718;
assign n_4607 = n_4594 ^ n_4595;
assign n_4608 = n_4596 ^ n_4254;
assign n_4609 = ~n_4271 & ~n_4597;
assign n_4610 = n_4599 ^ x294;
assign n_4611 = n_4601 ^ n_3619;
assign n_4612 = n_4602 ^ n_3097;
assign n_4613 = n_4603 & ~n_4580;
assign n_4614 = n_4580 ^ n_4603;
assign n_4615 = n_4604 ^ x284;
assign n_4616 = n_4605 ^ n_4595;
assign n_4617 = n_4606 & n_4607;
assign n_4618 = n_4608 & n_4270;
assign n_4619 = n_4490 ^ n_4608;
assign n_4620 = n_4609 ^ n_3434;
assign n_4621 = n_4611 ^ n_3677;
assign n_4622 = n_4612 ^ n_4588;
assign n_4623 = n_4612 ^ n_4598;
assign n_4624 = n_4614 ^ n_4611;
assign n_4625 = n_4615 ^ n_4616;
assign n_4626 = n_4616 ^ x283;
assign n_4627 = n_4617 ^ n_2718;
assign n_4628 = n_4618 ^ n_3515;
assign n_4629 = n_4620 ^ n_4296;
assign n_4630 = n_4614 ^ n_4621;
assign n_4631 = n_4598 & n_4622;
assign n_4632 = n_4623 ^ n_4599;
assign n_4633 = n_4623 ^ n_4610;
assign n_4634 = n_4621 & ~n_4624;
assign n_4635 = n_4625 ^ x283;
assign n_4636 = n_4625 & ~n_4626;
assign n_4637 = n_4627 ^ n_2761;
assign n_4638 = n_4628 ^ n_2761;
assign n_4639 = n_4627 ^ n_4628;
assign n_4640 = n_4629 ^ n_3476;
assign n_4641 = ~n_4629 & ~n_4313;
assign n_4642 = ~n_3664 & n_4630;
assign n_4643 = n_4631 ^ n_2567;
assign n_4644 = n_4610 & n_4632;
assign n_4645 = n_4600 & n_4633;
assign n_4646 = n_4633 ^ n_4600;
assign n_4647 = n_4634 ^ n_3677;
assign n_4648 = ~n_4635 & ~n_4613;
assign n_4649 = n_4613 ^ n_4635;
assign n_4650 = n_4636 ^ x283;
assign n_4651 = n_4637 ^ n_4628;
assign n_4652 = ~n_4638 & n_4639;
assign n_4653 = ~n_4640 & n_4312;
assign n_4654 = n_4640 ^ n_4296;
assign n_4655 = n_4511 ^ n_4640;
assign n_4656 = n_4641 ^ n_3476;
assign n_4657 = n_4642 ^ n_3137;
assign n_4658 = n_4644 ^ x294;
assign n_4659 = n_4647 ^ n_3713;
assign n_4660 = n_4649 ^ n_3713;
assign n_4661 = n_4647 ^ n_4649;
assign n_4662 = n_4650 ^ n_4651;
assign n_4663 = n_4651 ^ x282;
assign n_4664 = n_4652 ^ n_2761;
assign n_4665 = n_4653 ^ n_3556;
assign n_4666 = n_4656 ^ n_4367;
assign n_4667 = n_4643 ^ n_4657;
assign n_4668 = n_4657 ^ n_2610;
assign n_4669 = n_4659 ^ n_4649;
assign n_4670 = ~n_4660 & ~n_4661;
assign n_4671 = n_4662 ^ x282;
assign n_4672 = n_4662 & ~n_4663;
assign n_4673 = n_4664 ^ n_2803;
assign n_4674 = n_4665 ^ n_2803;
assign n_4675 = n_4665 ^ n_4664;
assign n_4676 = ~n_4666 & n_4355;
assign n_4677 = n_4531 ^ n_4666;
assign n_4678 = n_4666 ^ n_4339;
assign n_4679 = n_4667 ^ n_2610;
assign n_4680 = n_4667 & ~n_4668;
assign n_4681 = n_3703 & ~n_4669;
assign n_4682 = n_4670 ^ n_3713;
assign n_4683 = n_4671 & ~n_4648;
assign n_4684 = n_4648 ^ n_4671;
assign n_4685 = n_4672 ^ x282;
assign n_4686 = n_4665 ^ n_4673;
assign n_4687 = ~n_4674 & ~n_4675;
assign n_4688 = n_4676 ^ n_3587;
assign n_4689 = n_4658 ^ n_4679;
assign n_4690 = n_4679 ^ x293;
assign n_4691 = n_4680 ^ n_2610;
assign n_4692 = n_4681 ^ n_3178;
assign n_4693 = n_4682 ^ n_3751;
assign n_4694 = n_4684 ^ n_3751;
assign n_4695 = n_4682 ^ n_4684;
assign n_4696 = n_4685 ^ n_4686;
assign n_4697 = n_4686 ^ x281;
assign n_4698 = n_4687 ^ n_2803;
assign n_4699 = n_4688 ^ n_2833;
assign n_4700 = n_4689 ^ x293;
assign n_4701 = n_4689 & ~n_4690;
assign n_4702 = n_4691 ^ n_2647;
assign n_4703 = n_4692 ^ n_2647;
assign n_4704 = n_4691 ^ n_4692;
assign n_4705 = n_4693 ^ n_4684;
assign n_4706 = ~n_4694 & n_4695;
assign n_4707 = n_4696 ^ x281;
assign n_4708 = n_4696 & ~n_4697;
assign n_4709 = n_4698 ^ x280;
assign n_4710 = n_4700 & n_4645;
assign n_4711 = n_4645 ^ n_4700;
assign n_4712 = n_4701 ^ x293;
assign n_4713 = n_4702 ^ n_4692;
assign n_4714 = ~n_4703 & n_4704;
assign n_4715 = n_3740 & n_4705;
assign n_4716 = n_4706 ^ n_3751;
assign n_4717 = n_4707 & n_4683;
assign n_4718 = n_4683 ^ n_4707;
assign n_4719 = n_4708 ^ x281;
assign n_4720 = n_4709 ^ n_4699;
assign n_4721 = n_4712 ^ n_4713;
assign n_4722 = n_4713 ^ x292;
assign n_4723 = n_4714 ^ n_2647;
assign n_4724 = n_4715 ^ n_3218;
assign n_4725 = n_4716 ^ n_3787;
assign n_4726 = n_4718 ^ n_3787;
assign n_4727 = n_4716 ^ n_4718;
assign n_4728 = n_4719 ^ n_4720;
assign n_4729 = n_4721 ^ x292;
assign n_4730 = n_4721 & ~n_4722;
assign n_4731 = n_4723 ^ n_2688;
assign n_4732 = n_4724 ^ n_4723;
assign n_4733 = n_4725 ^ n_4718;
assign n_4734 = ~n_4726 & ~n_4727;
assign n_4735 = n_4728 ^ n_4717;
assign n_4736 = n_4710 & n_4729;
assign n_4737 = n_4729 ^ n_4710;
assign n_4738 = n_4730 ^ x292;
assign n_4739 = n_4724 ^ n_4731;
assign n_4740 = ~n_4731 & n_4732;
assign n_4741 = n_3776 & n_4733;
assign n_4742 = n_4734 ^ n_3787;
assign n_4743 = n_4735 ^ n_3824;
assign n_4744 = n_4738 ^ n_4739;
assign n_4745 = n_4739 ^ x291;
assign n_4746 = n_4740 ^ n_2688;
assign n_4747 = n_4741 ^ n_3260;
assign n_4748 = n_4742 ^ n_4735;
assign n_4749 = n_4742 ^ n_3824;
assign n_4750 = n_4744 ^ x291;
assign n_4751 = ~n_4744 & n_4745;
assign n_4752 = n_4746 ^ n_2727;
assign n_4753 = n_4747 ^ n_2727;
assign n_4754 = n_4746 ^ n_4747;
assign n_4755 = n_4743 & n_4748;
assign n_4756 = n_4749 ^ n_4735;
assign n_4757 = ~n_4736 & n_4750;
assign n_4758 = n_4750 ^ n_4736;
assign n_4759 = n_4751 ^ x291;
assign n_4760 = n_4752 ^ n_4747;
assign n_4761 = n_4753 & n_4754;
assign n_4762 = n_4755 ^ n_3824;
assign n_4763 = ~n_3814 & n_4756;
assign n_4764 = n_4759 ^ n_4760;
assign n_4765 = n_4760 ^ x290;
assign n_4766 = n_4761 ^ n_2727;
assign n_4767 = n_4762 ^ n_3866;
assign n_4768 = n_4763 ^ n_3299;
assign n_4769 = n_4764 ^ x290;
assign n_4770 = n_4764 & ~n_4765;
assign n_4771 = n_4766 ^ n_2770;
assign n_4772 = n_4767 & n_3881;
assign n_4773 = n_3634 ^ n_4767;
assign n_4774 = n_4768 ^ n_2770;
assign n_4775 = n_4766 ^ n_4768;
assign n_4776 = n_4769 & ~n_4757;
assign n_4777 = n_4757 ^ n_4769;
assign n_4778 = n_4770 ^ x290;
assign n_4779 = n_4771 ^ n_4768;
assign n_4780 = n_4772 ^ n_3634;
assign n_4781 = ~n_3854 & ~n_4773;
assign n_4782 = n_4773 ^ n_3866;
assign n_4783 = ~n_4774 & ~n_4775;
assign n_4784 = n_4778 ^ n_4779;
assign n_4785 = n_4779 ^ x289;
assign n_4786 = n_4780 ^ n_3907;
assign n_4787 = n_4781 ^ n_3342;
assign n_4788 = n_4783 ^ n_2770;
assign n_4789 = n_4784 ^ x289;
assign n_4790 = n_4784 & ~n_4785;
assign n_4791 = n_4786 & ~n_3922;
assign n_4792 = n_3675 ^ n_4786;
assign n_4793 = n_4787 ^ n_2812;
assign n_4794 = n_4788 ^ n_4787;
assign n_4795 = n_4788 ^ n_2812;
assign n_4796 = ~n_4776 & ~n_4789;
assign n_4797 = n_4789 ^ n_4776;
assign n_4798 = n_4790 ^ x289;
assign n_4799 = n_4791 ^ n_3675;
assign n_4800 = ~n_3896 & ~n_4792;
assign n_4801 = n_4792 ^ n_3907;
assign n_4802 = n_4793 & ~n_4794;
assign n_4803 = n_4795 ^ n_4787;
assign n_4804 = n_4799 ^ n_3949;
assign n_4805 = n_4800 ^ n_3382;
assign n_4806 = n_4802 ^ n_2812;
assign n_4807 = n_4798 ^ n_4803;
assign n_4808 = n_4803 ^ x288;
assign n_4809 = n_4804 & n_3964;
assign n_4810 = n_3734 ^ n_4804;
assign n_4811 = n_4805 ^ n_2855;
assign n_4812 = n_4806 ^ n_4805;
assign n_4813 = n_4806 ^ n_2855;
assign n_4814 = n_4807 ^ x288;
assign n_4815 = n_4807 & ~n_4808;
assign n_4816 = n_4809 ^ n_3734;
assign n_4817 = ~n_3938 & n_4810;
assign n_4818 = n_4810 ^ n_3949;
assign n_4819 = ~n_4811 & n_4812;
assign n_4820 = n_4813 ^ n_4805;
assign n_4821 = ~n_4796 & n_4814;
assign n_4822 = n_4814 ^ n_4796;
assign n_4823 = n_4815 ^ x288;
assign n_4824 = n_4816 ^ n_3992;
assign n_4825 = n_4816 ^ n_4007;
assign n_4826 = n_4817 ^ n_3424;
assign n_4827 = n_4819 ^ n_2855;
assign n_4828 = n_4820 ^ x303;
assign n_4829 = n_4823 ^ n_4820;
assign n_4830 = n_4007 & ~n_4824;
assign n_4831 = n_3981 & ~n_4825;
assign n_4832 = n_4825 ^ n_3992;
assign n_4833 = n_4826 ^ n_2890;
assign n_4834 = n_4827 ^ n_4826;
assign n_4835 = n_4827 ^ n_2890;
assign n_4836 = ~n_4829 & n_4828;
assign n_4837 = n_4829 ^ x303;
assign n_4838 = n_4830 ^ n_3782;
assign n_4839 = n_4831 ^ n_3466;
assign n_4840 = n_4833 & n_4834;
assign n_4841 = n_4835 ^ n_4826;
assign n_4842 = n_4836 ^ x303;
assign n_4843 = n_4821 & ~n_4837;
assign n_4844 = n_4837 ^ n_4821;
assign n_4845 = n_4838 ^ n_4035;
assign n_4846 = n_4840 ^ n_2890;
assign n_4847 = n_4841 ^ x302;
assign n_4848 = n_4842 ^ n_4841;
assign n_4849 = n_3834 ^ n_4845;
assign n_4850 = ~n_4845 & n_4052;
assign n_4851 = n_4846 ^ n_2918;
assign n_4852 = n_4839 ^ n_4846;
assign n_4853 = n_4848 & ~n_4847;
assign n_4854 = n_4848 ^ x302;
assign n_4855 = ~n_4024 & ~n_4849;
assign n_4856 = n_4849 ^ n_4035;
assign n_4857 = n_4850 ^ n_3834;
assign n_4858 = n_4839 ^ n_4851;
assign n_4859 = n_4851 & n_4852;
assign n_4860 = n_4853 ^ x302;
assign n_4861 = n_4843 & n_4854;
assign n_4862 = n_4854 ^ n_4843;
assign n_4863 = n_4855 ^ n_3508;
assign n_4864 = n_4857 ^ n_4079;
assign n_4865 = n_4858 ^ x301;
assign n_4866 = n_4859 ^ n_2918;
assign n_4867 = n_4860 ^ n_4858;
assign n_4868 = n_4863 ^ n_2940;
assign n_4869 = n_3876 ^ n_4864;
assign n_4870 = n_4864 & n_4092;
assign n_4871 = n_4866 ^ n_4863;
assign n_4872 = n_4866 ^ n_2940;
assign n_4873 = n_4867 & ~n_4865;
assign n_4874 = n_4867 ^ x301;
assign n_4875 = ~n_4067 & ~n_4869;
assign n_4876 = n_4600 ^ n_4869;
assign n_4877 = n_4869 ^ n_4079;
assign n_4878 = n_4870 ^ n_3876;
assign n_4879 = ~n_4868 & ~n_4871;
assign n_4880 = n_4872 ^ n_4863;
assign n_4881 = n_4873 ^ x301;
assign n_4882 = n_4861 & n_4874;
assign n_4883 = n_4874 ^ n_4861;
assign n_4884 = n_4875 ^ n_3550;
assign n_4885 = n_4878 ^ n_4120;
assign n_4886 = n_4879 ^ n_2940;
assign n_4887 = n_4881 ^ n_4880;
assign n_4888 = n_4881 ^ x300;
assign n_4889 = n_4884 ^ n_2959;
assign n_4890 = n_3917 ^ n_4885;
assign n_4891 = n_4885 & n_4135;
assign n_4892 = n_4886 ^ n_2959;
assign n_4893 = n_4886 ^ n_4884;
assign n_4894 = n_4887 ^ x300;
assign n_4895 = n_4887 & n_4888;
assign n_4896 = n_4107 & n_4890;
assign n_4897 = n_4890 ^ n_4120;
assign n_4898 = n_4646 ^ n_4890;
assign n_4899 = n_4891 ^ n_3917;
assign n_4900 = n_4892 ^ n_4884;
assign n_4901 = ~n_4889 & ~n_4893;
assign n_4902 = ~n_4882 & ~n_4894;
assign n_4903 = n_4894 ^ n_4882;
assign n_4904 = n_4895 ^ x300;
assign n_4905 = n_4896 ^ n_3595;
assign n_4906 = n_4899 ^ n_4162;
assign n_4907 = n_4900 ^ x299;
assign n_4908 = n_4901 ^ n_2959;
assign n_4909 = n_4904 ^ n_4900;
assign n_4910 = n_4904 ^ x299;
assign n_4911 = n_4905 ^ n_2980;
assign n_4912 = n_3959 ^ n_4906;
assign n_4913 = n_4906 & n_4176;
assign n_4914 = n_4908 ^ n_2980;
assign n_4915 = n_4908 ^ n_4905;
assign n_4916 = n_4907 & ~n_4909;
assign n_4917 = n_4910 ^ n_4900;
assign n_4918 = ~n_4151 & ~n_4912;
assign n_4919 = n_4912 ^ n_4162;
assign n_4920 = n_4711 ^ n_4912;
assign n_4921 = n_4913 ^ n_3959;
assign n_4922 = n_4914 ^ n_4905;
assign n_4923 = ~n_4911 & n_4915;
assign n_4924 = n_4916 ^ x299;
assign n_4925 = ~n_4902 & ~n_4917;
assign n_4926 = n_4917 ^ n_4902;
assign n_4927 = n_4918 ^ n_3643;
assign n_4928 = n_4921 ^ n_4204;
assign n_4929 = n_4922 ^ x298;
assign n_4930 = n_4923 ^ n_2980;
assign n_4931 = n_4924 ^ n_4922;
assign n_4932 = n_4927 ^ n_2999;
assign n_4933 = n_4002 ^ n_4928;
assign n_4934 = n_4928 & ~n_4219;
assign n_4935 = n_4930 ^ n_2999;
assign n_4936 = n_4930 ^ n_4927;
assign n_4937 = n_4931 & ~n_4929;
assign n_4938 = n_4931 ^ x298;
assign n_4939 = n_4193 & ~n_4933;
assign n_4940 = n_4933 ^ n_4204;
assign n_4941 = n_4737 ^ n_4933;
assign n_4942 = n_4934 ^ n_4002;
assign n_4943 = n_4935 ^ n_4927;
assign n_4944 = ~n_4932 & n_4936;
assign n_4945 = n_4937 ^ x298;
assign n_4946 = n_4938 & n_4925;
assign n_4947 = n_4925 ^ n_4938;
assign n_4948 = n_4939 ^ n_3684;
assign n_4949 = n_4942 ^ n_4247;
assign n_4950 = n_4943 ^ x297;
assign n_4951 = n_4944 ^ n_2999;
assign n_4952 = n_4945 ^ n_4943;
assign n_4953 = n_4948 ^ n_3019;
assign n_4954 = n_4047 ^ n_4949;
assign n_4955 = ~n_4949 & n_4262;
assign n_4956 = n_4951 ^ n_3019;
assign n_4957 = n_4951 ^ n_4948;
assign n_4958 = n_4952 & ~n_4950;
assign n_4959 = n_4952 ^ x297;
assign n_4960 = ~n_4236 & n_4954;
assign n_4961 = n_4954 ^ n_4247;
assign n_4962 = n_4758 ^ n_4954;
assign n_4963 = n_4955 ^ n_4047;
assign n_4964 = n_4956 ^ n_4948;
assign n_4965 = ~n_4953 & n_4957;
assign n_4966 = n_4958 ^ x297;
assign n_4967 = n_4946 & n_4959;
assign n_4968 = n_4959 ^ n_4946;
assign n_4969 = n_4960 ^ n_3720;
assign n_4970 = n_4963 ^ n_4087;
assign n_4971 = n_4963 ^ n_4289;
assign n_4972 = n_4964 ^ x296;
assign n_4973 = n_4965 ^ n_3019;
assign n_4974 = n_4966 ^ n_4964;
assign n_4975 = n_4969 ^ n_3033;
assign n_4976 = n_4970 ^ n_4289;
assign n_4977 = ~n_4304 & ~n_4971;
assign n_4978 = n_4973 ^ n_3033;
assign n_4979 = n_4973 ^ n_4969;
assign n_4980 = n_4974 & ~n_4972;
assign n_4981 = n_4974 ^ x296;
assign n_4982 = ~n_4279 & ~n_4976;
assign n_4983 = n_4777 ^ n_4976;
assign n_4984 = n_4977 ^ n_4087;
assign n_4985 = n_4978 ^ n_4969;
assign n_4986 = n_4975 & n_4979;
assign n_4987 = n_4980 ^ x296;
assign n_4988 = n_4981 & n_4967;
assign n_4989 = n_4967 ^ n_4981;
assign n_4990 = n_4982 ^ n_3745;
assign n_4991 = n_4984 ^ n_4332;
assign n_4992 = n_4985 ^ x311;
assign n_4993 = n_4986 ^ n_3033;
assign n_4994 = n_4987 ^ n_4985;
assign n_4995 = n_4990 ^ n_3059;
assign n_4996 = n_4130 ^ n_4991;
assign n_4997 = ~n_4991 & ~n_4346;
assign n_4998 = n_4993 ^ n_4990;
assign n_4999 = ~n_4994 & n_4992;
assign n_5000 = n_4994 ^ x311;
assign n_5001 = ~n_4321 & n_4996;
assign n_5002 = n_4996 ^ n_4332;
assign n_5003 = n_4797 ^ n_4996;
assign n_5004 = n_4997 ^ n_4130;
assign n_5005 = n_4998 ^ n_3059;
assign n_5006 = ~n_4998 & ~n_4995;
assign n_5007 = n_4999 ^ x311;
assign n_5008 = ~n_4988 & n_5000;
assign n_5009 = n_5000 ^ n_4988;
assign n_5010 = n_5001 ^ n_3793;
assign n_5011 = n_5004 ^ n_4373;
assign n_5012 = n_5005 ^ x310;
assign n_5013 = n_5006 ^ n_3059;
assign n_5014 = n_5007 ^ n_5005;
assign n_5015 = n_5010 ^ n_3083;
assign n_5016 = n_4171 ^ n_5011;
assign n_5017 = n_5011 & ~n_4384;
assign n_5018 = n_5013 ^ n_3083;
assign n_5019 = n_5013 ^ n_5010;
assign n_5020 = n_5014 ^ x310;
assign n_5021 = ~n_5014 & n_5012;
assign n_5022 = n_4362 & ~n_5016;
assign n_5023 = n_5016 ^ n_4373;
assign n_5024 = n_4822 ^ n_5016;
assign n_5025 = n_5017 ^ n_4171;
assign n_5026 = n_5018 ^ n_5010;
assign n_5027 = n_5015 & ~n_5019;
assign n_5028 = n_5020 & n_5008;
assign n_5029 = n_5008 ^ n_5020;
assign n_5030 = n_5021 ^ x310;
assign n_5031 = n_5022 ^ n_3831;
assign n_5032 = n_5025 ^ n_4403;
assign n_5033 = n_5026 ^ x309;
assign n_5034 = n_5027 ^ n_3083;
assign n_5035 = n_5030 ^ n_5026;
assign n_5036 = n_5031 ^ n_3113;
assign n_5037 = n_4214 ^ n_5032;
assign n_5038 = ~n_5032 & n_4412;
assign n_5039 = n_5034 ^ n_3113;
assign n_5040 = n_5034 ^ n_5031;
assign n_5041 = n_5035 ^ x309;
assign n_5042 = ~n_5035 & n_5033;
assign n_5043 = n_4395 & n_5037;
assign n_5044 = n_5037 ^ n_4403;
assign n_5045 = n_4844 ^ n_5037;
assign n_5046 = n_5038 ^ n_4214;
assign n_5047 = n_5039 ^ n_5031;
assign n_5048 = n_5036 & n_5040;
assign n_5049 = ~n_5028 & ~n_5041;
assign n_5050 = n_5041 ^ n_5028;
assign n_5051 = n_5042 ^ x309;
assign n_5052 = n_5043 ^ n_3873;
assign n_5053 = n_5046 ^ n_4426;
assign n_5054 = n_5047 ^ x308;
assign n_5055 = n_5048 ^ n_3113;
assign n_5056 = n_5051 ^ n_5047;
assign n_5057 = n_5052 ^ n_3147;
assign n_5058 = n_4257 ^ n_5053;
assign n_5059 = ~n_5053 & ~n_4434;
assign n_5060 = n_5055 ^ n_3147;
assign n_5061 = n_5055 ^ n_5052;
assign n_5062 = n_5056 ^ x308;
assign n_5063 = ~n_5056 & n_5054;
assign n_5064 = ~n_4420 & ~n_5058;
assign n_5065 = n_5058 ^ n_4426;
assign n_5066 = n_4862 ^ n_5058;
assign n_5067 = n_5059 ^ n_4257;
assign n_5068 = n_5060 ^ n_5052;
assign n_5069 = n_5057 & n_5061;
assign n_5070 = ~n_5049 & n_5062;
assign n_5071 = n_5063 ^ x308;
assign n_5072 = n_5064 ^ n_3914;
assign n_5073 = n_5067 ^ n_4440;
assign n_5074 = n_5068 ^ x307;
assign n_5075 = n_5069 ^ n_3147;
assign n_5076 = n_5071 ^ n_5068;
assign n_5077 = n_5072 ^ n_3185;
assign n_5078 = n_4299 ^ n_5073;
assign n_5079 = n_5073 & ~n_4449;
assign n_5080 = n_5075 ^ n_3185;
assign n_5081 = n_5075 ^ n_5072;
assign n_5082 = n_5076 ^ x307;
assign n_5083 = n_5076 & ~n_5074;
assign n_5084 = n_5078 & ~n_4448;
assign n_5085 = n_5078 ^ n_4440;
assign n_5086 = n_4883 ^ n_5078;
assign n_5087 = n_5079 ^ n_4299;
assign n_5088 = n_5080 ^ n_5072;
assign n_5089 = ~n_5077 & n_5081;
assign n_5090 = n_5070 ^ n_5082;
assign n_5091 = ~n_5082 & n_5070;
assign n_5092 = n_5083 ^ x307;
assign n_5093 = n_5084 ^ n_3956;
assign n_5094 = n_5087 ^ n_4466;
assign n_5095 = n_5088 ^ x306;
assign n_5096 = n_5089 ^ n_3185;
assign n_5097 = n_4562 & ~n_5090;
assign n_5098 = n_5090 ^ n_4562;
assign n_5099 = n_5092 ^ n_5088;
assign n_5100 = n_5093 ^ n_3225;
assign n_5101 = n_4341 ^ n_5094;
assign n_5102 = n_5094 & ~n_4475;
assign n_5103 = n_5096 ^ n_3225;
assign n_5104 = n_5096 ^ n_5093;
assign n_5105 = n_5097 ^ n_4591;
assign n_5106 = ~n_4554 & ~n_5098;
assign n_5107 = n_5099 ^ x306;
assign n_5108 = n_5099 & ~n_5095;
assign n_5109 = n_5101 & ~n_4474;
assign n_5110 = n_5101 ^ n_4466;
assign n_5111 = n_4903 ^ n_5101;
assign n_5112 = n_5102 ^ n_4341;
assign n_5113 = n_5103 ^ n_5093;
assign n_5114 = n_5100 & n_5104;
assign n_5115 = n_5106 ^ n_3574;
assign n_5116 = n_5091 ^ n_5107;
assign n_5117 = ~n_5107 & n_5091;
assign n_5118 = n_5108 ^ x306;
assign n_5119 = n_5109 ^ n_3999;
assign n_5120 = n_5112 ^ n_4487;
assign n_5121 = n_5113 ^ x305;
assign n_5122 = n_5114 ^ n_3225;
assign n_5123 = ~n_3070 & ~n_5115;
assign n_5124 = n_5115 ^ n_3070;
assign n_5125 = n_5105 ^ n_5116;
assign n_5126 = n_5097 ^ n_5116;
assign n_5127 = n_5118 ^ n_5113;
assign n_5128 = n_5119 ^ n_3267;
assign n_5129 = n_4379 ^ n_5120;
assign n_5130 = n_5120 & ~n_4496;
assign n_5131 = n_5122 ^ n_3267;
assign n_5132 = n_5122 ^ n_5119;
assign n_5133 = n_5123 ^ n_3097;
assign n_5134 = x327 & n_5124;
assign n_5135 = n_5124 ^ x327;
assign n_5136 = n_4590 & ~n_5125;
assign n_5137 = n_5126 & n_5105;
assign n_5138 = n_5127 ^ x305;
assign n_5139 = ~n_5127 & n_5121;
assign n_5140 = n_5129 & ~n_4495;
assign n_5141 = n_5129 ^ n_4487;
assign n_5142 = n_4926 ^ n_5129;
assign n_5143 = n_5130 ^ n_4379;
assign n_5144 = n_5131 ^ n_5119;
assign n_5145 = ~n_5128 & ~n_5132;
assign n_5146 = n_5134 ^ x326;
assign n_5147 = n_5136 ^ n_3619;
assign n_5148 = n_5137 ^ n_4591;
assign n_5149 = n_5117 ^ n_5138;
assign n_5150 = ~n_5138 & ~n_5117;
assign n_5151 = n_5139 ^ x305;
assign n_5152 = n_5140 ^ n_4029;
assign n_5153 = n_5143 ^ n_4407;
assign n_5154 = n_5143 ^ n_4508;
assign n_5155 = n_5144 ^ x304;
assign n_5156 = n_5145 ^ n_3267;
assign n_5157 = n_5147 ^ n_5133;
assign n_5158 = n_5147 ^ n_5123;
assign n_5159 = n_5148 ^ n_4630;
assign n_5160 = n_5149 ^ n_4630;
assign n_5161 = n_5148 ^ n_5149;
assign n_5162 = n_5151 ^ n_5144;
assign n_5163 = n_5152 ^ n_3306;
assign n_5164 = n_5153 ^ n_4508;
assign n_5165 = n_4516 & ~n_5154;
assign n_5166 = n_5152 ^ n_5156;
assign n_5167 = n_5157 ^ n_5134;
assign n_5168 = ~n_5133 & ~n_5158;
assign n_5169 = n_5159 ^ n_5149;
assign n_5170 = ~n_5160 & n_5161;
assign n_5171 = n_5162 ^ x304;
assign n_5172 = ~n_5162 & n_5155;
assign n_5173 = n_4502 & ~n_5164;
assign n_5174 = n_4947 ^ n_5164;
assign n_5175 = n_5165 ^ n_4407;
assign n_5176 = n_5166 ^ n_3306;
assign n_5177 = n_5166 & n_5163;
assign n_5178 = n_5167 & n_5146;
assign n_5179 = n_5167 ^ x326;
assign n_5180 = n_5168 ^ n_3097;
assign n_5181 = n_4624 & ~n_5169;
assign n_5182 = n_5170 ^ n_4630;
assign n_5183 = n_5171 ^ n_5150;
assign n_5184 = ~n_5150 & n_5171;
assign n_5185 = n_5172 ^ x304;
assign n_5186 = n_5173 ^ n_4084;
assign n_5187 = n_5175 ^ n_4528;
assign n_5188 = n_5176 ^ x319;
assign n_5189 = n_5177 ^ n_3306;
assign n_5190 = n_5178 ^ x326;
assign n_5191 = n_5135 & ~n_5179;
assign n_5192 = n_5179 ^ n_5135;
assign n_5193 = n_5180 ^ n_3137;
assign n_5194 = n_5181 ^ n_3677;
assign n_5195 = n_5182 ^ n_4669;
assign n_5196 = n_5183 ^ n_4669;
assign n_5197 = n_5182 ^ n_5183;
assign n_5198 = n_5185 ^ n_5176;
assign n_5199 = n_5186 ^ n_3348;
assign n_5200 = n_4429 ^ n_5187;
assign n_5201 = n_5187 & n_4537;
assign n_5202 = n_5189 ^ n_3348;
assign n_5203 = n_5189 ^ n_5186;
assign n_5204 = n_5190 ^ x325;
assign n_5205 = n_5193 ^ n_5194;
assign n_5206 = n_5194 ^ n_3137;
assign n_5207 = n_5180 ^ n_5194;
assign n_5208 = n_5195 ^ n_5183;
assign n_5209 = n_5196 & n_5197;
assign n_5210 = n_5198 ^ x319;
assign n_5211 = ~n_5198 & n_5188;
assign n_5212 = ~n_5200 & n_4536;
assign n_5213 = n_5200 ^ n_4528;
assign n_5214 = n_4968 ^ n_5200;
assign n_5215 = n_5201 ^ n_4429;
assign n_5216 = n_5202 ^ n_5186;
assign n_5217 = n_5199 & ~n_5203;
assign n_5218 = n_5190 ^ n_5205;
assign n_5219 = ~n_5206 & n_5207;
assign n_5220 = n_4661 & n_5208;
assign n_5221 = n_5209 ^ n_4669;
assign n_5222 = n_5184 ^ n_5210;
assign n_5223 = ~n_5210 & ~n_5184;
assign n_5224 = n_5211 ^ x319;
assign n_5225 = n_5212 ^ n_4127;
assign n_5226 = n_5215 ^ n_4452;
assign n_5227 = n_5215 ^ n_4551;
assign n_5228 = n_5216 ^ x318;
assign n_5229 = n_5217 ^ n_3348;
assign n_5230 = ~n_5218 & n_5204;
assign n_5231 = n_5218 ^ x325;
assign n_5232 = n_5219 ^ n_3137;
assign n_5233 = n_5220 ^ n_3713;
assign n_5234 = n_5221 ^ n_5222;
assign n_5235 = n_5222 ^ n_4705;
assign n_5236 = n_5224 ^ n_5216;
assign n_5237 = n_5225 ^ n_3389;
assign n_5238 = n_5226 ^ n_4551;
assign n_5239 = ~n_4559 & ~n_5227;
assign n_5240 = n_5229 ^ n_3389;
assign n_5241 = n_5229 ^ n_5225;
assign n_5242 = n_5230 ^ x325;
assign n_5243 = n_5231 & n_5191;
assign n_5244 = n_5191 ^ n_5231;
assign n_5245 = n_5232 ^ n_3178;
assign n_5246 = n_5233 ^ n_3178;
assign n_5247 = n_5232 ^ n_5233;
assign n_5248 = n_5234 ^ n_4705;
assign n_5249 = ~n_5234 & ~n_5235;
assign n_5250 = n_5236 ^ x318;
assign n_5251 = n_5236 & ~n_5228;
assign n_5252 = ~n_4544 & ~n_5238;
assign n_5253 = n_4989 ^ n_5238;
assign n_5254 = n_5239 ^ n_4452;
assign n_5255 = n_5240 ^ n_5225;
assign n_5256 = ~n_5237 & n_5241;
assign n_5257 = n_5242 ^ x324;
assign n_5258 = n_5245 ^ n_5233;
assign n_5259 = n_5246 & ~n_5247;
assign n_5260 = ~n_4695 & n_5248;
assign n_5261 = n_5249 ^ n_4705;
assign n_5262 = n_5223 ^ n_5250;
assign n_5263 = n_5250 & n_5223;
assign n_5264 = n_5251 ^ x318;
assign n_5265 = n_5252 ^ n_4168;
assign n_5266 = n_5254 ^ n_4576;
assign n_5267 = n_5255 ^ x317;
assign n_5268 = n_5256 ^ n_3389;
assign n_5269 = n_5242 ^ n_5258;
assign n_5270 = n_5259 ^ n_3178;
assign n_5271 = n_5260 ^ n_3751;
assign n_5272 = n_5261 ^ n_4733;
assign n_5273 = n_5262 ^ n_4733;
assign n_5274 = n_5261 ^ n_5262;
assign n_5275 = n_5264 ^ n_5255;
assign n_5276 = n_5265 ^ n_3431;
assign n_5277 = n_4469 ^ n_5266;
assign n_5278 = ~n_5266 & ~n_4586;
assign n_5279 = n_5268 ^ n_3431;
assign n_5280 = n_5268 ^ n_5265;
assign n_5281 = n_5269 & n_5257;
assign n_5282 = n_5269 ^ x324;
assign n_5283 = n_5270 ^ n_3218;
assign n_5284 = n_5271 ^ n_3218;
assign n_5285 = n_5270 ^ n_5271;
assign n_5286 = n_5272 ^ n_5262;
assign n_5287 = ~n_5273 & n_5274;
assign n_5288 = n_5275 ^ x317;
assign n_5289 = ~n_5275 & n_5267;
assign n_5290 = n_5277 & n_4585;
assign n_5291 = n_5277 ^ n_4576;
assign n_5292 = n_5009 ^ n_5277;
assign n_5293 = n_5278 ^ n_4469;
assign n_5294 = n_5279 ^ n_5265;
assign n_5295 = n_5276 & ~n_5280;
assign n_5296 = n_5281 ^ x324;
assign n_5297 = n_5243 & ~n_5282;
assign n_5298 = n_5282 ^ n_5243;
assign n_5299 = n_5283 ^ n_5271;
assign n_5300 = n_5284 & ~n_5285;
assign n_5301 = n_4727 & ~n_5286;
assign n_5302 = n_5287 ^ n_4733;
assign n_5303 = n_5263 ^ n_5288;
assign n_5304 = n_5288 & ~n_5263;
assign n_5305 = n_5289 ^ x317;
assign n_5306 = n_5290 ^ n_4211;
assign n_5307 = n_5293 ^ n_4608;
assign n_5308 = n_5294 ^ x316;
assign n_5309 = n_5295 ^ n_3431;
assign n_5310 = n_5296 ^ n_5299;
assign n_5311 = n_5299 ^ x323;
assign n_5312 = n_5300 ^ n_3218;
assign n_5313 = n_5301 ^ n_3787;
assign n_5314 = n_5302 ^ n_4756;
assign n_5315 = n_5303 ^ n_5302;
assign n_5316 = n_5303 ^ n_4756;
assign n_5317 = n_5305 ^ n_5294;
assign n_5318 = n_5306 ^ n_3473;
assign n_5319 = n_5307 ^ n_4490;
assign n_5320 = ~n_5307 & ~n_4619;
assign n_5321 = n_5309 ^ n_3473;
assign n_5322 = n_5309 ^ n_5306;
assign n_5323 = n_5310 ^ x323;
assign n_5324 = n_5310 & ~n_5311;
assign n_5325 = n_5312 ^ n_3260;
assign n_5326 = n_5313 ^ n_3260;
assign n_5327 = n_5312 ^ n_5313;
assign n_5328 = n_5314 ^ n_5303;
assign n_5329 = n_5315 & ~n_5316;
assign n_5330 = n_5317 ^ x316;
assign n_5331 = n_5317 & ~n_5308;
assign n_5332 = ~n_4596 & ~n_5319;
assign n_5333 = n_5319 ^ n_4608;
assign n_5334 = n_5029 ^ n_5319;
assign n_5335 = n_5320 ^ n_4490;
assign n_5336 = n_5321 ^ n_5306;
assign n_5337 = ~n_5318 & ~n_5322;
assign n_5338 = ~n_5297 & n_5323;
assign n_5339 = n_5323 ^ n_5297;
assign n_5340 = n_5324 ^ x323;
assign n_5341 = n_5325 ^ n_5313;
assign n_5342 = n_5326 & n_5327;
assign n_5343 = ~n_4748 & ~n_5328;
assign n_5344 = n_5329 ^ n_4756;
assign n_5345 = n_5330 ^ n_5304;
assign n_5346 = ~n_5304 & n_5330;
assign n_5347 = n_5331 ^ x316;
assign n_5348 = n_5332 ^ n_4254;
assign n_5349 = n_5335 ^ n_4640;
assign n_5350 = n_5336 ^ x315;
assign n_5351 = n_5337 ^ n_3473;
assign n_5352 = n_5340 ^ n_5341;
assign n_5353 = n_5341 ^ x322;
assign n_5354 = n_5342 ^ n_3260;
assign n_5355 = n_5343 ^ n_3824;
assign n_5356 = n_5344 ^ n_4773;
assign n_5357 = n_5345 ^ n_4773;
assign n_5358 = n_5344 ^ n_5345;
assign n_5359 = n_5347 ^ n_5336;
assign n_5360 = n_5348 ^ n_3515;
assign n_5361 = n_5349 ^ n_4511;
assign n_5362 = ~n_5349 & ~n_4655;
assign n_5363 = n_5351 ^ n_3515;
assign n_5364 = n_5351 ^ n_5348;
assign n_5365 = n_5352 ^ x322;
assign n_5366 = n_5352 & ~n_5353;
assign n_5367 = n_5354 ^ n_3299;
assign n_5368 = n_5355 ^ n_3299;
assign n_5369 = n_5354 ^ n_5355;
assign n_5370 = n_5356 ^ n_5345;
assign n_5371 = ~n_5357 & ~n_5358;
assign n_5372 = n_5359 ^ x315;
assign n_5373 = ~n_5359 & n_5350;
assign n_5374 = n_5361 & ~n_4654;
assign n_5375 = n_5361 ^ n_4640;
assign n_5376 = n_5050 ^ n_5361;
assign n_5377 = n_5362 ^ n_4511;
assign n_5378 = n_5363 ^ n_5348;
assign n_5379 = n_5360 & n_5364;
assign n_5380 = n_5338 & n_5365;
assign n_5381 = n_5365 ^ n_5338;
assign n_5382 = n_5366 ^ x322;
assign n_5383 = n_5367 ^ n_5355;
assign n_5384 = ~n_5368 & n_5369;
assign n_5385 = ~n_5370 & ~n_4782;
assign n_5386 = n_5371 ^ n_4773;
assign n_5387 = n_5372 ^ n_5346;
assign n_5388 = ~n_5346 & n_5372;
assign n_5389 = n_5373 ^ x315;
assign n_5390 = n_5374 ^ n_4296;
assign n_5391 = n_5377 ^ n_4677;
assign n_5392 = n_5378 ^ x314;
assign n_5393 = n_5379 ^ n_3515;
assign n_5394 = n_5382 ^ n_5383;
assign n_5395 = n_5383 ^ x321;
assign n_5396 = n_5384 ^ n_3299;
assign n_5397 = n_5385 ^ n_3866;
assign n_5398 = n_5386 ^ n_4792;
assign n_5399 = n_5387 ^ n_4792;
assign n_5400 = n_5386 ^ n_5387;
assign n_5401 = n_5389 ^ n_5378;
assign n_5402 = n_5390 ^ n_3556;
assign n_5403 = ~n_5391 & ~n_4678;
assign n_5404 = n_5391 ^ n_5049;
assign n_5405 = n_5391 ^ n_4666;
assign n_5406 = n_5393 ^ n_3556;
assign n_5407 = n_5390 ^ n_5393;
assign n_5408 = n_5394 ^ x321;
assign n_5409 = n_5394 & ~n_5395;
assign n_5410 = n_5396 ^ n_3342;
assign n_5411 = n_5397 ^ n_3342;
assign n_5412 = n_5396 ^ n_5397;
assign n_5413 = n_5398 ^ n_5387;
assign n_5414 = n_5399 & ~n_5400;
assign n_5415 = n_5401 ^ x314;
assign n_5416 = ~n_5401 & n_5392;
assign n_5417 = n_5403 ^ n_4339;
assign n_5418 = n_5404 ^ n_5062;
assign n_5419 = n_5390 ^ n_5406;
assign n_5420 = n_5402 & n_5407;
assign n_5421 = ~n_5380 & ~n_5408;
assign n_5422 = n_5408 ^ n_5380;
assign n_5423 = n_5409 ^ x321;
assign n_5424 = n_5410 ^ n_5397;
assign n_5425 = ~n_5411 & ~n_5412;
assign n_5426 = ~n_5413 & n_4801;
assign n_5427 = n_5414 ^ n_4792;
assign n_5428 = n_5415 ^ n_5388;
assign n_5429 = n_5388 & n_5415;
assign n_5430 = n_5416 ^ x314;
assign n_5431 = n_5417 ^ n_3587;
assign n_5432 = n_5419 ^ x313;
assign n_5433 = n_5420 ^ n_3556;
assign n_5434 = n_5423 ^ n_5424;
assign n_5435 = n_5424 ^ x320;
assign n_5436 = n_5425 ^ n_3342;
assign n_5437 = n_5426 ^ n_3907;
assign n_5438 = n_5427 ^ n_4810;
assign n_5439 = n_5428 ^ n_4810;
assign n_5440 = n_5427 ^ n_5428;
assign n_5441 = n_5430 ^ n_5419;
assign n_5442 = n_5433 ^ x312;
assign n_5443 = n_5434 ^ x320;
assign n_5444 = n_5434 & ~n_5435;
assign n_5445 = n_5436 ^ n_3382;
assign n_5446 = n_5437 ^ n_3382;
assign n_5447 = n_5436 ^ n_5437;
assign n_5448 = n_5438 ^ n_5428;
assign n_5449 = n_5439 & n_5440;
assign n_5450 = n_5441 ^ x313;
assign n_5451 = n_5441 & ~n_5432;
assign n_5452 = n_5442 ^ n_5431;
assign n_5453 = ~n_5421 & n_5443;
assign n_5454 = n_5443 ^ n_5421;
assign n_5455 = n_5444 ^ x320;
assign n_5456 = n_5445 ^ n_5437;
assign n_5457 = ~n_5446 & ~n_5447;
assign n_5458 = ~n_5448 & ~n_4818;
assign n_5459 = n_5449 ^ n_4810;
assign n_5460 = n_5429 ^ n_5450;
assign n_5461 = ~n_5450 & n_5429;
assign n_5462 = n_5451 ^ x313;
assign n_5463 = n_5455 ^ n_5456;
assign n_5464 = n_5456 ^ x335;
assign n_5465 = n_5457 ^ n_3382;
assign n_5466 = n_5458 ^ n_3949;
assign n_5467 = n_5459 ^ n_4825;
assign n_5468 = n_5459 ^ n_5460;
assign n_5469 = n_5460 ^ n_4825;
assign n_5470 = n_5462 ^ n_5452;
assign n_5471 = n_5463 ^ x335;
assign n_5472 = ~n_5463 & n_5464;
assign n_5473 = n_5465 ^ n_3424;
assign n_5474 = n_5466 ^ n_3424;
assign n_5475 = n_5465 ^ n_5466;
assign n_5476 = n_5467 ^ n_5460;
assign n_5477 = n_5468 & n_5469;
assign n_5478 = n_5470 ^ n_5461;
assign n_5479 = ~n_5471 & n_5453;
assign n_5480 = n_5453 ^ n_5471;
assign n_5481 = n_5472 ^ x335;
assign n_5482 = n_5473 ^ n_5466;
assign n_5483 = ~n_5474 & n_5475;
assign n_5484 = n_5476 & n_4832;
assign n_5485 = n_5477 ^ n_4825;
assign n_5486 = n_5478 ^ n_4849;
assign n_5487 = n_5481 ^ n_5482;
assign n_5488 = n_5482 ^ x334;
assign n_5489 = n_5483 ^ n_3424;
assign n_5490 = n_5484 ^ n_3992;
assign n_5491 = n_5485 ^ n_4849;
assign n_5492 = n_5485 ^ n_5478;
assign n_5493 = n_5487 ^ x334;
assign n_5494 = n_5487 & ~n_5488;
assign n_5495 = n_5489 ^ n_3466;
assign n_5496 = n_5490 ^ n_3466;
assign n_5497 = n_5489 ^ n_5490;
assign n_5498 = n_5491 ^ n_5478;
assign n_5499 = n_5486 & ~n_5492;
assign n_5500 = n_5479 & n_5493;
assign n_5501 = n_5493 ^ n_5479;
assign n_5502 = n_5494 ^ x334;
assign n_5503 = n_5495 ^ n_5490;
assign n_5504 = n_5496 & n_5497;
assign n_5505 = ~n_5498 & n_4856;
assign n_5506 = n_5499 ^ n_4849;
assign n_5507 = n_5502 ^ n_5503;
assign n_5508 = n_5503 ^ x333;
assign n_5509 = n_5504 ^ n_3466;
assign n_5510 = n_5505 ^ n_4035;
assign n_5511 = n_5506 ^ n_4876;
assign n_5512 = n_5506 ^ n_4600;
assign n_5513 = n_5507 ^ x333;
assign n_5514 = ~n_5507 & n_5508;
assign n_5515 = n_5509 ^ n_3508;
assign n_5516 = n_5510 ^ n_3508;
assign n_5517 = n_5509 ^ n_5510;
assign n_5518 = n_5511 & ~n_4877;
assign n_5519 = ~n_4876 & n_5512;
assign n_5520 = ~n_5500 & n_5513;
assign n_5521 = n_5513 ^ n_5500;
assign n_5522 = n_5514 ^ x333;
assign n_5523 = n_5515 ^ n_5510;
assign n_5524 = ~n_5516 & ~n_5517;
assign n_5525 = n_5518 ^ n_4079;
assign n_5526 = n_5519 ^ n_4869;
assign n_5527 = n_5522 ^ n_5523;
assign n_5528 = n_5523 ^ x332;
assign n_5529 = n_5524 ^ n_3508;
assign n_5530 = n_5526 ^ n_4646;
assign n_5531 = n_5526 ^ n_4890;
assign n_5532 = n_5527 ^ x332;
assign n_5533 = ~n_5527 & n_5528;
assign n_5534 = n_5529 ^ n_3550;
assign n_5535 = n_5525 ^ n_5529;
assign n_5536 = n_5530 ^ n_4890;
assign n_5537 = ~n_4898 & n_5531;
assign n_5538 = ~n_5520 & ~n_5532;
assign n_5539 = n_5532 ^ n_5520;
assign n_5540 = n_5533 ^ x332;
assign n_5541 = n_5525 ^ n_5534;
assign n_5542 = ~n_5534 & ~n_5535;
assign n_5543 = n_5536 & ~n_4897;
assign n_5544 = n_5537 ^ n_4646;
assign n_5545 = n_5540 ^ n_5541;
assign n_5546 = n_5541 ^ x331;
assign n_5547 = n_5542 ^ n_3550;
assign n_5548 = n_5543 ^ n_4120;
assign n_5549 = n_5544 ^ n_4912;
assign n_5550 = n_5545 ^ x331;
assign n_5551 = n_5545 & ~n_5546;
assign n_5552 = n_5547 ^ n_3595;
assign n_5553 = n_5548 ^ n_3595;
assign n_5554 = n_5547 ^ n_5548;
assign n_5555 = n_4711 ^ n_5549;
assign n_5556 = ~n_5549 & n_4920;
assign n_5557 = n_5538 & n_5550;
assign n_5558 = n_5550 ^ n_5538;
assign n_5559 = n_5551 ^ x331;
assign n_5560 = n_5552 ^ n_5548;
assign n_5561 = n_5553 & ~n_5554;
assign n_5562 = ~n_5555 & ~n_4919;
assign n_5563 = n_5555 ^ n_4912;
assign n_5564 = n_5556 ^ n_4711;
assign n_5565 = n_5559 ^ x330;
assign n_5566 = n_5559 ^ n_5560;
assign n_5567 = n_5561 ^ n_3595;
assign n_5568 = n_5562 ^ n_4162;
assign n_5569 = n_5564 ^ n_4933;
assign n_5570 = n_5566 & n_5565;
assign n_5571 = n_5566 ^ x330;
assign n_5572 = n_5567 ^ n_3643;
assign n_5573 = n_5568 ^ n_3643;
assign n_5574 = n_5567 ^ n_5568;
assign n_5575 = n_4737 ^ n_5569;
assign n_5576 = ~n_5569 & n_4941;
assign n_5577 = n_5570 ^ x330;
assign n_5578 = ~n_5557 & ~n_5571;
assign n_5579 = n_5571 ^ n_5557;
assign n_5580 = n_5572 ^ n_5568;
assign n_5581 = ~n_5573 & n_5574;
assign n_5582 = ~n_5575 & n_4940;
assign n_5583 = n_5575 ^ n_4933;
assign n_5584 = n_5576 ^ n_4737;
assign n_5585 = n_5577 ^ n_5580;
assign n_5586 = n_5580 ^ x329;
assign n_5587 = n_5581 ^ n_3643;
assign n_5588 = n_5582 ^ n_4204;
assign n_5589 = n_5584 ^ n_4954;
assign n_5590 = n_5585 ^ x329;
assign n_5591 = ~n_5585 & n_5586;
assign n_5592 = n_5587 ^ n_3684;
assign n_5593 = n_5588 ^ n_3684;
assign n_5594 = n_5587 ^ n_5588;
assign n_5595 = n_4758 ^ n_5589;
assign n_5596 = n_5589 & ~n_4962;
assign n_5597 = ~n_5578 & ~n_5590;
assign n_5598 = n_5590 ^ n_5578;
assign n_5599 = n_5591 ^ x329;
assign n_5600 = n_5592 ^ n_5588;
assign n_5601 = n_5593 & ~n_5594;
assign n_5602 = n_5595 & n_4961;
assign n_5603 = n_5595 ^ n_4954;
assign n_5604 = n_5596 ^ n_4758;
assign n_5605 = n_5599 ^ n_5600;
assign n_5606 = n_5600 ^ x328;
assign n_5607 = n_5601 ^ n_3684;
assign n_5608 = n_5602 ^ n_4247;
assign n_5609 = n_5604 ^ n_4777;
assign n_5610 = n_5604 ^ n_4976;
assign n_5611 = n_5605 ^ x328;
assign n_5612 = n_5605 & ~n_5606;
assign n_5613 = n_5608 ^ n_3720;
assign n_5614 = n_5607 ^ n_5608;
assign n_5615 = n_5609 ^ n_4976;
assign n_5616 = ~n_4983 & ~n_5610;
assign n_5617 = n_5611 ^ n_5597;
assign n_5618 = ~n_5597 & ~n_5611;
assign n_5619 = n_5612 ^ x328;
assign n_5620 = n_5607 ^ n_5613;
assign n_5621 = ~n_5613 & n_5614;
assign n_5622 = ~n_4970 & n_5615;
assign n_5623 = n_5135 ^ n_5615;
assign n_5624 = n_5616 ^ n_4777;
assign n_5625 = n_5617 ^ n_5098;
assign n_5626 = ~n_5098 & n_5617;
assign n_5627 = n_5619 ^ x343;
assign n_5628 = n_5620 ^ n_5619;
assign n_5629 = n_5621 ^ n_3720;
assign n_5630 = n_5622 ^ n_4289;
assign n_5631 = n_5624 ^ n_4996;
assign n_5632 = ~n_5090 & ~n_5625;
assign n_5633 = n_5626 ^ n_5125;
assign n_5634 = n_5628 ^ x343;
assign n_5635 = ~n_5628 & n_5627;
assign n_5636 = n_5629 ^ n_5630;
assign n_5637 = n_5630 ^ n_3745;
assign n_5638 = n_4797 ^ n_5631;
assign n_5639 = ~n_5631 & n_5003;
assign n_5640 = n_5632 ^ n_4562;
assign n_5641 = n_5618 ^ n_5634;
assign n_5642 = ~n_5634 & ~n_5618;
assign n_5643 = n_5635 ^ x343;
assign n_5644 = n_5636 ^ n_3745;
assign n_5645 = n_5636 & ~n_5637;
assign n_5646 = n_5638 & ~n_5002;
assign n_5647 = n_5638 ^ n_4996;
assign n_5648 = n_5192 ^ n_5638;
assign n_5649 = n_5639 ^ n_4797;
assign n_5650 = n_5640 ^ n_3574;
assign n_5651 = ~n_3574 & n_5640;
assign n_5652 = n_5641 ^ n_5633;
assign n_5653 = n_5641 ^ n_5626;
assign n_5654 = n_5643 ^ n_5644;
assign n_5655 = n_5644 ^ x342;
assign n_5656 = n_5645 ^ n_3745;
assign n_5657 = n_5646 ^ n_4332;
assign n_5658 = n_5649 ^ n_5016;
assign n_5659 = x359 & ~n_5650;
assign n_5660 = n_5650 ^ x359;
assign n_5661 = n_5651 ^ n_3619;
assign n_5662 = ~n_5126 & n_5652;
assign n_5663 = ~n_5633 & n_5653;
assign n_5664 = n_5654 ^ x342;
assign n_5665 = ~n_5654 & n_5655;
assign n_5666 = n_5656 ^ n_3793;
assign n_5667 = n_5657 ^ n_3793;
assign n_5668 = n_5656 ^ n_5657;
assign n_5669 = n_4822 ^ n_5658;
assign n_5670 = n_5658 & ~n_5024;
assign n_5671 = n_5659 ^ x358;
assign n_5672 = n_5662 ^ n_4591;
assign n_5673 = n_5663 ^ n_5125;
assign n_5674 = n_5642 ^ n_5664;
assign n_5675 = ~n_5664 & n_5642;
assign n_5676 = n_5665 ^ x342;
assign n_5677 = n_5666 ^ n_5657;
assign n_5678 = ~n_5667 & ~n_5668;
assign n_5679 = ~n_5669 & n_5023;
assign n_5680 = n_5669 ^ n_5016;
assign n_5681 = n_5244 ^ n_5669;
assign n_5682 = n_5670 ^ n_4822;
assign n_5683 = n_5672 ^ n_5661;
assign n_5684 = n_5672 ^ n_5651;
assign n_5685 = n_5673 ^ n_5169;
assign n_5686 = n_5674 ^ n_5169;
assign n_5687 = n_5673 ^ n_5674;
assign n_5688 = n_5676 ^ n_5677;
assign n_5689 = n_5677 ^ x341;
assign n_5690 = n_5678 ^ n_3793;
assign n_5691 = n_5679 ^ n_4373;
assign n_5692 = n_5682 ^ n_5037;
assign n_5693 = n_5683 ^ n_5659;
assign n_5694 = n_5683 ^ n_5671;
assign n_5695 = n_5661 & ~n_5684;
assign n_5696 = n_5685 ^ n_5674;
assign n_5697 = ~n_5686 & n_5687;
assign n_5698 = n_5688 ^ x341;
assign n_5699 = ~n_5688 & n_5689;
assign n_5700 = n_5690 ^ n_3831;
assign n_5701 = n_5691 ^ n_3831;
assign n_5702 = n_5690 ^ n_5691;
assign n_5703 = n_4844 ^ n_5692;
assign n_5704 = ~n_5692 & n_5045;
assign n_5705 = n_5671 & ~n_5693;
assign n_5706 = n_5695 ^ n_3619;
assign n_5707 = ~n_5161 & n_5696;
assign n_5708 = n_5697 ^ n_5169;
assign n_5709 = n_5675 ^ n_5698;
assign n_5710 = ~n_5698 & n_5675;
assign n_5711 = n_5699 ^ x341;
assign n_5712 = n_5700 ^ n_5691;
assign n_5713 = n_5701 & n_5702;
assign n_5714 = n_5703 & n_5044;
assign n_5715 = n_5703 ^ n_5037;
assign n_5716 = n_5298 ^ n_5703;
assign n_5717 = n_5704 ^ n_4844;
assign n_5718 = n_5705 ^ x358;
assign n_5719 = n_5706 ^ n_3677;
assign n_5720 = n_5707 ^ n_4630;
assign n_5721 = n_5708 ^ n_5208;
assign n_5722 = n_5709 ^ n_5208;
assign n_5723 = n_5708 ^ n_5709;
assign n_5724 = n_5711 ^ n_5712;
assign n_5725 = n_5712 ^ x340;
assign n_5726 = n_5713 ^ n_3831;
assign n_5727 = n_5714 ^ n_4403;
assign n_5728 = n_5717 ^ n_5058;
assign n_5729 = n_5719 ^ n_5720;
assign n_5730 = n_5720 ^ n_3677;
assign n_5731 = n_5706 ^ n_5720;
assign n_5732 = n_5721 ^ n_5709;
assign n_5733 = n_5722 & n_5723;
assign n_5734 = n_5724 ^ x340;
assign n_5735 = ~n_5724 & n_5725;
assign n_5736 = n_5726 ^ n_3873;
assign n_5737 = n_5727 ^ n_3873;
assign n_5738 = n_5726 ^ n_5727;
assign n_5739 = n_4862 ^ n_5728;
assign n_5740 = n_5728 & n_5066;
assign n_5741 = n_5718 ^ n_5729;
assign n_5742 = n_5729 ^ x357;
assign n_5743 = n_5730 & ~n_5731;
assign n_5744 = ~n_5197 & ~n_5732;
assign n_5745 = n_5733 ^ n_5208;
assign n_5746 = n_5710 ^ n_5734;
assign n_5747 = ~n_5734 & n_5710;
assign n_5748 = n_5735 ^ x340;
assign n_5749 = n_5736 ^ n_5727;
assign n_5750 = n_5737 & n_5738;
assign n_5751 = n_5739 & ~n_5065;
assign n_5752 = n_5739 ^ n_5058;
assign n_5753 = n_5339 ^ n_5739;
assign n_5754 = n_5740 ^ n_4862;
assign n_5755 = n_5741 ^ x357;
assign n_5756 = ~n_5741 & n_5742;
assign n_5757 = n_5743 ^ n_3677;
assign n_5758 = n_5744 ^ n_4669;
assign n_5759 = n_5745 ^ n_5248;
assign n_5760 = n_5746 ^ n_5248;
assign n_5761 = n_5745 ^ n_5746;
assign n_5762 = n_5748 ^ n_5749;
assign n_5763 = n_5749 ^ x339;
assign n_5764 = n_5750 ^ n_3873;
assign n_5765 = n_5751 ^ n_4426;
assign n_5766 = n_5754 ^ n_5078;
assign n_5767 = ~n_5694 & ~n_5755;
assign n_5768 = n_5755 ^ n_5694;
assign n_5769 = n_5756 ^ x357;
assign n_5770 = n_5757 ^ n_3713;
assign n_5771 = n_5758 ^ n_3713;
assign n_5772 = n_5757 ^ n_5758;
assign n_5773 = n_5759 ^ n_5746;
assign n_5774 = n_5760 & ~n_5761;
assign n_5775 = n_5762 ^ x339;
assign n_5776 = n_5762 & ~n_5763;
assign n_5777 = n_5764 ^ n_3914;
assign n_5778 = n_5765 ^ n_3914;
assign n_5779 = n_5764 ^ n_5765;
assign n_5780 = n_4883 ^ n_5766;
assign n_5781 = n_5766 & ~n_5086;
assign n_5782 = n_5770 ^ n_5758;
assign n_5783 = n_5771 & n_5772;
assign n_5784 = n_5234 & n_5773;
assign n_5785 = n_5774 ^ n_5248;
assign n_5786 = n_5747 ^ n_5775;
assign n_5787 = n_5775 & n_5747;
assign n_5788 = n_5776 ^ x339;
assign n_5789 = n_5777 ^ n_5765;
assign n_5790 = ~n_5778 & ~n_5779;
assign n_5791 = n_5780 & n_5085;
assign n_5792 = n_5780 ^ n_5078;
assign n_5793 = n_5381 ^ n_5780;
assign n_5794 = n_5781 ^ n_4883;
assign n_5795 = n_5769 ^ n_5782;
assign n_5796 = n_5782 ^ x356;
assign n_5797 = n_5783 ^ n_3713;
assign n_5798 = n_5784 ^ n_4705;
assign n_5799 = n_5785 ^ n_5286;
assign n_5800 = n_5786 ^ n_5286;
assign n_5801 = n_5785 ^ n_5786;
assign n_5802 = n_5788 ^ n_5789;
assign n_5803 = n_5789 ^ x338;
assign n_5804 = n_5790 ^ n_3914;
assign n_5805 = n_5791 ^ n_4440;
assign n_5806 = n_5794 ^ n_5101;
assign n_5807 = n_5795 ^ x356;
assign n_5808 = ~n_5795 & n_5796;
assign n_5809 = n_5797 ^ n_3751;
assign n_5810 = n_5798 ^ n_3751;
assign n_5811 = n_5797 ^ n_5798;
assign n_5812 = n_5799 ^ n_5786;
assign n_5813 = n_5800 & n_5801;
assign n_5814 = n_5802 ^ x338;
assign n_5815 = n_5802 & ~n_5803;
assign n_5816 = n_5804 ^ n_3956;
assign n_5817 = n_5805 ^ n_3956;
assign n_5818 = n_5804 ^ n_5805;
assign n_5819 = n_4903 ^ n_5806;
assign n_5820 = n_5806 & n_5111;
assign n_5821 = n_5767 & ~n_5807;
assign n_5822 = n_5807 ^ n_5767;
assign n_5823 = n_5808 ^ x356;
assign n_5824 = n_5809 ^ n_5798;
assign n_5825 = ~n_5810 & n_5811;
assign n_5826 = ~n_5274 & n_5812;
assign n_5827 = n_5813 ^ n_5286;
assign n_5828 = n_5814 ^ n_5787;
assign n_5829 = n_5787 & n_5814;
assign n_5830 = n_5815 ^ x338;
assign n_5831 = n_5816 ^ n_5805;
assign n_5832 = ~n_5817 & n_5818;
assign n_5833 = ~n_5819 & n_5110;
assign n_5834 = n_5819 ^ n_5101;
assign n_5835 = n_5422 ^ n_5819;
assign n_5836 = n_5820 ^ n_4903;
assign n_5837 = n_5823 ^ n_5824;
assign n_5838 = n_5824 ^ x355;
assign n_5839 = n_5825 ^ n_3751;
assign n_5840 = n_5826 ^ n_4733;
assign n_5841 = n_5827 ^ n_5328;
assign n_5842 = n_5828 ^ n_5328;
assign n_5843 = n_5828 ^ n_5827;
assign n_5844 = n_5830 ^ n_5831;
assign n_5845 = n_5831 ^ x337;
assign n_5846 = n_5832 ^ n_3956;
assign n_5847 = n_5833 ^ n_4466;
assign n_5848 = n_5836 ^ n_5129;
assign n_5849 = n_5837 ^ x355;
assign n_5850 = ~n_5837 & n_5838;
assign n_5851 = n_5839 ^ n_3787;
assign n_5852 = n_5840 ^ n_3787;
assign n_5853 = n_5839 ^ n_5840;
assign n_5854 = n_5828 ^ n_5841;
assign n_5855 = n_5842 & ~n_5843;
assign n_5856 = n_5844 ^ x337;
assign n_5857 = ~n_5844 & n_5845;
assign n_5858 = n_5846 ^ n_3999;
assign n_5859 = n_5847 ^ n_3999;
assign n_5860 = n_5846 ^ n_5847;
assign n_5861 = n_4926 ^ n_5848;
assign n_5862 = ~n_5848 & ~n_5142;
assign n_5863 = n_5821 & ~n_5849;
assign n_5864 = n_5849 ^ n_5821;
assign n_5865 = n_5850 ^ x355;
assign n_5866 = n_5851 ^ n_5840;
assign n_5867 = n_5852 & n_5853;
assign n_5868 = ~n_5315 & ~n_5854;
assign n_5869 = n_5855 ^ n_5328;
assign n_5870 = n_5856 ^ n_5829;
assign n_5871 = n_5829 & ~n_5856;
assign n_5872 = n_5857 ^ x337;
assign n_5873 = n_5858 ^ n_5847;
assign n_5874 = ~n_5859 & n_5860;
assign n_5875 = ~n_5861 & n_5141;
assign n_5876 = n_5861 ^ n_5129;
assign n_5877 = n_5454 ^ n_5861;
assign n_5878 = n_5862 ^ n_4926;
assign n_5879 = n_5865 ^ n_5866;
assign n_5880 = n_5866 ^ x354;
assign n_5881 = n_5867 ^ n_3787;
assign n_5882 = n_5868 ^ n_4756;
assign n_5883 = n_5869 ^ n_5370;
assign n_5884 = n_5870 ^ n_5370;
assign n_5885 = n_5870 ^ n_5869;
assign n_5886 = n_5872 ^ n_5873;
assign n_5887 = n_5873 ^ x336;
assign n_5888 = n_5874 ^ n_3999;
assign n_5889 = n_5875 ^ n_4487;
assign n_5890 = n_5878 ^ n_4947;
assign n_5891 = n_5878 ^ n_5164;
assign n_5892 = n_5879 ^ x354;
assign n_5893 = n_5879 & ~n_5880;
assign n_5894 = n_5881 ^ n_3824;
assign n_5895 = n_5882 ^ n_3824;
assign n_5896 = n_5881 ^ n_5882;
assign n_5897 = n_5870 ^ n_5883;
assign n_5898 = ~n_5884 & n_5885;
assign n_5899 = n_5886 ^ x336;
assign n_5900 = ~n_5886 & n_5887;
assign n_5901 = n_5888 ^ n_5889;
assign n_5902 = n_5889 ^ n_4029;
assign n_5903 = n_5890 ^ n_5164;
assign n_5904 = n_5174 & ~n_5891;
assign n_5905 = n_5892 & n_5863;
assign n_5906 = n_5863 ^ n_5892;
assign n_5907 = n_5893 ^ x354;
assign n_5908 = n_5894 ^ n_5882;
assign n_5909 = ~n_5895 & ~n_5896;
assign n_5910 = n_5358 & n_5897;
assign n_5911 = n_5898 ^ n_5370;
assign n_5912 = n_5871 ^ n_5899;
assign n_5913 = ~n_5899 & n_5871;
assign n_5914 = n_5900 ^ x336;
assign n_5915 = n_5901 ^ n_4029;
assign n_5916 = n_5901 & ~n_5902;
assign n_5917 = n_5153 & ~n_5903;
assign n_5918 = n_5480 ^ n_5903;
assign n_5919 = n_5904 ^ n_4947;
assign n_5920 = n_5907 ^ n_5908;
assign n_5921 = n_5908 ^ x353;
assign n_5922 = n_5909 ^ n_3824;
assign n_5923 = n_5910 ^ n_4773;
assign n_5924 = n_5911 ^ n_5413;
assign n_5925 = n_5912 ^ n_5413;
assign n_5926 = n_5911 ^ n_5912;
assign n_5927 = n_5914 ^ n_5915;
assign n_5928 = n_5915 ^ x351;
assign n_5929 = n_5916 ^ n_4029;
assign n_5930 = n_5917 ^ n_4508;
assign n_5931 = n_5919 ^ n_5200;
assign n_5932 = n_5920 ^ x353;
assign n_5933 = n_5920 & ~n_5921;
assign n_5934 = n_5922 ^ n_3866;
assign n_5935 = n_5923 ^ n_3866;
assign n_5936 = n_5923 ^ n_5922;
assign n_5937 = n_5924 ^ n_5912;
assign n_5938 = ~n_5925 & n_5926;
assign n_5939 = n_5927 ^ x351;
assign n_5940 = ~n_5927 & n_5928;
assign n_5941 = n_5929 ^ n_5930;
assign n_5942 = n_5930 ^ n_4084;
assign n_5943 = n_4968 ^ n_5931;
assign n_5944 = ~n_5931 & n_5214;
assign n_5945 = ~n_5905 & ~n_5932;
assign n_5946 = n_5932 ^ n_5905;
assign n_5947 = n_5933 ^ x353;
assign n_5948 = n_5923 ^ n_5934;
assign n_5949 = ~n_5935 & ~n_5936;
assign n_5950 = n_5400 & n_5937;
assign n_5951 = n_5938 ^ n_5413;
assign n_5952 = n_5913 ^ n_5939;
assign n_5953 = ~n_5939 & n_5913;
assign n_5954 = n_5940 ^ x351;
assign n_5955 = n_5941 ^ n_4084;
assign n_5956 = ~n_5941 & n_5942;
assign n_5957 = ~n_5943 & ~n_5213;
assign n_5958 = n_5943 ^ n_5200;
assign n_5959 = n_5501 ^ n_5943;
assign n_5960 = n_5944 ^ n_4968;
assign n_5961 = n_5947 ^ n_5948;
assign n_5962 = n_5948 ^ x352;
assign n_5963 = n_5949 ^ n_3866;
assign n_5964 = n_5950 ^ n_4792;
assign n_5965 = n_5951 ^ n_5448;
assign n_5966 = n_5952 ^ n_5448;
assign n_5967 = n_5951 ^ n_5952;
assign n_5968 = n_5954 ^ n_5955;
assign n_5969 = n_5955 ^ x350;
assign n_5970 = n_5956 ^ n_4084;
assign n_5971 = n_5957 ^ n_4528;
assign n_5972 = n_5960 ^ n_4989;
assign n_5973 = n_5960 ^ n_5238;
assign n_5974 = n_5961 ^ x352;
assign n_5975 = ~n_5961 & n_5962;
assign n_5976 = n_5963 ^ n_3907;
assign n_5977 = n_5964 ^ n_3907;
assign n_5978 = n_5963 ^ n_5964;
assign n_5979 = n_5965 ^ n_5952;
assign n_5980 = ~n_5966 & n_5967;
assign n_5981 = n_5968 ^ x350;
assign n_5982 = n_5968 & ~n_5969;
assign n_5983 = n_5970 ^ n_5971;
assign n_5984 = n_5971 ^ n_4127;
assign n_5985 = n_5972 ^ n_5238;
assign n_5986 = n_5253 & ~n_5973;
assign n_5987 = ~n_5974 & ~n_5945;
assign n_5988 = n_5945 ^ n_5974;
assign n_5989 = n_5975 ^ x352;
assign n_5990 = n_5976 ^ n_5964;
assign n_5991 = n_5977 & n_5978;
assign n_5992 = ~n_5440 & n_5979;
assign n_5993 = n_5980 ^ n_5448;
assign n_5994 = n_5981 ^ n_5953;
assign n_5995 = n_5953 & n_5981;
assign n_5996 = n_5982 ^ x350;
assign n_5997 = n_5983 ^ n_4127;
assign n_5998 = n_5983 & n_5984;
assign n_5999 = ~n_5226 & ~n_5985;
assign n_6000 = n_5521 ^ n_5985;
assign n_6001 = n_5986 ^ n_4989;
assign n_6002 = n_5989 ^ n_5990;
assign n_6003 = n_5990 ^ x367;
assign n_6004 = n_5991 ^ n_3907;
assign n_6005 = n_5992 ^ n_4810;
assign n_6006 = n_5993 ^ n_5476;
assign n_6007 = n_5994 ^ n_5993;
assign n_6008 = n_5994 ^ n_5476;
assign n_6009 = n_5996 ^ n_5997;
assign n_6010 = n_5997 ^ x349;
assign n_6011 = n_5998 ^ n_4127;
assign n_6012 = n_5999 ^ n_4551;
assign n_6013 = n_6001 ^ n_5277;
assign n_6014 = n_6002 ^ x367;
assign n_6015 = ~n_6002 & n_6003;
assign n_6016 = n_6004 ^ n_3949;
assign n_6017 = n_6005 ^ n_3949;
assign n_6018 = n_6004 ^ n_6005;
assign n_6019 = n_6006 ^ n_5994;
assign n_6020 = ~n_6007 & ~n_6008;
assign n_6021 = n_6009 ^ x349;
assign n_6022 = n_6009 & ~n_6010;
assign n_6023 = n_6011 ^ n_4168;
assign n_6024 = n_6012 ^ n_4168;
assign n_6025 = n_6011 ^ n_6012;
assign n_6026 = n_5009 ^ n_6013;
assign n_6027 = n_6013 & ~n_5292;
assign n_6028 = n_5987 & ~n_6014;
assign n_6029 = n_6014 ^ n_5987;
assign n_6030 = n_6015 ^ x367;
assign n_6031 = n_6016 ^ n_6005;
assign n_6032 = ~n_6017 & n_6018;
assign n_6033 = ~n_5468 & n_6019;
assign n_6034 = n_6020 ^ n_5476;
assign n_6035 = n_5995 ^ n_6021;
assign n_6036 = n_6021 & n_5995;
assign n_6037 = n_6022 ^ x349;
assign n_6038 = n_6023 ^ n_6012;
assign n_6039 = ~n_6024 & ~n_6025;
assign n_6040 = n_6026 & ~n_5291;
assign n_6041 = n_6026 ^ n_5277;
assign n_6042 = n_5539 ^ n_6026;
assign n_6043 = n_6027 ^ n_5009;
assign n_6044 = n_6030 ^ n_6031;
assign n_6045 = n_6031 ^ x366;
assign n_6046 = n_6032 ^ n_3949;
assign n_6047 = n_6033 ^ n_4825;
assign n_6048 = n_6034 ^ n_5498;
assign n_6049 = n_6035 ^ n_5498;
assign n_6050 = n_6034 ^ n_6035;
assign n_6051 = n_6037 ^ n_6038;
assign n_6052 = n_6038 ^ x348;
assign n_6053 = n_6039 ^ n_4168;
assign n_6054 = n_6040 ^ n_4576;
assign n_6055 = n_6043 ^ n_5319;
assign n_6056 = n_6044 ^ x366;
assign n_6057 = ~n_6044 & n_6045;
assign n_6058 = n_6046 ^ n_3992;
assign n_6059 = n_6047 ^ n_3992;
assign n_6060 = n_6046 ^ n_6047;
assign n_6061 = n_6048 ^ n_6035;
assign n_6062 = n_6049 & n_6050;
assign n_6063 = n_6051 ^ x348;
assign n_6064 = n_6051 & ~n_6052;
assign n_6065 = n_6053 ^ n_4211;
assign n_6066 = n_6054 ^ n_4211;
assign n_6067 = n_6053 ^ n_6054;
assign n_6068 = n_6055 ^ n_5029;
assign n_6069 = ~n_6055 & ~n_5334;
assign n_6070 = n_6028 & ~n_6056;
assign n_6071 = n_6056 ^ n_6028;
assign n_6072 = n_6057 ^ x366;
assign n_6073 = n_6058 ^ n_6047;
assign n_6074 = n_6059 & ~n_6060;
assign n_6075 = n_5492 & n_6061;
assign n_6076 = n_6062 ^ n_5498;
assign n_6077 = n_6036 ^ n_6063;
assign n_6078 = n_6063 & n_6036;
assign n_6079 = n_6064 ^ x348;
assign n_6080 = n_6065 ^ n_6054;
assign n_6081 = n_6066 & ~n_6067;
assign n_6082 = n_6068 & ~n_5333;
assign n_6083 = n_6068 ^ n_5319;
assign n_6084 = n_5558 ^ n_6068;
assign n_6085 = n_6069 ^ n_5029;
assign n_6086 = n_6072 ^ n_6073;
assign n_6087 = n_6073 ^ x365;
assign n_6088 = n_6074 ^ n_3992;
assign n_6089 = n_6075 ^ n_4849;
assign n_6090 = n_6076 ^ n_5511;
assign n_6091 = n_6077 ^ n_5511;
assign n_6092 = n_6076 ^ n_6077;
assign n_6093 = n_6079 ^ n_6080;
assign n_6094 = n_6080 ^ x347;
assign n_6095 = n_6081 ^ n_4211;
assign n_6096 = n_6082 ^ n_4608;
assign n_6097 = n_6085 ^ n_5361;
assign n_6098 = n_6086 ^ x365;
assign n_6099 = n_6086 & ~n_6087;
assign n_6100 = n_6089 ^ n_4035;
assign n_6101 = n_6088 ^ n_6089;
assign n_6102 = n_6090 ^ n_6077;
assign n_6103 = ~n_6091 & ~n_6092;
assign n_6104 = n_6093 ^ x347;
assign n_6105 = n_6093 & ~n_6094;
assign n_6106 = n_6095 ^ n_4254;
assign n_6107 = n_6096 ^ n_4254;
assign n_6108 = n_6095 ^ n_6096;
assign n_6109 = n_6097 ^ n_5050;
assign n_6110 = ~n_6097 & ~n_5376;
assign n_6111 = n_6098 ^ n_6070;
assign n_6112 = n_6070 & n_6098;
assign n_6113 = n_6099 ^ x365;
assign n_6114 = n_6088 ^ n_6100;
assign n_6115 = n_6100 & ~n_6101;
assign n_6116 = ~n_5512 & n_6102;
assign n_6117 = n_6103 ^ n_5511;
assign n_6118 = n_6078 ^ n_6104;
assign n_6119 = n_6104 & n_6078;
assign n_6120 = n_6105 ^ x347;
assign n_6121 = n_6106 ^ n_6096;
assign n_6122 = ~n_6107 & n_6108;
assign n_6123 = ~n_6109 & ~n_5375;
assign n_6124 = n_6109 ^ n_5361;
assign n_6125 = n_5579 ^ n_6109;
assign n_6126 = n_6110 ^ n_5050;
assign n_6127 = n_6111 ^ n_5625;
assign n_6128 = ~n_5625 & ~n_6111;
assign n_6129 = n_6113 ^ n_6114;
assign n_6130 = n_6114 ^ x364;
assign n_6131 = n_6115 ^ n_4035;
assign n_6132 = n_6116 ^ n_4869;
assign n_6133 = n_6117 ^ n_5536;
assign n_6134 = n_6118 ^ n_5536;
assign n_6135 = n_6117 ^ n_6118;
assign n_6136 = n_6120 ^ n_6121;
assign n_6137 = n_6121 ^ x346;
assign n_6138 = n_6122 ^ n_4254;
assign n_6139 = n_6123 ^ n_4640;
assign n_6140 = n_6126 ^ n_5418;
assign n_6141 = n_5617 & n_6127;
assign n_6142 = n_6128 ^ n_5652;
assign n_6143 = n_6129 ^ x364;
assign n_6144 = n_6129 & ~n_6130;
assign n_6145 = n_6131 ^ n_6132;
assign n_6146 = n_6132 ^ n_4079;
assign n_6147 = n_6133 ^ n_6118;
assign n_6148 = ~n_6134 & n_6135;
assign n_6149 = n_6136 ^ x346;
assign n_6150 = ~n_6136 & n_6137;
assign n_6151 = n_6138 ^ n_4296;
assign n_6152 = n_6139 ^ n_4296;
assign n_6153 = n_6139 ^ n_6138;
assign n_6154 = ~n_6140 & n_5405;
assign n_6155 = n_6140 ^ n_5391;
assign n_6156 = n_6141 ^ n_5098;
assign n_6157 = n_6143 ^ n_6112;
assign n_6158 = ~n_6112 & ~n_6143;
assign n_6159 = n_6144 ^ x364;
assign n_6160 = n_6145 ^ n_4079;
assign n_6161 = ~n_6145 & ~n_6146;
assign n_6162 = n_5530 & ~n_6147;
assign n_6163 = n_6148 ^ n_5536;
assign n_6164 = n_6149 ^ n_6119;
assign n_6165 = n_6119 & ~n_6149;
assign n_6166 = n_6150 ^ x346;
assign n_6167 = n_6139 ^ n_6151;
assign n_6168 = ~n_6152 & ~n_6153;
assign n_6169 = n_6154 ^ n_4666;
assign n_6170 = n_6156 ^ n_4562;
assign n_6171 = n_4562 & ~n_6156;
assign n_6172 = n_6157 ^ n_6142;
assign n_6173 = n_6157 ^ n_6128;
assign n_6174 = n_6159 ^ n_6160;
assign n_6175 = n_6160 ^ x363;
assign n_6176 = n_6161 ^ n_4079;
assign n_6177 = n_6162 ^ n_4890;
assign n_6178 = n_6163 ^ n_5555;
assign n_6179 = n_6164 ^ n_5555;
assign n_6180 = n_6163 ^ n_6164;
assign n_6181 = n_6166 ^ n_6167;
assign n_6182 = n_6167 ^ x345;
assign n_6183 = n_6168 ^ n_4296;
assign n_6184 = n_6169 ^ n_4339;
assign n_6185 = x391 & ~n_6170;
assign n_6186 = n_6170 ^ x391;
assign n_6187 = n_6171 ^ n_4591;
assign n_6188 = ~n_5653 & n_6172;
assign n_6189 = n_6142 & ~n_6173;
assign n_6190 = n_6174 ^ x363;
assign n_6191 = ~n_6174 & n_6175;
assign n_6192 = n_6176 ^ n_4120;
assign n_6193 = n_6177 ^ n_4120;
assign n_6194 = n_6176 ^ n_6177;
assign n_6195 = n_6178 ^ n_6164;
assign n_6196 = ~n_6179 & ~n_6180;
assign n_6197 = n_6181 ^ x345;
assign n_6198 = ~n_6181 & n_6182;
assign n_6199 = n_6183 ^ x344;
assign n_6200 = n_6185 ^ x390;
assign n_6201 = n_6188 ^ n_5125;
assign n_6202 = n_6189 ^ n_5652;
assign n_6203 = n_6190 ^ n_6158;
assign n_6204 = ~n_6158 & ~n_6190;
assign n_6205 = n_6191 ^ x363;
assign n_6206 = n_6192 ^ n_6177;
assign n_6207 = ~n_6193 & ~n_6194;
assign n_6208 = ~n_6195 & n_5563;
assign n_6209 = n_6196 ^ n_5555;
assign n_6210 = n_6197 ^ n_6165;
assign n_6211 = n_6165 & ~n_6197;
assign n_6212 = n_6198 ^ x345;
assign n_6213 = n_6199 ^ n_6184;
assign n_6214 = n_6201 ^ n_6187;
assign n_6215 = n_6201 ^ n_6171;
assign n_6216 = n_6202 ^ n_5696;
assign n_6217 = n_6203 ^ n_5696;
assign n_6218 = n_6202 ^ n_6203;
assign n_6219 = n_6205 ^ n_6206;
assign n_6220 = n_6206 ^ x362;
assign n_6221 = n_6207 ^ n_4120;
assign n_6222 = n_6208 ^ n_4912;
assign n_6223 = n_6209 ^ n_5575;
assign n_6224 = n_6210 ^ n_5575;
assign n_6225 = n_6209 ^ n_6210;
assign n_6226 = n_6212 ^ n_6213;
assign n_6227 = n_6214 ^ n_6185;
assign n_6228 = n_6214 ^ n_6200;
assign n_6229 = n_6187 & n_6215;
assign n_6230 = n_6216 ^ n_6203;
assign n_6231 = ~n_6217 & n_6218;
assign n_6232 = n_6219 ^ x362;
assign n_6233 = n_6219 & ~n_6220;
assign n_6234 = n_6221 ^ n_4162;
assign n_6235 = n_6222 ^ n_4162;
assign n_6236 = n_6221 ^ n_6222;
assign n_6237 = n_6223 ^ n_6210;
assign n_6238 = ~n_6224 & n_6225;
assign n_6239 = n_6226 ^ n_6211;
assign n_6240 = n_6200 & n_6227;
assign n_6241 = n_6229 ^ n_4591;
assign n_6242 = ~n_5687 & ~n_6230;
assign n_6243 = n_6231 ^ n_5696;
assign n_6244 = n_6232 ^ n_6204;
assign n_6245 = ~n_6204 & ~n_6232;
assign n_6246 = n_6233 ^ x362;
assign n_6247 = n_6234 ^ n_6222;
assign n_6248 = ~n_6235 & ~n_6236;
assign n_6249 = n_6237 & n_5583;
assign n_6250 = n_6238 ^ n_5575;
assign n_6251 = n_6239 ^ n_5595;
assign n_6252 = n_6240 ^ x390;
assign n_6253 = n_6241 ^ n_4630;
assign n_6254 = n_6242 ^ n_5169;
assign n_6255 = n_6243 ^ n_5732;
assign n_6256 = n_6244 ^ n_5732;
assign n_6257 = n_6243 ^ n_6244;
assign n_6258 = n_6246 ^ x361;
assign n_6259 = n_6247 ^ x361;
assign n_6260 = n_6246 ^ n_6247;
assign n_6261 = n_6248 ^ n_4162;
assign n_6262 = n_6249 ^ n_4933;
assign n_6263 = n_6250 ^ n_6239;
assign n_6264 = n_6253 ^ n_6254;
assign n_6265 = n_6254 ^ n_4630;
assign n_6266 = n_6241 ^ n_6254;
assign n_6267 = n_6255 ^ n_6244;
assign n_6268 = ~n_6256 & ~n_6257;
assign n_6269 = n_6258 ^ n_6247;
assign n_6270 = n_6259 & ~n_6260;
assign n_6271 = n_6261 ^ n_4204;
assign n_6272 = n_6262 ^ n_4204;
assign n_6273 = n_6261 ^ n_6262;
assign n_6274 = n_6263 ^ n_5595;
assign n_6275 = ~n_6263 & ~n_6251;
assign n_6276 = n_6252 ^ n_6264;
assign n_6277 = n_6264 ^ x389;
assign n_6278 = ~n_6265 & n_6266;
assign n_6279 = ~n_5723 & ~n_6267;
assign n_6280 = n_6268 ^ n_5732;
assign n_6281 = n_6269 ^ n_6245;
assign n_6282 = ~n_6245 & ~n_6269;
assign n_6283 = n_6270 ^ x361;
assign n_6284 = n_6271 ^ n_6262;
assign n_6285 = n_6272 & n_6273;
assign n_6286 = n_6274 & n_5603;
assign n_6287 = n_6275 ^ n_5595;
assign n_6288 = n_6276 ^ x389;
assign n_6289 = n_6276 & ~n_6277;
assign n_6290 = n_6278 ^ n_4630;
assign n_6291 = n_6279 ^ n_5208;
assign n_6292 = n_6280 ^ n_5773;
assign n_6293 = n_6281 ^ n_5773;
assign n_6294 = n_6280 ^ n_6281;
assign n_6295 = n_6283 ^ n_6284;
assign n_6296 = n_6284 ^ x360;
assign n_6297 = n_6285 ^ n_4204;
assign n_6298 = n_6286 ^ n_4954;
assign n_6299 = n_6287 ^ n_5135;
assign n_6300 = n_6287 ^ n_5615;
assign n_6301 = ~n_6288 & ~n_6228;
assign n_6302 = n_6228 ^ n_6288;
assign n_6303 = n_6289 ^ x389;
assign n_6304 = n_6290 ^ n_4669;
assign n_6305 = n_6291 ^ n_4669;
assign n_6306 = n_6290 ^ n_6291;
assign n_6307 = n_6292 ^ n_6281;
assign n_6308 = ~n_6293 & ~n_6294;
assign n_6309 = n_6295 ^ x360;
assign n_6310 = ~n_6295 & n_6296;
assign n_6311 = n_6297 ^ n_6298;
assign n_6312 = n_6298 ^ n_4247;
assign n_6313 = n_6299 ^ n_5615;
assign n_6314 = ~n_5623 & ~n_6300;
assign n_6315 = n_6304 ^ n_6291;
assign n_6316 = ~n_6305 & ~n_6306;
assign n_6317 = n_5761 & n_6307;
assign n_6318 = n_6308 ^ n_5773;
assign n_6319 = n_6309 ^ n_6282;
assign n_6320 = n_6282 & ~n_6309;
assign n_6321 = n_6310 ^ x360;
assign n_6322 = n_6311 ^ n_4247;
assign n_6323 = n_6311 & n_6312;
assign n_6324 = ~n_5609 & ~n_6313;
assign n_6325 = n_6314 ^ n_5135;
assign n_6326 = n_6303 ^ n_6315;
assign n_6327 = n_6315 ^ x388;
assign n_6328 = n_6316 ^ n_4669;
assign n_6329 = n_6317 ^ n_5248;
assign n_6330 = n_6318 ^ n_5812;
assign n_6331 = n_6319 ^ n_5812;
assign n_6332 = n_6318 ^ n_6319;
assign n_6333 = n_6321 ^ n_6322;
assign n_6334 = n_6322 ^ x375;
assign n_6335 = n_6323 ^ n_4247;
assign n_6336 = n_6324 ^ n_4976;
assign n_6337 = n_6325 ^ n_5192;
assign n_6338 = n_6325 ^ n_5638;
assign n_6339 = n_6326 ^ x388;
assign n_6340 = n_6326 & ~n_6327;
assign n_6341 = n_6328 ^ n_4705;
assign n_6342 = n_6329 ^ n_4705;
assign n_6343 = n_6328 ^ n_6329;
assign n_6344 = n_6330 ^ n_6319;
assign n_6345 = n_6331 & ~n_6332;
assign n_6346 = n_6333 ^ x375;
assign n_6347 = n_6333 & ~n_6334;
assign n_6348 = n_6335 ^ n_6336;
assign n_6349 = n_6336 ^ n_4289;
assign n_6350 = n_6337 ^ n_5638;
assign n_6351 = ~n_5648 & n_6338;
assign n_6352 = n_6301 & ~n_6339;
assign n_6353 = n_6339 ^ n_6301;
assign n_6354 = n_6340 ^ x388;
assign n_6355 = n_6341 ^ n_6329;
assign n_6356 = n_6342 & n_6343;
assign n_6357 = ~n_5801 & n_6344;
assign n_6358 = n_6345 ^ n_5812;
assign n_6359 = n_6320 ^ n_6346;
assign n_6360 = ~n_6346 & ~n_6320;
assign n_6361 = n_6347 ^ x375;
assign n_6362 = n_6348 ^ n_4289;
assign n_6363 = n_6348 & ~n_6349;
assign n_6364 = n_6350 & n_5647;
assign n_6365 = n_6351 ^ n_5192;
assign n_6366 = n_6354 ^ n_6355;
assign n_6367 = n_6355 ^ x387;
assign n_6368 = n_6356 ^ n_4705;
assign n_6369 = n_6357 ^ n_5286;
assign n_6370 = n_6358 ^ n_5854;
assign n_6371 = n_6359 ^ n_6358;
assign n_6372 = n_6359 ^ n_5854;
assign n_6373 = n_6361 ^ n_6362;
assign n_6374 = n_6362 ^ x374;
assign n_6375 = n_6363 ^ n_4289;
assign n_6376 = n_6364 ^ n_4996;
assign n_6377 = n_6365 ^ n_5669;
assign n_6378 = n_6366 ^ x387;
assign n_6379 = n_6366 & ~n_6367;
assign n_6380 = n_6368 ^ n_4733;
assign n_6381 = n_6369 ^ n_4733;
assign n_6382 = n_6368 ^ n_6369;
assign n_6383 = n_6370 ^ n_6359;
assign n_6384 = ~n_6371 & ~n_6372;
assign n_6385 = n_6373 ^ x374;
assign n_6386 = n_6373 & ~n_6374;
assign n_6387 = n_6375 ^ n_4332;
assign n_6388 = n_6376 ^ n_4332;
assign n_6389 = n_6375 ^ n_6376;
assign n_6390 = n_5244 ^ n_6377;
assign n_6391 = ~n_6377 & ~n_5681;
assign n_6392 = ~n_6378 & n_6352;
assign n_6393 = n_6352 ^ n_6378;
assign n_6394 = n_6379 ^ x387;
assign n_6395 = n_6380 ^ n_6369;
assign n_6396 = ~n_6381 & n_6382;
assign n_6397 = n_5843 & ~n_6383;
assign n_6398 = n_6384 ^ n_5854;
assign n_6399 = n_6385 ^ n_6360;
assign n_6400 = n_6360 & ~n_6385;
assign n_6401 = n_6386 ^ x374;
assign n_6402 = n_6387 ^ n_6376;
assign n_6403 = ~n_6388 & ~n_6389;
assign n_6404 = n_6390 & n_5680;
assign n_6405 = n_6390 ^ n_5669;
assign n_6406 = n_6391 ^ n_5244;
assign n_6407 = n_6394 ^ n_6395;
assign n_6408 = n_6395 ^ x386;
assign n_6409 = n_6396 ^ n_4733;
assign n_6410 = n_6397 ^ n_5328;
assign n_6411 = n_6398 ^ n_5897;
assign n_6412 = n_6399 ^ n_5897;
assign n_6413 = n_6398 ^ n_6399;
assign n_6414 = n_6401 ^ n_6402;
assign n_6415 = n_6402 ^ x373;
assign n_6416 = n_6403 ^ n_4332;
assign n_6417 = n_6404 ^ n_5016;
assign n_6418 = n_6406 ^ n_5298;
assign n_6419 = n_6406 ^ n_5703;
assign n_6420 = n_6407 ^ x386;
assign n_6421 = n_6407 & ~n_6408;
assign n_6422 = n_6409 ^ n_4756;
assign n_6423 = n_6410 ^ n_4756;
assign n_6424 = n_6409 ^ n_6410;
assign n_6425 = n_6411 ^ n_6399;
assign n_6426 = ~n_6412 & ~n_6413;
assign n_6427 = n_6414 ^ x373;
assign n_6428 = n_6414 & ~n_6415;
assign n_6429 = n_6416 ^ n_4373;
assign n_6430 = n_6417 ^ n_4373;
assign n_6431 = n_6416 ^ n_6417;
assign n_6432 = n_6418 ^ n_5703;
assign n_6433 = ~n_5716 & ~n_6419;
assign n_6434 = ~n_6392 & n_6420;
assign n_6435 = n_6420 ^ n_6392;
assign n_6436 = n_6421 ^ x386;
assign n_6437 = n_6422 ^ n_6410;
assign n_6438 = ~n_6423 & n_6424;
assign n_6439 = ~n_5885 & n_6425;
assign n_6440 = n_6186 ^ n_6425;
assign n_6441 = n_6426 ^ n_5897;
assign n_6442 = n_6400 ^ n_6427;
assign n_6443 = n_6427 & ~n_6400;
assign n_6444 = n_6428 ^ x373;
assign n_6445 = n_6429 ^ n_6417;
assign n_6446 = n_6430 & ~n_6431;
assign n_6447 = ~n_6432 & n_5715;
assign n_6448 = n_6433 ^ n_5298;
assign n_6449 = n_6436 ^ n_6437;
assign n_6450 = n_6437 ^ x385;
assign n_6451 = n_6438 ^ n_4756;
assign n_6452 = n_6439 ^ n_5370;
assign n_6453 = n_6441 ^ n_5937;
assign n_6454 = n_6441 ^ n_6442;
assign n_6455 = n_6442 ^ n_5937;
assign n_6456 = n_6444 ^ n_6445;
assign n_6457 = n_6445 ^ x372;
assign n_6458 = n_6446 ^ n_4373;
assign n_6459 = n_6447 ^ n_5037;
assign n_6460 = n_6448 ^ n_5739;
assign n_6461 = n_6449 ^ x385;
assign n_6462 = n_6449 & ~n_6450;
assign n_6463 = n_6451 ^ n_4773;
assign n_6464 = n_6452 ^ n_4773;
assign n_6465 = n_6451 ^ n_6452;
assign n_6466 = n_6453 ^ n_6442;
assign n_6467 = ~n_6454 & n_6455;
assign n_6468 = n_6456 ^ x372;
assign n_6469 = n_6456 & ~n_6457;
assign n_6470 = n_6458 ^ n_4403;
assign n_6471 = n_6459 ^ n_4403;
assign n_6472 = n_6458 ^ n_6459;
assign n_6473 = n_5339 ^ n_6460;
assign n_6474 = n_6460 & n_5753;
assign n_6475 = ~n_6434 & ~n_6461;
assign n_6476 = n_6461 ^ n_6434;
assign n_6477 = n_6462 ^ x385;
assign n_6478 = n_6463 ^ n_6452;
assign n_6479 = n_6464 & n_6465;
assign n_6480 = ~n_5926 & n_6466;
assign n_6481 = n_6228 ^ n_6466;
assign n_6482 = n_6467 ^ n_5937;
assign n_6483 = n_6468 ^ n_6443;
assign n_6484 = n_6443 & n_6468;
assign n_6485 = n_6469 ^ x372;
assign n_6486 = n_6470 ^ n_6459;
assign n_6487 = n_6471 & n_6472;
assign n_6488 = ~n_6473 & ~n_5752;
assign n_6489 = n_6473 ^ n_5739;
assign n_6490 = n_6474 ^ n_5339;
assign n_6491 = n_6477 ^ n_6478;
assign n_6492 = n_6478 ^ x384;
assign n_6493 = n_6479 ^ n_4773;
assign n_6494 = n_6480 ^ n_5413;
assign n_6495 = n_6482 ^ n_5979;
assign n_6496 = n_6483 ^ n_5979;
assign n_6497 = n_6482 ^ n_6483;
assign n_6498 = n_6485 ^ n_6486;
assign n_6499 = n_6486 ^ x371;
assign n_6500 = n_6487 ^ n_4403;
assign n_6501 = n_6488 ^ n_5058;
assign n_6502 = n_6490 ^ n_5780;
assign n_6503 = n_6491 ^ x384;
assign n_6504 = ~n_6491 & n_6492;
assign n_6505 = n_6493 ^ n_4792;
assign n_6506 = n_6494 ^ n_4792;
assign n_6507 = n_6493 ^ n_6494;
assign n_6508 = n_6495 ^ n_6483;
assign n_6509 = ~n_6496 & n_6497;
assign n_6510 = n_6498 ^ x371;
assign n_6511 = n_6498 & ~n_6499;
assign n_6512 = n_6500 ^ n_6501;
assign n_6513 = n_6501 ^ n_4426;
assign n_6514 = n_5381 ^ n_6502;
assign n_6515 = ~n_6502 & ~n_5793;
assign n_6516 = n_6503 & n_6475;
assign n_6517 = n_6475 ^ n_6503;
assign n_6518 = n_6504 ^ x384;
assign n_6519 = n_6505 ^ n_6494;
assign n_6520 = n_6506 & ~n_6507;
assign n_6521 = ~n_5967 & ~n_6508;
assign n_6522 = n_6302 ^ n_6508;
assign n_6523 = n_6509 ^ n_5979;
assign n_6524 = n_6484 ^ n_6510;
assign n_6525 = n_6510 & n_6484;
assign n_6526 = n_6511 ^ x371;
assign n_6527 = n_6512 ^ n_4426;
assign n_6528 = n_6512 & ~n_6513;
assign n_6529 = ~n_6514 & n_5792;
assign n_6530 = n_6514 ^ n_5780;
assign n_6531 = n_5660 ^ n_6514;
assign n_6532 = n_6515 ^ n_5381;
assign n_6533 = n_6518 ^ n_6519;
assign n_6534 = n_6519 ^ x399;
assign n_6535 = n_6520 ^ n_4792;
assign n_6536 = n_6521 ^ n_5448;
assign n_6537 = n_6523 ^ n_6019;
assign n_6538 = n_6524 ^ n_6019;
assign n_6539 = n_6523 ^ n_6524;
assign n_6540 = n_6526 ^ n_6527;
assign n_6541 = n_6527 ^ x370;
assign n_6542 = n_6528 ^ n_4426;
assign n_6543 = n_6529 ^ n_5078;
assign n_6544 = n_6532 ^ n_5819;
assign n_6545 = n_6533 ^ x399;
assign n_6546 = n_6533 & ~n_6534;
assign n_6547 = n_6535 ^ n_4810;
assign n_6548 = n_6536 ^ n_4810;
assign n_6549 = n_6535 ^ n_6536;
assign n_6550 = n_6537 ^ n_6524;
assign n_6551 = ~n_6538 & n_6539;
assign n_6552 = n_6540 ^ x370;
assign n_6553 = n_6540 & ~n_6541;
assign n_6554 = n_6542 ^ n_4440;
assign n_6555 = n_6543 ^ n_4440;
assign n_6556 = n_6542 ^ n_6543;
assign n_6557 = n_5422 ^ n_6544;
assign n_6558 = ~n_6544 & ~n_5835;
assign n_6559 = n_6545 & ~n_6516;
assign n_6560 = n_6516 ^ n_6545;
assign n_6561 = n_6546 ^ x399;
assign n_6562 = n_6547 ^ n_6536;
assign n_6563 = ~n_6548 & ~n_6549;
assign n_6564 = n_6007 & ~n_6550;
assign n_6565 = n_6353 ^ n_6550;
assign n_6566 = n_6551 ^ n_6019;
assign n_6567 = n_6525 ^ n_6552;
assign n_6568 = ~n_6552 & ~n_6525;
assign n_6569 = n_6553 ^ x370;
assign n_6570 = n_6554 ^ n_6543;
assign n_6571 = n_6555 & ~n_6556;
assign n_6572 = n_6557 & ~n_5834;
assign n_6573 = n_6557 ^ n_5819;
assign n_6574 = n_6557 ^ n_5694;
assign n_6575 = n_6558 ^ n_5422;
assign n_6576 = n_6561 ^ n_6562;
assign n_6577 = n_6562 ^ x398;
assign n_6578 = n_6563 ^ n_4810;
assign n_6579 = n_6564 ^ n_5476;
assign n_6580 = n_6566 ^ n_6061;
assign n_6581 = n_6567 ^ n_6061;
assign n_6582 = n_6566 ^ n_6567;
assign n_6583 = n_6569 ^ n_6570;
assign n_6584 = n_6570 ^ x369;
assign n_6585 = n_6571 ^ n_4440;
assign n_6586 = n_6572 ^ n_5101;
assign n_6587 = n_6575 ^ n_5861;
assign n_6588 = n_6576 ^ x398;
assign n_6589 = ~n_6576 & n_6577;
assign n_6590 = n_6578 ^ n_4825;
assign n_6591 = n_6579 ^ n_4825;
assign n_6592 = n_6578 ^ n_6579;
assign n_6593 = n_6580 ^ n_6567;
assign n_6594 = n_6581 & ~n_6582;
assign n_6595 = n_6583 ^ x369;
assign n_6596 = ~n_6583 & n_6584;
assign n_6597 = n_6585 ^ n_6586;
assign n_6598 = n_6586 ^ n_4466;
assign n_6599 = n_5454 ^ n_6587;
assign n_6600 = n_6587 & ~n_5877;
assign n_6601 = ~n_6559 & n_6588;
assign n_6602 = n_6588 ^ n_6559;
assign n_6603 = n_6589 ^ x398;
assign n_6604 = n_6590 ^ n_6579;
assign n_6605 = ~n_6591 & ~n_6592;
assign n_6606 = ~n_6050 & n_6593;
assign n_6607 = n_6393 ^ n_6593;
assign n_6608 = n_6594 ^ n_6061;
assign n_6609 = n_6595 ^ n_6568;
assign n_6610 = ~n_6568 & ~n_6595;
assign n_6611 = n_6596 ^ x369;
assign n_6612 = n_6597 ^ n_4466;
assign n_6613 = ~n_6597 & n_6598;
assign n_6614 = ~n_6599 & ~n_5876;
assign n_6615 = n_6599 ^ n_5768;
assign n_6616 = n_6599 ^ n_5861;
assign n_6617 = n_6600 ^ n_5454;
assign n_6618 = n_6603 ^ n_6604;
assign n_6619 = n_6604 ^ x397;
assign n_6620 = n_6605 ^ n_4825;
assign n_6621 = n_6606 ^ n_5498;
assign n_6622 = n_6608 ^ n_6102;
assign n_6623 = n_6609 ^ n_6102;
assign n_6624 = n_6608 ^ n_6609;
assign n_6625 = n_6611 ^ n_6612;
assign n_6626 = n_6612 ^ x368;
assign n_6627 = n_6613 ^ n_4466;
assign n_6628 = n_6614 ^ n_5129;
assign n_6629 = n_6617 ^ n_5480;
assign n_6630 = n_6617 ^ n_5903;
assign n_6631 = n_6618 ^ x397;
assign n_6632 = n_6618 & ~n_6619;
assign n_6633 = n_6620 ^ n_4849;
assign n_6634 = n_6621 ^ n_4849;
assign n_6635 = n_6620 ^ n_6621;
assign n_6636 = n_6622 ^ n_6609;
assign n_6637 = ~n_6623 & n_6624;
assign n_6638 = n_6625 ^ x368;
assign n_6639 = ~n_6625 & n_6626;
assign n_6640 = n_6627 ^ n_6628;
assign n_6641 = n_6628 ^ n_4487;
assign n_6642 = n_6629 ^ n_5903;
assign n_6643 = ~n_5918 & n_6630;
assign n_6644 = ~n_6631 & n_6601;
assign n_6645 = n_6601 ^ n_6631;
assign n_6646 = n_6632 ^ x397;
assign n_6647 = n_6633 ^ n_6621;
assign n_6648 = n_6634 & ~n_6635;
assign n_6649 = n_6092 & ~n_6636;
assign n_6650 = n_6435 ^ n_6636;
assign n_6651 = n_6637 ^ n_6102;
assign n_6652 = n_6638 ^ n_6610;
assign n_6653 = ~n_6610 & n_6638;
assign n_6654 = n_6639 ^ x368;
assign n_6655 = n_6640 ^ n_4487;
assign n_6656 = ~n_6640 & n_6641;
assign n_6657 = n_5890 & ~n_6642;
assign n_6658 = n_5822 ^ n_6642;
assign n_6659 = n_6643 ^ n_5480;
assign n_6660 = n_6646 ^ n_6647;
assign n_6661 = n_6647 ^ x396;
assign n_6662 = n_6648 ^ n_4849;
assign n_6663 = n_6649 ^ n_5511;
assign n_6664 = n_6651 ^ n_6147;
assign n_6665 = n_6652 ^ n_6147;
assign n_6666 = n_6651 ^ n_6652;
assign n_6667 = n_6654 ^ n_6655;
assign n_6668 = n_6655 ^ x383;
assign n_6669 = n_6656 ^ n_4487;
assign n_6670 = n_6657 ^ n_5164;
assign n_6671 = n_6659 ^ n_5943;
assign n_6672 = n_6660 ^ x396;
assign n_6673 = n_6660 & ~n_6661;
assign n_6674 = n_6662 ^ n_4869;
assign n_6675 = n_6663 ^ n_4869;
assign n_6676 = n_6662 ^ n_6663;
assign n_6677 = n_6664 ^ n_6652;
assign n_6678 = n_6665 & n_6666;
assign n_6679 = n_6667 ^ x383;
assign n_6680 = ~n_6667 & n_6668;
assign n_6681 = n_6669 ^ n_6670;
assign n_6682 = n_6670 ^ n_4508;
assign n_6683 = n_5501 ^ n_6671;
assign n_6684 = n_6671 & n_5959;
assign n_6685 = n_6644 & ~n_6672;
assign n_6686 = n_6672 ^ n_6644;
assign n_6687 = n_6673 ^ x396;
assign n_6688 = n_6674 ^ n_6663;
assign n_6689 = ~n_6675 & n_6676;
assign n_6690 = ~n_6135 & n_6677;
assign n_6691 = n_6476 ^ n_6677;
assign n_6692 = n_6678 ^ n_6147;
assign n_6693 = n_6679 ^ n_6653;
assign n_6694 = ~n_6653 & ~n_6679;
assign n_6695 = n_6680 ^ x383;
assign n_6696 = n_6681 ^ n_4508;
assign n_6697 = n_6681 & n_6682;
assign n_6698 = n_6683 & n_5958;
assign n_6699 = n_6683 ^ n_5943;
assign n_6700 = n_5864 ^ n_6683;
assign n_6701 = n_6684 ^ n_5501;
assign n_6702 = n_6687 ^ n_6688;
assign n_6703 = n_6688 ^ x395;
assign n_6704 = n_6689 ^ n_4869;
assign n_6705 = n_6690 ^ n_5536;
assign n_6706 = n_6692 ^ n_6195;
assign n_6707 = n_6693 ^ n_6195;
assign n_6708 = n_6692 ^ n_6693;
assign n_6709 = n_6695 ^ n_6696;
assign n_6710 = n_6696 ^ x382;
assign n_6711 = n_6697 ^ n_4508;
assign n_6712 = n_6698 ^ n_5200;
assign n_6713 = n_6701 ^ n_5985;
assign n_6714 = n_6702 ^ x395;
assign n_6715 = ~n_6702 & n_6703;
assign n_6716 = n_6704 ^ n_4890;
assign n_6717 = n_6705 ^ n_4890;
assign n_6718 = n_6704 ^ n_6705;
assign n_6719 = n_6706 ^ n_6693;
assign n_6720 = n_6707 & ~n_6708;
assign n_6721 = n_6709 ^ x382;
assign n_6722 = ~n_6709 & n_6710;
assign n_6723 = n_6711 ^ n_6712;
assign n_6724 = n_6712 ^ n_4528;
assign n_6725 = n_5521 ^ n_6713;
assign n_6726 = ~n_6713 & n_6000;
assign n_6727 = ~n_6685 & ~n_6714;
assign n_6728 = n_6714 ^ n_6685;
assign n_6729 = n_6715 ^ x395;
assign n_6730 = n_6716 ^ n_6705;
assign n_6731 = n_6717 & n_6718;
assign n_6732 = n_6180 & ~n_6719;
assign n_6733 = n_6517 ^ n_6719;
assign n_6734 = n_6720 ^ n_6195;
assign n_6735 = n_6694 ^ n_6721;
assign n_6736 = n_6721 & ~n_6694;
assign n_6737 = n_6722 ^ x382;
assign n_6738 = n_6723 ^ n_4528;
assign n_6739 = ~n_6723 & ~n_6724;
assign n_6740 = n_5972 & ~n_6725;
assign n_6741 = n_6725 ^ n_5985;
assign n_6742 = n_5906 ^ n_6725;
assign n_6743 = n_6726 ^ n_5521;
assign n_6744 = n_6729 ^ n_6730;
assign n_6745 = n_6730 ^ x394;
assign n_6746 = n_6731 ^ n_4890;
assign n_6747 = n_6732 ^ n_5555;
assign n_6748 = n_6734 ^ n_6237;
assign n_6749 = n_6734 ^ n_6735;
assign n_6750 = n_6735 ^ n_6237;
assign n_6751 = n_6737 ^ n_6738;
assign n_6752 = n_6738 ^ x381;
assign n_6753 = n_6739 ^ n_4528;
assign n_6754 = n_6740 ^ n_5238;
assign n_6755 = n_6743 ^ n_6026;
assign n_6756 = n_6744 ^ x394;
assign n_6757 = n_6744 & ~n_6745;
assign n_6758 = n_6746 ^ n_4912;
assign n_6759 = n_6747 ^ n_4912;
assign n_6760 = n_6746 ^ n_6747;
assign n_6761 = n_6748 ^ n_6735;
assign n_6762 = ~n_6749 & ~n_6750;
assign n_6763 = n_6751 ^ x381;
assign n_6764 = ~n_6751 & n_6752;
assign n_6765 = n_6753 ^ n_6754;
assign n_6766 = n_6754 ^ n_4551;
assign n_6767 = n_5539 ^ n_6755;
assign n_6768 = n_6755 & ~n_6042;
assign n_6769 = ~n_6727 & ~n_6756;
assign n_6770 = n_6756 ^ n_6727;
assign n_6771 = n_6757 ^ x394;
assign n_6772 = n_6758 ^ n_6747;
assign n_6773 = n_6759 & n_6760;
assign n_6774 = ~n_6225 & n_6761;
assign n_6775 = n_6560 ^ n_6761;
assign n_6776 = n_6762 ^ n_6237;
assign n_6777 = n_6763 ^ n_6736;
assign n_6778 = n_6736 & n_6763;
assign n_6779 = n_6764 ^ x381;
assign n_6780 = n_6765 ^ n_4551;
assign n_6781 = n_6765 & ~n_6766;
assign n_6782 = n_6767 & n_6041;
assign n_6783 = n_6767 ^ n_6026;
assign n_6784 = n_5946 ^ n_6767;
assign n_6785 = n_6768 ^ n_5539;
assign n_6786 = n_6771 ^ n_6772;
assign n_6787 = n_6772 ^ x393;
assign n_6788 = n_6773 ^ n_4912;
assign n_6789 = n_6774 ^ n_5575;
assign n_6790 = n_6776 ^ n_6274;
assign n_6791 = n_6777 ^ n_6274;
assign n_6792 = n_6776 ^ n_6777;
assign n_6793 = n_6779 ^ n_6780;
assign n_6794 = n_6780 ^ x380;
assign n_6795 = n_6781 ^ n_4551;
assign n_6796 = n_6782 ^ n_5277;
assign n_6797 = n_6785 ^ n_6068;
assign n_6798 = n_6786 ^ x393;
assign n_6799 = ~n_6786 & n_6787;
assign n_6800 = n_6788 ^ n_4933;
assign n_6801 = n_6789 ^ n_4933;
assign n_6802 = n_6788 ^ n_6789;
assign n_6803 = n_6790 ^ n_6777;
assign n_6804 = n_6791 & ~n_6792;
assign n_6805 = n_6793 ^ x380;
assign n_6806 = n_6793 & ~n_6794;
assign n_6807 = n_6795 ^ n_4576;
assign n_6808 = n_6796 ^ n_4576;
assign n_6809 = n_6795 ^ n_6796;
assign n_6810 = n_6797 ^ n_5558;
assign n_6811 = n_6797 & ~n_6084;
assign n_6812 = n_6769 & n_6798;
assign n_6813 = n_6798 ^ n_6769;
assign n_6814 = n_6799 ^ x393;
assign n_6815 = n_6800 ^ n_6789;
assign n_6816 = n_6801 & ~n_6802;
assign n_6817 = n_6263 & n_6803;
assign n_6818 = n_6602 ^ n_6803;
assign n_6819 = n_6804 ^ n_6274;
assign n_6820 = n_6778 ^ n_6805;
assign n_6821 = n_6805 & ~n_6778;
assign n_6822 = n_6806 ^ x380;
assign n_6823 = n_6807 ^ n_6796;
assign n_6824 = ~n_6808 & ~n_6809;
assign n_6825 = n_6810 & ~n_6083;
assign n_6826 = n_6810 ^ n_6068;
assign n_6827 = n_6810 ^ n_5988;
assign n_6828 = n_6811 ^ n_5558;
assign n_6829 = n_6814 ^ n_6815;
assign n_6830 = n_6815 ^ x392;
assign n_6831 = n_6816 ^ n_4933;
assign n_6832 = n_6817 ^ n_5595;
assign n_6833 = n_6819 ^ n_6313;
assign n_6834 = n_6820 ^ n_6313;
assign n_6835 = n_6819 ^ n_6820;
assign n_6836 = n_6822 ^ n_6823;
assign n_6837 = n_6823 ^ x379;
assign n_6838 = n_6824 ^ n_4576;
assign n_6839 = n_6825 ^ n_5319;
assign n_6840 = n_6828 ^ n_6109;
assign n_6841 = n_6829 ^ x392;
assign n_6842 = n_6829 & ~n_6830;
assign n_6843 = n_6831 ^ n_6832;
assign n_6844 = n_6832 ^ n_4954;
assign n_6845 = n_6833 ^ n_6820;
assign n_6846 = ~n_6834 & ~n_6835;
assign n_6847 = n_6836 ^ x379;
assign n_6848 = n_6836 & ~n_6837;
assign n_6849 = n_6838 ^ n_4608;
assign n_6850 = n_6839 ^ n_4608;
assign n_6851 = n_6838 ^ n_6839;
assign n_6852 = n_6840 ^ n_5579;
assign n_6853 = ~n_6840 & ~n_6125;
assign n_6854 = n_6812 & ~n_6841;
assign n_6855 = n_6841 ^ n_6812;
assign n_6856 = n_6842 ^ x392;
assign n_6857 = n_6843 ^ n_4954;
assign n_6858 = n_6843 & n_6844;
assign n_6859 = ~n_6299 & ~n_6845;
assign n_6860 = n_6645 ^ n_6845;
assign n_6861 = n_6846 ^ n_6313;
assign n_6862 = n_6847 ^ n_6821;
assign n_6863 = ~n_6821 & ~n_6847;
assign n_6864 = n_6848 ^ x379;
assign n_6865 = n_6849 ^ n_6839;
assign n_6866 = ~n_6850 & ~n_6851;
assign n_6867 = n_6852 & ~n_6124;
assign n_6868 = n_6852 ^ n_6109;
assign n_6869 = n_6029 ^ n_6852;
assign n_6870 = n_6853 ^ n_5579;
assign n_6871 = n_6856 ^ n_6857;
assign n_6872 = n_6857 ^ x407;
assign n_6873 = n_6858 ^ n_4954;
assign n_6874 = n_6859 ^ n_5615;
assign n_6875 = n_6861 ^ n_6350;
assign n_6876 = n_6862 ^ n_6350;
assign n_6877 = n_6861 ^ n_6862;
assign n_6878 = n_6864 ^ n_6865;
assign n_6879 = n_6865 ^ x378;
assign n_6880 = n_6866 ^ n_4608;
assign n_6881 = n_6867 ^ n_5361;
assign n_6882 = n_6870 ^ n_6140;
assign n_6883 = n_6871 ^ x407;
assign n_6884 = n_6871 & ~n_6872;
assign n_6885 = n_6873 ^ n_6874;
assign n_6886 = n_6874 ^ n_4976;
assign n_6887 = n_6875 ^ n_6862;
assign n_6888 = n_6876 & n_6877;
assign n_6889 = n_6878 ^ x378;
assign n_6890 = ~n_6878 & n_6879;
assign n_6891 = n_6880 ^ n_4640;
assign n_6892 = n_6881 ^ n_4640;
assign n_6893 = n_6881 ^ n_6880;
assign n_6894 = n_6882 ^ n_5598;
assign n_6895 = n_6854 & ~n_6883;
assign n_6896 = n_6883 ^ n_6854;
assign n_6897 = n_6884 ^ x407;
assign n_6898 = n_6885 ^ n_4976;
assign n_6899 = ~n_6885 & ~n_6886;
assign n_6900 = n_6337 & ~n_6887;
assign n_6901 = n_6686 ^ n_6887;
assign n_6902 = n_6888 ^ n_6350;
assign n_6903 = n_6889 ^ n_6863;
assign n_6904 = n_6863 & n_6889;
assign n_6905 = n_6890 ^ x378;
assign n_6906 = n_6881 ^ n_6891;
assign n_6907 = ~n_6892 & ~n_6893;
assign n_6908 = n_6894 & n_6155;
assign n_6909 = n_6071 ^ n_6894;
assign n_6910 = n_6894 ^ n_6140;
assign n_6911 = n_6897 ^ n_6898;
assign n_6912 = n_6898 ^ x406;
assign n_6913 = n_6899 ^ n_4976;
assign n_6914 = n_6900 ^ n_5638;
assign n_6915 = n_6902 ^ n_6390;
assign n_6916 = n_6903 ^ n_6390;
assign n_6917 = n_6902 ^ n_6903;
assign n_6918 = n_6905 ^ n_6906;
assign n_6919 = n_6906 ^ x377;
assign n_6920 = n_6907 ^ n_4640;
assign n_6921 = n_6908 ^ n_5391;
assign n_6922 = n_6911 ^ x406;
assign n_6923 = n_6911 & ~n_6912;
assign n_6924 = n_6913 ^ n_4996;
assign n_6925 = n_6914 ^ n_6913;
assign n_6926 = n_6915 ^ n_6903;
assign n_6927 = n_6916 & ~n_6917;
assign n_6928 = n_6918 ^ x377;
assign n_6929 = n_6918 & ~n_6919;
assign n_6930 = n_6920 ^ x376;
assign n_6931 = n_6921 ^ n_4666;
assign n_6932 = n_6895 & ~n_6922;
assign n_6933 = n_6922 ^ n_6895;
assign n_6934 = n_6923 ^ x406;
assign n_6935 = n_6914 ^ n_6924;
assign n_6936 = ~n_6924 & n_6925;
assign n_6937 = n_6926 & ~n_6405;
assign n_6938 = n_6728 ^ n_6926;
assign n_6939 = n_6927 ^ n_6390;
assign n_6940 = n_6928 ^ n_6904;
assign n_6941 = n_6904 & ~n_6928;
assign n_6942 = n_6929 ^ x377;
assign n_6943 = n_6930 ^ n_6931;
assign n_6944 = n_6934 ^ n_6935;
assign n_6945 = n_6935 ^ x405;
assign n_6946 = n_6936 ^ n_4996;
assign n_6947 = n_6937 ^ n_5669;
assign n_6948 = n_6939 ^ n_6432;
assign n_6949 = n_6940 ^ n_6432;
assign n_6950 = n_6939 ^ n_6940;
assign n_6951 = n_6942 ^ n_6943;
assign n_6952 = n_6944 ^ x405;
assign n_6953 = n_6944 & ~n_6945;
assign n_6954 = n_6946 ^ n_5016;
assign n_6955 = n_6947 ^ n_5016;
assign n_6956 = n_6946 ^ n_6947;
assign n_6957 = n_6948 ^ n_6940;
assign n_6958 = n_6949 & n_6950;
assign n_6959 = n_6951 ^ n_6941;
assign n_6960 = n_6932 & ~n_6952;
assign n_6961 = n_6952 ^ n_6932;
assign n_6962 = n_6953 ^ x405;
assign n_6963 = n_6954 ^ n_6947;
assign n_6964 = n_6955 & n_6956;
assign n_6965 = ~n_6418 & n_6957;
assign n_6966 = n_6770 ^ n_6957;
assign n_6967 = n_6958 ^ n_6432;
assign n_6968 = n_6959 ^ n_6473;
assign n_6969 = n_6962 ^ n_6963;
assign n_6970 = n_6963 ^ x404;
assign n_6971 = n_6964 ^ n_5016;
assign n_6972 = n_6965 ^ n_5703;
assign n_6973 = n_6967 ^ n_6473;
assign n_6974 = n_6967 ^ n_6959;
assign n_6975 = n_6969 ^ x404;
assign n_6976 = ~n_6969 & n_6970;
assign n_6977 = n_6971 ^ n_5037;
assign n_6978 = n_6972 ^ n_5037;
assign n_6979 = n_6971 ^ n_6972;
assign n_6980 = n_6973 ^ n_6959;
assign n_6981 = ~n_6968 & n_6974;
assign n_6982 = n_6960 & n_6975;
assign n_6983 = n_6975 ^ n_6960;
assign n_6984 = n_6976 ^ x404;
assign n_6985 = n_6977 ^ n_6972;
assign n_6986 = n_6978 & n_6979;
assign n_6987 = n_6980 & ~n_6489;
assign n_6988 = n_6813 ^ n_6980;
assign n_6989 = n_6981 ^ n_6473;
assign n_6990 = n_6984 ^ n_6985;
assign n_6991 = n_6985 ^ x403;
assign n_6992 = n_6986 ^ n_5037;
assign n_6993 = n_6987 ^ n_5739;
assign n_6994 = n_6989 ^ n_6514;
assign n_6995 = n_6990 ^ x403;
assign n_6996 = n_6990 & ~n_6991;
assign n_6997 = n_6992 ^ n_5058;
assign n_6998 = n_6993 ^ n_5058;
assign n_6999 = n_6992 ^ n_6993;
assign n_7000 = n_5660 ^ n_6994;
assign n_7001 = ~n_6994 & n_6531;
assign n_7002 = ~n_6982 & n_6995;
assign n_7003 = n_6995 ^ n_6982;
assign n_7004 = n_6996 ^ x403;
assign n_7005 = n_6997 ^ n_6993;
assign n_7006 = ~n_6998 & ~n_6999;
assign n_7007 = ~n_7000 & ~n_6530;
assign n_7008 = n_7000 ^ n_6514;
assign n_7009 = n_6855 ^ n_7000;
assign n_7010 = n_7001 ^ n_5660;
assign n_7011 = n_7004 ^ n_7005;
assign n_7012 = n_7005 ^ x402;
assign n_7013 = n_7006 ^ n_5058;
assign n_7014 = n_7007 ^ n_5780;
assign n_7015 = n_7010 ^ n_6557;
assign n_7016 = n_7011 ^ x402;
assign n_7017 = n_7011 & ~n_7012;
assign n_7018 = n_7013 ^ n_5078;
assign n_7019 = n_7014 ^ n_5078;
assign n_7020 = n_7013 ^ n_7014;
assign n_7021 = n_7015 ^ n_5694;
assign n_7022 = n_7015 & ~n_6574;
assign n_7023 = ~n_7002 & ~n_7016;
assign n_7024 = n_7016 ^ n_7002;
assign n_7025 = n_7017 ^ x402;
assign n_7026 = n_7018 ^ n_7014;
assign n_7027 = n_7019 & n_7020;
assign n_7028 = n_7021 & ~n_6573;
assign n_7029 = n_7021 ^ n_6557;
assign n_7030 = n_6896 ^ n_7021;
assign n_7031 = n_7022 ^ n_5694;
assign n_7032 = n_7025 ^ n_7026;
assign n_7033 = n_7026 ^ x401;
assign n_7034 = n_7027 ^ n_5078;
assign n_7035 = n_7028 ^ n_5819;
assign n_7036 = n_7031 ^ n_6615;
assign n_7037 = n_7031 ^ n_6599;
assign n_7038 = n_7032 ^ x401;
assign n_7039 = n_7032 & ~n_7033;
assign n_7040 = n_7034 ^ n_5101;
assign n_7041 = n_7035 ^ n_7034;
assign n_7042 = ~n_7036 & n_6616;
assign n_7043 = n_7036 ^ n_6599;
assign n_7044 = n_6933 ^ n_7036;
assign n_7045 = n_6615 & ~n_7037;
assign n_7046 = n_7023 & ~n_7038;
assign n_7047 = n_7038 ^ n_7023;
assign n_7048 = n_7039 ^ x401;
assign n_7049 = n_7035 ^ n_7040;
assign n_7050 = n_7040 & n_7041;
assign n_7051 = n_7042 ^ n_5861;
assign n_7052 = n_7045 ^ n_5768;
assign n_7053 = n_7048 ^ n_7049;
assign n_7054 = n_7049 ^ x400;
assign n_7055 = n_7050 ^ n_5101;
assign n_7056 = n_7051 ^ n_5129;
assign n_7057 = n_7052 ^ n_6642;
assign n_7058 = n_7053 ^ x400;
assign n_7059 = n_7053 & ~n_7054;
assign n_7060 = n_7055 ^ n_7051;
assign n_7061 = n_5822 ^ n_7057;
assign n_7062 = ~n_7057 & ~n_6658;
assign n_7063 = ~n_7046 & n_7058;
assign n_7064 = n_7058 ^ n_7046;
assign n_7065 = n_7059 ^ x400;
assign n_7066 = n_7060 ^ n_5129;
assign n_7067 = n_7060 & ~n_7056;
assign n_7068 = n_6629 & n_7061;
assign n_7069 = n_7061 ^ n_6642;
assign n_7070 = n_6961 ^ n_7061;
assign n_7071 = n_7062 ^ n_5822;
assign n_7072 = n_7065 ^ x415;
assign n_7073 = n_7065 ^ n_7066;
assign n_7074 = n_7067 ^ n_5129;
assign n_7075 = n_7068 ^ n_5903;
assign n_7076 = n_7071 ^ n_6683;
assign n_7077 = n_7073 ^ x415;
assign n_7078 = n_7073 & n_7072;
assign n_7079 = n_7074 ^ n_7075;
assign n_7080 = n_7075 ^ n_5164;
assign n_7081 = n_5864 ^ n_7076;
assign n_7082 = ~n_7076 & n_6700;
assign n_7083 = n_7063 & n_7077;
assign n_7084 = n_7077 ^ n_7063;
assign n_7085 = n_7078 ^ x415;
assign n_7086 = n_7079 ^ n_5164;
assign n_7087 = n_7079 & n_7080;
assign n_7088 = n_7081 & ~n_6699;
assign n_7089 = n_7081 ^ n_6683;
assign n_7090 = n_6983 ^ n_7081;
assign n_7091 = n_7082 ^ n_5864;
assign n_7092 = n_7085 ^ n_7086;
assign n_7093 = n_7086 ^ x414;
assign n_7094 = n_7087 ^ n_5164;
assign n_7095 = n_7088 ^ n_5943;
assign n_7096 = n_7091 ^ n_6725;
assign n_7097 = n_7092 ^ x414;
assign n_7098 = ~n_7092 & n_7093;
assign n_7099 = n_7094 ^ n_5200;
assign n_7100 = n_7095 ^ n_5200;
assign n_7101 = n_7094 ^ n_7095;
assign n_7102 = n_5906 ^ n_7096;
assign n_7103 = n_7096 & n_6742;
assign n_7104 = n_7083 ^ n_7097;
assign n_7105 = ~n_7097 & n_7083;
assign n_7106 = n_7098 ^ x414;
assign n_7107 = n_7099 ^ n_7095;
assign n_7108 = n_7100 & ~n_7101;
assign n_7109 = n_7102 & n_6741;
assign n_7110 = n_7102 ^ n_6725;
assign n_7111 = n_7003 ^ n_7102;
assign n_7112 = n_7103 ^ n_5906;
assign n_7113 = n_6127 & n_7104;
assign n_7114 = n_7104 ^ n_6127;
assign n_7115 = n_7106 ^ n_7107;
assign n_7116 = n_7107 ^ x413;
assign n_7117 = n_7108 ^ n_5200;
assign n_7118 = n_7109 ^ n_5985;
assign n_7119 = n_7112 ^ n_6767;
assign n_7120 = n_7113 ^ n_6172;
assign n_7121 = ~n_6111 & n_7114;
assign n_7122 = n_7115 ^ x413;
assign n_7123 = n_7115 & ~n_7116;
assign n_7124 = n_7117 ^ n_5238;
assign n_7125 = n_7118 ^ n_5238;
assign n_7126 = n_7117 ^ n_7118;
assign n_7127 = n_5946 ^ n_7119;
assign n_7128 = n_7119 & n_6784;
assign n_7129 = n_7121 ^ n_5625;
assign n_7130 = ~n_7105 & ~n_7122;
assign n_7131 = n_7122 ^ n_7105;
assign n_7132 = n_7123 ^ x413;
assign n_7133 = n_7124 ^ n_7118;
assign n_7134 = n_7125 & ~n_7126;
assign n_7135 = ~n_7127 & n_6783;
assign n_7136 = n_7127 ^ n_6767;
assign n_7137 = n_7024 ^ n_7127;
assign n_7138 = n_7128 ^ n_5946;
assign n_7139 = ~n_5098 & ~n_7129;
assign n_7140 = n_7129 ^ n_5098;
assign n_7141 = n_7131 ^ n_7113;
assign n_7142 = n_7131 ^ n_7120;
assign n_7143 = n_7132 ^ n_7133;
assign n_7144 = n_7133 ^ x412;
assign n_7145 = n_7134 ^ n_5238;
assign n_7146 = n_7135 ^ n_6026;
assign n_7147 = n_7138 ^ n_6810;
assign n_7148 = n_7139 ^ n_5125;
assign n_7149 = x423 & n_7140;
assign n_7150 = n_7140 ^ x423;
assign n_7151 = n_7120 & ~n_7141;
assign n_7152 = n_6173 & n_7142;
assign n_7153 = n_7143 ^ x412;
assign n_7154 = n_7143 & ~n_7144;
assign n_7155 = n_7145 ^ n_5277;
assign n_7156 = n_7146 ^ n_5277;
assign n_7157 = n_7145 ^ n_7146;
assign n_7158 = n_7147 ^ n_5988;
assign n_7159 = ~n_7147 & ~n_6827;
assign n_7160 = n_7149 ^ x422;
assign n_7161 = n_7151 ^ n_6172;
assign n_7162 = n_7152 ^ n_5652;
assign n_7163 = n_7153 & ~n_7130;
assign n_7164 = n_7130 ^ n_7153;
assign n_7165 = n_7154 ^ x412;
assign n_7166 = n_7155 ^ n_7146;
assign n_7167 = n_7156 & n_7157;
assign n_7168 = ~n_7158 & n_6826;
assign n_7169 = n_7158 ^ n_6810;
assign n_7170 = n_7047 ^ n_7158;
assign n_7171 = n_7159 ^ n_5988;
assign n_7172 = n_7161 ^ n_6230;
assign n_7173 = n_7162 ^ n_7139;
assign n_7174 = n_7162 ^ n_7148;
assign n_7175 = n_7164 ^ n_7161;
assign n_7176 = n_7164 ^ n_6230;
assign n_7177 = n_7165 ^ n_7166;
assign n_7178 = n_7166 ^ x411;
assign n_7179 = n_7167 ^ n_5277;
assign n_7180 = n_7168 ^ n_6068;
assign n_7181 = n_7171 ^ n_6852;
assign n_7182 = n_7172 ^ n_7164;
assign n_7183 = ~n_7148 & ~n_7173;
assign n_7184 = n_7174 ^ n_7149;
assign n_7185 = n_7174 ^ n_7160;
assign n_7186 = ~n_7175 & ~n_7176;
assign n_7187 = n_7177 ^ x411;
assign n_7188 = n_7177 & ~n_7178;
assign n_7189 = n_7179 ^ n_5319;
assign n_7190 = n_7180 ^ n_5319;
assign n_7191 = n_7179 ^ n_7180;
assign n_7192 = n_7181 ^ n_6029;
assign n_7193 = n_7181 & n_6869;
assign n_7194 = ~n_6218 & ~n_7182;
assign n_7195 = n_7183 ^ n_5125;
assign n_7196 = n_7160 & n_7184;
assign n_7197 = ~n_7150 & n_7185;
assign n_7198 = n_7185 ^ n_7150;
assign n_7199 = n_7186 ^ n_6230;
assign n_7200 = ~n_7187 & ~n_7163;
assign n_7201 = n_7163 ^ n_7187;
assign n_7202 = n_7188 ^ x411;
assign n_7203 = n_7189 ^ n_7180;
assign n_7204 = ~n_7190 & ~n_7191;
assign n_7205 = ~n_7192 & ~n_6868;
assign n_7206 = n_7192 ^ n_6852;
assign n_7207 = n_7064 ^ n_7192;
assign n_7208 = n_7193 ^ n_6029;
assign n_7209 = n_7194 ^ n_5696;
assign n_7210 = n_7195 ^ n_5169;
assign n_7211 = n_7196 ^ x422;
assign n_7212 = n_7199 ^ n_6267;
assign n_7213 = n_7201 ^ n_6267;
assign n_7214 = n_7199 ^ n_7201;
assign n_7215 = n_7202 ^ n_7203;
assign n_7216 = n_7203 ^ x410;
assign n_7217 = n_7204 ^ n_5319;
assign n_7218 = n_7205 ^ n_6109;
assign n_7219 = n_7208 ^ n_6909;
assign n_7220 = n_7209 ^ n_5169;
assign n_7221 = n_7195 ^ n_7209;
assign n_7222 = n_7210 ^ n_7209;
assign n_7223 = n_7212 ^ n_7201;
assign n_7224 = ~n_7213 & n_7214;
assign n_7225 = n_7215 ^ x410;
assign n_7226 = n_7215 & ~n_7216;
assign n_7227 = n_7217 ^ n_5361;
assign n_7228 = n_7218 ^ n_5361;
assign n_7229 = n_7218 ^ n_7217;
assign n_7230 = n_7219 & ~n_6910;
assign n_7231 = n_7084 ^ n_7219;
assign n_7232 = n_7219 ^ n_6894;
assign n_7233 = ~n_7220 & n_7221;
assign n_7234 = n_7211 ^ n_7222;
assign n_7235 = n_7222 ^ x421;
assign n_7236 = n_6257 & n_7223;
assign n_7237 = n_7224 ^ n_6267;
assign n_7238 = n_7225 & ~n_7200;
assign n_7239 = n_7200 ^ n_7225;
assign n_7240 = n_7226 ^ x410;
assign n_7241 = n_7218 ^ n_7227;
assign n_7242 = ~n_7228 & ~n_7229;
assign n_7243 = n_7230 ^ n_6140;
assign n_7244 = n_7233 ^ n_5169;
assign n_7245 = n_7234 ^ x421;
assign n_7246 = ~n_7234 & n_7235;
assign n_7247 = n_7236 ^ n_5732;
assign n_7248 = n_7237 ^ n_6307;
assign n_7249 = n_7239 ^ n_6307;
assign n_7250 = n_7237 ^ n_7239;
assign n_7251 = n_7240 ^ n_7241;
assign n_7252 = n_7241 ^ x409;
assign n_7253 = n_7242 ^ n_5361;
assign n_7254 = n_7243 ^ n_5391;
assign n_7255 = n_7244 ^ n_5208;
assign n_7256 = n_7245 & ~n_7197;
assign n_7257 = n_7197 ^ n_7245;
assign n_7258 = n_7246 ^ x421;
assign n_7259 = n_7247 ^ n_5208;
assign n_7260 = n_7244 ^ n_7247;
assign n_7261 = n_7248 ^ n_7239;
assign n_7262 = n_7249 & n_7250;
assign n_7263 = n_7251 ^ x409;
assign n_7264 = ~n_7251 & n_7252;
assign n_7265 = n_7253 ^ x408;
assign n_7266 = n_7255 ^ n_7247;
assign n_7267 = ~n_7259 & ~n_7260;
assign n_7268 = n_6294 & ~n_7261;
assign n_7269 = n_7262 ^ n_6307;
assign n_7270 = n_7238 & ~n_7263;
assign n_7271 = n_7263 ^ n_7238;
assign n_7272 = n_7264 ^ x409;
assign n_7273 = n_7265 ^ n_7254;
assign n_7274 = n_7258 ^ n_7266;
assign n_7275 = n_7266 ^ x420;
assign n_7276 = n_7267 ^ n_5208;
assign n_7277 = n_7268 ^ n_5773;
assign n_7278 = n_7269 ^ n_6344;
assign n_7279 = n_7271 ^ n_7269;
assign n_7280 = n_7271 ^ n_6344;
assign n_7281 = n_7272 ^ n_7273;
assign n_7282 = n_7274 ^ x420;
assign n_7283 = ~n_7274 & n_7275;
assign n_7284 = n_7276 ^ n_5248;
assign n_7285 = n_7277 ^ n_5248;
assign n_7286 = n_7276 ^ n_7277;
assign n_7287 = n_7278 ^ n_7271;
assign n_7288 = ~n_7279 & n_7280;
assign n_7289 = n_7281 ^ n_7270;
assign n_7290 = n_7256 & n_7282;
assign n_7291 = n_7282 ^ n_7256;
assign n_7292 = n_7283 ^ x420;
assign n_7293 = n_7284 ^ n_7277;
assign n_7294 = n_7285 & ~n_7286;
assign n_7295 = n_6332 & n_7287;
assign n_7296 = n_7288 ^ n_6344;
assign n_7297 = n_7289 ^ n_6383;
assign n_7298 = n_7292 ^ n_7293;
assign n_7299 = n_7293 ^ x419;
assign n_7300 = n_7294 ^ n_5248;
assign n_7301 = n_7295 ^ n_5812;
assign n_7302 = n_7296 ^ n_7289;
assign n_7303 = n_7296 ^ n_7297;
assign n_7304 = n_7298 ^ x419;
assign n_7305 = ~n_7298 & n_7299;
assign n_7306 = n_7300 ^ n_5286;
assign n_7307 = n_7301 ^ n_5286;
assign n_7308 = n_7300 ^ n_7301;
assign n_7309 = n_7297 & n_7302;
assign n_7310 = n_6371 & n_7303;
assign n_7311 = ~n_7290 & ~n_7304;
assign n_7312 = n_7304 ^ n_7290;
assign n_7313 = n_7305 ^ x419;
assign n_7314 = n_7306 ^ n_7301;
assign n_7315 = ~n_7307 & ~n_7308;
assign n_7316 = n_7309 ^ n_6383;
assign n_7317 = n_7310 ^ n_5854;
assign n_7318 = n_7313 ^ n_7314;
assign n_7319 = n_7314 ^ x418;
assign n_7320 = n_7315 ^ n_5286;
assign n_7321 = n_7316 ^ n_6425;
assign n_7322 = n_7317 ^ n_5328;
assign n_7323 = n_7318 ^ x418;
assign n_7324 = n_7318 & ~n_7319;
assign n_7325 = n_7320 ^ n_7317;
assign n_7326 = n_7320 ^ n_5328;
assign n_7327 = n_7321 & ~n_6440;
assign n_7328 = n_6186 ^ n_7321;
assign n_7329 = ~n_7311 & ~n_7323;
assign n_7330 = n_7323 ^ n_7311;
assign n_7331 = n_7324 ^ x418;
assign n_7332 = n_7322 & ~n_7325;
assign n_7333 = n_7326 ^ n_7317;
assign n_7334 = n_7327 ^ n_6186;
assign n_7335 = n_6413 & n_7328;
assign n_7336 = n_7328 ^ n_6425;
assign n_7337 = n_7332 ^ n_5328;
assign n_7338 = n_7331 ^ n_7333;
assign n_7339 = n_7333 ^ x417;
assign n_7340 = n_7334 ^ n_6466;
assign n_7341 = n_7334 ^ n_6228;
assign n_7342 = n_7335 ^ n_5897;
assign n_7343 = n_7337 ^ n_5370;
assign n_7344 = n_7338 ^ x417;
assign n_7345 = n_7338 & ~n_7339;
assign n_7346 = n_7340 ^ n_6228;
assign n_7347 = n_7341 & n_6481;
assign n_7348 = n_7342 ^ n_5370;
assign n_7349 = n_7337 ^ n_7342;
assign n_7350 = n_7343 ^ n_7342;
assign n_7351 = n_7329 & ~n_7344;
assign n_7352 = n_7344 ^ n_7329;
assign n_7353 = n_7345 ^ x417;
assign n_7354 = n_6454 & ~n_7346;
assign n_7355 = n_7347 ^ n_6466;
assign n_7356 = ~n_7348 & n_7349;
assign n_7357 = n_7350 ^ x416;
assign n_7358 = n_7353 ^ n_7350;
assign n_7359 = n_7354 ^ n_5937;
assign n_7360 = n_7355 ^ n_6508;
assign n_7361 = n_7356 ^ n_5370;
assign n_7362 = ~n_7358 & n_7357;
assign n_7363 = n_7358 ^ x416;
assign n_7364 = n_6302 ^ n_7360;
assign n_7365 = n_7360 & ~n_6522;
assign n_7366 = n_7361 ^ n_5413;
assign n_7367 = n_7359 ^ n_7361;
assign n_7368 = n_7362 ^ x416;
assign n_7369 = ~n_7351 & ~n_7363;
assign n_7370 = n_7363 ^ n_7351;
assign n_7371 = ~n_6497 & ~n_7364;
assign n_7372 = n_7364 ^ n_6508;
assign n_7373 = n_7365 ^ n_6302;
assign n_7374 = n_7359 ^ n_7366;
assign n_7375 = n_7366 & n_7367;
assign n_7376 = n_7371 ^ n_5979;
assign n_7377 = n_7373 ^ n_6550;
assign n_7378 = n_7374 ^ x431;
assign n_7379 = n_7368 ^ n_7374;
assign n_7380 = n_7375 ^ n_5413;
assign n_7381 = n_7376 ^ n_5448;
assign n_7382 = n_6353 ^ n_7377;
assign n_7383 = n_7377 & n_6565;
assign n_7384 = n_7368 ^ n_7378;
assign n_7385 = n_7378 & ~n_7379;
assign n_7386 = n_7380 ^ n_5448;
assign n_7387 = n_7380 ^ n_7376;
assign n_7388 = ~n_6539 & n_7382;
assign n_7389 = n_7382 ^ n_6550;
assign n_7390 = n_7383 ^ n_6353;
assign n_7391 = ~n_7384 & n_7369;
assign n_7392 = n_7369 ^ n_7384;
assign n_7393 = n_7385 ^ x431;
assign n_7394 = n_7386 ^ n_7376;
assign n_7395 = ~n_7381 & n_7387;
assign n_7396 = n_7388 ^ n_6019;
assign n_7397 = n_7390 ^ n_6393;
assign n_7398 = n_7390 ^ n_6593;
assign n_7399 = n_7393 ^ n_7394;
assign n_7400 = n_7394 ^ x430;
assign n_7401 = n_7395 ^ n_5448;
assign n_7402 = n_7396 ^ n_5476;
assign n_7403 = n_7397 ^ n_6593;
assign n_7404 = ~n_6607 & n_7398;
assign n_7405 = n_7399 ^ x430;
assign n_7406 = ~n_7399 & n_7400;
assign n_7407 = n_7401 ^ n_5476;
assign n_7408 = n_7401 ^ n_7396;
assign n_7409 = n_6582 & n_7403;
assign n_7410 = n_7404 ^ n_6393;
assign n_7411 = ~n_7391 & n_7405;
assign n_7412 = n_7405 ^ n_7391;
assign n_7413 = n_7406 ^ x430;
assign n_7414 = n_7407 ^ n_7396;
assign n_7415 = n_7402 & n_7408;
assign n_7416 = n_7409 ^ n_6061;
assign n_7417 = n_7410 ^ n_6636;
assign n_7418 = n_7413 ^ n_7414;
assign n_7419 = n_7414 ^ x429;
assign n_7420 = n_7415 ^ n_5476;
assign n_7421 = n_7416 ^ n_5498;
assign n_7422 = n_6435 ^ n_7417;
assign n_7423 = ~n_7417 & ~n_6650;
assign n_7424 = n_7418 ^ x429;
assign n_7425 = n_7418 & ~n_7419;
assign n_7426 = n_7420 ^ n_7416;
assign n_7427 = ~n_6624 & n_7422;
assign n_7428 = n_7150 ^ n_7422;
assign n_7429 = n_7422 ^ n_6636;
assign n_7430 = n_7423 ^ n_6435;
assign n_7431 = n_7411 & ~n_7424;
assign n_7432 = n_7424 ^ n_7411;
assign n_7433 = n_7425 ^ x429;
assign n_7434 = n_7426 ^ n_5498;
assign n_7435 = ~n_7426 & ~n_7421;
assign n_7436 = n_7427 ^ n_6102;
assign n_7437 = n_7430 ^ n_6677;
assign n_7438 = n_7433 ^ n_7434;
assign n_7439 = n_7434 ^ x428;
assign n_7440 = n_7435 ^ n_5498;
assign n_7441 = n_7436 ^ n_5511;
assign n_7442 = n_6476 ^ n_7437;
assign n_7443 = ~n_7437 & n_6691;
assign n_7444 = n_7438 ^ x428;
assign n_7445 = n_7438 & ~n_7439;
assign n_7446 = n_7440 ^ n_5511;
assign n_7447 = n_7440 ^ n_7436;
assign n_7448 = ~n_6666 & n_7442;
assign n_7449 = n_7442 ^ n_6677;
assign n_7450 = n_7198 ^ n_7442;
assign n_7451 = n_7443 ^ n_6476;
assign n_7452 = n_7431 & ~n_7444;
assign n_7453 = n_7444 ^ n_7431;
assign n_7454 = n_7445 ^ x428;
assign n_7455 = n_7446 ^ n_7436;
assign n_7456 = n_7441 & n_7447;
assign n_7457 = n_7448 ^ n_6147;
assign n_7458 = n_7451 ^ n_6719;
assign n_7459 = n_7454 ^ n_7455;
assign n_7460 = n_7455 ^ x427;
assign n_7461 = n_7456 ^ n_5511;
assign n_7462 = n_7457 ^ n_5536;
assign n_7463 = n_6517 ^ n_7458;
assign n_7464 = n_7458 & ~n_6733;
assign n_7465 = n_7459 ^ x427;
assign n_7466 = n_7459 & ~n_7460;
assign n_7467 = n_7461 ^ n_5536;
assign n_7468 = n_7461 ^ n_7457;
assign n_7469 = n_6708 & ~n_7463;
assign n_7470 = n_7463 ^ n_6719;
assign n_7471 = n_7257 ^ n_7463;
assign n_7472 = n_7464 ^ n_6517;
assign n_7473 = ~n_7452 & n_7465;
assign n_7474 = n_7465 ^ n_7452;
assign n_7475 = n_7466 ^ x427;
assign n_7476 = n_7467 ^ n_7457;
assign n_7477 = ~n_7462 & n_7468;
assign n_7478 = n_7469 ^ n_6195;
assign n_7479 = n_7472 ^ n_6761;
assign n_7480 = n_7475 ^ n_7476;
assign n_7481 = n_7476 ^ x426;
assign n_7482 = n_7477 ^ n_5536;
assign n_7483 = n_7478 ^ n_5555;
assign n_7484 = n_6560 ^ n_7479;
assign n_7485 = ~n_7479 & n_6775;
assign n_7486 = n_7480 ^ x426;
assign n_7487 = n_7480 & ~n_7481;
assign n_7488 = n_7482 ^ n_7478;
assign n_7489 = n_6749 & n_7484;
assign n_7490 = n_7484 ^ n_6761;
assign n_7491 = n_7291 ^ n_7484;
assign n_7492 = n_7485 ^ n_6560;
assign n_7493 = n_7473 & n_7486;
assign n_7494 = n_7486 ^ n_7473;
assign n_7495 = n_7487 ^ x426;
assign n_7496 = n_7488 ^ n_5555;
assign n_7497 = n_7488 & n_7483;
assign n_7498 = n_7489 ^ n_6237;
assign n_7499 = n_7492 ^ n_6803;
assign n_7500 = n_7495 ^ n_7496;
assign n_7501 = n_7496 ^ x425;
assign n_7502 = n_7497 ^ n_5555;
assign n_7503 = n_7498 ^ n_5575;
assign n_7504 = n_6602 ^ n_7499;
assign n_7505 = ~n_7499 & ~n_6818;
assign n_7506 = n_7500 ^ x425;
assign n_7507 = ~n_7500 & n_7501;
assign n_7508 = n_7502 ^ n_5575;
assign n_7509 = n_7502 ^ n_7498;
assign n_7510 = n_6792 & ~n_7504;
assign n_7511 = n_7504 ^ n_6803;
assign n_7512 = n_7312 ^ n_7504;
assign n_7513 = n_7505 ^ n_6602;
assign n_7514 = n_7493 & ~n_7506;
assign n_7515 = n_7506 ^ n_7493;
assign n_7516 = n_7507 ^ x425;
assign n_7517 = n_7508 ^ n_7498;
assign n_7518 = ~n_7503 & n_7509;
assign n_7519 = n_7510 ^ n_6274;
assign n_7520 = n_7513 ^ n_6645;
assign n_7521 = n_7513 ^ n_6845;
assign n_7522 = n_7516 ^ n_7517;
assign n_7523 = n_7517 ^ x424;
assign n_7524 = n_7518 ^ n_5575;
assign n_7525 = n_7519 ^ n_5595;
assign n_7526 = n_7520 ^ n_6845;
assign n_7527 = n_6860 & ~n_7521;
assign n_7528 = n_7522 ^ x424;
assign n_7529 = ~n_7522 & n_7523;
assign n_7530 = n_7524 ^ n_7519;
assign n_7531 = n_6835 & ~n_7526;
assign n_7532 = n_7330 ^ n_7526;
assign n_7533 = n_7527 ^ n_6645;
assign n_7534 = n_7528 & ~n_7514;
assign n_7535 = n_7514 ^ n_7528;
assign n_7536 = n_7529 ^ x424;
assign n_7537 = n_7530 ^ n_5595;
assign n_7538 = n_7530 & n_7525;
assign n_7539 = n_7531 ^ n_6313;
assign n_7540 = n_7533 ^ n_6887;
assign n_7541 = n_7536 ^ n_7537;
assign n_7542 = n_7537 ^ x439;
assign n_7543 = n_7538 ^ n_5595;
assign n_7544 = n_7539 ^ n_5615;
assign n_7545 = n_6686 ^ n_7540;
assign n_7546 = ~n_7540 & n_6901;
assign n_7547 = n_7541 ^ x439;
assign n_7548 = n_7541 & ~n_7542;
assign n_7549 = n_7543 ^ n_5615;
assign n_7550 = n_7543 ^ n_7539;
assign n_7551 = ~n_6877 & ~n_7545;
assign n_7552 = n_7545 ^ n_6887;
assign n_7553 = n_7352 ^ n_7545;
assign n_7554 = n_7546 ^ n_6686;
assign n_7555 = n_7534 & ~n_7547;
assign n_7556 = n_7547 ^ n_7534;
assign n_7557 = n_7548 ^ x439;
assign n_7558 = n_7549 ^ n_7539;
assign n_7559 = ~n_7544 & n_7550;
assign n_7560 = n_7551 ^ n_6350;
assign n_7561 = n_7554 ^ n_6926;
assign n_7562 = n_7557 ^ n_7558;
assign n_7563 = n_7558 ^ x438;
assign n_7564 = n_7559 ^ n_5615;
assign n_7565 = n_7560 ^ n_5638;
assign n_7566 = n_6728 ^ n_7561;
assign n_7567 = n_7561 & ~n_6938;
assign n_7568 = n_7562 ^ x438;
assign n_7569 = n_7562 & ~n_7563;
assign n_7570 = n_7564 ^ n_7560;
assign n_7571 = n_6917 & n_7566;
assign n_7572 = n_7566 ^ n_6926;
assign n_7573 = n_7370 ^ n_7566;
assign n_7574 = n_7567 ^ n_6728;
assign n_7575 = n_7555 & ~n_7568;
assign n_7576 = n_7568 ^ n_7555;
assign n_7577 = n_7569 ^ x438;
assign n_7578 = n_7570 ^ n_5638;
assign n_7579 = ~n_7570 & n_7565;
assign n_7580 = n_7571 ^ n_6390;
assign n_7581 = n_7574 ^ n_6957;
assign n_7582 = n_7577 ^ n_7578;
assign n_7583 = n_7578 ^ x437;
assign n_7584 = n_7579 ^ n_5638;
assign n_7585 = n_7580 ^ n_5669;
assign n_7586 = n_6770 ^ n_7581;
assign n_7587 = n_7581 & n_6966;
assign n_7588 = n_7582 ^ x437;
assign n_7589 = ~n_7582 & n_7583;
assign n_7590 = n_7584 ^ n_5669;
assign n_7591 = n_7584 ^ n_7580;
assign n_7592 = ~n_6950 & ~n_7586;
assign n_7593 = n_7586 ^ n_6957;
assign n_7594 = n_7392 ^ n_7586;
assign n_7595 = n_7587 ^ n_6770;
assign n_7596 = n_7575 & n_7588;
assign n_7597 = n_7588 ^ n_7575;
assign n_7598 = n_7589 ^ x437;
assign n_7599 = n_7590 ^ n_7580;
assign n_7600 = ~n_7585 & ~n_7591;
assign n_7601 = n_7592 ^ n_6432;
assign n_7602 = n_7595 ^ n_6980;
assign n_7603 = n_7598 ^ n_7599;
assign n_7604 = n_7599 ^ x436;
assign n_7605 = n_7600 ^ n_5669;
assign n_7606 = n_7601 ^ n_5703;
assign n_7607 = n_6813 ^ n_7602;
assign n_7608 = ~n_7602 & n_6988;
assign n_7609 = n_7603 ^ x436;
assign n_7610 = n_7603 & ~n_7604;
assign n_7611 = n_7605 ^ n_5703;
assign n_7612 = n_7605 ^ n_7601;
assign n_7613 = ~n_6974 & n_7607;
assign n_7614 = n_7607 ^ n_6980;
assign n_7615 = n_7412 ^ n_7607;
assign n_7616 = n_7608 ^ n_6813;
assign n_7617 = ~n_7596 & n_7609;
assign n_7618 = n_7609 ^ n_7596;
assign n_7619 = n_7610 ^ x436;
assign n_7620 = n_7611 ^ n_7601;
assign n_7621 = ~n_7606 & ~n_7612;
assign n_7622 = n_7613 ^ n_6473;
assign n_7623 = n_7616 ^ n_7000;
assign n_7624 = n_7619 ^ n_7620;
assign n_7625 = n_7620 ^ x435;
assign n_7626 = n_7621 ^ n_5703;
assign n_7627 = n_7622 ^ n_5739;
assign n_7628 = n_6855 ^ n_7623;
assign n_7629 = n_7623 & n_7009;
assign n_7630 = n_7624 ^ x435;
assign n_7631 = ~n_7624 & n_7625;
assign n_7632 = n_7626 ^ n_5739;
assign n_7633 = n_7626 ^ n_7622;
assign n_7634 = n_7628 & n_7008;
assign n_7635 = n_7628 ^ n_7000;
assign n_7636 = n_7432 ^ n_7628;
assign n_7637 = n_7629 ^ n_6855;
assign n_7638 = n_7617 ^ n_7630;
assign n_7639 = ~n_7630 & n_7617;
assign n_7640 = n_7631 ^ x435;
assign n_7641 = n_7632 ^ n_7622;
assign n_7642 = ~n_7627 & n_7633;
assign n_7643 = n_7634 ^ n_6514;
assign n_7644 = n_7637 ^ n_7021;
assign n_7645 = n_7638 ^ n_7114;
assign n_7646 = n_7114 & n_7638;
assign n_7647 = n_7640 ^ n_7641;
assign n_7648 = n_7641 ^ x434;
assign n_7649 = n_7642 ^ n_5739;
assign n_7650 = n_7643 ^ n_5780;
assign n_7651 = n_6896 ^ n_7644;
assign n_7652 = n_7644 & ~n_7030;
assign n_7653 = n_7104 & n_7645;
assign n_7654 = n_7646 ^ n_7142;
assign n_7655 = n_7647 ^ x434;
assign n_7656 = n_7647 & ~n_7648;
assign n_7657 = n_7649 ^ n_5780;
assign n_7658 = n_7649 ^ n_7643;
assign n_7659 = n_7651 & n_7029;
assign n_7660 = n_7651 ^ n_7021;
assign n_7661 = n_7453 ^ n_7651;
assign n_7662 = n_7652 ^ n_6896;
assign n_7663 = n_7653 ^ n_6127;
assign n_7664 = n_7639 ^ n_7655;
assign n_7665 = ~n_7655 & ~n_7639;
assign n_7666 = n_7656 ^ x434;
assign n_7667 = n_7657 ^ n_7643;
assign n_7668 = ~n_7650 & n_7658;
assign n_7669 = n_7659 ^ n_6557;
assign n_7670 = n_7662 ^ n_7036;
assign n_7671 = n_7663 ^ n_5625;
assign n_7672 = ~n_5625 & n_7663;
assign n_7673 = n_7664 ^ n_7654;
assign n_7674 = n_7664 ^ n_7646;
assign n_7675 = n_7666 ^ n_7667;
assign n_7676 = n_7667 ^ x433;
assign n_7677 = n_7668 ^ n_5780;
assign n_7678 = n_7669 ^ n_5819;
assign n_7679 = n_6933 ^ n_7670;
assign n_7680 = ~n_7670 & n_7044;
assign n_7681 = x455 & ~n_7671;
assign n_7682 = n_7671 ^ x455;
assign n_7683 = n_7672 ^ n_5652;
assign n_7684 = n_7141 & n_7673;
assign n_7685 = n_7654 & ~n_7674;
assign n_7686 = n_7675 ^ x433;
assign n_7687 = n_7675 & ~n_7676;
assign n_7688 = n_7677 ^ n_5819;
assign n_7689 = n_7677 ^ n_7669;
assign n_7690 = ~n_7679 & n_7043;
assign n_7691 = n_7679 ^ n_7036;
assign n_7692 = n_7474 ^ n_7679;
assign n_7693 = n_7680 ^ n_6933;
assign n_7694 = n_7681 ^ x454;
assign n_7695 = n_7684 ^ n_6172;
assign n_7696 = n_7685 ^ n_7142;
assign n_7697 = n_7686 ^ n_7665;
assign n_7698 = n_7665 & ~n_7686;
assign n_7699 = n_7687 ^ x433;
assign n_7700 = n_7688 ^ n_7669;
assign n_7701 = ~n_7678 & ~n_7689;
assign n_7702 = n_7690 ^ n_6599;
assign n_7703 = n_7693 ^ n_6961;
assign n_7704 = n_7693 ^ n_7061;
assign n_7705 = n_7695 ^ n_7683;
assign n_7706 = n_7695 ^ n_7672;
assign n_7707 = n_7696 ^ n_7182;
assign n_7708 = n_7697 ^ n_7182;
assign n_7709 = n_7696 ^ n_7697;
assign n_7710 = n_7699 ^ n_7700;
assign n_7711 = n_7700 ^ x432;
assign n_7712 = n_7701 ^ n_5819;
assign n_7713 = n_7702 ^ n_5861;
assign n_7714 = n_7703 ^ n_7061;
assign n_7715 = ~n_7070 & n_7704;
assign n_7716 = n_7705 ^ n_7681;
assign n_7717 = n_7705 ^ n_7694;
assign n_7718 = n_7683 & ~n_7706;
assign n_7719 = n_7707 ^ n_7697;
assign n_7720 = n_7708 & n_7709;
assign n_7721 = n_7710 ^ x432;
assign n_7722 = n_7710 & ~n_7711;
assign n_7723 = n_7712 ^ n_7702;
assign n_7724 = n_7714 & ~n_7069;
assign n_7725 = n_7494 ^ n_7714;
assign n_7726 = n_7715 ^ n_6961;
assign n_7727 = n_7694 & ~n_7716;
assign n_7728 = n_7718 ^ n_5652;
assign n_7729 = n_7175 & n_7719;
assign n_7730 = n_7720 ^ n_7182;
assign n_7731 = n_7721 ^ n_7698;
assign n_7732 = ~n_7698 & n_7721;
assign n_7733 = n_7722 ^ x432;
assign n_7734 = n_7723 ^ n_5861;
assign n_7735 = ~n_7723 & n_7713;
assign n_7736 = n_7724 ^ n_6642;
assign n_7737 = n_7726 ^ n_7081;
assign n_7738 = n_7727 ^ x454;
assign n_7739 = n_7728 ^ n_5696;
assign n_7740 = n_7729 ^ n_6230;
assign n_7741 = n_7730 ^ n_7223;
assign n_7742 = n_7731 ^ n_7223;
assign n_7743 = n_7730 ^ n_7731;
assign n_7744 = n_7733 ^ n_7734;
assign n_7745 = n_7734 ^ x447;
assign n_7746 = n_7735 ^ n_5861;
assign n_7747 = n_7736 ^ n_5903;
assign n_7748 = n_6983 ^ n_7737;
assign n_7749 = n_7737 & n_7090;
assign n_7750 = n_7739 ^ n_7740;
assign n_7751 = n_7740 ^ n_5696;
assign n_7752 = n_7728 ^ n_7740;
assign n_7753 = n_7741 ^ n_7731;
assign n_7754 = n_7742 & n_7743;
assign n_7755 = n_7744 ^ x447;
assign n_7756 = n_7744 & ~n_7745;
assign n_7757 = n_7746 ^ n_5903;
assign n_7758 = n_7746 ^ n_7736;
assign n_7759 = ~n_7748 & n_7089;
assign n_7760 = n_7748 ^ n_7081;
assign n_7761 = n_7515 ^ n_7748;
assign n_7762 = n_7749 ^ n_6983;
assign n_7763 = n_7738 ^ n_7750;
assign n_7764 = n_7750 ^ x453;
assign n_7765 = ~n_7751 & n_7752;
assign n_7766 = ~n_7214 & ~n_7753;
assign n_7767 = n_7754 ^ n_7223;
assign n_7768 = n_7755 ^ n_7732;
assign n_7769 = n_7732 & n_7755;
assign n_7770 = n_7756 ^ x447;
assign n_7771 = n_7757 ^ n_7736;
assign n_7772 = n_7747 & ~n_7758;
assign n_7773 = n_7759 ^ n_6683;
assign n_7774 = n_7762 ^ n_7102;
assign n_7775 = n_7763 ^ x453;
assign n_7776 = n_7763 & ~n_7764;
assign n_7777 = n_7765 ^ n_5696;
assign n_7778 = n_7766 ^ n_6267;
assign n_7779 = n_7767 ^ n_7261;
assign n_7780 = n_7768 ^ n_7261;
assign n_7781 = n_7767 ^ n_7768;
assign n_7782 = n_7770 ^ n_7771;
assign n_7783 = n_7771 ^ x446;
assign n_7784 = n_7772 ^ n_5903;
assign n_7785 = n_7773 ^ n_5943;
assign n_7786 = n_7003 ^ n_7774;
assign n_7787 = ~n_7774 & n_7111;
assign n_7788 = n_7775 & ~n_7717;
assign n_7789 = n_7717 ^ n_7775;
assign n_7790 = n_7776 ^ x453;
assign n_7791 = n_7777 ^ n_5732;
assign n_7792 = n_7778 ^ n_5732;
assign n_7793 = n_7777 ^ n_7778;
assign n_7794 = n_7779 ^ n_7768;
assign n_7795 = n_7780 & n_7781;
assign n_7796 = n_7782 ^ x446;
assign n_7797 = n_7782 & ~n_7783;
assign n_7798 = n_7784 ^ n_5943;
assign n_7799 = n_7784 ^ n_7773;
assign n_7800 = n_7786 & ~n_7110;
assign n_7801 = n_7786 ^ n_7102;
assign n_7802 = n_7535 ^ n_7786;
assign n_7803 = n_7787 ^ n_7003;
assign n_7804 = n_7791 ^ n_7778;
assign n_7805 = n_7792 & n_7793;
assign n_7806 = ~n_7250 & n_7794;
assign n_7807 = n_7795 ^ n_7261;
assign n_7808 = n_7796 ^ n_7769;
assign n_7809 = ~n_7769 & ~n_7796;
assign n_7810 = n_7797 ^ x446;
assign n_7811 = n_7798 ^ n_7773;
assign n_7812 = ~n_7785 & n_7799;
assign n_7813 = n_7800 ^ n_6725;
assign n_7814 = n_7803 ^ n_7127;
assign n_7815 = n_7790 ^ n_7804;
assign n_7816 = n_7804 ^ x452;
assign n_7817 = n_7805 ^ n_5732;
assign n_7818 = n_7806 ^ n_6307;
assign n_7819 = n_7807 ^ n_7287;
assign n_7820 = n_7808 ^ n_7287;
assign n_7821 = n_7807 ^ n_7808;
assign n_7822 = n_7810 ^ n_7811;
assign n_7823 = n_7811 ^ x445;
assign n_7824 = n_7812 ^ n_5943;
assign n_7825 = n_7813 ^ n_5985;
assign n_7826 = n_7024 ^ n_7814;
assign n_7827 = n_7814 & ~n_7137;
assign n_7828 = n_7815 ^ x452;
assign n_7829 = ~n_7815 & n_7816;
assign n_7830 = n_7817 ^ n_5773;
assign n_7831 = n_7818 ^ n_5773;
assign n_7832 = n_7817 ^ n_7818;
assign n_7833 = n_7819 ^ n_7808;
assign n_7834 = n_7820 & n_7821;
assign n_7835 = n_7822 ^ x445;
assign n_7836 = ~n_7822 & n_7823;
assign n_7837 = n_7824 ^ n_5985;
assign n_7838 = n_7824 ^ n_7813;
assign n_7839 = ~n_7826 & ~n_7136;
assign n_7840 = n_7826 ^ n_7127;
assign n_7841 = n_7556 ^ n_7826;
assign n_7842 = n_7827 ^ n_7024;
assign n_7843 = n_7788 & ~n_7828;
assign n_7844 = n_7828 ^ n_7788;
assign n_7845 = n_7829 ^ x452;
assign n_7846 = n_7830 ^ n_7818;
assign n_7847 = n_7831 & n_7832;
assign n_7848 = n_7279 & ~n_7833;
assign n_7849 = n_7834 ^ n_7287;
assign n_7850 = n_7809 ^ n_7835;
assign n_7851 = ~n_7835 & ~n_7809;
assign n_7852 = n_7836 ^ x445;
assign n_7853 = n_7837 ^ n_7813;
assign n_7854 = n_7825 & ~n_7838;
assign n_7855 = n_7839 ^ n_6767;
assign n_7856 = n_7842 ^ n_7158;
assign n_7857 = n_7845 ^ n_7846;
assign n_7858 = n_7846 ^ x451;
assign n_7859 = n_7847 ^ n_5773;
assign n_7860 = n_7848 ^ n_6344;
assign n_7861 = n_7850 ^ n_7303;
assign n_7862 = n_7849 ^ n_7850;
assign n_7863 = n_7852 ^ n_7853;
assign n_7864 = n_7853 ^ x444;
assign n_7865 = n_7854 ^ n_5985;
assign n_7866 = n_7855 ^ n_6026;
assign n_7867 = n_7856 ^ n_7047;
assign n_7868 = n_7856 & n_7170;
assign n_7869 = n_7857 ^ x451;
assign n_7870 = n_7857 & ~n_7858;
assign n_7871 = n_7859 ^ n_5812;
assign n_7872 = n_7860 ^ n_5812;
assign n_7873 = n_7859 ^ n_7860;
assign n_7874 = n_7849 ^ n_7861;
assign n_7875 = ~n_7861 & n_7862;
assign n_7876 = n_7863 ^ x444;
assign n_7877 = n_7863 & ~n_7864;
assign n_7878 = n_7865 ^ n_6026;
assign n_7879 = n_7865 ^ n_7855;
assign n_7880 = n_7867 & ~n_7169;
assign n_7881 = n_7867 ^ n_7158;
assign n_7882 = n_7576 ^ n_7867;
assign n_7883 = n_7868 ^ n_7047;
assign n_7884 = ~n_7843 & ~n_7869;
assign n_7885 = n_7869 ^ n_7843;
assign n_7886 = n_7870 ^ x451;
assign n_7887 = n_7871 ^ n_7860;
assign n_7888 = n_7872 & ~n_7873;
assign n_7889 = ~n_7302 & ~n_7874;
assign n_7890 = n_7875 ^ n_7303;
assign n_7891 = n_7851 ^ n_7876;
assign n_7892 = n_7876 & n_7851;
assign n_7893 = n_7877 ^ x444;
assign n_7894 = n_7878 ^ n_7855;
assign n_7895 = n_7866 & n_7879;
assign n_7896 = n_7880 ^ n_6810;
assign n_7897 = n_7883 ^ n_7192;
assign n_7898 = n_7886 ^ n_7887;
assign n_7899 = n_7887 ^ x450;
assign n_7900 = n_7888 ^ n_5812;
assign n_7901 = n_7889 ^ n_6383;
assign n_7902 = n_7890 ^ n_7328;
assign n_7903 = n_7891 ^ n_7328;
assign n_7904 = n_7890 ^ n_7891;
assign n_7905 = n_7893 ^ n_7894;
assign n_7906 = n_7894 ^ x443;
assign n_7907 = n_7895 ^ n_6026;
assign n_7908 = n_7896 ^ n_6068;
assign n_7909 = n_7897 ^ n_7064;
assign n_7910 = ~n_7897 & ~n_7207;
assign n_7911 = n_7898 ^ x450;
assign n_7912 = ~n_7898 & n_7899;
assign n_7913 = n_7900 ^ n_5854;
assign n_7914 = n_7901 ^ n_7900;
assign n_7915 = n_7902 ^ n_7891;
assign n_7916 = ~n_7903 & n_7904;
assign n_7917 = n_7905 ^ x443;
assign n_7918 = n_7905 & ~n_7906;
assign n_7919 = n_7907 ^ n_6068;
assign n_7920 = n_7907 ^ n_7896;
assign n_7921 = n_7909 & ~n_7206;
assign n_7922 = n_7909 ^ n_7192;
assign n_7923 = n_7597 ^ n_7909;
assign n_7924 = n_7910 ^ n_7064;
assign n_7925 = n_7911 & n_7884;
assign n_7926 = n_7884 ^ n_7911;
assign n_7927 = n_7912 ^ x450;
assign n_7928 = n_7901 ^ n_7913;
assign n_7929 = ~n_7913 & n_7914;
assign n_7930 = ~n_7915 & n_7336;
assign n_7931 = n_7916 ^ n_7328;
assign n_7932 = n_7892 ^ n_7917;
assign n_7933 = n_7917 & n_7892;
assign n_7934 = n_7918 ^ x443;
assign n_7935 = n_7919 ^ n_7896;
assign n_7936 = n_7908 & ~n_7920;
assign n_7937 = n_7921 ^ n_6852;
assign n_7938 = n_7924 ^ n_7231;
assign n_7939 = n_7927 ^ n_7928;
assign n_7940 = n_7928 ^ x449;
assign n_7941 = n_7929 ^ n_5854;
assign n_7942 = n_7930 ^ n_6425;
assign n_7943 = n_7931 ^ n_7346;
assign n_7944 = n_7932 ^ n_7346;
assign n_7945 = n_7931 ^ n_7932;
assign n_7946 = n_7934 ^ n_7935;
assign n_7947 = n_7935 ^ x442;
assign n_7948 = n_7936 ^ n_6068;
assign n_7949 = n_7937 ^ n_6109;
assign n_7950 = ~n_7938 & n_7232;
assign n_7951 = n_7618 ^ n_7938;
assign n_7952 = n_7938 ^ n_7219;
assign n_7953 = n_7939 ^ x449;
assign n_7954 = ~n_7939 & n_7940;
assign n_7955 = n_7941 ^ n_5897;
assign n_7956 = n_7942 ^ n_5897;
assign n_7957 = n_7941 ^ n_7942;
assign n_7958 = n_7943 ^ n_7932;
assign n_7959 = n_7944 & n_7945;
assign n_7960 = n_7946 ^ x442;
assign n_7961 = ~n_7946 & n_7947;
assign n_7962 = n_7948 ^ n_6109;
assign n_7963 = n_7937 ^ n_7948;
assign n_7964 = n_7950 ^ n_6894;
assign n_7965 = n_7925 & n_7953;
assign n_7966 = n_7953 ^ n_7925;
assign n_7967 = n_7954 ^ x449;
assign n_7968 = n_7955 ^ n_7942;
assign n_7969 = n_7956 & n_7957;
assign n_7970 = ~n_7341 & n_7958;
assign n_7971 = n_7959 ^ n_7346;
assign n_7972 = n_7960 ^ n_7933;
assign n_7973 = n_7933 & ~n_7960;
assign n_7974 = n_7961 ^ x442;
assign n_7975 = n_7937 ^ n_7962;
assign n_7976 = ~n_7949 & ~n_7963;
assign n_7977 = n_7964 ^ n_6140;
assign n_7978 = n_7967 ^ n_7968;
assign n_7979 = n_7968 ^ x448;
assign n_7980 = n_7969 ^ n_5897;
assign n_7981 = n_7970 ^ n_6466;
assign n_7982 = n_7971 ^ n_7364;
assign n_7983 = n_7972 ^ n_7364;
assign n_7984 = n_7971 ^ n_7972;
assign n_7985 = n_7974 ^ n_7975;
assign n_7986 = n_7975 ^ x441;
assign n_7987 = n_7976 ^ n_6109;
assign n_7988 = n_7978 ^ x448;
assign n_7989 = n_7978 & ~n_7979;
assign n_7990 = n_7980 ^ n_5937;
assign n_7991 = n_7981 ^ n_5937;
assign n_7992 = n_7980 ^ n_7981;
assign n_7993 = n_7982 ^ n_7972;
assign n_7994 = ~n_7983 & n_7984;
assign n_7995 = n_7985 ^ x441;
assign n_7996 = n_7985 & ~n_7986;
assign n_7997 = n_7987 ^ x440;
assign n_7998 = ~n_7965 & n_7988;
assign n_7999 = n_7988 ^ n_7965;
assign n_8000 = n_7989 ^ x448;
assign n_8001 = n_7990 ^ n_7981;
assign n_8002 = n_7991 & ~n_7992;
assign n_8003 = n_7993 & n_7372;
assign n_8004 = n_7994 ^ n_7364;
assign n_8005 = n_7995 ^ n_7973;
assign n_8006 = n_7973 & n_7995;
assign n_8007 = n_7996 ^ x441;
assign n_8008 = n_7997 ^ n_7977;
assign n_8009 = n_8000 ^ n_8001;
assign n_8010 = n_8001 ^ x463;
assign n_8011 = n_8002 ^ n_5937;
assign n_8012 = n_8003 ^ n_6508;
assign n_8013 = n_8004 ^ n_7382;
assign n_8014 = n_8005 ^ n_7382;
assign n_8015 = n_8004 ^ n_8005;
assign n_8016 = n_8007 ^ n_8008;
assign n_8017 = n_8009 ^ x463;
assign n_8018 = ~n_8009 & n_8010;
assign n_8019 = n_8011 ^ n_5979;
assign n_8020 = n_8012 ^ n_5979;
assign n_8021 = n_8011 ^ n_8012;
assign n_8022 = n_8013 ^ n_8005;
assign n_8023 = ~n_8014 & ~n_8015;
assign n_8024 = n_8016 ^ n_8006;
assign n_8025 = n_7998 & ~n_8017;
assign n_8026 = n_8017 ^ n_7998;
assign n_8027 = n_8018 ^ x463;
assign n_8028 = n_8019 ^ n_8012;
assign n_8029 = ~n_8020 & n_8021;
assign n_8030 = n_8022 & ~n_7389;
assign n_8031 = n_8023 ^ n_7382;
assign n_8032 = n_8024 ^ n_7403;
assign n_8033 = n_8027 ^ n_8028;
assign n_8034 = n_8028 ^ x462;
assign n_8035 = n_8029 ^ n_5979;
assign n_8036 = n_8030 ^ n_6550;
assign n_8037 = n_8031 ^ n_7403;
assign n_8038 = n_8031 ^ n_8024;
assign n_8039 = n_8033 ^ x462;
assign n_8040 = n_8033 & ~n_8034;
assign n_8041 = n_8035 ^ n_6019;
assign n_8042 = n_8036 ^ n_6019;
assign n_8043 = n_8035 ^ n_8036;
assign n_8044 = n_8037 ^ n_8024;
assign n_8045 = n_8032 & ~n_8038;
assign n_8046 = n_8025 & n_8039;
assign n_8047 = n_8039 ^ n_8025;
assign n_8048 = n_8040 ^ x462;
assign n_8049 = n_8041 ^ n_8036;
assign n_8050 = ~n_8042 & n_8043;
assign n_8051 = n_7397 & n_8044;
assign n_8052 = n_8045 ^ n_7403;
assign n_8053 = n_8048 ^ n_8049;
assign n_8054 = n_8049 ^ x461;
assign n_8055 = n_8050 ^ n_6019;
assign n_8056 = n_8051 ^ n_6593;
assign n_8057 = n_8052 ^ n_7428;
assign n_8058 = n_8052 ^ n_7150;
assign n_8059 = n_8053 ^ x461;
assign n_8060 = n_8053 & ~n_8054;
assign n_8061 = n_8055 ^ n_6061;
assign n_8062 = n_8056 ^ n_6061;
assign n_8063 = n_8055 ^ n_8056;
assign n_8064 = ~n_8057 & ~n_7429;
assign n_8065 = ~n_7428 & n_8058;
assign n_8066 = ~n_8046 & ~n_8059;
assign n_8067 = n_8059 ^ n_8046;
assign n_8068 = n_8060 ^ x461;
assign n_8069 = n_8061 ^ n_8056;
assign n_8070 = n_8062 & ~n_8063;
assign n_8071 = n_8064 ^ n_6636;
assign n_8072 = n_8065 ^ n_7422;
assign n_8073 = n_8068 ^ n_8069;
assign n_8074 = n_8069 ^ x460;
assign n_8075 = n_8070 ^ n_6061;
assign n_8076 = n_8072 ^ n_7442;
assign n_8077 = n_8073 ^ x460;
assign n_8078 = ~n_8073 & n_8074;
assign n_8079 = n_8075 ^ n_6102;
assign n_8080 = n_8071 ^ n_8075;
assign n_8081 = n_7198 ^ n_8076;
assign n_8082 = ~n_8076 & n_7450;
assign n_8083 = n_8066 & n_8077;
assign n_8084 = n_8077 ^ n_8066;
assign n_8085 = n_8078 ^ x460;
assign n_8086 = n_8071 ^ n_8079;
assign n_8087 = n_8079 & n_8080;
assign n_8088 = n_8081 & n_7449;
assign n_8089 = n_8081 ^ n_7442;
assign n_8090 = n_8082 ^ n_7198;
assign n_8091 = n_8085 ^ n_8086;
assign n_8092 = n_8086 ^ x459;
assign n_8093 = n_8087 ^ n_6102;
assign n_8094 = n_8088 ^ n_6677;
assign n_8095 = n_8090 ^ n_7463;
assign n_8096 = n_8091 ^ x459;
assign n_8097 = n_8091 & ~n_8092;
assign n_8098 = n_8093 ^ n_6147;
assign n_8099 = n_8094 ^ n_6147;
assign n_8100 = n_8093 ^ n_8094;
assign n_8101 = n_7257 ^ n_8095;
assign n_8102 = n_8095 & n_7471;
assign n_8103 = n_8083 & ~n_8096;
assign n_8104 = n_8096 ^ n_8083;
assign n_8105 = n_8097 ^ x459;
assign n_8106 = n_8098 ^ n_8094;
assign n_8107 = ~n_8099 & ~n_8100;
assign n_8108 = n_8101 & n_7470;
assign n_8109 = n_8101 ^ n_7463;
assign n_8110 = n_8102 ^ n_7257;
assign n_8111 = n_8105 ^ n_8106;
assign n_8112 = n_8106 ^ x458;
assign n_8113 = n_8107 ^ n_6147;
assign n_8114 = n_8108 ^ n_6719;
assign n_8115 = n_8110 ^ n_7291;
assign n_8116 = n_8110 ^ n_7484;
assign n_8117 = n_8111 ^ x458;
assign n_8118 = n_8111 & ~n_8112;
assign n_8119 = n_8113 ^ n_6195;
assign n_8120 = n_8114 ^ n_6195;
assign n_8121 = n_8113 ^ n_8114;
assign n_8122 = n_8115 ^ n_7484;
assign n_8123 = n_7491 & n_8116;
assign n_8124 = n_8103 & ~n_8117;
assign n_8125 = n_8117 ^ n_8103;
assign n_8126 = n_8118 ^ x458;
assign n_8127 = n_8119 ^ n_8114;
assign n_8128 = n_8120 & ~n_8121;
assign n_8129 = ~n_8122 & n_7490;
assign n_8130 = n_8123 ^ n_7291;
assign n_8131 = n_8126 ^ n_8127;
assign n_8132 = n_8127 ^ x457;
assign n_8133 = n_8128 ^ n_6195;
assign n_8134 = n_8129 ^ n_6761;
assign n_8135 = n_8130 ^ n_7504;
assign n_8136 = n_8131 ^ x457;
assign n_8137 = n_8131 & ~n_8132;
assign n_8138 = n_8133 ^ n_6237;
assign n_8139 = n_8134 ^ n_6237;
assign n_8140 = n_8133 ^ n_8134;
assign n_8141 = n_7312 ^ n_8135;
assign n_8142 = n_8135 & n_7512;
assign n_8143 = ~n_8124 & n_8136;
assign n_8144 = n_8136 ^ n_8124;
assign n_8145 = n_8137 ^ x457;
assign n_8146 = n_8138 ^ n_8134;
assign n_8147 = n_8139 & n_8140;
assign n_8148 = n_8141 & ~n_7511;
assign n_8149 = n_8141 ^ n_7504;
assign n_8150 = n_8142 ^ n_7312;
assign n_8151 = n_8145 ^ n_8146;
assign n_8152 = n_8146 ^ x456;
assign n_8153 = n_8147 ^ n_6237;
assign n_8154 = n_8148 ^ n_6803;
assign n_8155 = n_8150 ^ n_7330;
assign n_8156 = n_8150 ^ n_7526;
assign n_8157 = n_8151 ^ x456;
assign n_8158 = n_8151 & ~n_8152;
assign n_8159 = n_8153 ^ n_8154;
assign n_8160 = n_8154 ^ n_6274;
assign n_8161 = n_8155 ^ n_7526;
assign n_8162 = ~n_7532 & ~n_8156;
assign n_8163 = n_8143 ^ n_8157;
assign n_8164 = ~n_8157 & ~n_8143;
assign n_8165 = n_8158 ^ x456;
assign n_8166 = n_8159 ^ n_6274;
assign n_8167 = ~n_8159 & n_8160;
assign n_8168 = n_7520 & n_8161;
assign n_8169 = n_8161 ^ n_7682;
assign n_8170 = n_8162 ^ n_7330;
assign n_8171 = n_8163 ^ n_7645;
assign n_8172 = n_8163 ^ n_7114;
assign n_8173 = n_7645 & n_8163;
assign n_8174 = n_8165 ^ n_8166;
assign n_8175 = n_8166 ^ x471;
assign n_8176 = n_8167 ^ n_6274;
assign n_8177 = n_8168 ^ n_6845;
assign n_8178 = n_8170 ^ n_7545;
assign n_8179 = n_7638 & ~n_8172;
assign n_8180 = n_8173 ^ n_7673;
assign n_8181 = n_8174 ^ x471;
assign n_8182 = ~n_8174 & n_8175;
assign n_8183 = n_8176 ^ n_6313;
assign n_8184 = n_8177 ^ n_6313;
assign n_8185 = n_8176 ^ n_8177;
assign n_8186 = n_7352 ^ n_8178;
assign n_8187 = n_8178 & n_7553;
assign n_8188 = n_8179 ^ n_7114;
assign n_8189 = n_8164 ^ n_8181;
assign n_8190 = ~n_8181 & ~n_8164;
assign n_8191 = n_8182 ^ x471;
assign n_8192 = n_8183 ^ n_8177;
assign n_8193 = n_8184 & n_8185;
assign n_8194 = n_8186 & n_7552;
assign n_8195 = n_8186 ^ n_7717;
assign n_8196 = n_8186 ^ n_7545;
assign n_8197 = n_8187 ^ n_7352;
assign n_8198 = n_8188 ^ n_6127;
assign n_8199 = n_6127 & n_8188;
assign n_8200 = n_8189 ^ n_8180;
assign n_8201 = n_8189 ^ n_8173;
assign n_8202 = n_8191 ^ n_8192;
assign n_8203 = n_8192 ^ x470;
assign n_8204 = n_8193 ^ n_6313;
assign n_8205 = n_8194 ^ n_6887;
assign n_8206 = n_8197 ^ n_7566;
assign n_8207 = x487 & n_8198;
assign n_8208 = n_8198 ^ x487;
assign n_8209 = n_8199 ^ n_6172;
assign n_8210 = n_7674 & ~n_8200;
assign n_8211 = n_8180 & n_8201;
assign n_8212 = n_8202 ^ x470;
assign n_8213 = ~n_8202 & n_8203;
assign n_8214 = n_8204 ^ n_8205;
assign n_8215 = n_8205 ^ n_6350;
assign n_8216 = n_7370 ^ n_8206;
assign n_8217 = n_8206 & ~n_7573;
assign n_8218 = n_8207 ^ x486;
assign n_8219 = n_8210 ^ n_7142;
assign n_8220 = n_8211 ^ n_7673;
assign n_8221 = n_8212 ^ n_8190;
assign n_8222 = ~n_8190 & n_8212;
assign n_8223 = n_8213 ^ x470;
assign n_8224 = n_8214 ^ n_6350;
assign n_8225 = ~n_8214 & ~n_8215;
assign n_8226 = n_8216 & n_7572;
assign n_8227 = n_7789 ^ n_8216;
assign n_8228 = n_8216 ^ n_7566;
assign n_8229 = n_8217 ^ n_7370;
assign n_8230 = n_8219 ^ n_8209;
assign n_8231 = n_8219 ^ n_8199;
assign n_8232 = n_8220 ^ n_7719;
assign n_8233 = n_8221 ^ n_7719;
assign n_8234 = n_8220 ^ n_8221;
assign n_8235 = n_8223 ^ n_8224;
assign n_8236 = n_8224 ^ x469;
assign n_8237 = n_8225 ^ n_6350;
assign n_8238 = n_8226 ^ n_6926;
assign n_8239 = n_8229 ^ n_7586;
assign n_8240 = n_8230 ^ n_8207;
assign n_8241 = n_8230 ^ n_8218;
assign n_8242 = n_8209 & ~n_8231;
assign n_8243 = n_8232 ^ n_8221;
assign n_8244 = ~n_8233 & n_8234;
assign n_8245 = n_8235 ^ x469;
assign n_8246 = ~n_8235 & n_8236;
assign n_8247 = n_8237 ^ n_6390;
assign n_8248 = n_8238 ^ n_6390;
assign n_8249 = n_8237 ^ n_8238;
assign n_8250 = n_7392 ^ n_8239;
assign n_8251 = ~n_8239 & ~n_7594;
assign n_8252 = n_8218 & ~n_8240;
assign n_8253 = n_8208 & n_8241;
assign n_8254 = n_8241 ^ n_8208;
assign n_8255 = n_8242 ^ n_6172;
assign n_8256 = ~n_7709 & ~n_8243;
assign n_8257 = n_8244 ^ n_7719;
assign n_8258 = n_8245 ^ n_8222;
assign n_8259 = n_8222 & n_8245;
assign n_8260 = n_8246 ^ x469;
assign n_8261 = n_8247 ^ n_8238;
assign n_8262 = n_8248 & ~n_8249;
assign n_8263 = n_8250 & ~n_7593;
assign n_8264 = n_8250 ^ n_7844;
assign n_8265 = n_8250 ^ n_7586;
assign n_8266 = n_8251 ^ n_7392;
assign n_8267 = n_8252 ^ x486;
assign n_8268 = n_8255 ^ n_6230;
assign n_8269 = n_8256 ^ n_7182;
assign n_8270 = n_8257 ^ n_7753;
assign n_8271 = n_8258 ^ n_7753;
assign n_8272 = n_8257 ^ n_8258;
assign n_8273 = n_8260 ^ n_8261;
assign n_8274 = n_8261 ^ x468;
assign n_8275 = n_8262 ^ n_6390;
assign n_8276 = n_8263 ^ n_6957;
assign n_8277 = n_8266 ^ n_7607;
assign n_8278 = n_8268 ^ n_8269;
assign n_8279 = n_8269 ^ n_6230;
assign n_8280 = n_8255 ^ n_8269;
assign n_8281 = n_8270 ^ n_8258;
assign n_8282 = ~n_8271 & ~n_8272;
assign n_8283 = n_8273 ^ x468;
assign n_8284 = ~n_8273 & n_8274;
assign n_8285 = n_8275 ^ n_6432;
assign n_8286 = n_8276 ^ n_6432;
assign n_8287 = n_8275 ^ n_8276;
assign n_8288 = n_7412 ^ n_8277;
assign n_8289 = ~n_8277 & ~n_7615;
assign n_8290 = n_8267 ^ n_8278;
assign n_8291 = n_8278 ^ x485;
assign n_8292 = n_8279 & n_8280;
assign n_8293 = ~n_7743 & ~n_8281;
assign n_8294 = n_8282 ^ n_7753;
assign n_8295 = n_8283 ^ n_8259;
assign n_8296 = ~n_8259 & ~n_8283;
assign n_8297 = n_8284 ^ x468;
assign n_8298 = n_8285 ^ n_8276;
assign n_8299 = ~n_8286 & ~n_8287;
assign n_8300 = ~n_8288 & n_7614;
assign n_8301 = n_7885 ^ n_8288;
assign n_8302 = n_8288 ^ n_7607;
assign n_8303 = n_8289 ^ n_7412;
assign n_8304 = n_8290 ^ x485;
assign n_8305 = ~n_8290 & n_8291;
assign n_8306 = n_8292 ^ n_6230;
assign n_8307 = n_8293 ^ n_7223;
assign n_8308 = n_8294 ^ n_7794;
assign n_8309 = n_8295 ^ n_7794;
assign n_8310 = n_8294 ^ n_8295;
assign n_8311 = n_8297 ^ n_8298;
assign n_8312 = n_8298 ^ x467;
assign n_8313 = n_8299 ^ n_6432;
assign n_8314 = n_8300 ^ n_6980;
assign n_8315 = n_8303 ^ n_7628;
assign n_8316 = n_8253 & n_8304;
assign n_8317 = n_8304 ^ n_8253;
assign n_8318 = n_8305 ^ x485;
assign n_8319 = n_8306 ^ n_6267;
assign n_8320 = n_8307 ^ n_6267;
assign n_8321 = n_8306 ^ n_8307;
assign n_8322 = n_8308 ^ n_8295;
assign n_8323 = ~n_8309 & ~n_8310;
assign n_8324 = n_8311 ^ x467;
assign n_8325 = n_8311 & ~n_8312;
assign n_8326 = n_8313 ^ n_6473;
assign n_8327 = n_8314 ^ n_6473;
assign n_8328 = n_8313 ^ n_8314;
assign n_8329 = n_7432 ^ n_8315;
assign n_8330 = n_8315 & ~n_7636;
assign n_8331 = n_8319 ^ n_8307;
assign n_8332 = ~n_8320 & n_8321;
assign n_8333 = ~n_7781 & n_8322;
assign n_8334 = n_8323 ^ n_7794;
assign n_8335 = n_8324 ^ n_8296;
assign n_8336 = n_8296 & n_8324;
assign n_8337 = n_8325 ^ x467;
assign n_8338 = n_8326 ^ n_8314;
assign n_8339 = ~n_8327 & n_8328;
assign n_8340 = n_8329 & ~n_7635;
assign n_8341 = n_8329 ^ n_7628;
assign n_8342 = n_8329 ^ n_7926;
assign n_8343 = n_8330 ^ n_7432;
assign n_8344 = n_8318 ^ n_8331;
assign n_8345 = n_8331 ^ x484;
assign n_8346 = n_8332 ^ n_6267;
assign n_8347 = n_8333 ^ n_7261;
assign n_8348 = n_8334 ^ n_7833;
assign n_8349 = n_8335 ^ n_7833;
assign n_8350 = n_8334 ^ n_8335;
assign n_8351 = n_8337 ^ n_8338;
assign n_8352 = n_8338 ^ x466;
assign n_8353 = n_8339 ^ n_6473;
assign n_8354 = n_8340 ^ n_7000;
assign n_8355 = n_8343 ^ n_7651;
assign n_8356 = n_8344 ^ x484;
assign n_8357 = ~n_8344 & n_8345;
assign n_8358 = n_8346 ^ n_6307;
assign n_8359 = n_8347 ^ n_6307;
assign n_8360 = n_8346 ^ n_8347;
assign n_8361 = n_8348 ^ n_8335;
assign n_8362 = n_8349 & n_8350;
assign n_8363 = n_8351 ^ x466;
assign n_8364 = ~n_8351 & n_8352;
assign n_8365 = n_8353 ^ n_6514;
assign n_8366 = n_8354 ^ n_6514;
assign n_8367 = n_8353 ^ n_8354;
assign n_8368 = n_7453 ^ n_8355;
assign n_8369 = n_8355 & ~n_7661;
assign n_8370 = n_8356 & n_8316;
assign n_8371 = n_8316 ^ n_8356;
assign n_8372 = n_8357 ^ x484;
assign n_8373 = n_8358 ^ n_8347;
assign n_8374 = ~n_8359 & ~n_8360;
assign n_8375 = ~n_7821 & n_8361;
assign n_8376 = n_8362 ^ n_7833;
assign n_8377 = n_8363 ^ n_8336;
assign n_8378 = n_8336 & ~n_8363;
assign n_8379 = n_8364 ^ x466;
assign n_8380 = n_8365 ^ n_8354;
assign n_8381 = n_8366 & ~n_8367;
assign n_8382 = n_8368 & n_7660;
assign n_8383 = n_8368 ^ n_7651;
assign n_8384 = n_7966 ^ n_8368;
assign n_8385 = n_8369 ^ n_7453;
assign n_8386 = n_8372 ^ n_8373;
assign n_8387 = n_8373 ^ x483;
assign n_8388 = n_8374 ^ n_6307;
assign n_8389 = n_8375 ^ n_7287;
assign n_8390 = n_8376 ^ n_7874;
assign n_8391 = n_8377 ^ n_7874;
assign n_8392 = n_8376 ^ n_8377;
assign n_8393 = n_8379 ^ n_8380;
assign n_8394 = n_8380 ^ x465;
assign n_8395 = n_8381 ^ n_6514;
assign n_8396 = n_8382 ^ n_7021;
assign n_8397 = n_8385 ^ n_7679;
assign n_8398 = n_8386 ^ x483;
assign n_8399 = ~n_8386 & n_8387;
assign n_8400 = n_8388 ^ n_6344;
assign n_8401 = n_8389 ^ n_6344;
assign n_8402 = n_8388 ^ n_8389;
assign n_8403 = n_8390 ^ n_8377;
assign n_8404 = ~n_8391 & n_8392;
assign n_8405 = n_8393 ^ x465;
assign n_8406 = n_8393 & ~n_8394;
assign n_8407 = n_8395 ^ n_6557;
assign n_8408 = n_8396 ^ n_6557;
assign n_8409 = n_8395 ^ n_8396;
assign n_8410 = n_7474 ^ n_8397;
assign n_8411 = ~n_8397 & ~n_7692;
assign n_8412 = n_8370 & n_8398;
assign n_8413 = n_8398 ^ n_8370;
assign n_8414 = n_8399 ^ x483;
assign n_8415 = n_8400 ^ n_8389;
assign n_8416 = n_8401 & ~n_8402;
assign n_8417 = ~n_7862 & n_8403;
assign n_8418 = n_8404 ^ n_7874;
assign n_8419 = n_8405 ^ n_8378;
assign n_8420 = n_8378 & n_8405;
assign n_8421 = n_8406 ^ x465;
assign n_8422 = n_8407 ^ n_8396;
assign n_8423 = n_8408 & n_8409;
assign n_8424 = n_8410 & n_7691;
assign n_8425 = n_8410 ^ n_7999;
assign n_8426 = n_8410 ^ n_7679;
assign n_8427 = n_8411 ^ n_7474;
assign n_8428 = n_8414 ^ n_8415;
assign n_8429 = n_8415 ^ x482;
assign n_8430 = n_8416 ^ n_6344;
assign n_8431 = n_8417 ^ n_7303;
assign n_8432 = n_8418 ^ n_7915;
assign n_8433 = n_8419 ^ n_7915;
assign n_8434 = n_8418 ^ n_8419;
assign n_8435 = n_8421 ^ n_8422;
assign n_8436 = n_8422 ^ x464;
assign n_8437 = n_8423 ^ n_6557;
assign n_8438 = n_8424 ^ n_7036;
assign n_8439 = n_8427 ^ n_7494;
assign n_8440 = n_8427 ^ n_7714;
assign n_8441 = n_8428 ^ x482;
assign n_8442 = ~n_8428 & n_8429;
assign n_8443 = n_8430 ^ n_6383;
assign n_8444 = n_8431 ^ n_6383;
assign n_8445 = n_8430 ^ n_8431;
assign n_8446 = n_8432 ^ n_8419;
assign n_8447 = n_8433 & ~n_8434;
assign n_8448 = n_8435 ^ x464;
assign n_8449 = n_8435 & ~n_8436;
assign n_8450 = n_8438 ^ n_6599;
assign n_8451 = n_8437 ^ n_8438;
assign n_8452 = n_8439 ^ n_7714;
assign n_8453 = ~n_7725 & ~n_8440;
assign n_8454 = ~n_8412 & ~n_8441;
assign n_8455 = n_8441 ^ n_8412;
assign n_8456 = n_8442 ^ x482;
assign n_8457 = n_8443 ^ n_8431;
assign n_8458 = ~n_8444 & ~n_8445;
assign n_8459 = ~n_7904 & ~n_8446;
assign n_8460 = n_8447 ^ n_7915;
assign n_8461 = n_8448 ^ n_8420;
assign n_8462 = ~n_8420 & ~n_8448;
assign n_8463 = n_8449 ^ x464;
assign n_8464 = n_8437 ^ n_8450;
assign n_8465 = n_8450 & n_8451;
assign n_8466 = n_7703 & ~n_8452;
assign n_8467 = n_8452 ^ n_8026;
assign n_8468 = n_8453 ^ n_7494;
assign n_8469 = n_8456 ^ n_8457;
assign n_8470 = n_8457 ^ x481;
assign n_8471 = n_8458 ^ n_6383;
assign n_8472 = n_8459 ^ n_7328;
assign n_8473 = n_8460 ^ n_7958;
assign n_8474 = n_8461 ^ n_7958;
assign n_8475 = n_8460 ^ n_8461;
assign n_8476 = n_8463 ^ x479;
assign n_8477 = n_8464 ^ n_8463;
assign n_8478 = n_8465 ^ n_6599;
assign n_8479 = n_8466 ^ n_7061;
assign n_8480 = n_8468 ^ n_7748;
assign n_8481 = n_8469 ^ x481;
assign n_8482 = n_8469 & ~n_8470;
assign n_8483 = n_8471 ^ n_6425;
assign n_8484 = n_8472 ^ n_6425;
assign n_8485 = n_8471 ^ n_8472;
assign n_8486 = n_8473 ^ n_8461;
assign n_8487 = n_8474 & n_8475;
assign n_8488 = n_8477 ^ x479;
assign n_8489 = ~n_8477 & n_8476;
assign n_8490 = n_8478 ^ n_6642;
assign n_8491 = n_8479 ^ n_6642;
assign n_8492 = n_8478 ^ n_8479;
assign n_8493 = n_7515 ^ n_8480;
assign n_8494 = ~n_8480 & ~n_7761;
assign n_8495 = ~n_8454 & ~n_8481;
assign n_8496 = n_8481 ^ n_8454;
assign n_8497 = n_8482 ^ x481;
assign n_8498 = n_8483 ^ n_8472;
assign n_8499 = n_8484 & n_8485;
assign n_8500 = ~n_7945 & ~n_8486;
assign n_8501 = n_8487 ^ n_7958;
assign n_8502 = n_8488 ^ n_8462;
assign n_8503 = n_8462 & n_8488;
assign n_8504 = n_8489 ^ x479;
assign n_8505 = n_8490 ^ n_8479;
assign n_8506 = ~n_8491 & n_8492;
assign n_8507 = n_8493 & ~n_7760;
assign n_8508 = n_8493 ^ n_7748;
assign n_8509 = n_8047 ^ n_8493;
assign n_8510 = n_8494 ^ n_7515;
assign n_8511 = n_8497 ^ n_8498;
assign n_8512 = n_8498 ^ x480;
assign n_8513 = n_8499 ^ n_6425;
assign n_8514 = n_8500 ^ n_7346;
assign n_8515 = n_8501 ^ n_7993;
assign n_8516 = n_8502 ^ n_7993;
assign n_8517 = n_8501 ^ n_8502;
assign n_8518 = n_8504 ^ n_8505;
assign n_8519 = n_8505 ^ x478;
assign n_8520 = n_8506 ^ n_6642;
assign n_8521 = n_8507 ^ n_7081;
assign n_8522 = n_8510 ^ n_7786;
assign n_8523 = n_8511 ^ x480;
assign n_8524 = n_8511 & ~n_8512;
assign n_8525 = n_8513 ^ n_6466;
assign n_8526 = n_8514 ^ n_6466;
assign n_8527 = n_8513 ^ n_8514;
assign n_8528 = n_8515 ^ n_8502;
assign n_8529 = n_8516 & ~n_8517;
assign n_8530 = n_8518 ^ x478;
assign n_8531 = ~n_8518 & n_8519;
assign n_8532 = n_8520 ^ n_6683;
assign n_8533 = n_8521 ^ n_6683;
assign n_8534 = n_8520 ^ n_8521;
assign n_8535 = n_7535 ^ n_8522;
assign n_8536 = ~n_8522 & ~n_7802;
assign n_8537 = n_8495 & ~n_8523;
assign n_8538 = n_8523 ^ n_8495;
assign n_8539 = n_8524 ^ x480;
assign n_8540 = n_8525 ^ n_8514;
assign n_8541 = ~n_8526 & n_8527;
assign n_8542 = ~n_7984 & n_8528;
assign n_8543 = n_8529 ^ n_7993;
assign n_8544 = n_8530 ^ n_8503;
assign n_8545 = ~n_8503 & ~n_8530;
assign n_8546 = n_8531 ^ x478;
assign n_8547 = n_8532 ^ n_8521;
assign n_8548 = n_8533 & n_8534;
assign n_8549 = ~n_8535 & n_7801;
assign n_8550 = n_8535 ^ n_7786;
assign n_8551 = n_8067 ^ n_8535;
assign n_8552 = n_8536 ^ n_7535;
assign n_8553 = n_8539 ^ n_8540;
assign n_8554 = n_8540 ^ x495;
assign n_8555 = n_8541 ^ n_6466;
assign n_8556 = n_8542 ^ n_7364;
assign n_8557 = n_8543 ^ n_8022;
assign n_8558 = n_8544 ^ n_8543;
assign n_8559 = n_8546 ^ n_8547;
assign n_8560 = n_8547 ^ x477;
assign n_8561 = n_8548 ^ n_6683;
assign n_8562 = n_8549 ^ n_7102;
assign n_8563 = n_8552 ^ n_7826;
assign n_8564 = n_8553 ^ x495;
assign n_8565 = n_8553 & ~n_8554;
assign n_8566 = n_8555 ^ n_6508;
assign n_8567 = n_8556 ^ n_6508;
assign n_8568 = n_8555 ^ n_8556;
assign n_8569 = n_8544 ^ n_8557;
assign n_8570 = n_8557 & n_8558;
assign n_8571 = n_8559 ^ x477;
assign n_8572 = n_8559 & ~n_8560;
assign n_8573 = n_8561 ^ n_6725;
assign n_8574 = n_8562 ^ n_6725;
assign n_8575 = n_8561 ^ n_8562;
assign n_8576 = n_7556 ^ n_8563;
assign n_8577 = ~n_8563 & n_7841;
assign n_8578 = n_8537 & ~n_8564;
assign n_8579 = n_8564 ^ n_8537;
assign n_8580 = n_8565 ^ x495;
assign n_8581 = n_8566 ^ n_8556;
assign n_8582 = n_8567 & n_8568;
assign n_8583 = n_8015 & ~n_8569;
assign n_8584 = n_8570 ^ n_8022;
assign n_8585 = n_8545 ^ n_8571;
assign n_8586 = n_8571 & n_8545;
assign n_8587 = n_8572 ^ x477;
assign n_8588 = n_8573 ^ n_8562;
assign n_8589 = ~n_8574 & ~n_8575;
assign n_8590 = ~n_8576 & n_7840;
assign n_8591 = n_8576 ^ n_7826;
assign n_8592 = n_8084 ^ n_8576;
assign n_8593 = n_8577 ^ n_7556;
assign n_8594 = n_8580 ^ n_8581;
assign n_8595 = n_8581 ^ x494;
assign n_8596 = n_8582 ^ n_6508;
assign n_8597 = n_8583 ^ n_7382;
assign n_8598 = n_8584 ^ n_8044;
assign n_8599 = n_8585 ^ n_8044;
assign n_8600 = n_8584 ^ n_8585;
assign n_8601 = n_8587 ^ n_8588;
assign n_8602 = n_8588 ^ x476;
assign n_8603 = n_8589 ^ n_6725;
assign n_8604 = n_8590 ^ n_7127;
assign n_8605 = n_8593 ^ n_7576;
assign n_8606 = n_8593 ^ n_7867;
assign n_8607 = n_8594 ^ x494;
assign n_8608 = ~n_8594 & n_8595;
assign n_8609 = n_8596 ^ n_6550;
assign n_8610 = n_8597 ^ n_6550;
assign n_8611 = n_8596 ^ n_8597;
assign n_8612 = n_8598 ^ n_8585;
assign n_8613 = ~n_8599 & n_8600;
assign n_8614 = n_8601 ^ x476;
assign n_8615 = n_8601 & ~n_8602;
assign n_8616 = n_8603 ^ n_6767;
assign n_8617 = n_8604 ^ n_6767;
assign n_8618 = n_8603 ^ n_8604;
assign n_8619 = n_8605 ^ n_7867;
assign n_8620 = ~n_7882 & n_8606;
assign n_8621 = n_8578 & n_8607;
assign n_8622 = n_8607 ^ n_8578;
assign n_8623 = n_8608 ^ x494;
assign n_8624 = n_8609 ^ n_8597;
assign n_8625 = ~n_8610 & n_8611;
assign n_8626 = n_8038 & ~n_8612;
assign n_8627 = n_8613 ^ n_8044;
assign n_8628 = n_8586 ^ n_8614;
assign n_8629 = ~n_8614 & ~n_8586;
assign n_8630 = n_8615 ^ x476;
assign n_8631 = n_8616 ^ n_8604;
assign n_8632 = ~n_8617 & ~n_8618;
assign n_8633 = n_8619 & ~n_7881;
assign n_8634 = n_8104 ^ n_8619;
assign n_8635 = n_8620 ^ n_7576;
assign n_8636 = n_8623 ^ n_8624;
assign n_8637 = n_8624 ^ x493;
assign n_8638 = n_8625 ^ n_6550;
assign n_8639 = n_8626 ^ n_7403;
assign n_8640 = n_8627 ^ n_8057;
assign n_8641 = n_8628 ^ n_8057;
assign n_8642 = n_8627 ^ n_8628;
assign n_8643 = n_8630 ^ n_8631;
assign n_8644 = n_8631 ^ x475;
assign n_8645 = n_8632 ^ n_6767;
assign n_8646 = n_8633 ^ n_7158;
assign n_8647 = n_8635 ^ n_7909;
assign n_8648 = n_8636 ^ x493;
assign n_8649 = ~n_8636 & n_8637;
assign n_8650 = n_8638 ^ n_6593;
assign n_8651 = n_8639 ^ n_8638;
assign n_8652 = n_8640 ^ n_8628;
assign n_8653 = ~n_8641 & ~n_8642;
assign n_8654 = n_8643 ^ x475;
assign n_8655 = ~n_8643 & n_8644;
assign n_8656 = n_8645 ^ n_6810;
assign n_8657 = n_8646 ^ n_6810;
assign n_8658 = n_8645 ^ n_8646;
assign n_8659 = n_8647 ^ n_7597;
assign n_8660 = n_8647 & n_7923;
assign n_8661 = n_8621 ^ n_8648;
assign n_8662 = n_8648 & n_8621;
assign n_8663 = n_8649 ^ x493;
assign n_8664 = n_8639 ^ n_8650;
assign n_8665 = ~n_8650 & n_8651;
assign n_8666 = ~n_8058 & ~n_8652;
assign n_8667 = n_8653 ^ n_8057;
assign n_8668 = n_8654 ^ n_8629;
assign n_8669 = n_8629 & n_8654;
assign n_8670 = n_8655 ^ x475;
assign n_8671 = n_8656 ^ n_8646;
assign n_8672 = ~n_8657 & n_8658;
assign n_8673 = ~n_8659 & ~n_7922;
assign n_8674 = n_8659 ^ n_7909;
assign n_8675 = n_8125 ^ n_8659;
assign n_8676 = n_8660 ^ n_7597;
assign n_8677 = n_8171 ^ n_8661;
assign n_8678 = n_8661 & n_8171;
assign n_8679 = n_8663 ^ n_8664;
assign n_8680 = n_8664 ^ x492;
assign n_8681 = n_8665 ^ n_6593;
assign n_8682 = n_8666 ^ n_7422;
assign n_8683 = n_8667 ^ n_8081;
assign n_8684 = n_8668 ^ n_8081;
assign n_8685 = n_8667 ^ n_8668;
assign n_8686 = n_8670 ^ n_8671;
assign n_8687 = n_8671 ^ x474;
assign n_8688 = n_8672 ^ n_6810;
assign n_8689 = n_8673 ^ n_7192;
assign n_8690 = n_8676 ^ n_7951;
assign n_8691 = n_8677 ^ n_8163;
assign n_8692 = n_8678 ^ n_8200;
assign n_8693 = n_8679 ^ x492;
assign n_8694 = n_8679 & ~n_8680;
assign n_8695 = n_8681 ^ n_6636;
assign n_8696 = n_8682 ^ n_6636;
assign n_8697 = n_8681 ^ n_8682;
assign n_8698 = n_8683 ^ n_8668;
assign n_8699 = n_8684 & n_8685;
assign n_8700 = n_8686 ^ x474;
assign n_8701 = n_8686 & ~n_8687;
assign n_8702 = n_8688 ^ n_6852;
assign n_8703 = n_8689 ^ n_6852;
assign n_8704 = n_8689 ^ n_8688;
assign n_8705 = ~n_8690 & ~n_7952;
assign n_8706 = n_8690 ^ n_7938;
assign n_8707 = n_7645 & n_8691;
assign n_8708 = n_8693 & ~n_8662;
assign n_8709 = n_8662 ^ n_8693;
assign n_8710 = n_8694 ^ x492;
assign n_8711 = n_8695 ^ n_8682;
assign n_8712 = ~n_8696 & ~n_8697;
assign n_8713 = ~n_8698 & n_8089;
assign n_8714 = n_8699 ^ n_8081;
assign n_8715 = n_8700 ^ n_8669;
assign n_8716 = ~n_8669 & n_8700;
assign n_8717 = n_8701 ^ x474;
assign n_8718 = n_8689 ^ n_8702;
assign n_8719 = ~n_8703 & n_8704;
assign n_8720 = n_8705 ^ n_7219;
assign n_8721 = n_8707 ^ n_8163;
assign n_8722 = n_8678 ^ n_8709;
assign n_8723 = n_8692 ^ n_8709;
assign n_8724 = n_8710 ^ n_8711;
assign n_8725 = n_8711 ^ x491;
assign n_8726 = n_8712 ^ n_6636;
assign n_8727 = n_8713 ^ n_7442;
assign n_8728 = n_8714 ^ n_8101;
assign n_8729 = n_8715 ^ n_8101;
assign n_8730 = n_8714 ^ n_8715;
assign n_8731 = n_8717 ^ n_8718;
assign n_8732 = n_8718 ^ x473;
assign n_8733 = n_8719 ^ n_6852;
assign n_8734 = n_8720 ^ n_6894;
assign n_8735 = n_8721 ^ n_7114;
assign n_8736 = n_7114 & n_8721;
assign n_8737 = ~n_8722 & ~n_8692;
assign n_8738 = n_7673 & n_8722;
assign n_8739 = n_8724 ^ x491;
assign n_8740 = n_8724 & ~n_8725;
assign n_8741 = n_8726 ^ n_6677;
assign n_8742 = n_8727 ^ n_6677;
assign n_8743 = n_8726 ^ n_8727;
assign n_8744 = n_8728 ^ n_8715;
assign n_8745 = n_8729 & ~n_8730;
assign n_8746 = n_8731 ^ x473;
assign n_8747 = n_8731 & ~n_8732;
assign n_8748 = n_8733 ^ x472;
assign n_8749 = n_8735 ^ x39;
assign n_8750 = x39 & n_8735;
assign n_8751 = n_8736 ^ n_7142;
assign n_8752 = n_8737 ^ n_8200;
assign n_8753 = n_8738 ^ n_8200;
assign n_8754 = ~n_8708 & ~n_8739;
assign n_8755 = n_8739 ^ n_8708;
assign n_8756 = n_8740 ^ x491;
assign n_8757 = n_8741 ^ n_8727;
assign n_8758 = n_8742 & n_8743;
assign n_8759 = n_8744 & ~n_8109;
assign n_8760 = n_8745 ^ n_8101;
assign n_8761 = n_8746 ^ n_8716;
assign n_8762 = ~n_8716 & ~n_8746;
assign n_8763 = n_8747 ^ x473;
assign n_8764 = n_8748 ^ n_8734;
assign n_8765 = n_8750 ^ x38;
assign n_8766 = n_8752 ^ n_8243;
assign n_8767 = n_8753 ^ n_8736;
assign n_8768 = n_8753 ^ n_8751;
assign n_8769 = n_8755 ^ n_8752;
assign n_8770 = n_8755 ^ n_8243;
assign n_8771 = n_8756 ^ n_8757;
assign n_8772 = n_8757 ^ x490;
assign n_8773 = n_8758 ^ n_6677;
assign n_8774 = n_8759 ^ n_7463;
assign n_8775 = n_8760 ^ n_8122;
assign n_8776 = n_8761 ^ n_8122;
assign n_8777 = n_8760 ^ n_8761;
assign n_8778 = n_8763 ^ n_8764;
assign n_8779 = n_8766 ^ n_8755;
assign n_8780 = n_8751 & n_8767;
assign n_8781 = n_8768 ^ n_8750;
assign n_8782 = n_8768 ^ n_8765;
assign n_8783 = n_7719 & ~n_8769;
assign n_8784 = n_8769 & ~n_8770;
assign n_8785 = n_8771 ^ x490;
assign n_8786 = n_8771 & ~n_8772;
assign n_8787 = n_8773 ^ n_6719;
assign n_8788 = n_8774 ^ n_6719;
assign n_8789 = n_8773 ^ n_8774;
assign n_8790 = n_8775 ^ n_8761;
assign n_8791 = ~n_8776 & ~n_8777;
assign n_8792 = n_8778 ^ n_8762;
assign n_8793 = n_8780 ^ n_7142;
assign n_8794 = n_8765 & n_8781;
assign n_8795 = n_8783 ^ n_8243;
assign n_8796 = n_8784 ^ n_8243;
assign n_8797 = n_8754 & ~n_8785;
assign n_8798 = n_8785 ^ n_8754;
assign n_8799 = n_8786 ^ x490;
assign n_8800 = n_8787 ^ n_8774;
assign n_8801 = n_8788 & n_8789;
assign n_8802 = ~n_8115 & ~n_8790;
assign n_8803 = n_8791 ^ n_8122;
assign n_8804 = n_8792 ^ n_8141;
assign n_8805 = n_8793 ^ n_7182;
assign n_8806 = n_8794 ^ x38;
assign n_8807 = n_8795 ^ n_7182;
assign n_8808 = n_8793 ^ n_8795;
assign n_8809 = n_8796 ^ n_8281;
assign n_8810 = n_8798 ^ n_8796;
assign n_8811 = n_8798 ^ n_8281;
assign n_8812 = n_8799 ^ n_8800;
assign n_8813 = n_8800 ^ x489;
assign n_8814 = n_8801 ^ n_6719;
assign n_8815 = n_8802 ^ n_7484;
assign n_8816 = n_8803 ^ n_8792;
assign n_8817 = n_8803 ^ n_8141;
assign n_8818 = n_8805 ^ n_8795;
assign n_8819 = n_8807 & n_8808;
assign n_8820 = n_8809 ^ n_8798;
assign n_8821 = ~n_7753 & n_8810;
assign n_8822 = ~n_8810 & n_8811;
assign n_8823 = n_8812 ^ x489;
assign n_8824 = ~n_8812 & n_8813;
assign n_8825 = n_8814 ^ n_6761;
assign n_8826 = n_8815 ^ n_6761;
assign n_8827 = n_8814 ^ n_8815;
assign n_8828 = ~n_8804 & ~n_8816;
assign n_8829 = n_8817 ^ n_8792;
assign n_8830 = n_8806 ^ n_8818;
assign n_8831 = n_8818 ^ x37;
assign n_8832 = n_8819 ^ n_7182;
assign n_8833 = n_8821 ^ n_8281;
assign n_8834 = n_8822 ^ n_8281;
assign n_8835 = n_8823 ^ n_8797;
assign n_8836 = n_8797 & n_8823;
assign n_8837 = n_8824 ^ x489;
assign n_8838 = n_8825 ^ n_8815;
assign n_8839 = n_8826 & n_8827;
assign n_8840 = n_8828 ^ n_8141;
assign n_8841 = n_8829 & ~n_8149;
assign n_8842 = n_8830 ^ x37;
assign n_8843 = ~n_8830 & n_8831;
assign n_8844 = n_8832 ^ n_7223;
assign n_8845 = n_8833 ^ n_7223;
assign n_8846 = n_8832 ^ n_8833;
assign n_8847 = n_8834 ^ n_8322;
assign n_8848 = n_8835 ^ n_8834;
assign n_8849 = n_8835 ^ n_8322;
assign n_8850 = n_8837 ^ n_8838;
assign n_8851 = n_8838 ^ x488;
assign n_8852 = n_8839 ^ n_6761;
assign n_8853 = n_8840 ^ n_8161;
assign n_8854 = n_8840 ^ n_7682;
assign n_8855 = n_8841 ^ n_7504;
assign n_8856 = n_8842 & ~n_8782;
assign n_8857 = n_8782 ^ n_8842;
assign n_8858 = n_8843 ^ x37;
assign n_8859 = n_8844 ^ n_8833;
assign n_8860 = ~n_8845 & ~n_8846;
assign n_8861 = n_8847 ^ n_8835;
assign n_8862 = n_7794 & ~n_8848;
assign n_8863 = n_8848 & n_8849;
assign n_8864 = n_8850 ^ x488;
assign n_8865 = n_8850 & ~n_8851;
assign n_8866 = n_8852 ^ n_6803;
assign n_8867 = ~n_8169 & ~n_8853;
assign n_8868 = n_8854 ^ n_7526;
assign n_8869 = n_8854 ^ n_8161;
assign n_8870 = n_8855 ^ n_6803;
assign n_8871 = n_8855 ^ n_8852;
assign n_8872 = n_8858 ^ n_8859;
assign n_8873 = n_8859 ^ x36;
assign n_8874 = n_8860 ^ n_7223;
assign n_8875 = n_8862 ^ n_8322;
assign n_8876 = n_8863 ^ n_8322;
assign n_8877 = n_8864 ^ n_8836;
assign n_8878 = n_8836 & ~n_8864;
assign n_8879 = n_8865 ^ x488;
assign n_8880 = n_8867 ^ n_7682;
assign n_8881 = ~n_8155 & ~n_8868;
assign n_8882 = n_8870 ^ n_8852;
assign n_8883 = n_8866 & n_8871;
assign n_8884 = n_8872 ^ x36;
assign n_8885 = ~n_8872 & n_8873;
assign n_8886 = n_8874 ^ n_7261;
assign n_8887 = n_8875 ^ n_7261;
assign n_8888 = n_8874 ^ n_8875;
assign n_8889 = n_8876 ^ n_8361;
assign n_8890 = n_8877 ^ n_8876;
assign n_8891 = n_8877 ^ n_8361;
assign n_8892 = n_8879 ^ x503;
assign n_8893 = n_8880 ^ n_8186;
assign n_8894 = n_8881 ^ n_7526;
assign n_8895 = n_8882 ^ n_8879;
assign n_8896 = n_8883 ^ n_6803;
assign n_8897 = n_8856 & n_8884;
assign n_8898 = n_8884 ^ n_8856;
assign n_8899 = n_8885 ^ x36;
assign n_8900 = n_8886 ^ n_8875;
assign n_8901 = ~n_8887 & ~n_8888;
assign n_8902 = n_8889 ^ n_8877;
assign n_8903 = ~n_7833 & ~n_8890;
assign n_8904 = n_8890 & ~n_8891;
assign n_8905 = n_8882 ^ n_8892;
assign n_8906 = n_8893 & ~n_8195;
assign n_8907 = n_8893 ^ n_7717;
assign n_8908 = n_8894 ^ n_6845;
assign n_8909 = n_8892 & n_8895;
assign n_8910 = n_8896 ^ n_8894;
assign n_8911 = n_8899 ^ n_8900;
assign n_8912 = n_8900 ^ x35;
assign n_8913 = n_8901 ^ n_7261;
assign n_8914 = n_8749 ^ n_8902;
assign n_8915 = n_8903 ^ n_8361;
assign n_8916 = n_8904 ^ n_8361;
assign n_8917 = ~n_8905 & n_8878;
assign n_8918 = n_8878 ^ n_8905;
assign n_8919 = n_8906 ^ n_7717;
assign n_8920 = n_8907 & ~n_8196;
assign n_8921 = n_8909 ^ x503;
assign n_8922 = n_8910 ^ n_6845;
assign n_8923 = n_8910 & n_8908;
assign n_8924 = n_8911 ^ x35;
assign n_8925 = n_8911 & ~n_8912;
assign n_8926 = n_8913 ^ n_7287;
assign n_8927 = n_8915 ^ n_7287;
assign n_8928 = n_8913 ^ n_8915;
assign n_8929 = n_8916 ^ n_8403;
assign n_8930 = n_8918 ^ n_8916;
assign n_8931 = n_8918 ^ n_8403;
assign n_8932 = n_8919 ^ n_8216;
assign n_8933 = n_8920 ^ n_7545;
assign n_8934 = n_8921 ^ n_8922;
assign n_8935 = n_8922 ^ x502;
assign n_8936 = n_8923 ^ n_6845;
assign n_8937 = n_8897 & ~n_8924;
assign n_8938 = n_8924 ^ n_8897;
assign n_8939 = n_8925 ^ x35;
assign n_8940 = n_8926 ^ n_8915;
assign n_8941 = n_8927 & n_8928;
assign n_8942 = n_8929 ^ n_8918;
assign n_8943 = ~n_7874 & ~n_8930;
assign n_8944 = n_8930 & ~n_8931;
assign n_8945 = n_8932 & n_8227;
assign n_8946 = n_7789 ^ n_8932;
assign n_8947 = n_8934 ^ x502;
assign n_8948 = ~n_8934 & n_8935;
assign n_8949 = n_8936 ^ n_6887;
assign n_8950 = n_8933 ^ n_8936;
assign n_8951 = n_8939 ^ n_8940;
assign n_8952 = n_8940 ^ x34;
assign n_8953 = n_8941 ^ n_7287;
assign n_8954 = n_8942 ^ n_8782;
assign n_8955 = n_8943 ^ n_8403;
assign n_8956 = n_8944 ^ n_8403;
assign n_8957 = n_8945 ^ n_7789;
assign n_8958 = ~n_8946 & n_8228;
assign n_8959 = n_8917 & n_8947;
assign n_8960 = n_8947 ^ n_8917;
assign n_8961 = n_8948 ^ x502;
assign n_8962 = n_8933 ^ n_8949;
assign n_8963 = n_8949 & ~n_8950;
assign n_8964 = n_8951 ^ x34;
assign n_8965 = n_8951 & ~n_8952;
assign n_8966 = n_8953 ^ n_7303;
assign n_8967 = n_8955 ^ n_7303;
assign n_8968 = n_8953 ^ n_8955;
assign n_8969 = n_8956 ^ n_8446;
assign n_8970 = n_8957 ^ n_8250;
assign n_8971 = n_8957 ^ n_7844;
assign n_8972 = n_8958 ^ n_7566;
assign n_8973 = n_8956 ^ n_8960;
assign n_8974 = n_8961 ^ n_8962;
assign n_8975 = n_8962 ^ x501;
assign n_8976 = n_8963 ^ n_6887;
assign n_8977 = ~n_8937 & n_8964;
assign n_8978 = n_8964 ^ n_8937;
assign n_8979 = n_8965 ^ x34;
assign n_8980 = n_8966 ^ n_8955;
assign n_8981 = n_8967 & ~n_8968;
assign n_8982 = n_8264 & ~n_8970;
assign n_8983 = n_8971 ^ n_8250;
assign n_8984 = n_8972 ^ n_6926;
assign n_8985 = ~n_8973 & ~n_8969;
assign n_8986 = ~n_7915 & n_8973;
assign n_8987 = n_8973 ^ n_8446;
assign n_8988 = n_8974 ^ x501;
assign n_8989 = n_8974 & ~n_8975;
assign n_8990 = n_8976 ^ n_6926;
assign n_8991 = n_8976 ^ n_8972;
assign n_8992 = n_8979 ^ x33;
assign n_8993 = n_8980 ^ x33;
assign n_8994 = n_8979 ^ n_8980;
assign n_8995 = n_8981 ^ n_7303;
assign n_8996 = n_8982 ^ n_7844;
assign n_8997 = n_8983 & ~n_8265;
assign n_8998 = n_8985 ^ n_8446;
assign n_8999 = n_8986 ^ n_8446;
assign n_9000 = n_8857 ^ n_8987;
assign n_9001 = ~n_8959 & n_8988;
assign n_9002 = n_8988 ^ n_8959;
assign n_9003 = n_8989 ^ x501;
assign n_9004 = n_8990 ^ n_8972;
assign n_9005 = n_8984 & n_8991;
assign n_9006 = n_8992 ^ n_8980;
assign n_9007 = n_8993 & ~n_8994;
assign n_9008 = n_8995 ^ n_7328;
assign n_9009 = n_8996 ^ n_8288;
assign n_9010 = n_8997 ^ n_7586;
assign n_9011 = n_8998 ^ n_8486;
assign n_9012 = n_8999 ^ n_7328;
assign n_9013 = n_8995 ^ n_8999;
assign n_9014 = n_9002 ^ n_8998;
assign n_9015 = n_9002 ^ n_8486;
assign n_9016 = n_9003 ^ n_9004;
assign n_9017 = n_9004 ^ x500;
assign n_9018 = n_9005 ^ n_6926;
assign n_9019 = n_8977 & ~n_9006;
assign n_9020 = n_9006 ^ n_8977;
assign n_9021 = n_9007 ^ x33;
assign n_9022 = n_9008 ^ n_8999;
assign n_9023 = n_9009 & ~n_8301;
assign n_9024 = n_7885 ^ n_9009;
assign n_9025 = n_9010 ^ n_6957;
assign n_9026 = n_9011 ^ n_9002;
assign n_9027 = ~n_9012 & n_9013;
assign n_9028 = n_7958 & ~n_9014;
assign n_9029 = n_9014 & ~n_9015;
assign n_9030 = n_9016 ^ x500;
assign n_9031 = n_9016 & ~n_9017;
assign n_9032 = n_9018 ^ n_6957;
assign n_9033 = n_9018 ^ n_9010;
assign n_9034 = n_9021 ^ n_9022;
assign n_9035 = n_9022 ^ x32;
assign n_9036 = n_9023 ^ n_7885;
assign n_9037 = ~n_9024 & ~n_8302;
assign n_9038 = n_8898 ^ n_9026;
assign n_9039 = n_9027 ^ n_7328;
assign n_9040 = n_9028 ^ n_8486;
assign n_9041 = n_9029 ^ n_8486;
assign n_9042 = ~n_9001 & ~n_9030;
assign n_9043 = n_9030 ^ n_9001;
assign n_9044 = n_9031 ^ x500;
assign n_9045 = n_9032 ^ n_9010;
assign n_9046 = ~n_9025 & n_9033;
assign n_9047 = n_9034 ^ x32;
assign n_9048 = n_9034 & ~n_9035;
assign n_9049 = n_9036 ^ n_7926;
assign n_9050 = n_9036 ^ n_8329;
assign n_9051 = n_9037 ^ n_7607;
assign n_9052 = n_9039 ^ n_7346;
assign n_9053 = n_9040 ^ n_9039;
assign n_9054 = n_9041 ^ n_8528;
assign n_9055 = n_9043 ^ n_9041;
assign n_9056 = n_9043 ^ n_8528;
assign n_9057 = n_9044 ^ n_9045;
assign n_9058 = n_9045 ^ x499;
assign n_9059 = n_9046 ^ n_6957;
assign n_9060 = ~n_9019 & ~n_9047;
assign n_9061 = n_9047 ^ n_9019;
assign n_9062 = n_9048 ^ x32;
assign n_9063 = n_9049 ^ n_8329;
assign n_9064 = n_8342 & ~n_9050;
assign n_9065 = n_9051 ^ n_6980;
assign n_9066 = n_9040 ^ n_9052;
assign n_9067 = ~n_9052 & n_9053;
assign n_9068 = n_9054 ^ n_9043;
assign n_9069 = n_7993 & ~n_9055;
assign n_9070 = n_9055 & n_9056;
assign n_9071 = n_9057 ^ x499;
assign n_9072 = n_9057 & ~n_9058;
assign n_9073 = n_9059 ^ n_6980;
assign n_9074 = n_9059 ^ n_9051;
assign n_9075 = n_9063 ^ n_8208;
assign n_9076 = n_9063 & n_8341;
assign n_9077 = n_9064 ^ n_7926;
assign n_9078 = n_9062 ^ n_9066;
assign n_9079 = n_9066 ^ x47;
assign n_9080 = n_9067 ^ n_7346;
assign n_9081 = n_8938 ^ n_9068;
assign n_9082 = n_9069 ^ n_8528;
assign n_9083 = n_9070 ^ n_8528;
assign n_9084 = ~n_9042 & n_9071;
assign n_9085 = n_9071 ^ n_9042;
assign n_9086 = n_9072 ^ x499;
assign n_9087 = n_9073 ^ n_9051;
assign n_9088 = n_9065 & ~n_9074;
assign n_9089 = n_9076 ^ n_7628;
assign n_9090 = n_9077 ^ n_8368;
assign n_9091 = n_9078 ^ x47;
assign n_9092 = ~n_9078 & n_9079;
assign n_9093 = n_9080 ^ n_7364;
assign n_9094 = n_9082 ^ n_7364;
assign n_9095 = n_9080 ^ n_9082;
assign n_9096 = n_9083 ^ n_8569;
assign n_9097 = n_9085 ^ n_9083;
assign n_9098 = n_9085 ^ n_8569;
assign n_9099 = n_9086 ^ n_9087;
assign n_9100 = n_9087 ^ x498;
assign n_9101 = n_9088 ^ n_6980;
assign n_9102 = n_9089 ^ n_7000;
assign n_9103 = n_7966 ^ n_9090;
assign n_9104 = ~n_9090 & n_8384;
assign n_9105 = ~n_9060 & ~n_9091;
assign n_9106 = n_9091 ^ n_9060;
assign n_9107 = n_9092 ^ x47;
assign n_9108 = n_9093 ^ n_9082;
assign n_9109 = ~n_9094 & n_9095;
assign n_9110 = n_9096 ^ n_9085;
assign n_9111 = n_8022 & n_9097;
assign n_9112 = ~n_9097 & ~n_9098;
assign n_9113 = n_9099 ^ x498;
assign n_9114 = ~n_9099 & n_9100;
assign n_9115 = n_9101 ^ n_7000;
assign n_9116 = n_9101 ^ n_9089;
assign n_9117 = n_9103 & n_8383;
assign n_9118 = n_8254 ^ n_9103;
assign n_9119 = n_9104 ^ n_7966;
assign n_9120 = n_9107 ^ n_9108;
assign n_9121 = n_9108 ^ x46;
assign n_9122 = n_9109 ^ n_7364;
assign n_9123 = n_8978 ^ n_9110;
assign n_9124 = n_9111 ^ n_8569;
assign n_9125 = n_9112 ^ n_8569;
assign n_9126 = ~n_9113 & n_9084;
assign n_9127 = n_9084 ^ n_9113;
assign n_9128 = n_9114 ^ x498;
assign n_9129 = n_9115 ^ n_9089;
assign n_9130 = ~n_9102 & ~n_9116;
assign n_9131 = n_9117 ^ n_7651;
assign n_9132 = n_9119 ^ n_8425;
assign n_9133 = n_9119 ^ n_8410;
assign n_9134 = n_9120 ^ x46;
assign n_9135 = ~n_9120 & n_9121;
assign n_9136 = n_9122 ^ n_7382;
assign n_9137 = n_9124 ^ n_7382;
assign n_9138 = n_9122 ^ n_9124;
assign n_9139 = n_9125 ^ n_8612;
assign n_9140 = n_9127 ^ n_9125;
assign n_9141 = n_9127 ^ n_8612;
assign n_9142 = n_9128 ^ n_9129;
assign n_9143 = n_9129 ^ x497;
assign n_9144 = n_9130 ^ n_7000;
assign n_9145 = n_9131 ^ n_7021;
assign n_9146 = n_9132 & ~n_8426;
assign n_9147 = n_8317 ^ n_9132;
assign n_9148 = n_8425 & ~n_9133;
assign n_9149 = ~n_9105 & n_9134;
assign n_9150 = n_9134 ^ n_9105;
assign n_9151 = n_9135 ^ x46;
assign n_9152 = n_9136 ^ n_9124;
assign n_9153 = ~n_9137 & ~n_9138;
assign n_9154 = n_9139 ^ n_9127;
assign n_9155 = n_8044 & ~n_9140;
assign n_9156 = n_9140 & ~n_9141;
assign n_9157 = n_9142 ^ x497;
assign n_9158 = n_9142 & ~n_9143;
assign n_9159 = n_9144 ^ n_7021;
assign n_9160 = n_9144 ^ n_9131;
assign n_9161 = n_9146 ^ n_7679;
assign n_9162 = n_9148 ^ n_7999;
assign n_9163 = n_9151 ^ n_9152;
assign n_9164 = n_9152 ^ x45;
assign n_9165 = n_9153 ^ n_7382;
assign n_9166 = n_9020 ^ n_9154;
assign n_9167 = n_9155 ^ n_8612;
assign n_9168 = n_9156 ^ n_8612;
assign n_9169 = ~n_9157 & ~n_9126;
assign n_9170 = n_9126 ^ n_9157;
assign n_9171 = n_9158 ^ x497;
assign n_9172 = n_9159 ^ n_9131;
assign n_9173 = n_9145 & n_9160;
assign n_9174 = n_9161 ^ n_7036;
assign n_9175 = n_9162 ^ n_8026;
assign n_9176 = n_9162 ^ n_8452;
assign n_9177 = n_9163 ^ x45;
assign n_9178 = ~n_9163 & n_9164;
assign n_9179 = n_9165 ^ n_7403;
assign n_9180 = n_9167 ^ n_7403;
assign n_9181 = n_9165 ^ n_9167;
assign n_9182 = n_9168 ^ n_8652;
assign n_9183 = n_9170 ^ n_9168;
assign n_9184 = n_9170 ^ n_8652;
assign n_9185 = n_9171 ^ n_9172;
assign n_9186 = n_9172 ^ x496;
assign n_9187 = n_9173 ^ n_7021;
assign n_9188 = n_9175 ^ n_7714;
assign n_9189 = n_9175 ^ n_8452;
assign n_9190 = ~n_8467 & n_9176;
assign n_9191 = ~n_9177 & ~n_9149;
assign n_9192 = n_9149 ^ n_9177;
assign n_9193 = n_9178 ^ x45;
assign n_9194 = n_9179 ^ n_9167;
assign n_9195 = ~n_9180 & n_9181;
assign n_9196 = n_9182 ^ n_9170;
assign n_9197 = ~n_8057 & ~n_9183;
assign n_9198 = n_9183 & ~n_9184;
assign n_9199 = n_9185 ^ x496;
assign n_9200 = n_9185 & ~n_9186;
assign n_9201 = n_9187 ^ n_9161;
assign n_9202 = ~n_8439 & ~n_9188;
assign n_9203 = n_8371 ^ n_9189;
assign n_9204 = n_9190 ^ n_8026;
assign n_9205 = n_9193 ^ n_9194;
assign n_9206 = n_9194 ^ x44;
assign n_9207 = n_9195 ^ n_7403;
assign n_9208 = n_9061 ^ n_9196;
assign n_9209 = n_9197 ^ n_8652;
assign n_9210 = n_9198 ^ n_8652;
assign n_9211 = n_9199 & ~n_9169;
assign n_9212 = n_9169 ^ n_9199;
assign n_9213 = n_9200 ^ x496;
assign n_9214 = n_9201 ^ n_7036;
assign n_9215 = n_9201 & n_9174;
assign n_9216 = n_9202 ^ n_7714;
assign n_9217 = n_9204 ^ n_8493;
assign n_9218 = n_9205 ^ x44;
assign n_9219 = n_9205 & ~n_9206;
assign n_9220 = n_9207 ^ n_7422;
assign n_9221 = n_9209 ^ n_9207;
assign n_9222 = n_9210 ^ n_8698;
assign n_9223 = n_9212 ^ n_9210;
assign n_9224 = n_9212 ^ n_8698;
assign n_9225 = n_9213 ^ n_9214;
assign n_9226 = n_9214 ^ x511;
assign n_9227 = n_9215 ^ n_7036;
assign n_9228 = n_9216 ^ n_7061;
assign n_9229 = n_8047 ^ n_9217;
assign n_9230 = ~n_9217 & ~n_8509;
assign n_9231 = ~n_9191 & ~n_9218;
assign n_9232 = n_9218 ^ n_9191;
assign n_9233 = n_9219 ^ x44;
assign n_9234 = n_9209 ^ n_9220;
assign n_9235 = n_9220 & n_9221;
assign n_9236 = n_9222 ^ n_9212;
assign n_9237 = n_8081 & ~n_9223;
assign n_9238 = n_9223 & ~n_9224;
assign n_9239 = n_9225 ^ x511;
assign n_9240 = ~n_9225 & n_9226;
assign n_9241 = n_9227 ^ n_9216;
assign n_9242 = ~n_9229 & ~n_8508;
assign n_9243 = n_8413 ^ n_9229;
assign n_9244 = n_9230 ^ n_8047;
assign n_9245 = n_9233 ^ n_9234;
assign n_9246 = n_9234 ^ x43;
assign n_9247 = n_9235 ^ n_7422;
assign n_9248 = n_9106 ^ n_9236;
assign n_9249 = n_9237 ^ n_8698;
assign n_9250 = n_9238 ^ n_8698;
assign n_9251 = ~n_9239 & n_9211;
assign n_9252 = n_9211 ^ n_9239;
assign n_9253 = n_9240 ^ x511;
assign n_9254 = n_9241 ^ n_7061;
assign n_9255 = n_9241 & n_9228;
assign n_9256 = n_9242 ^ n_7748;
assign n_9257 = n_9244 ^ n_8535;
assign n_9258 = n_9245 ^ x43;
assign n_9259 = n_9245 & ~n_9246;
assign n_9260 = n_9247 ^ n_7442;
assign n_9261 = n_9249 ^ n_7442;
assign n_9262 = n_9247 ^ n_9249;
assign n_9263 = n_9250 ^ n_8744;
assign n_9264 = n_9250 ^ n_9252;
assign n_9265 = n_9252 ^ n_8744;
assign n_9266 = n_9253 ^ n_9254;
assign n_9267 = n_9254 ^ x510;
assign n_9268 = n_9255 ^ n_7061;
assign n_9269 = n_9256 ^ n_7081;
assign n_9270 = n_8067 ^ n_9257;
assign n_9271 = ~n_9257 & ~n_8551;
assign n_9272 = ~n_9258 & n_9231;
assign n_9273 = n_9231 ^ n_9258;
assign n_9274 = n_9259 ^ x43;
assign n_9275 = n_9260 ^ n_9249;
assign n_9276 = ~n_9261 & n_9262;
assign n_9277 = n_9263 ^ n_9252;
assign n_9278 = n_8101 & ~n_9264;
assign n_9279 = n_9264 & n_9265;
assign n_9280 = n_9266 ^ x510;
assign n_9281 = n_9266 & ~n_9267;
assign n_9282 = n_9268 ^ n_9256;
assign n_9283 = n_9270 & ~n_8550;
assign n_9284 = n_8455 ^ n_9270;
assign n_9285 = n_9271 ^ n_8067;
assign n_9286 = n_9274 ^ n_9275;
assign n_9287 = n_9275 ^ x42;
assign n_9288 = n_9276 ^ n_7442;
assign n_9289 = n_9150 ^ n_9277;
assign n_9290 = n_9278 ^ n_8744;
assign n_9291 = n_9279 ^ n_8744;
assign n_9292 = ~n_9280 & ~n_9251;
assign n_9293 = n_9251 ^ n_9280;
assign n_9294 = n_9281 ^ x510;
assign n_9295 = n_9282 ^ n_7081;
assign n_9296 = n_9282 & ~n_9269;
assign n_9297 = n_9283 ^ n_7786;
assign n_9298 = n_9285 ^ n_8576;
assign n_9299 = n_9286 ^ x42;
assign n_9300 = n_9286 & ~n_9287;
assign n_9301 = n_9288 ^ n_7463;
assign n_9302 = n_9290 ^ n_9288;
assign n_9303 = n_9291 ^ n_8790;
assign n_9304 = n_9291 ^ n_9293;
assign n_9305 = n_9293 ^ n_8790;
assign n_9306 = n_9294 ^ n_9295;
assign n_9307 = n_9295 ^ x509;
assign n_9308 = n_9296 ^ n_7081;
assign n_9309 = n_9297 ^ n_7102;
assign n_9310 = n_8084 ^ n_9298;
assign n_9311 = n_9298 & ~n_8592;
assign n_9312 = ~n_9272 & n_9299;
assign n_9313 = n_9299 ^ n_9272;
assign n_9314 = n_9300 ^ x42;
assign n_9315 = n_9290 ^ n_9301;
assign n_9316 = ~n_9301 & ~n_9302;
assign n_9317 = n_9303 ^ n_9293;
assign n_9318 = ~n_8122 & n_9304;
assign n_9319 = ~n_9304 & ~n_9305;
assign n_9320 = n_9306 ^ x509;
assign n_9321 = n_9306 & ~n_9307;
assign n_9322 = n_9308 ^ n_7102;
assign n_9323 = n_9308 ^ n_9297;
assign n_9324 = ~n_9310 & n_8591;
assign n_9325 = n_8496 ^ n_9310;
assign n_9326 = n_9311 ^ n_8084;
assign n_9327 = n_9314 ^ n_9315;
assign n_9328 = n_9315 ^ x41;
assign n_9329 = n_9316 ^ n_7463;
assign n_9330 = n_9192 ^ n_9317;
assign n_9331 = n_9318 ^ n_8790;
assign n_9332 = n_9319 ^ n_8790;
assign n_9333 = n_9292 & ~n_9320;
assign n_9334 = n_9320 ^ n_9292;
assign n_9335 = n_9321 ^ x509;
assign n_9336 = n_9322 ^ n_9297;
assign n_9337 = n_9309 & ~n_9323;
assign n_9338 = n_9324 ^ n_7826;
assign n_9339 = n_9326 ^ n_8619;
assign n_9340 = n_9327 ^ x41;
assign n_9341 = n_9327 & ~n_9328;
assign n_9342 = n_9329 ^ n_9331;
assign n_9343 = n_9331 ^ n_7484;
assign n_9344 = n_9332 ^ n_9334;
assign n_9345 = n_9334 ^ n_8829;
assign n_9346 = n_9335 ^ n_9336;
assign n_9347 = n_9336 ^ x508;
assign n_9348 = n_9337 ^ n_7102;
assign n_9349 = n_9338 ^ n_7127;
assign n_9350 = n_8104 ^ n_9339;
assign n_9351 = ~n_9339 & ~n_8634;
assign n_9352 = ~n_9312 & ~n_9340;
assign n_9353 = n_9340 ^ n_9312;
assign n_9354 = n_9341 ^ x41;
assign n_9355 = n_9342 ^ n_7484;
assign n_9356 = ~n_9342 & ~n_9343;
assign n_9357 = n_8141 & n_9344;
assign n_9358 = ~n_9344 & ~n_9345;
assign n_9359 = n_9345 ^ n_9332;
assign n_9360 = n_9346 ^ x508;
assign n_9361 = ~n_9346 & n_9347;
assign n_9362 = n_9348 ^ n_7127;
assign n_9363 = n_9348 ^ n_9338;
assign n_9364 = n_8605 & ~n_9350;
assign n_9365 = n_8538 ^ n_9350;
assign n_9366 = n_9351 ^ n_8104;
assign n_9367 = n_9354 ^ n_9355;
assign n_9368 = n_9355 ^ x40;
assign n_9369 = n_9356 ^ n_7484;
assign n_9370 = n_9357 ^ n_8829;
assign n_9371 = n_9358 ^ n_8829;
assign n_9372 = n_9232 ^ n_9359;
assign n_9373 = ~n_9333 & ~n_9360;
assign n_9374 = n_9360 ^ n_9333;
assign n_9375 = n_9361 ^ x508;
assign n_9376 = n_9362 ^ n_9338;
assign n_9377 = n_9349 & n_9363;
assign n_9378 = n_9364 ^ n_7867;
assign n_9379 = n_9366 ^ n_8659;
assign n_9380 = n_9367 ^ x40;
assign n_9381 = ~n_9367 & n_9368;
assign n_9382 = n_9369 ^ n_7504;
assign n_9383 = n_9370 ^ n_9369;
assign n_9384 = n_9370 ^ n_7504;
assign n_9385 = n_9371 ^ n_9374;
assign n_9386 = n_8869 ^ n_9374;
assign n_9387 = n_9375 ^ n_9376;
assign n_9388 = n_9376 ^ x507;
assign n_9389 = n_9377 ^ n_7127;
assign n_9390 = n_9378 ^ n_7158;
assign n_9391 = n_8125 ^ n_9379;
assign n_9392 = ~n_9379 & n_8675;
assign n_9393 = n_9352 & n_9380;
assign n_9394 = n_9380 ^ n_9352;
assign n_9395 = n_9381 ^ x40;
assign n_9396 = ~n_9382 & ~n_9383;
assign n_9397 = n_9384 ^ n_9369;
assign n_9398 = n_8869 ^ n_9385;
assign n_9399 = n_9385 & n_9386;
assign n_9400 = n_9387 ^ x507;
assign n_9401 = ~n_9387 & n_9388;
assign n_9402 = n_9389 ^ n_7158;
assign n_9403 = n_9389 ^ n_9378;
assign n_9404 = ~n_9391 & ~n_8674;
assign n_9405 = n_8579 ^ n_9391;
assign n_9406 = n_9392 ^ n_8125;
assign n_9407 = n_9395 ^ x55;
assign n_9408 = n_9396 ^ n_7504;
assign n_9409 = n_9397 ^ n_9395;
assign n_9410 = n_9398 ^ n_8854;
assign n_9411 = n_9398 ^ n_9273;
assign n_9412 = n_9399 ^ n_8869;
assign n_9413 = n_9400 & ~n_9373;
assign n_9414 = n_9373 ^ n_9400;
assign n_9415 = n_9401 ^ x507;
assign n_9416 = n_9402 ^ n_9378;
assign n_9417 = ~n_9390 & n_9403;
assign n_9418 = n_9404 ^ n_7909;
assign n_9419 = n_9406 ^ n_8690;
assign n_9420 = n_9397 ^ n_9407;
assign n_9421 = n_9407 & n_9409;
assign n_9422 = n_8161 & ~n_9410;
assign n_9423 = n_9412 ^ n_9414;
assign n_9424 = n_9414 ^ n_8907;
assign n_9425 = n_9415 ^ n_9416;
assign n_9426 = n_9416 ^ x506;
assign n_9427 = n_9417 ^ n_7158;
assign n_9428 = n_9418 ^ n_7192;
assign n_9429 = n_9419 ^ n_8144;
assign n_9430 = n_9393 & ~n_9420;
assign n_9431 = n_9420 ^ n_9393;
assign n_9432 = n_9421 ^ x55;
assign n_9433 = n_9422 ^ n_8854;
assign n_9434 = n_8186 & n_9423;
assign n_9435 = n_9423 ^ n_8907;
assign n_9436 = ~n_9423 & ~n_9424;
assign n_9437 = n_9425 ^ x506;
assign n_9438 = ~n_9425 & n_9426;
assign n_9439 = n_9427 ^ n_7192;
assign n_9440 = n_9427 ^ n_9418;
assign n_9441 = n_9429 & n_8706;
assign n_9442 = n_9408 ^ n_9433;
assign n_9443 = n_9433 ^ n_7526;
assign n_9444 = n_9434 ^ n_8907;
assign n_9445 = n_9313 ^ n_9435;
assign n_9446 = n_9436 ^ n_8907;
assign n_9447 = n_9413 & n_9437;
assign n_9448 = n_9437 ^ n_9413;
assign n_9449 = n_9438 ^ x506;
assign n_9450 = n_9439 ^ n_9418;
assign n_9451 = ~n_9428 & n_9440;
assign n_9452 = n_9441 ^ n_7938;
assign n_9453 = n_9442 ^ n_7526;
assign n_9454 = ~n_9442 & n_9443;
assign n_9455 = n_9444 ^ n_7545;
assign n_9456 = n_9446 ^ n_8946;
assign n_9457 = n_9448 ^ n_9446;
assign n_9458 = n_9448 ^ n_8946;
assign n_9459 = n_9449 ^ n_9450;
assign n_9460 = n_9450 ^ x505;
assign n_9461 = n_9451 ^ n_7192;
assign n_9462 = n_9452 ^ n_7219;
assign n_9463 = n_9432 ^ n_9453;
assign n_9464 = n_9453 ^ x54;
assign n_9465 = n_9454 ^ n_7526;
assign n_9466 = n_9456 ^ n_9448;
assign n_9467 = n_8216 & n_9457;
assign n_9468 = ~n_9457 & ~n_9458;
assign n_9469 = n_9459 ^ x505;
assign n_9470 = ~n_9459 & n_9460;
assign n_9471 = n_9461 ^ x504;
assign n_9472 = n_9463 ^ x54;
assign n_9473 = n_9463 & ~n_9464;
assign n_9474 = n_9465 ^ n_9444;
assign n_9475 = n_9465 ^ n_7545;
assign n_9476 = n_9353 ^ n_9466;
assign n_9477 = n_9467 ^ n_8946;
assign n_9478 = n_9468 ^ n_8946;
assign n_9479 = ~n_9469 & ~n_9447;
assign n_9480 = n_9447 ^ n_9469;
assign n_9481 = n_9470 ^ x505;
assign n_9482 = n_9471 ^ n_9462;
assign n_9483 = ~n_9430 & n_9472;
assign n_9484 = n_9472 ^ n_9430;
assign n_9485 = n_9473 ^ x54;
assign n_9486 = ~n_9455 & n_9474;
assign n_9487 = n_9475 ^ n_9444;
assign n_9488 = n_9477 ^ n_7566;
assign n_9489 = n_9478 ^ n_8983;
assign n_9490 = n_9480 ^ n_8983;
assign n_9491 = n_9478 ^ n_9480;
assign n_9492 = n_9481 ^ n_9479;
assign n_9493 = n_9486 ^ n_7545;
assign n_9494 = n_9485 ^ n_9487;
assign n_9495 = n_9487 ^ x53;
assign n_9496 = n_9489 ^ n_9480;
assign n_9497 = ~n_9490 & ~n_9491;
assign n_9498 = n_9492 ^ n_9482;
assign n_9499 = n_9493 ^ n_9477;
assign n_9500 = n_9493 ^ n_7566;
assign n_9501 = n_9494 ^ x53;
assign n_9502 = ~n_9494 & n_9495;
assign n_9503 = n_9496 ^ n_8971;
assign n_9504 = n_9394 ^ n_9496;
assign n_9505 = n_9497 ^ n_8983;
assign n_9506 = n_9498 ^ n_9024;
assign n_9507 = ~n_9488 & ~n_9499;
assign n_9508 = n_9500 ^ n_9477;
assign n_9509 = ~n_9501 & n_9483;
assign n_9510 = n_9483 ^ n_9501;
assign n_9511 = n_9502 ^ x53;
assign n_9512 = n_8250 & n_9503;
assign n_9513 = n_9498 ^ n_9505;
assign n_9514 = n_9505 ^ n_9024;
assign n_9515 = n_9507 ^ n_7566;
assign n_9516 = n_9508 ^ x52;
assign n_9517 = n_9511 ^ n_9508;
assign n_9518 = n_9512 ^ n_8971;
assign n_9519 = n_9513 & n_9506;
assign n_9520 = ~n_8288 & ~n_9513;
assign n_9521 = n_9514 ^ n_9498;
assign n_9522 = n_9515 ^ n_7586;
assign n_9523 = ~n_9517 & n_9516;
assign n_9524 = n_9517 ^ x52;
assign n_9525 = n_9518 ^ n_7586;
assign n_9526 = n_9515 ^ n_9518;
assign n_9527 = n_9519 ^ n_9024;
assign n_9528 = n_9520 ^ n_9024;
assign n_9529 = n_9431 ^ n_9521;
assign n_9530 = n_9522 ^ n_9518;
assign n_9531 = n_9523 ^ x52;
assign n_9532 = ~n_9524 & n_9509;
assign n_9533 = n_9509 ^ n_9524;
assign n_9534 = ~n_9525 & ~n_9526;
assign n_9535 = n_9527 ^ n_9063;
assign n_9536 = n_9527 ^ n_9075;
assign n_9537 = n_9528 ^ n_7607;
assign n_9538 = n_9530 ^ x51;
assign n_9539 = n_9531 ^ n_9530;
assign n_9540 = n_9534 ^ n_7586;
assign n_9541 = ~n_9075 & n_9535;
assign n_9542 = n_9536 ^ n_9049;
assign n_9543 = n_9484 ^ n_9536;
assign n_9544 = n_9539 & ~n_9538;
assign n_9545 = n_9539 ^ x51;
assign n_9546 = n_9540 ^ n_9528;
assign n_9547 = n_9540 ^ n_7607;
assign n_9548 = n_9541 ^ n_8208;
assign n_9549 = n_8329 & n_9542;
assign n_9550 = n_9544 ^ x51;
assign n_9551 = n_9532 & n_9545;
assign n_9552 = n_9545 ^ n_9532;
assign n_9553 = ~n_9537 & ~n_9546;
assign n_9554 = n_9547 ^ n_9528;
assign n_9555 = n_9548 ^ n_9103;
assign n_9556 = n_9549 ^ n_9049;
assign n_9557 = n_9553 ^ n_7607;
assign n_9558 = n_9550 ^ n_9554;
assign n_9559 = n_9554 ^ x50;
assign n_9560 = n_9555 & n_9118;
assign n_9561 = n_8254 ^ n_9555;
assign n_9562 = n_9557 ^ n_7628;
assign n_9563 = n_9556 ^ n_9557;
assign n_9564 = n_9558 ^ x50;
assign n_9565 = ~n_9558 & n_9559;
assign n_9566 = n_9560 ^ n_8254;
assign n_9567 = n_9561 ^ n_9103;
assign n_9568 = n_9510 ^ n_9561;
assign n_9569 = n_9556 ^ n_9562;
assign n_9570 = n_9562 & ~n_9563;
assign n_9571 = n_9564 & ~n_9551;
assign n_9572 = n_9551 ^ n_9564;
assign n_9573 = n_9565 ^ x50;
assign n_9574 = n_9566 ^ n_9132;
assign n_9575 = n_8368 & ~n_9567;
assign n_9576 = n_9569 ^ x49;
assign n_9577 = n_9570 ^ n_7628;
assign n_9578 = n_9573 ^ n_9569;
assign n_9579 = ~n_9574 & n_9147;
assign n_9580 = n_8317 ^ n_9574;
assign n_9581 = n_9575 ^ n_9103;
assign n_9582 = n_9577 ^ n_7651;
assign n_9583 = ~n_9578 & n_9576;
assign n_9584 = n_9578 ^ x49;
assign n_9585 = n_9579 ^ n_8317;
assign n_9586 = n_9580 ^ n_9132;
assign n_9587 = n_9533 ^ n_9580;
assign n_9588 = n_9581 ^ n_7651;
assign n_9589 = n_9577 ^ n_9581;
assign n_9590 = n_9582 ^ n_9581;
assign n_9591 = n_9583 ^ x49;
assign n_9592 = n_9571 & n_9584;
assign n_9593 = n_9584 ^ n_9571;
assign n_9594 = n_9585 ^ n_8371;
assign n_9595 = n_9585 ^ n_9189;
assign n_9596 = n_8410 & n_9586;
assign n_9597 = n_9588 & ~n_9589;
assign n_9598 = n_9590 ^ x48;
assign n_9599 = n_9591 ^ n_9590;
assign n_9600 = n_9594 ^ n_9189;
assign n_9601 = ~n_9203 & n_9595;
assign n_9602 = n_9596 ^ n_9132;
assign n_9603 = n_9597 ^ n_7651;
assign n_9604 = ~n_9599 & n_9598;
assign n_9605 = n_9599 ^ x48;
assign n_9606 = n_9600 ^ n_9175;
assign n_9607 = n_9552 ^ n_9600;
assign n_9608 = n_9601 ^ n_8371;
assign n_9609 = n_9602 ^ n_7679;
assign n_9610 = n_9603 ^ n_9602;
assign n_9611 = n_9604 ^ x48;
assign n_9612 = n_9592 & n_9605;
assign n_9613 = n_9605 ^ n_9592;
assign n_9614 = ~n_8452 & ~n_9606;
assign n_9615 = n_9608 ^ n_9229;
assign n_9616 = ~n_9610 & ~n_9609;
assign n_9617 = n_9610 ^ n_7679;
assign n_9618 = n_9611 ^ x63;
assign n_9619 = n_9614 ^ n_9175;
assign n_9620 = n_8413 ^ n_9615;
assign n_9621 = n_9615 & ~n_9243;
assign n_9622 = n_9616 ^ n_7679;
assign n_9623 = n_9617 ^ x63;
assign n_9624 = n_9611 ^ n_9617;
assign n_9625 = n_9618 ^ n_9617;
assign n_9626 = n_9619 ^ n_7714;
assign n_9627 = n_9620 ^ n_9229;
assign n_9628 = n_9572 ^ n_9620;
assign n_9629 = n_9621 ^ n_8413;
assign n_9630 = n_9622 ^ n_9619;
assign n_9631 = n_9622 ^ n_7714;
assign n_9632 = ~n_9623 & n_9624;
assign n_9633 = n_9612 & ~n_9625;
assign n_9634 = n_9625 ^ n_9612;
assign n_9635 = n_8493 & n_9627;
assign n_9636 = n_9629 ^ n_9270;
assign n_9637 = n_9626 & n_9630;
assign n_9638 = n_9631 ^ n_9619;
assign n_9639 = n_9632 ^ x63;
assign n_9640 = n_9635 ^ n_9229;
assign n_9641 = n_8455 ^ n_9636;
assign n_9642 = ~n_9636 & ~n_9284;
assign n_9643 = n_9637 ^ n_7714;
assign n_9644 = n_9638 ^ x62;
assign n_9645 = n_9639 ^ n_9638;
assign n_9646 = n_9640 ^ n_7748;
assign n_9647 = n_9641 ^ n_9270;
assign n_9648 = n_9593 ^ n_9641;
assign n_9649 = n_9642 ^ n_8455;
assign n_9650 = n_9643 ^ n_7748;
assign n_9651 = n_9643 ^ n_9640;
assign n_9652 = n_9645 & ~n_9644;
assign n_9653 = n_9645 ^ x62;
assign n_9654 = ~n_8535 & ~n_9647;
assign n_9655 = n_9649 ^ n_9310;
assign n_9656 = n_9650 ^ n_9640;
assign n_9657 = n_9646 & n_9651;
assign n_9658 = n_9652 ^ x62;
assign n_9659 = ~n_9633 & n_9653;
assign n_9660 = n_9653 ^ n_9633;
assign n_9661 = n_9654 ^ n_9270;
assign n_9662 = n_8496 ^ n_9655;
assign n_9663 = ~n_9655 & ~n_9325;
assign n_9664 = n_9656 ^ x61;
assign n_9665 = n_9657 ^ n_7748;
assign n_9666 = n_9658 ^ n_9656;
assign n_9667 = n_9658 ^ x61;
assign n_9668 = n_9661 ^ n_7786;
assign n_9669 = n_9662 ^ n_9310;
assign n_9670 = n_9613 ^ n_9662;
assign n_9671 = n_9663 ^ n_8496;
assign n_9672 = n_9665 ^ n_9661;
assign n_9673 = n_9664 & ~n_9666;
assign n_9674 = n_9667 ^ n_9656;
assign n_9675 = ~n_8576 & ~n_9669;
assign n_9676 = n_9671 ^ n_8538;
assign n_9677 = n_9671 ^ n_9350;
assign n_9678 = n_9672 ^ n_7786;
assign n_9679 = n_9672 & n_9668;
assign n_9680 = n_9673 ^ x61;
assign n_9681 = n_9659 & ~n_9674;
assign n_9682 = n_9674 ^ n_9659;
assign n_9683 = n_9675 ^ n_9310;
assign n_9684 = n_8619 & ~n_9676;
assign n_9685 = n_9676 ^ n_9350;
assign n_9686 = n_9365 & n_9677;
assign n_9687 = n_9678 ^ x60;
assign n_9688 = n_9679 ^ n_7786;
assign n_9689 = n_9680 ^ n_9678;
assign n_9690 = n_9683 ^ n_7826;
assign n_9691 = n_9684 ^ n_9350;
assign n_9692 = n_9634 ^ n_9685;
assign n_9693 = n_9686 ^ n_8538;
assign n_9694 = n_9688 ^ n_7826;
assign n_9695 = n_9688 ^ n_9683;
assign n_9696 = n_9689 & ~n_9687;
assign n_9697 = n_9689 ^ x60;
assign n_9698 = n_9691 ^ n_7867;
assign n_9699 = n_9693 ^ n_9391;
assign n_9700 = n_9694 ^ n_9683;
assign n_9701 = n_9690 & n_9695;
assign n_9702 = n_9696 ^ x60;
assign n_9703 = ~n_9681 & ~n_9697;
assign n_9704 = n_9697 ^ n_9681;
assign n_9705 = n_8579 ^ n_9699;
assign n_9706 = ~n_9699 & n_9405;
assign n_9707 = n_9700 ^ x59;
assign n_9708 = n_9701 ^ n_7826;
assign n_9709 = n_9702 ^ n_9700;
assign n_9710 = n_8677 & n_9704;
assign n_9711 = n_9704 ^ n_8677;
assign n_9712 = n_9705 ^ n_9391;
assign n_9713 = n_9660 ^ n_9705;
assign n_9714 = n_9706 ^ n_8579;
assign n_9715 = n_9708 ^ n_7867;
assign n_9716 = n_9708 ^ n_9691;
assign n_9717 = n_9709 ^ x59;
assign n_9718 = ~n_9709 & n_9707;
assign n_9719 = n_8723 ^ n_9710;
assign n_9720 = n_9711 ^ n_8661;
assign n_9721 = ~n_8659 & n_9712;
assign n_9722 = n_9714 ^ n_9429;
assign n_9723 = n_9715 ^ n_9691;
assign n_9724 = ~n_9698 & ~n_9716;
assign n_9725 = n_9717 ^ n_9703;
assign n_9726 = ~n_9703 & ~n_9717;
assign n_9727 = n_9718 ^ x59;
assign n_9728 = n_8171 & n_9720;
assign n_9729 = n_9721 ^ n_9391;
assign n_9730 = n_9722 ^ n_8622;
assign n_9731 = n_9723 ^ x58;
assign n_9732 = n_9724 ^ n_7867;
assign n_9733 = n_9725 ^ n_9710;
assign n_9734 = n_9719 ^ n_9725;
assign n_9735 = n_9727 ^ n_9723;
assign n_9736 = n_9728 ^ n_8661;
assign n_9737 = n_9729 ^ n_7909;
assign n_9738 = n_9730 ^ n_9429;
assign n_9739 = n_9732 ^ n_7909;
assign n_9740 = n_9732 ^ n_9729;
assign n_9741 = n_9733 & ~n_9719;
assign n_9742 = ~n_8200 & ~n_9733;
assign n_9743 = n_9735 ^ x58;
assign n_9744 = ~n_9735 & n_9731;
assign n_9745 = n_7645 & n_9736;
assign n_9746 = n_9736 ^ n_7645;
assign n_9747 = ~n_8690 & ~n_9738;
assign n_9748 = n_9739 ^ n_9729;
assign n_9749 = ~n_9737 & n_9740;
assign n_9750 = n_9741 ^ n_8723;
assign n_9751 = n_9742 ^ n_8723;
assign n_9752 = n_9726 ^ n_9743;
assign n_9753 = ~n_9743 & n_9726;
assign n_9754 = n_9744 ^ x58;
assign n_9755 = n_9745 ^ n_7673;
assign n_9756 = x199 & n_9746;
assign n_9757 = n_9746 ^ x199;
assign n_9758 = n_9747 ^ n_9429;
assign n_9759 = n_9748 ^ x57;
assign n_9760 = n_9749 ^ n_7909;
assign n_9761 = n_8779 ^ n_9750;
assign n_9762 = n_9751 ^ n_9745;
assign n_9763 = n_9750 ^ n_9752;
assign n_9764 = n_8779 ^ n_9752;
assign n_9765 = n_9754 ^ n_9748;
assign n_9766 = n_9751 ^ n_9755;
assign n_9767 = n_9756 ^ x198;
assign n_9768 = n_9758 ^ n_7938;
assign n_9769 = n_9760 ^ x56;
assign n_9770 = n_9761 ^ n_9752;
assign n_9771 = n_9755 & n_9762;
assign n_9772 = ~n_8243 & ~n_9763;
assign n_9773 = n_9763 & n_9764;
assign n_9774 = n_9765 ^ x57;
assign n_9775 = n_9765 & ~n_9759;
assign n_9776 = n_9766 ^ n_9756;
assign n_9777 = n_9766 ^ n_9767;
assign n_9778 = n_9769 ^ n_9768;
assign n_9779 = n_9771 ^ n_7673;
assign n_9780 = n_9772 ^ n_8779;
assign n_9781 = n_9773 ^ n_8779;
assign n_9782 = n_9753 ^ n_9774;
assign n_9783 = n_9774 & n_9753;
assign n_9784 = n_9775 ^ x57;
assign n_9785 = n_9767 & n_9776;
assign n_9786 = n_9779 ^ n_7719;
assign n_9787 = n_9780 ^ n_7719;
assign n_9788 = n_9779 ^ n_9780;
assign n_9789 = n_8820 ^ n_9781;
assign n_9790 = n_9781 ^ n_9782;
assign n_9791 = n_8820 ^ n_9782;
assign n_9792 = n_9784 ^ n_9783;
assign n_9793 = n_9785 ^ x198;
assign n_9794 = n_9786 ^ n_9780;
assign n_9795 = n_9787 & ~n_9788;
assign n_9796 = n_9789 ^ n_9782;
assign n_9797 = ~n_8281 & ~n_9790;
assign n_9798 = n_9790 & n_9791;
assign n_9799 = n_9792 ^ n_9778;
assign n_9800 = n_9793 ^ n_9794;
assign n_9801 = n_9794 ^ x197;
assign n_9802 = n_9795 ^ n_7719;
assign n_9803 = n_9797 ^ n_8820;
assign n_9804 = n_9798 ^ n_8820;
assign n_9805 = n_8861 ^ n_9799;
assign n_9806 = n_9800 ^ x197;
assign n_9807 = ~n_9800 & n_9801;
assign n_9808 = n_9802 ^ n_7753;
assign n_9809 = n_9803 ^ n_7753;
assign n_9810 = n_9802 ^ n_9803;
assign n_9811 = n_9804 ^ n_9799;
assign n_9812 = n_8861 ^ n_9804;
assign n_9813 = n_9807 ^ x197;
assign n_9814 = n_9808 ^ n_9803;
assign n_9815 = n_9809 & n_9810;
assign n_9816 = ~n_9811 & n_9805;
assign n_9817 = n_8322 & n_9811;
assign n_9818 = n_9812 ^ n_9799;
assign n_9819 = n_9813 ^ n_9814;
assign n_9820 = n_9814 ^ x196;
assign n_9821 = n_9815 ^ n_7753;
assign n_9822 = n_9816 ^ n_8861;
assign n_9823 = n_9817 ^ n_8861;
assign n_9824 = n_9819 ^ x196;
assign n_9825 = ~n_9819 & n_9820;
assign n_9826 = n_9821 ^ n_7794;
assign n_9827 = n_8902 ^ n_9822;
assign n_9828 = n_9823 ^ n_7794;
assign n_9829 = n_9821 ^ n_9823;
assign n_9830 = n_9825 ^ x196;
assign n_9831 = n_9826 ^ n_9823;
assign n_9832 = n_8749 ^ n_9827;
assign n_9833 = ~n_9827 & ~n_8914;
assign n_9834 = ~n_9828 & ~n_9829;
assign n_9835 = n_9830 ^ n_9831;
assign n_9836 = n_9831 ^ x195;
assign n_9837 = n_9832 ^ n_8902;
assign n_9838 = n_9833 ^ n_8749;
assign n_9839 = n_9834 ^ n_7794;
assign n_9840 = n_9835 ^ x195;
assign n_9841 = ~n_9835 & n_9836;
assign n_9842 = n_8361 & ~n_9837;
assign n_9843 = n_9838 ^ n_8782;
assign n_9844 = n_8942 ^ n_9838;
assign n_9845 = n_9839 ^ n_7833;
assign n_9846 = n_9841 ^ x195;
assign n_9847 = n_9842 ^ n_8902;
assign n_9848 = n_8403 & n_9843;
assign n_9849 = ~n_9843 & ~n_8954;
assign n_9850 = n_9844 ^ n_8782;
assign n_9851 = n_9847 ^ n_7833;
assign n_9852 = n_9839 ^ n_9847;
assign n_9853 = n_9845 ^ n_9847;
assign n_9854 = n_9848 ^ n_8942;
assign n_9855 = n_9849 ^ n_8942;
assign n_9856 = n_9851 & n_9852;
assign n_9857 = n_9846 ^ n_9853;
assign n_9858 = n_9853 ^ x194;
assign n_9859 = n_8987 ^ n_9855;
assign n_9860 = n_9856 ^ n_7833;
assign n_9861 = n_9857 ^ x194;
assign n_9862 = ~n_9857 & n_9858;
assign n_9863 = n_8857 ^ n_9859;
assign n_9864 = ~n_9859 & n_9000;
assign n_9865 = n_9860 ^ n_7874;
assign n_9866 = n_9854 ^ n_9860;
assign n_9867 = n_9862 ^ x194;
assign n_9868 = n_9863 ^ n_8973;
assign n_9869 = n_9864 ^ n_8857;
assign n_9870 = n_9854 ^ n_9865;
assign n_9871 = n_9865 & ~n_9866;
assign n_9872 = ~n_8446 & ~n_9868;
assign n_9873 = n_9026 ^ n_9869;
assign n_9874 = n_9867 ^ n_9870;
assign n_9875 = n_9870 ^ x193;
assign n_9876 = n_9871 ^ n_7874;
assign n_9877 = n_9872 ^ n_8973;
assign n_9878 = n_8898 ^ n_9873;
assign n_9879 = n_9873 & n_9038;
assign n_9880 = n_9874 ^ x193;
assign n_9881 = n_9874 & ~n_9875;
assign n_9882 = n_9876 ^ n_7915;
assign n_9883 = n_9877 ^ n_7915;
assign n_9884 = n_9876 ^ n_9877;
assign n_9885 = n_9878 ^ n_9026;
assign n_9886 = n_9879 ^ n_8898;
assign n_9887 = n_9881 ^ x193;
assign n_9888 = n_9882 ^ n_9877;
assign n_9889 = ~n_9883 & n_9884;
assign n_9890 = ~n_8486 & ~n_9885;
assign n_9891 = n_9886 ^ n_8938;
assign n_9892 = n_9886 ^ n_9068;
assign n_9893 = n_9888 ^ x192;
assign n_9894 = n_9887 ^ n_9888;
assign n_9895 = n_9889 ^ n_7915;
assign n_9896 = n_9890 ^ n_9026;
assign n_9897 = n_8528 & ~n_9891;
assign n_9898 = n_9891 ^ n_9068;
assign n_9899 = n_9081 & n_9892;
assign n_9900 = n_9887 ^ n_9893;
assign n_9901 = n_9893 & ~n_9894;
assign n_9902 = n_9895 ^ n_7958;
assign n_9903 = n_9896 ^ n_7958;
assign n_9904 = n_9895 ^ n_9896;
assign n_9905 = n_9897 ^ n_9068;
assign n_9906 = n_9757 ^ n_9898;
assign n_9907 = n_9899 ^ n_8938;
assign n_9908 = ~n_9880 & n_9900;
assign n_9909 = n_9900 ^ n_9880;
assign n_9910 = n_9901 ^ x192;
assign n_9911 = n_9902 ^ n_9896;
assign n_9912 = n_9903 & n_9904;
assign n_9913 = n_9905 ^ n_7993;
assign n_9914 = n_9110 ^ n_9907;
assign n_9915 = n_9910 ^ n_9911;
assign n_9916 = n_9911 ^ x207;
assign n_9917 = n_9912 ^ n_7958;
assign n_9918 = n_8978 ^ n_9914;
assign n_9919 = ~n_9914 & ~n_9123;
assign n_9920 = n_9915 ^ x207;
assign n_9921 = n_9915 & ~n_9916;
assign n_9922 = n_9917 ^ n_7993;
assign n_9923 = n_9917 ^ n_9905;
assign n_9924 = n_9918 ^ n_9110;
assign n_9925 = n_9777 ^ n_9918;
assign n_9926 = n_9919 ^ n_8978;
assign n_9927 = ~n_9908 & n_9920;
assign n_9928 = n_9920 ^ n_9908;
assign n_9929 = n_9921 ^ x207;
assign n_9930 = n_9922 ^ n_9905;
assign n_9931 = ~n_9913 & n_9923;
assign n_9932 = ~n_8569 & ~n_9924;
assign n_9933 = n_9154 ^ n_9926;
assign n_9934 = n_9929 ^ n_9930;
assign n_9935 = n_9930 ^ x206;
assign n_9936 = n_9931 ^ n_7993;
assign n_9937 = n_9932 ^ n_9110;
assign n_9938 = n_9020 ^ n_9933;
assign n_9939 = ~n_9933 & n_9166;
assign n_9940 = n_9934 ^ x206;
assign n_9941 = n_9934 & ~n_9935;
assign n_9942 = n_9936 ^ n_8022;
assign n_9943 = n_9937 ^ n_8022;
assign n_9944 = n_9936 ^ n_9937;
assign n_9945 = n_9938 ^ n_9154;
assign n_9946 = n_9806 ^ n_9938;
assign n_9947 = n_9939 ^ n_9020;
assign n_9948 = n_9927 & n_9940;
assign n_9949 = n_9940 ^ n_9927;
assign n_9950 = n_9941 ^ x206;
assign n_9951 = n_9942 ^ n_9937;
assign n_9952 = ~n_9943 & n_9944;
assign n_9953 = ~n_8612 & n_9945;
assign n_9954 = n_9196 ^ n_9947;
assign n_9955 = n_9950 ^ n_9951;
assign n_9956 = n_9951 ^ x205;
assign n_9957 = n_9952 ^ n_8022;
assign n_9958 = n_9953 ^ n_9154;
assign n_9959 = n_9061 ^ n_9954;
assign n_9960 = ~n_9954 & n_9208;
assign n_9961 = n_9955 ^ x205;
assign n_9962 = n_9955 & ~n_9956;
assign n_9963 = n_9957 ^ n_8044;
assign n_9964 = n_9958 ^ n_8044;
assign n_9965 = n_9957 ^ n_9958;
assign n_9966 = n_9959 ^ n_9196;
assign n_9967 = n_9824 ^ n_9959;
assign n_9968 = n_9960 ^ n_9061;
assign n_9969 = ~n_9948 & ~n_9961;
assign n_9970 = n_9961 ^ n_9948;
assign n_9971 = n_9962 ^ x205;
assign n_9972 = n_9963 ^ n_9958;
assign n_9973 = n_9964 & ~n_9965;
assign n_9974 = ~n_8652 & n_9966;
assign n_9975 = n_9236 ^ n_9968;
assign n_9976 = n_9971 ^ n_9972;
assign n_9977 = n_9972 ^ x204;
assign n_9978 = n_9973 ^ n_8044;
assign n_9979 = n_9974 ^ n_9196;
assign n_9980 = n_9106 ^ n_9975;
assign n_9981 = ~n_9975 & ~n_9248;
assign n_9982 = n_9976 ^ x204;
assign n_9983 = ~n_9976 & n_9977;
assign n_9984 = n_9978 ^ n_8057;
assign n_9985 = n_9979 ^ n_8057;
assign n_9986 = n_9978 ^ n_9979;
assign n_9987 = n_9980 ^ n_9236;
assign n_9988 = n_9840 ^ n_9980;
assign n_9989 = n_9981 ^ n_9106;
assign n_9990 = n_9969 & n_9982;
assign n_9991 = n_9982 ^ n_9969;
assign n_9992 = n_9983 ^ x204;
assign n_9993 = n_9984 ^ n_9979;
assign n_9994 = ~n_9985 & ~n_9986;
assign n_9995 = ~n_8698 & ~n_9987;
assign n_9996 = n_9277 ^ n_9989;
assign n_9997 = n_9992 ^ n_9993;
assign n_9998 = n_9993 ^ x203;
assign n_9999 = n_9994 ^ n_8057;
assign n_10000 = n_9995 ^ n_9236;
assign n_10001 = n_9150 ^ n_9996;
assign n_10002 = ~n_9996 & n_9289;
assign n_10003 = n_9997 ^ x203;
assign n_10004 = n_9997 & ~n_9998;
assign n_10005 = n_9999 ^ n_8081;
assign n_10006 = n_10000 ^ n_8081;
assign n_10007 = n_9999 ^ n_10000;
assign n_10008 = n_10001 ^ n_9277;
assign n_10009 = n_9861 ^ n_10001;
assign n_10010 = n_10002 ^ n_9150;
assign n_10011 = ~n_9990 & n_10003;
assign n_10012 = n_10003 ^ n_9990;
assign n_10013 = n_10004 ^ x203;
assign n_10014 = n_10005 ^ n_10000;
assign n_10015 = n_10006 & n_10007;
assign n_10016 = n_8744 & n_10008;
assign n_10017 = n_9317 ^ n_10010;
assign n_10018 = n_10013 ^ n_10014;
assign n_10019 = n_10014 ^ x202;
assign n_10020 = n_10015 ^ n_8081;
assign n_10021 = n_10016 ^ n_9277;
assign n_10022 = n_9192 ^ n_10017;
assign n_10023 = ~n_10017 & n_9330;
assign n_10024 = n_10018 ^ x202;
assign n_10025 = n_10018 & ~n_10019;
assign n_10026 = n_10020 ^ n_8101;
assign n_10027 = n_10021 ^ n_8101;
assign n_10028 = n_10020 ^ n_10021;
assign n_10029 = n_10022 ^ n_9317;
assign n_10030 = n_9880 ^ n_10022;
assign n_10031 = n_10023 ^ n_9192;
assign n_10032 = n_10024 & n_10011;
assign n_10033 = n_10011 ^ n_10024;
assign n_10034 = n_10025 ^ x202;
assign n_10035 = n_10026 ^ n_10021;
assign n_10036 = ~n_10027 & n_10028;
assign n_10037 = ~n_8790 & n_10029;
assign n_10038 = n_10031 ^ n_9232;
assign n_10039 = n_10031 ^ n_9359;
assign n_10040 = n_10034 ^ n_10035;
assign n_10041 = n_10035 ^ x201;
assign n_10042 = n_10036 ^ n_8101;
assign n_10043 = n_10037 ^ n_9317;
assign n_10044 = n_8829 & ~n_10038;
assign n_10045 = n_10038 ^ n_9359;
assign n_10046 = n_9372 & n_10039;
assign n_10047 = n_10040 ^ x201;
assign n_10048 = n_10040 & ~n_10041;
assign n_10049 = n_10042 ^ n_8122;
assign n_10050 = n_10043 ^ n_8122;
assign n_10051 = n_10042 ^ n_10043;
assign n_10052 = n_10044 ^ n_9359;
assign n_10053 = n_9909 ^ n_10045;
assign n_10054 = n_10046 ^ n_9232;
assign n_10055 = ~n_10047 & ~n_10032;
assign n_10056 = n_10032 ^ n_10047;
assign n_10057 = n_10048 ^ x201;
assign n_10058 = n_10049 ^ n_10043;
assign n_10059 = n_10050 & n_10051;
assign n_10060 = n_10052 ^ n_8141;
assign n_10061 = n_10054 ^ n_9273;
assign n_10062 = n_10054 ^ n_9398;
assign n_10063 = n_10057 ^ n_10058;
assign n_10064 = n_10058 ^ x200;
assign n_10065 = n_10059 ^ n_8122;
assign n_10066 = n_10061 ^ n_9398;
assign n_10067 = ~n_9411 & ~n_10062;
assign n_10068 = n_10063 ^ x200;
assign n_10069 = ~n_10063 & n_10064;
assign n_10070 = n_10065 ^ n_10060;
assign n_10071 = n_10065 ^ n_10052;
assign n_10072 = n_10066 ^ n_9385;
assign n_10073 = n_9928 ^ n_10066;
assign n_10074 = n_10067 ^ n_9273;
assign n_10075 = ~n_10055 & ~n_10068;
assign n_10076 = n_10068 ^ n_10055;
assign n_10077 = n_10069 ^ x200;
assign n_10078 = n_10060 & n_10071;
assign n_10079 = ~n_8869 & n_10072;
assign n_10080 = n_9435 ^ n_10074;
assign n_10081 = n_10077 ^ x215;
assign n_10082 = n_10070 ^ n_10077;
assign n_10083 = n_10078 ^ n_8141;
assign n_10084 = n_10079 ^ n_9385;
assign n_10085 = n_9313 ^ n_10080;
assign n_10086 = n_10080 & n_9445;
assign n_10087 = n_10070 ^ n_10081;
assign n_10088 = n_10081 & n_10082;
assign n_10089 = n_10083 ^ n_10084;
assign n_10090 = n_10084 ^ n_8161;
assign n_10091 = n_10085 ^ n_9423;
assign n_10092 = n_9949 ^ n_10085;
assign n_10093 = n_10086 ^ n_9313;
assign n_10094 = ~n_10087 & ~n_10075;
assign n_10095 = n_10075 ^ n_10087;
assign n_10096 = n_10088 ^ x215;
assign n_10097 = n_10089 ^ n_8161;
assign n_10098 = n_10089 & ~n_10090;
assign n_10099 = n_8907 & ~n_10091;
assign n_10100 = n_9466 ^ n_10093;
assign n_10101 = n_10096 ^ n_10097;
assign n_10102 = n_10097 ^ x214;
assign n_10103 = n_10098 ^ n_8161;
assign n_10104 = n_10099 ^ n_9423;
assign n_10105 = n_9353 ^ n_10100;
assign n_10106 = n_10100 & ~n_9476;
assign n_10107 = n_10101 ^ x214;
assign n_10108 = n_10101 & ~n_10102;
assign n_10109 = n_10103 ^ n_8186;
assign n_10110 = n_10104 ^ n_8186;
assign n_10111 = n_10103 ^ n_10104;
assign n_10112 = n_10105 ^ n_9466;
assign n_10113 = n_9970 ^ n_10105;
assign n_10114 = n_10106 ^ n_9353;
assign n_10115 = n_10094 & ~n_10107;
assign n_10116 = n_10107 ^ n_10094;
assign n_10117 = n_10108 ^ x214;
assign n_10118 = n_10109 ^ n_10104;
assign n_10119 = n_10110 & ~n_10111;
assign n_10120 = ~n_8946 & n_10112;
assign n_10121 = n_10114 ^ n_9496;
assign n_10122 = n_10117 ^ n_10118;
assign n_10123 = n_10118 ^ x213;
assign n_10124 = n_10119 ^ n_8186;
assign n_10125 = n_10120 ^ n_9466;
assign n_10126 = n_9394 ^ n_10121;
assign n_10127 = ~n_10121 & n_9504;
assign n_10128 = n_10122 ^ x213;
assign n_10129 = ~n_10122 & n_10123;
assign n_10130 = n_10124 ^ n_8216;
assign n_10131 = n_10125 ^ n_8216;
assign n_10132 = n_10124 ^ n_10125;
assign n_10133 = n_10126 ^ n_9496;
assign n_10134 = n_9991 ^ n_10126;
assign n_10135 = n_10127 ^ n_9394;
assign n_10136 = n_10128 & n_10115;
assign n_10137 = n_10115 ^ n_10128;
assign n_10138 = n_10129 ^ x213;
assign n_10139 = n_10130 ^ n_10125;
assign n_10140 = ~n_10131 & n_10132;
assign n_10141 = n_8983 & n_10133;
assign n_10142 = n_9521 ^ n_10135;
assign n_10143 = n_10138 ^ n_10139;
assign n_10144 = n_10139 ^ x212;
assign n_10145 = n_10140 ^ n_8216;
assign n_10146 = n_10141 ^ n_9496;
assign n_10147 = n_9431 ^ n_10142;
assign n_10148 = ~n_10142 & ~n_9529;
assign n_10149 = n_10143 ^ x212;
assign n_10150 = n_10143 & ~n_10144;
assign n_10151 = n_10145 ^ n_8250;
assign n_10152 = n_10146 ^ n_8250;
assign n_10153 = n_10145 ^ n_10146;
assign n_10154 = n_10147 ^ n_9521;
assign n_10155 = n_10012 ^ n_10147;
assign n_10156 = n_10148 ^ n_9431;
assign n_10157 = n_10136 & ~n_10149;
assign n_10158 = n_10149 ^ n_10136;
assign n_10159 = n_10150 ^ x212;
assign n_10160 = n_10151 ^ n_10146;
assign n_10161 = n_10152 & ~n_10153;
assign n_10162 = ~n_9024 & ~n_10154;
assign n_10163 = n_10156 ^ n_9536;
assign n_10164 = n_10159 ^ n_10160;
assign n_10165 = n_10160 ^ x211;
assign n_10166 = n_10161 ^ n_8250;
assign n_10167 = n_10162 ^ n_9521;
assign n_10168 = n_9484 ^ n_10163;
assign n_10169 = n_10163 & n_9543;
assign n_10170 = n_10164 ^ x211;
assign n_10171 = ~n_10164 & n_10165;
assign n_10172 = n_10166 ^ n_8288;
assign n_10173 = n_10167 ^ n_8288;
assign n_10174 = n_10166 ^ n_10167;
assign n_10175 = n_10168 ^ n_9536;
assign n_10176 = n_10033 ^ n_10168;
assign n_10177 = n_10169 ^ n_9484;
assign n_10178 = n_10157 & n_10170;
assign n_10179 = n_10170 ^ n_10157;
assign n_10180 = n_10171 ^ x211;
assign n_10181 = n_10172 ^ n_10167;
assign n_10182 = ~n_10173 & ~n_10174;
assign n_10183 = n_9063 & ~n_10175;
assign n_10184 = n_10177 ^ n_9561;
assign n_10185 = n_10180 ^ n_10181;
assign n_10186 = n_10181 ^ x210;
assign n_10187 = n_10182 ^ n_8288;
assign n_10188 = n_10183 ^ n_9536;
assign n_10189 = n_9510 ^ n_10184;
assign n_10190 = n_10184 & ~n_9568;
assign n_10191 = n_10185 ^ x210;
assign n_10192 = n_10185 & ~n_10186;
assign n_10193 = n_10187 ^ n_8329;
assign n_10194 = n_10188 ^ n_8329;
assign n_10195 = n_10187 ^ n_10188;
assign n_10196 = n_10189 ^ n_9561;
assign n_10197 = n_10056 ^ n_10189;
assign n_10198 = n_10190 ^ n_9510;
assign n_10199 = n_10178 & ~n_10191;
assign n_10200 = n_10191 ^ n_10178;
assign n_10201 = n_10192 ^ x210;
assign n_10202 = n_10193 ^ n_10188;
assign n_10203 = n_10194 & n_10195;
assign n_10204 = n_9103 & n_10196;
assign n_10205 = n_10198 ^ n_9533;
assign n_10206 = n_10198 ^ n_9580;
assign n_10207 = n_10201 ^ n_10202;
assign n_10208 = n_10202 ^ x209;
assign n_10209 = n_10203 ^ n_8329;
assign n_10210 = n_10204 ^ n_9561;
assign n_10211 = n_9132 & n_10205;
assign n_10212 = n_10205 ^ n_9580;
assign n_10213 = n_9587 & ~n_10206;
assign n_10214 = n_10207 ^ x209;
assign n_10215 = n_10207 & ~n_10208;
assign n_10216 = n_10209 ^ n_8368;
assign n_10217 = n_10210 ^ n_8368;
assign n_10218 = n_10209 ^ n_10210;
assign n_10219 = n_10211 ^ n_9580;
assign n_10220 = n_10076 ^ n_10212;
assign n_10221 = n_10213 ^ n_9533;
assign n_10222 = ~n_10199 & n_10214;
assign n_10223 = n_10214 ^ n_10199;
assign n_10224 = n_10215 ^ x209;
assign n_10225 = n_10216 ^ n_10210;
assign n_10226 = ~n_10217 & n_10218;
assign n_10227 = n_10219 ^ n_8410;
assign n_10228 = n_10221 ^ n_9600;
assign n_10229 = n_10224 ^ n_10225;
assign n_10230 = n_10225 ^ x208;
assign n_10231 = n_10226 ^ n_8368;
assign n_10232 = n_9552 ^ n_10228;
assign n_10233 = n_10228 & n_9607;
assign n_10234 = n_10229 ^ x208;
assign n_10235 = n_10229 & ~n_10230;
assign n_10236 = n_10231 ^ n_10219;
assign n_10237 = n_10232 ^ n_9594;
assign n_10238 = n_10232 ^ n_10095;
assign n_10239 = n_10233 ^ n_9552;
assign n_10240 = n_10234 ^ n_10222;
assign n_10241 = ~n_10222 & ~n_10234;
assign n_10242 = n_10235 ^ x208;
assign n_10243 = n_10236 ^ n_8410;
assign n_10244 = ~n_10236 & n_10227;
assign n_10245 = ~n_9189 & n_10237;
assign n_10246 = n_10239 ^ n_9572;
assign n_10247 = n_10239 ^ n_9620;
assign n_10248 = n_10240 ^ n_9711;
assign n_10249 = n_9711 & n_10240;
assign n_10250 = n_10242 ^ x223;
assign n_10251 = n_10243 ^ x223;
assign n_10252 = n_10243 ^ n_10242;
assign n_10253 = n_10244 ^ n_8410;
assign n_10254 = n_10245 ^ n_9594;
assign n_10255 = ~n_9229 & n_10246;
assign n_10256 = n_10246 ^ n_9620;
assign n_10257 = n_9628 & ~n_10247;
assign n_10258 = n_10248 ^ n_9704;
assign n_10259 = n_9734 ^ n_10249;
assign n_10260 = n_10243 ^ n_10250;
assign n_10261 = n_10251 & ~n_10252;
assign n_10262 = n_10253 ^ n_8452;
assign n_10263 = n_10254 ^ n_8452;
assign n_10264 = n_10253 ^ n_10254;
assign n_10265 = n_10255 ^ n_9620;
assign n_10266 = n_10116 ^ n_10256;
assign n_10267 = n_10257 ^ n_9572;
assign n_10268 = n_8677 & n_10258;
assign n_10269 = n_10241 & n_10260;
assign n_10270 = n_10260 ^ n_10241;
assign n_10271 = n_10261 ^ x223;
assign n_10272 = n_10262 ^ n_10254;
assign n_10273 = ~n_10263 & ~n_10264;
assign n_10274 = n_10265 ^ n_8493;
assign n_10275 = n_10267 ^ n_9641;
assign n_10276 = n_10268 ^ n_9704;
assign n_10277 = n_10249 ^ n_10270;
assign n_10278 = n_10259 ^ n_10270;
assign n_10279 = n_10271 ^ x222;
assign n_10280 = n_10271 ^ n_10272;
assign n_10281 = n_10273 ^ n_8452;
assign n_10282 = n_9593 ^ n_10275;
assign n_10283 = ~n_10275 & ~n_9648;
assign n_10284 = n_10276 ^ n_8171;
assign n_10285 = n_8171 & n_10276;
assign n_10286 = ~n_10277 & n_10259;
assign n_10287 = ~n_8723 & n_10277;
assign n_10288 = n_10280 & n_10279;
assign n_10289 = n_10280 ^ x222;
assign n_10290 = n_10281 ^ n_10265;
assign n_10291 = n_10282 ^ n_9641;
assign n_10292 = n_10282 ^ n_10137;
assign n_10293 = n_10283 ^ n_9593;
assign n_10294 = n_10284 ^ x359;
assign n_10295 = x359 & n_10284;
assign n_10296 = n_10285 ^ n_8200;
assign n_10297 = n_10286 ^ n_9734;
assign n_10298 = n_10287 ^ n_9734;
assign n_10299 = n_10288 ^ x222;
assign n_10300 = n_10269 & ~n_10289;
assign n_10301 = n_10289 ^ n_10269;
assign n_10302 = n_10290 ^ n_8493;
assign n_10303 = ~n_10290 & ~n_10274;
assign n_10304 = n_9270 & ~n_10291;
assign n_10305 = n_10293 ^ n_9662;
assign n_10306 = n_10295 ^ x358;
assign n_10307 = n_9770 ^ n_10297;
assign n_10308 = n_10298 ^ n_10285;
assign n_10309 = n_10298 ^ n_10296;
assign n_10310 = n_10301 ^ n_10297;
assign n_10311 = n_9770 ^ n_10301;
assign n_10312 = n_10299 ^ n_10302;
assign n_10313 = n_10302 ^ x221;
assign n_10314 = n_10303 ^ n_8493;
assign n_10315 = n_10304 ^ n_9641;
assign n_10316 = n_9613 ^ n_10305;
assign n_10317 = ~n_10305 & n_9670;
assign n_10318 = n_10307 ^ n_10301;
assign n_10319 = ~n_10296 & ~n_10308;
assign n_10320 = n_10295 ^ n_10309;
assign n_10321 = n_8779 & ~n_10310;
assign n_10322 = n_10310 & n_10311;
assign n_10323 = n_10312 ^ x221;
assign n_10324 = ~n_10312 & n_10313;
assign n_10325 = n_10314 ^ n_8535;
assign n_10326 = n_10315 ^ n_8535;
assign n_10327 = n_10314 ^ n_10315;
assign n_10328 = n_10316 ^ n_9662;
assign n_10329 = n_10158 ^ n_10316;
assign n_10330 = n_10317 ^ n_9613;
assign n_10331 = n_10319 ^ n_8200;
assign n_10332 = n_10320 & n_10306;
assign n_10333 = n_10320 ^ x358;
assign n_10334 = n_10321 ^ n_9770;
assign n_10335 = n_10322 ^ n_9770;
assign n_10336 = n_10300 & n_10323;
assign n_10337 = n_10323 ^ n_10300;
assign n_10338 = n_10324 ^ x221;
assign n_10339 = n_10325 ^ n_10315;
assign n_10340 = n_10326 & n_10327;
assign n_10341 = ~n_9310 & n_10328;
assign n_10342 = n_9685 ^ n_10330;
assign n_10343 = n_10331 ^ n_8243;
assign n_10344 = n_10332 ^ x358;
assign n_10345 = n_10294 & ~n_10333;
assign n_10346 = n_10333 ^ n_10294;
assign n_10347 = n_10334 ^ n_8243;
assign n_10348 = n_10331 ^ n_10334;
assign n_10349 = n_9796 ^ n_10335;
assign n_10350 = n_10337 ^ n_10335;
assign n_10351 = n_9796 ^ n_10337;
assign n_10352 = n_10338 ^ n_10339;
assign n_10353 = n_10339 ^ x220;
assign n_10354 = n_10340 ^ n_8535;
assign n_10355 = n_10341 ^ n_9662;
assign n_10356 = n_9634 ^ n_10342;
assign n_10357 = ~n_10342 & ~n_9692;
assign n_10358 = n_10343 ^ n_10334;
assign n_10359 = n_10347 & ~n_10348;
assign n_10360 = n_10349 ^ n_10337;
assign n_10361 = ~n_8820 & ~n_10350;
assign n_10362 = n_10350 & n_10351;
assign n_10363 = n_10352 ^ x220;
assign n_10364 = ~n_10352 & n_10353;
assign n_10365 = n_10354 ^ n_8576;
assign n_10366 = n_10355 ^ n_8576;
assign n_10367 = n_10354 ^ n_10355;
assign n_10368 = n_10356 ^ n_9676;
assign n_10369 = n_10179 ^ n_10356;
assign n_10370 = n_10357 ^ n_9634;
assign n_10371 = n_10344 ^ n_10358;
assign n_10372 = n_10358 ^ x357;
assign n_10373 = n_10359 ^ n_8243;
assign n_10374 = n_10361 ^ n_9796;
assign n_10375 = n_10362 ^ n_9796;
assign n_10376 = n_10336 & n_10363;
assign n_10377 = n_10363 ^ n_10336;
assign n_10378 = n_10364 ^ x220;
assign n_10379 = n_10365 ^ n_10355;
assign n_10380 = ~n_10366 & n_10367;
assign n_10381 = ~n_9350 & n_10368;
assign n_10382 = n_10370 ^ n_9705;
assign n_10383 = n_10371 ^ x357;
assign n_10384 = n_10371 & ~n_10372;
assign n_10385 = n_10373 ^ n_8281;
assign n_10386 = n_10374 ^ n_10373;
assign n_10387 = n_10375 ^ n_9818;
assign n_10388 = n_9818 ^ n_10377;
assign n_10389 = n_10375 ^ n_10377;
assign n_10390 = n_10378 ^ n_10379;
assign n_10391 = n_10379 ^ x219;
assign n_10392 = n_10380 ^ n_8576;
assign n_10393 = n_10381 ^ n_9676;
assign n_10394 = n_9660 ^ n_10382;
assign n_10395 = ~n_10382 & ~n_9713;
assign n_10396 = n_10345 & ~n_10383;
assign n_10397 = n_10383 ^ n_10345;
assign n_10398 = n_10384 ^ x357;
assign n_10399 = n_10374 ^ n_10385;
assign n_10400 = n_10385 & n_10386;
assign n_10401 = n_10387 ^ n_10377;
assign n_10402 = ~n_10388 & ~n_10389;
assign n_10403 = ~n_8861 & n_10389;
assign n_10404 = n_10390 ^ x219;
assign n_10405 = ~n_10390 & n_10391;
assign n_10406 = n_10392 ^ n_8619;
assign n_10407 = n_10393 ^ n_8619;
assign n_10408 = n_10392 ^ n_10393;
assign n_10409 = n_10394 ^ n_9705;
assign n_10410 = n_10200 ^ n_10394;
assign n_10411 = n_10395 ^ n_9660;
assign n_10412 = n_10398 ^ n_10399;
assign n_10413 = n_10399 ^ x356;
assign n_10414 = n_10400 ^ n_8281;
assign n_10415 = n_10402 ^ n_9818;
assign n_10416 = n_10403 ^ n_9818;
assign n_10417 = n_10376 & n_10404;
assign n_10418 = n_10404 ^ n_10376;
assign n_10419 = n_10405 ^ x219;
assign n_10420 = n_10406 ^ n_10393;
assign n_10421 = ~n_10407 & ~n_10408;
assign n_10422 = ~n_9391 & ~n_10409;
assign n_10423 = n_10411 ^ n_9730;
assign n_10424 = n_10412 ^ x356;
assign n_10425 = ~n_10412 & n_10413;
assign n_10426 = n_10414 ^ n_8322;
assign n_10427 = n_10415 ^ n_9832;
assign n_10428 = n_10416 ^ n_8322;
assign n_10429 = n_10414 ^ n_10416;
assign n_10430 = n_10418 ^ n_10415;
assign n_10431 = n_10419 ^ n_10420;
assign n_10432 = n_10420 ^ x218;
assign n_10433 = n_10421 ^ n_8619;
assign n_10434 = n_10422 ^ n_9705;
assign n_10435 = n_10423 ^ n_9682;
assign n_10436 = n_10396 & n_10424;
assign n_10437 = n_10424 ^ n_10396;
assign n_10438 = n_10425 ^ x356;
assign n_10439 = n_10426 ^ n_10416;
assign n_10440 = n_10418 ^ n_10427;
assign n_10441 = ~n_10428 & ~n_10429;
assign n_10442 = ~n_10427 & n_10430;
assign n_10443 = ~n_8902 & ~n_10430;
assign n_10444 = n_10431 ^ x218;
assign n_10445 = ~n_10431 & n_10432;
assign n_10446 = n_10433 ^ n_8659;
assign n_10447 = n_10434 ^ n_8659;
assign n_10448 = n_10433 ^ n_10434;
assign n_10449 = n_10435 ^ n_9730;
assign n_10450 = n_10223 ^ n_10435;
assign n_10451 = n_10438 ^ n_10439;
assign n_10452 = n_10439 ^ x355;
assign n_10453 = n_10441 ^ n_8322;
assign n_10454 = n_10442 ^ n_9832;
assign n_10455 = n_10443 ^ n_9832;
assign n_10456 = n_10417 & n_10444;
assign n_10457 = n_10444 ^ n_10417;
assign n_10458 = n_10445 ^ x218;
assign n_10459 = n_10446 ^ n_10434;
assign n_10460 = n_10447 & n_10448;
assign n_10461 = n_9429 & n_10449;
assign n_10462 = n_10451 ^ x355;
assign n_10463 = ~n_10451 & n_10452;
assign n_10464 = n_10453 ^ n_8361;
assign n_10465 = n_10454 ^ n_9850;
assign n_10466 = n_10455 ^ n_8361;
assign n_10467 = n_10453 ^ n_10455;
assign n_10468 = n_9850 ^ n_10457;
assign n_10469 = n_10454 ^ n_10457;
assign n_10470 = n_10458 ^ n_10459;
assign n_10471 = n_10459 ^ x217;
assign n_10472 = n_10460 ^ n_8659;
assign n_10473 = n_10461 ^ n_9730;
assign n_10474 = ~n_10436 & ~n_10462;
assign n_10475 = n_10462 ^ n_10436;
assign n_10476 = n_10463 ^ x355;
assign n_10477 = n_10464 ^ n_10455;
assign n_10478 = n_10465 ^ n_10457;
assign n_10479 = n_10466 & ~n_10467;
assign n_10480 = ~n_10468 & ~n_10469;
assign n_10481 = ~n_8942 & n_10469;
assign n_10482 = n_10470 ^ x217;
assign n_10483 = ~n_10470 & n_10471;
assign n_10484 = n_10472 ^ x216;
assign n_10485 = n_10473 ^ n_8690;
assign n_10486 = n_10476 ^ n_10477;
assign n_10487 = n_10477 ^ x354;
assign n_10488 = n_10479 ^ n_8361;
assign n_10489 = n_10480 ^ n_9850;
assign n_10490 = n_10481 ^ n_9850;
assign n_10491 = ~n_10456 & ~n_10482;
assign n_10492 = n_10482 ^ n_10456;
assign n_10493 = n_10483 ^ x217;
assign n_10494 = n_10484 ^ n_10485;
assign n_10495 = n_10486 ^ x354;
assign n_10496 = ~n_10486 & n_10487;
assign n_10497 = n_10488 ^ n_8403;
assign n_10498 = n_10489 ^ n_9863;
assign n_10499 = n_10490 ^ n_8403;
assign n_10500 = n_10488 ^ n_10490;
assign n_10501 = n_10492 ^ n_9863;
assign n_10502 = n_10489 ^ n_10492;
assign n_10503 = n_10493 ^ n_10491;
assign n_10504 = ~n_10474 & n_10495;
assign n_10505 = n_10495 ^ n_10474;
assign n_10506 = n_10496 ^ x354;
assign n_10507 = n_10497 ^ n_10490;
assign n_10508 = n_10498 ^ n_10492;
assign n_10509 = ~n_10499 & n_10500;
assign n_10510 = n_10501 & ~n_10502;
assign n_10511 = ~n_8987 & n_10502;
assign n_10512 = n_10503 ^ n_10494;
assign n_10513 = n_10506 ^ n_10507;
assign n_10514 = n_10507 ^ x353;
assign n_10515 = n_10509 ^ n_8403;
assign n_10516 = n_10510 ^ n_9863;
assign n_10517 = n_10511 ^ n_9863;
assign n_10518 = n_10512 ^ n_9878;
assign n_10519 = n_10513 ^ x353;
assign n_10520 = n_10513 & ~n_10514;
assign n_10521 = n_10515 ^ n_8446;
assign n_10522 = n_10516 ^ n_10512;
assign n_10523 = n_10516 ^ n_9878;
assign n_10524 = n_10517 ^ n_10515;
assign n_10525 = ~n_10504 & n_10519;
assign n_10526 = n_10519 ^ n_10504;
assign n_10527 = n_10520 ^ x353;
assign n_10528 = n_10517 ^ n_10521;
assign n_10529 = n_10518 & ~n_10522;
assign n_10530 = n_9026 & n_10522;
assign n_10531 = n_10523 ^ n_10512;
assign n_10532 = ~n_10521 & n_10524;
assign n_10533 = n_10527 ^ n_10528;
assign n_10534 = n_10528 ^ x352;
assign n_10535 = n_10529 ^ n_9878;
assign n_10536 = n_10530 ^ n_9878;
assign n_10537 = n_10532 ^ n_8446;
assign n_10538 = n_10533 ^ x352;
assign n_10539 = ~n_10533 & n_10534;
assign n_10540 = n_9898 ^ n_10535;
assign n_10541 = n_10536 ^ n_8486;
assign n_10542 = n_10537 ^ n_10536;
assign n_10543 = n_10537 ^ n_8486;
assign n_10544 = ~n_10525 & n_10538;
assign n_10545 = n_10538 ^ n_10525;
assign n_10546 = n_10539 ^ x352;
assign n_10547 = n_10540 & n_9906;
assign n_10548 = n_9757 ^ n_10540;
assign n_10549 = n_10541 & ~n_10542;
assign n_10550 = n_10543 ^ n_10536;
assign n_10551 = n_10547 ^ n_9757;
assign n_10552 = n_10548 ^ n_9891;
assign n_10553 = n_10549 ^ n_8486;
assign n_10554 = n_10546 ^ n_10550;
assign n_10555 = n_10550 ^ x367;
assign n_10556 = n_10551 ^ n_9918;
assign n_10557 = ~n_9068 & n_10552;
assign n_10558 = n_10553 ^ n_8528;
assign n_10559 = n_10554 ^ x367;
assign n_10560 = n_10554 & ~n_10555;
assign n_10561 = ~n_10556 & ~n_9925;
assign n_10562 = n_9777 ^ n_10556;
assign n_10563 = n_10557 ^ n_9891;
assign n_10564 = n_10544 & ~n_10559;
assign n_10565 = n_10559 ^ n_10544;
assign n_10566 = n_10560 ^ x367;
assign n_10567 = n_10561 ^ n_9777;
assign n_10568 = n_10562 ^ n_9918;
assign n_10569 = n_10563 ^ n_8528;
assign n_10570 = n_10553 ^ n_10563;
assign n_10571 = n_10558 ^ n_10563;
assign n_10572 = n_10567 ^ n_9938;
assign n_10573 = ~n_9110 & ~n_10568;
assign n_10574 = ~n_10569 & ~n_10570;
assign n_10575 = n_10566 ^ n_10571;
assign n_10576 = n_10571 ^ x366;
assign n_10577 = n_10572 & n_9946;
assign n_10578 = n_9806 ^ n_10572;
assign n_10579 = n_10573 ^ n_9918;
assign n_10580 = n_10574 ^ n_8528;
assign n_10581 = n_10575 ^ x366;
assign n_10582 = ~n_10575 & n_10576;
assign n_10583 = n_10577 ^ n_9806;
assign n_10584 = n_10578 ^ n_9938;
assign n_10585 = n_10579 ^ n_8569;
assign n_10586 = n_10580 ^ n_10579;
assign n_10587 = n_10580 ^ n_8569;
assign n_10588 = ~n_10581 & ~n_10564;
assign n_10589 = n_10564 ^ n_10581;
assign n_10590 = n_10582 ^ x366;
assign n_10591 = n_10583 ^ n_9959;
assign n_10592 = n_9154 & ~n_10584;
assign n_10593 = ~n_10585 & ~n_10586;
assign n_10594 = n_10587 ^ n_10579;
assign n_10595 = ~n_10591 & n_9967;
assign n_10596 = n_9824 ^ n_10591;
assign n_10597 = n_10592 ^ n_9938;
assign n_10598 = n_10593 ^ n_8569;
assign n_10599 = n_10590 ^ n_10594;
assign n_10600 = n_10594 ^ x365;
assign n_10601 = n_10595 ^ n_9824;
assign n_10602 = n_10596 ^ n_9959;
assign n_10603 = n_10597 ^ n_8612;
assign n_10604 = n_10598 ^ n_10597;
assign n_10605 = n_10598 ^ n_8612;
assign n_10606 = n_10599 ^ x365;
assign n_10607 = n_10599 & ~n_10600;
assign n_10608 = n_10601 ^ n_9980;
assign n_10609 = n_9196 & n_10602;
assign n_10610 = ~n_10603 & n_10604;
assign n_10611 = n_10605 ^ n_10597;
assign n_10612 = ~n_10588 & ~n_10606;
assign n_10613 = n_10606 ^ n_10588;
assign n_10614 = n_10607 ^ x365;
assign n_10615 = n_10608 & ~n_9988;
assign n_10616 = n_9840 ^ n_10608;
assign n_10617 = n_10609 ^ n_9959;
assign n_10618 = n_10610 ^ n_8612;
assign n_10619 = n_10611 ^ x364;
assign n_10620 = n_10614 ^ n_10611;
assign n_10621 = n_10615 ^ n_9840;
assign n_10622 = n_10616 ^ n_9980;
assign n_10623 = n_10617 ^ n_8652;
assign n_10624 = n_10618 ^ n_10617;
assign n_10625 = n_10618 ^ n_8652;
assign n_10626 = ~n_10620 & n_10619;
assign n_10627 = n_10620 ^ x364;
assign n_10628 = n_10621 ^ n_10001;
assign n_10629 = n_9236 & n_10622;
assign n_10630 = ~n_10623 & n_10624;
assign n_10631 = n_10625 ^ n_10617;
assign n_10632 = n_10626 ^ x364;
assign n_10633 = ~n_10627 & ~n_10612;
assign n_10634 = n_10612 ^ n_10627;
assign n_10635 = n_9861 ^ n_10628;
assign n_10636 = n_10628 & ~n_10009;
assign n_10637 = n_10629 ^ n_9980;
assign n_10638 = n_10630 ^ n_8652;
assign n_10639 = n_10631 ^ x363;
assign n_10640 = n_10632 ^ n_10631;
assign n_10641 = n_10294 ^ n_10635;
assign n_10642 = n_10635 ^ n_10001;
assign n_10643 = n_10636 ^ n_9861;
assign n_10644 = n_10637 ^ n_8698;
assign n_10645 = n_10638 ^ n_10637;
assign n_10646 = n_10638 ^ n_8698;
assign n_10647 = ~n_10640 & n_10639;
assign n_10648 = n_10640 ^ x363;
assign n_10649 = ~n_9277 & n_10642;
assign n_10650 = n_10643 ^ n_10022;
assign n_10651 = n_10643 ^ n_10030;
assign n_10652 = n_10644 & ~n_10645;
assign n_10653 = n_10646 ^ n_10637;
assign n_10654 = n_10647 ^ x363;
assign n_10655 = n_10633 & ~n_10648;
assign n_10656 = n_10648 ^ n_10633;
assign n_10657 = n_10649 ^ n_10001;
assign n_10658 = ~n_10030 & n_10650;
assign n_10659 = n_10651 ^ n_10022;
assign n_10660 = n_10346 ^ n_10651;
assign n_10661 = n_10652 ^ n_8698;
assign n_10662 = n_10653 ^ x362;
assign n_10663 = n_10654 ^ n_10653;
assign n_10664 = n_10657 ^ n_8744;
assign n_10665 = n_10658 ^ n_9880;
assign n_10666 = ~n_9317 & n_10659;
assign n_10667 = n_10661 ^ n_10657;
assign n_10668 = n_10661 ^ n_8744;
assign n_10669 = n_10663 & ~n_10662;
assign n_10670 = n_10663 ^ x362;
assign n_10671 = n_10665 ^ n_10045;
assign n_10672 = n_10665 ^ n_9909;
assign n_10673 = n_10666 ^ n_10022;
assign n_10674 = ~n_10664 & ~n_10667;
assign n_10675 = n_10668 ^ n_10657;
assign n_10676 = n_10669 ^ x362;
assign n_10677 = ~n_10655 & ~n_10670;
assign n_10678 = n_10670 ^ n_10655;
assign n_10679 = n_10053 & n_10671;
assign n_10680 = n_9359 & ~n_10672;
assign n_10681 = n_10672 ^ n_10045;
assign n_10682 = n_10674 ^ n_8744;
assign n_10683 = n_10676 ^ n_10675;
assign n_10684 = n_10676 ^ x361;
assign n_10685 = n_10679 ^ n_9909;
assign n_10686 = n_10680 ^ n_10045;
assign n_10687 = n_10681 ^ n_10397;
assign n_10688 = n_10682 ^ n_8790;
assign n_10689 = n_10673 ^ n_10682;
assign n_10690 = n_10683 ^ x361;
assign n_10691 = ~n_10683 & n_10684;
assign n_10692 = n_10685 ^ n_10066;
assign n_10693 = n_10685 ^ n_9928;
assign n_10694 = n_10686 ^ n_8829;
assign n_10695 = n_10673 ^ n_10688;
assign n_10696 = ~n_10688 & n_10689;
assign n_10697 = ~n_10690 & ~n_10677;
assign n_10698 = n_10677 ^ n_10690;
assign n_10699 = n_10691 ^ x361;
assign n_10700 = ~n_10073 & ~n_10692;
assign n_10701 = n_10693 ^ n_10066;
assign n_10702 = n_10695 ^ x360;
assign n_10703 = n_10696 ^ n_8790;
assign n_10704 = n_10699 ^ n_10695;
assign n_10705 = n_10700 ^ n_9928;
assign n_10706 = n_10701 ^ n_10061;
assign n_10707 = n_10437 ^ n_10701;
assign n_10708 = n_10703 ^ n_10686;
assign n_10709 = ~n_10704 & n_10702;
assign n_10710 = n_10704 ^ x360;
assign n_10711 = n_10705 ^ n_10085;
assign n_10712 = n_9398 & ~n_10706;
assign n_10713 = ~n_10708 & ~n_10694;
assign n_10714 = n_10708 ^ n_8829;
assign n_10715 = n_10709 ^ x360;
assign n_10716 = ~n_10697 & n_10710;
assign n_10717 = n_10710 ^ n_10697;
assign n_10718 = n_10711 & n_10092;
assign n_10719 = n_9949 ^ n_10711;
assign n_10720 = n_10712 ^ n_10061;
assign n_10721 = n_10713 ^ n_8829;
assign n_10722 = n_10714 ^ x375;
assign n_10723 = n_10715 ^ n_10714;
assign n_10724 = n_10715 ^ x375;
assign n_10725 = n_10718 ^ n_9949;
assign n_10726 = n_10719 ^ n_10085;
assign n_10727 = n_10475 ^ n_10719;
assign n_10728 = n_10720 ^ n_8869;
assign n_10729 = n_10721 ^ n_10720;
assign n_10730 = n_10722 & ~n_10723;
assign n_10731 = n_10724 ^ n_10714;
assign n_10732 = n_10725 ^ n_10105;
assign n_10733 = n_9435 & ~n_10726;
assign n_10734 = n_10729 & n_10728;
assign n_10735 = n_10729 ^ n_8869;
assign n_10736 = n_10730 ^ x375;
assign n_10737 = n_10716 & n_10731;
assign n_10738 = n_10731 ^ n_10716;
assign n_10739 = ~n_10732 & ~n_10113;
assign n_10740 = n_9970 ^ n_10732;
assign n_10741 = n_10733 ^ n_10085;
assign n_10742 = n_10734 ^ n_8869;
assign n_10743 = n_10735 ^ x374;
assign n_10744 = n_10735 ^ n_10736;
assign n_10745 = n_10739 ^ n_9970;
assign n_10746 = n_10740 ^ n_10105;
assign n_10747 = n_10505 ^ n_10740;
assign n_10748 = n_10741 ^ n_8907;
assign n_10749 = n_10742 ^ n_10741;
assign n_10750 = n_10742 ^ n_8907;
assign n_10751 = ~n_10744 & n_10743;
assign n_10752 = n_10744 ^ x374;
assign n_10753 = n_10745 ^ n_10126;
assign n_10754 = ~n_9466 & ~n_10746;
assign n_10755 = ~n_10748 & ~n_10749;
assign n_10756 = n_10750 ^ n_10741;
assign n_10757 = n_10751 ^ x374;
assign n_10758 = ~n_10752 & ~n_10737;
assign n_10759 = n_10737 ^ n_10752;
assign n_10760 = ~n_10753 & n_10134;
assign n_10761 = n_9991 ^ n_10753;
assign n_10762 = n_10754 ^ n_10105;
assign n_10763 = n_10755 ^ n_8907;
assign n_10764 = n_10756 ^ x373;
assign n_10765 = n_10757 ^ n_10756;
assign n_10766 = n_10760 ^ n_9991;
assign n_10767 = n_10761 ^ n_10126;
assign n_10768 = n_10526 ^ n_10761;
assign n_10769 = n_10762 ^ n_8946;
assign n_10770 = n_10763 ^ n_10762;
assign n_10771 = n_10763 ^ n_8946;
assign n_10772 = ~n_10765 & n_10764;
assign n_10773 = n_10765 ^ x373;
assign n_10774 = n_10766 ^ n_10147;
assign n_10775 = n_9496 & n_10767;
assign n_10776 = n_10769 & n_10770;
assign n_10777 = n_10771 ^ n_10762;
assign n_10778 = n_10772 ^ x373;
assign n_10779 = ~n_10773 & n_10758;
assign n_10780 = n_10758 ^ n_10773;
assign n_10781 = n_10774 & ~n_10155;
assign n_10782 = n_10012 ^ n_10774;
assign n_10783 = n_10775 ^ n_10126;
assign n_10784 = n_10776 ^ n_8946;
assign n_10785 = n_10777 ^ x372;
assign n_10786 = n_10778 ^ n_10777;
assign n_10787 = n_10248 & n_10780;
assign n_10788 = n_10780 ^ n_10248;
assign n_10789 = n_10781 ^ n_10012;
assign n_10790 = n_10782 ^ n_10147;
assign n_10791 = n_10545 ^ n_10782;
assign n_10792 = n_10783 ^ n_8983;
assign n_10793 = n_10784 ^ n_10783;
assign n_10794 = n_10784 ^ n_8983;
assign n_10795 = ~n_10786 & n_10785;
assign n_10796 = n_10786 ^ x372;
assign n_10797 = n_10278 ^ n_10787;
assign n_10798 = n_10788 ^ n_10240;
assign n_10799 = n_10789 ^ n_10168;
assign n_10800 = n_9521 & n_10790;
assign n_10801 = n_10792 & n_10793;
assign n_10802 = n_10794 ^ n_10783;
assign n_10803 = n_10795 ^ x372;
assign n_10804 = n_10779 & ~n_10796;
assign n_10805 = n_10796 ^ n_10779;
assign n_10806 = n_9711 & n_10798;
assign n_10807 = n_10799 & n_10176;
assign n_10808 = n_10033 ^ n_10799;
assign n_10809 = n_10800 ^ n_10147;
assign n_10810 = n_10801 ^ n_8983;
assign n_10811 = n_10802 ^ x371;
assign n_10812 = n_10803 ^ n_10802;
assign n_10813 = n_10805 ^ n_10787;
assign n_10814 = n_10797 ^ n_10805;
assign n_10815 = n_10806 ^ n_10240;
assign n_10816 = n_10807 ^ n_10033;
assign n_10817 = n_10808 ^ n_10168;
assign n_10818 = n_10565 ^ n_10808;
assign n_10819 = n_10809 ^ n_9024;
assign n_10820 = n_10810 ^ n_10809;
assign n_10821 = n_10810 ^ n_9024;
assign n_10822 = n_10812 & ~n_10811;
assign n_10823 = n_10812 ^ x371;
assign n_10824 = ~n_10813 & n_10797;
assign n_10825 = n_9734 & n_10813;
assign n_10826 = n_8677 & n_10815;
assign n_10827 = n_10815 ^ n_8677;
assign n_10828 = n_10816 ^ n_10189;
assign n_10829 = n_9536 & ~n_10817;
assign n_10830 = n_10819 & n_10820;
assign n_10831 = n_10821 ^ n_10809;
assign n_10832 = n_10822 ^ x371;
assign n_10833 = n_10804 & n_10823;
assign n_10834 = n_10823 ^ n_10804;
assign n_10835 = n_10824 ^ n_10278;
assign n_10836 = n_10825 ^ n_10278;
assign n_10837 = n_10826 ^ n_8723;
assign n_10838 = x7 & n_10827;
assign n_10839 = n_10827 ^ x7;
assign n_10840 = n_10056 ^ n_10828;
assign n_10841 = ~n_10828 & ~n_10197;
assign n_10842 = n_10829 ^ n_10168;
assign n_10843 = n_10830 ^ n_9024;
assign n_10844 = n_10832 ^ n_10831;
assign n_10845 = n_10832 ^ x370;
assign n_10846 = n_10318 ^ n_10834;
assign n_10847 = n_10835 ^ n_10834;
assign n_10848 = n_10318 ^ n_10835;
assign n_10849 = n_10836 ^ n_10826;
assign n_10850 = n_10836 ^ n_10837;
assign n_10851 = n_10838 ^ x6;
assign n_10852 = n_10840 ^ n_10189;
assign n_10853 = n_10589 ^ n_10840;
assign n_10854 = n_10841 ^ n_10056;
assign n_10855 = n_10842 ^ n_9063;
assign n_10856 = n_10843 ^ n_10842;
assign n_10857 = n_10843 ^ n_9063;
assign n_10858 = n_10844 ^ x370;
assign n_10859 = ~n_10844 & n_10845;
assign n_10860 = n_10847 & ~n_10846;
assign n_10861 = ~n_9770 & ~n_10847;
assign n_10862 = n_10848 ^ n_10834;
assign n_10863 = ~n_10837 & ~n_10849;
assign n_10864 = n_10850 ^ n_10838;
assign n_10865 = n_10850 ^ n_10851;
assign n_10866 = ~n_9561 & ~n_10852;
assign n_10867 = n_10212 ^ n_10854;
assign n_10868 = ~n_10855 & ~n_10856;
assign n_10869 = n_10857 ^ n_10842;
assign n_10870 = ~n_10833 & n_10858;
assign n_10871 = n_10858 ^ n_10833;
assign n_10872 = n_10859 ^ x370;
assign n_10873 = n_10860 ^ n_10318;
assign n_10874 = n_10861 ^ n_10318;
assign n_10875 = n_10863 ^ n_8723;
assign n_10876 = n_10851 & n_10864;
assign n_10877 = n_10866 ^ n_10189;
assign n_10878 = n_10076 ^ n_10867;
assign n_10879 = ~n_10867 & ~n_10220;
assign n_10880 = n_10868 ^ n_9063;
assign n_10881 = n_10869 ^ x369;
assign n_10882 = n_10360 ^ n_10871;
assign n_10883 = n_10872 ^ n_10869;
assign n_10884 = n_10873 ^ n_10871;
assign n_10885 = n_10360 ^ n_10873;
assign n_10886 = n_10874 ^ n_8779;
assign n_10887 = n_10875 ^ n_10874;
assign n_10888 = n_10875 ^ n_8779;
assign n_10889 = n_10876 ^ x6;
assign n_10890 = n_10877 ^ n_9103;
assign n_10891 = n_10878 ^ n_10205;
assign n_10892 = n_10613 ^ n_10878;
assign n_10893 = n_10879 ^ n_10076;
assign n_10894 = n_10880 ^ n_10877;
assign n_10895 = n_10880 ^ n_9103;
assign n_10896 = ~n_10883 & n_10881;
assign n_10897 = n_10883 ^ x369;
assign n_10898 = n_10884 & n_10882;
assign n_10899 = n_9796 & ~n_10884;
assign n_10900 = n_10885 ^ n_10871;
assign n_10901 = n_10886 & n_10887;
assign n_10902 = n_10888 ^ n_10874;
assign n_10903 = n_9580 & ~n_10891;
assign n_10904 = n_10893 ^ n_10095;
assign n_10905 = n_10893 ^ n_10232;
assign n_10906 = ~n_10890 & n_10894;
assign n_10907 = n_10895 ^ n_10877;
assign n_10908 = n_10896 ^ x369;
assign n_10909 = ~n_10870 & ~n_10897;
assign n_10910 = n_10897 ^ n_10870;
assign n_10911 = n_10898 ^ n_10360;
assign n_10912 = n_10899 ^ n_10360;
assign n_10913 = n_10901 ^ n_8779;
assign n_10914 = n_10889 ^ n_10902;
assign n_10915 = n_10902 ^ x5;
assign n_10916 = n_10903 ^ n_10205;
assign n_10917 = ~n_9600 & ~n_10904;
assign n_10918 = n_10904 ^ n_10232;
assign n_10919 = n_10238 & n_10905;
assign n_10920 = n_10906 ^ n_9103;
assign n_10921 = n_10907 ^ x368;
assign n_10922 = n_10908 ^ n_10907;
assign n_10923 = n_10910 ^ n_10911;
assign n_10924 = n_10401 ^ n_10911;
assign n_10925 = n_10912 ^ n_8820;
assign n_10926 = n_10913 ^ n_10912;
assign n_10927 = n_10913 ^ n_8820;
assign n_10928 = n_10914 ^ x5;
assign n_10929 = n_10914 & ~n_10915;
assign n_10930 = n_10916 ^ n_9132;
assign n_10931 = n_10917 ^ n_10232;
assign n_10932 = n_10634 ^ n_10918;
assign n_10933 = n_10919 ^ n_10095;
assign n_10934 = n_10920 ^ n_10916;
assign n_10935 = n_10922 & ~n_10921;
assign n_10936 = n_10922 ^ x368;
assign n_10937 = ~n_9818 & n_10923;
assign n_10938 = ~n_10923 & n_10924;
assign n_10939 = n_10924 ^ n_10910;
assign n_10940 = n_10925 & n_10926;
assign n_10941 = n_10927 ^ n_10912;
assign n_10942 = ~n_10928 & ~n_10865;
assign n_10943 = n_10865 ^ n_10928;
assign n_10944 = n_10929 ^ x5;
assign n_10945 = n_10931 ^ n_9189;
assign n_10946 = n_10256 ^ n_10933;
assign n_10947 = ~n_10934 & n_10930;
assign n_10948 = n_10934 ^ n_9132;
assign n_10949 = n_10935 ^ x368;
assign n_10950 = ~n_10936 & ~n_10909;
assign n_10951 = n_10909 ^ n_10936;
assign n_10952 = n_10937 ^ n_10401;
assign n_10953 = n_10938 ^ n_10401;
assign n_10954 = n_10940 ^ n_8820;
assign n_10955 = n_10941 ^ x4;
assign n_10956 = n_10944 ^ n_10941;
assign n_10957 = n_10116 ^ n_10946;
assign n_10958 = n_10946 & n_10266;
assign n_10959 = n_10947 ^ n_9132;
assign n_10960 = n_10948 ^ x383;
assign n_10961 = n_10949 ^ n_10948;
assign n_10962 = n_10949 ^ x383;
assign n_10963 = n_10440 ^ n_10951;
assign n_10964 = n_10952 ^ n_8861;
assign n_10965 = n_10951 ^ n_10953;
assign n_10966 = n_10440 ^ n_10953;
assign n_10967 = n_10954 ^ n_10952;
assign n_10968 = n_10954 ^ n_8861;
assign n_10969 = ~n_10956 & n_10955;
assign n_10970 = n_10956 ^ x4;
assign n_10971 = n_10957 ^ n_10246;
assign n_10972 = n_10656 ^ n_10957;
assign n_10973 = n_10958 ^ n_10116;
assign n_10974 = n_10959 ^ n_9189;
assign n_10975 = n_10959 ^ n_10931;
assign n_10976 = n_10960 & ~n_10961;
assign n_10977 = n_10962 ^ n_10948;
assign n_10978 = n_10965 & ~n_10963;
assign n_10979 = n_9832 & ~n_10965;
assign n_10980 = n_10966 ^ n_10951;
assign n_10981 = n_10964 & ~n_10967;
assign n_10982 = n_10968 ^ n_10952;
assign n_10983 = n_10969 ^ x4;
assign n_10984 = ~n_10942 & ~n_10970;
assign n_10985 = n_10970 ^ n_10942;
assign n_10986 = ~n_9620 & n_10971;
assign n_10987 = n_10973 ^ n_10137;
assign n_10988 = n_10973 ^ n_10282;
assign n_10989 = n_10974 ^ n_10931;
assign n_10990 = ~n_10945 & ~n_10975;
assign n_10991 = n_10976 ^ x383;
assign n_10992 = n_10977 & n_10950;
assign n_10993 = n_10950 ^ n_10977;
assign n_10994 = n_10978 ^ n_10440;
assign n_10995 = n_10979 ^ n_10440;
assign n_10996 = n_10981 ^ n_8861;
assign n_10997 = n_10982 ^ x3;
assign n_10998 = n_10983 ^ n_10982;
assign n_10999 = n_10986 ^ n_10246;
assign n_11000 = ~n_9641 & ~n_10987;
assign n_11001 = n_10987 ^ n_10282;
assign n_11002 = n_10292 & n_10988;
assign n_11003 = n_10990 ^ n_9189;
assign n_11004 = n_10989 ^ n_10991;
assign n_11005 = n_10991 ^ x382;
assign n_11006 = n_10478 ^ n_10993;
assign n_11007 = n_10994 ^ n_10993;
assign n_11008 = n_10478 ^ n_10994;
assign n_11009 = n_10995 ^ n_8902;
assign n_11010 = n_10996 ^ n_10995;
assign n_11011 = n_10996 ^ n_8902;
assign n_11012 = n_10998 & ~n_10997;
assign n_11013 = n_10998 ^ x3;
assign n_11014 = n_10999 ^ n_9229;
assign n_11015 = n_11000 ^ n_10282;
assign n_11016 = n_10678 ^ n_11001;
assign n_11017 = n_11002 ^ n_10137;
assign n_11018 = n_11003 ^ n_9229;
assign n_11019 = n_11003 ^ n_10999;
assign n_11020 = n_11004 ^ x382;
assign n_11021 = n_11004 & n_11005;
assign n_11022 = n_11007 & ~n_11006;
assign n_11023 = ~n_9850 & ~n_11007;
assign n_11024 = n_11008 ^ n_10993;
assign n_11025 = n_11009 & ~n_11010;
assign n_11026 = n_11011 ^ n_10995;
assign n_11027 = n_11012 ^ x3;
assign n_11028 = ~n_10984 & ~n_11013;
assign n_11029 = n_11013 ^ n_10984;
assign n_11030 = n_11015 ^ n_9270;
assign n_11031 = n_11017 ^ n_10316;
assign n_11032 = n_11018 ^ n_10999;
assign n_11033 = ~n_11014 & n_11019;
assign n_11034 = n_11020 & ~n_10992;
assign n_11035 = n_10992 ^ n_11020;
assign n_11036 = n_11021 ^ x382;
assign n_11037 = n_11022 ^ n_10478;
assign n_11038 = n_11023 ^ n_10478;
assign n_11039 = n_11025 ^ n_8902;
assign n_11040 = n_11026 ^ x2;
assign n_11041 = n_11027 ^ n_11026;
assign n_11042 = n_10158 ^ n_11031;
assign n_11043 = ~n_11031 & ~n_10329;
assign n_11044 = n_11032 ^ x381;
assign n_11045 = n_11033 ^ n_9229;
assign n_11046 = n_10508 ^ n_11035;
assign n_11047 = n_11036 ^ n_11032;
assign n_11048 = n_11037 ^ n_11035;
assign n_11049 = n_10508 ^ n_11037;
assign n_11050 = n_11038 ^ n_8942;
assign n_11051 = n_11039 ^ n_11038;
assign n_11052 = n_11039 ^ n_8942;
assign n_11053 = n_11041 & ~n_11040;
assign n_11054 = n_11041 ^ x2;
assign n_11055 = n_11042 ^ n_10316;
assign n_11056 = n_10698 ^ n_11042;
assign n_11057 = n_11043 ^ n_10158;
assign n_11058 = n_11045 ^ n_9270;
assign n_11059 = n_11045 ^ n_11015;
assign n_11060 = ~n_11047 & n_11044;
assign n_11061 = n_11047 ^ x381;
assign n_11062 = n_11048 & ~n_11046;
assign n_11063 = ~n_9863 & ~n_11048;
assign n_11064 = n_11049 ^ n_11035;
assign n_11065 = n_11050 & ~n_11051;
assign n_11066 = n_11052 ^ n_11038;
assign n_11067 = n_11053 ^ x2;
assign n_11068 = ~n_11028 & n_11054;
assign n_11069 = n_11054 ^ n_11028;
assign n_11070 = n_9662 & ~n_11055;
assign n_11071 = n_11057 ^ n_10179;
assign n_11072 = n_11057 ^ n_10356;
assign n_11073 = n_11058 ^ n_11015;
assign n_11074 = n_11030 & n_11059;
assign n_11075 = n_11060 ^ x381;
assign n_11076 = ~n_11061 & n_11034;
assign n_11077 = n_11034 ^ n_11061;
assign n_11078 = n_11062 ^ n_10508;
assign n_11079 = n_11063 ^ n_10508;
assign n_11080 = n_11065 ^ n_8942;
assign n_11081 = n_11066 ^ x1;
assign n_11082 = n_11067 ^ n_11066;
assign n_11083 = n_11070 ^ n_10316;
assign n_11084 = n_9685 & ~n_11071;
assign n_11085 = n_11071 ^ n_10356;
assign n_11086 = ~n_10369 & ~n_11072;
assign n_11087 = n_11073 ^ x380;
assign n_11088 = n_11074 ^ n_9270;
assign n_11089 = n_11075 ^ n_11073;
assign n_11090 = n_10531 ^ n_11077;
assign n_11091 = n_11078 ^ n_11077;
assign n_11092 = n_10531 ^ n_11078;
assign n_11093 = n_11080 ^ n_8987;
assign n_11094 = n_11079 ^ n_11080;
assign n_11095 = n_11082 & ~n_11081;
assign n_11096 = n_11082 ^ x1;
assign n_11097 = n_11083 ^ n_9310;
assign n_11098 = n_11084 ^ n_10356;
assign n_11099 = n_10717 ^ n_11085;
assign n_11100 = n_11086 ^ n_10179;
assign n_11101 = n_11088 ^ n_9310;
assign n_11102 = n_11088 ^ n_11083;
assign n_11103 = n_11089 & ~n_11087;
assign n_11104 = n_11089 ^ x380;
assign n_11105 = n_11091 & ~n_11090;
assign n_11106 = ~n_9878 & ~n_11091;
assign n_11107 = n_11092 ^ n_11077;
assign n_11108 = n_11079 ^ n_11093;
assign n_11109 = n_11093 & ~n_11094;
assign n_11110 = n_11095 ^ x1;
assign n_11111 = ~n_11068 & ~n_11096;
assign n_11112 = n_11096 ^ n_11068;
assign n_11113 = n_11098 ^ n_9350;
assign n_11114 = n_11100 ^ n_10394;
assign n_11115 = n_11101 ^ n_11083;
assign n_11116 = ~n_11097 & ~n_11102;
assign n_11117 = n_11103 ^ x380;
assign n_11118 = ~n_11076 & ~n_11104;
assign n_11119 = n_11104 ^ n_11076;
assign n_11120 = n_11105 ^ n_10531;
assign n_11121 = n_11106 ^ n_10531;
assign n_11122 = n_11108 ^ x0;
assign n_11123 = n_11109 ^ n_8987;
assign n_11124 = n_11110 ^ n_11108;
assign n_11125 = n_11114 ^ n_10200;
assign n_11126 = ~n_11114 & ~n_10410;
assign n_11127 = n_11115 ^ x379;
assign n_11128 = n_11116 ^ n_9310;
assign n_11129 = n_11117 ^ n_11115;
assign n_11130 = n_11119 ^ n_10548;
assign n_11131 = n_11120 ^ n_11119;
assign n_11132 = n_11120 ^ n_10548;
assign n_11133 = n_11121 ^ n_9026;
assign n_11134 = n_11123 ^ n_11121;
assign n_11135 = n_11123 ^ n_9026;
assign n_11136 = n_11124 & ~n_11122;
assign n_11137 = n_11124 ^ x0;
assign n_11138 = n_11125 ^ n_10394;
assign n_11139 = n_10738 ^ n_11125;
assign n_11140 = n_11126 ^ n_10200;
assign n_11141 = n_11128 ^ n_9350;
assign n_11142 = n_11128 ^ n_11098;
assign n_11143 = n_11129 ^ x379;
assign n_11144 = n_11129 & ~n_11127;
assign n_11145 = n_11131 & ~n_11130;
assign n_11146 = n_9898 & ~n_11131;
assign n_11147 = n_11132 ^ n_11119;
assign n_11148 = ~n_11133 & ~n_11134;
assign n_11149 = n_11135 ^ n_11121;
assign n_11150 = n_11136 ^ x0;
assign n_11151 = ~n_11111 & n_11137;
assign n_11152 = n_11137 ^ n_11111;
assign n_11153 = ~n_9705 & ~n_11138;
assign n_11154 = n_11140 ^ n_10450;
assign n_11155 = n_11141 ^ n_11098;
assign n_11156 = n_11113 & ~n_11142;
assign n_11157 = ~n_11143 & n_11118;
assign n_11158 = n_11118 ^ n_11143;
assign n_11159 = n_11144 ^ x379;
assign n_11160 = n_11145 ^ n_10548;
assign n_11161 = n_11146 ^ n_10548;
assign n_11162 = n_11148 ^ n_9026;
assign n_11163 = n_11149 ^ x15;
assign n_11164 = n_11150 ^ n_11149;
assign n_11165 = n_11153 ^ n_10394;
assign n_11166 = n_11154 ^ n_10435;
assign n_11167 = n_11155 ^ x378;
assign n_11168 = n_11156 ^ n_9350;
assign n_11169 = n_11158 ^ n_10562;
assign n_11170 = n_11159 ^ n_11155;
assign n_11171 = n_11160 ^ n_11158;
assign n_11172 = n_11160 ^ n_10562;
assign n_11173 = n_11161 ^ n_9068;
assign n_11174 = n_11162 ^ n_11161;
assign n_11175 = n_11162 ^ n_9068;
assign n_11176 = ~n_11164 & n_11163;
assign n_11177 = n_11164 ^ x15;
assign n_11178 = n_11165 ^ n_9391;
assign n_11179 = ~n_9730 & ~n_11166;
assign n_11180 = n_11168 ^ n_9391;
assign n_11181 = n_11165 ^ n_11168;
assign n_11182 = n_11170 ^ x378;
assign n_11183 = n_11170 & ~n_11167;
assign n_11184 = ~n_11171 & n_11169;
assign n_11185 = n_9918 & n_11171;
assign n_11186 = n_11172 ^ n_11158;
assign n_11187 = n_11173 & n_11174;
assign n_11188 = n_11175 ^ n_11161;
assign n_11189 = n_11176 ^ x15;
assign n_11190 = ~n_11177 & n_11151;
assign n_11191 = n_11151 ^ n_11177;
assign n_11192 = n_11179 ^ n_10435;
assign n_11193 = n_11165 ^ n_11180;
assign n_11194 = ~n_11178 & n_11181;
assign n_11195 = n_11157 ^ n_11182;
assign n_11196 = n_11182 & ~n_11157;
assign n_11197 = n_11183 ^ x378;
assign n_11198 = n_11184 ^ n_10562;
assign n_11199 = n_11185 ^ n_10562;
assign n_11200 = n_11187 ^ n_9068;
assign n_11201 = n_11188 ^ x14;
assign n_11202 = n_11189 ^ n_11188;
assign n_11203 = n_11192 ^ n_9429;
assign n_11204 = n_11193 ^ x377;
assign n_11205 = n_11194 ^ n_9391;
assign n_11206 = n_11195 ^ n_10578;
assign n_11207 = n_11197 ^ n_11193;
assign n_11208 = n_11195 ^ n_11198;
assign n_11209 = n_11198 ^ n_10578;
assign n_11210 = n_11200 ^ n_9110;
assign n_11211 = n_11199 ^ n_11200;
assign n_11212 = ~n_11202 & n_11201;
assign n_11213 = n_11202 ^ x14;
assign n_11214 = n_11205 ^ x376;
assign n_11215 = n_11207 ^ x377;
assign n_11216 = ~n_11207 & n_11204;
assign n_11217 = n_11208 & ~n_11206;
assign n_11218 = n_9938 & ~n_11208;
assign n_11219 = n_11195 ^ n_11209;
assign n_11220 = n_11199 ^ n_11210;
assign n_11221 = n_11210 & ~n_11211;
assign n_11222 = n_11212 ^ x14;
assign n_11223 = n_11190 & ~n_11213;
assign n_11224 = n_11213 ^ n_11190;
assign n_11225 = n_11214 ^ n_11203;
assign n_11226 = n_11196 ^ n_11215;
assign n_11227 = n_11215 & ~n_11196;
assign n_11228 = n_11216 ^ x377;
assign n_11229 = n_11217 ^ n_10578;
assign n_11230 = n_11218 ^ n_10578;
assign n_11231 = n_11220 ^ x13;
assign n_11232 = n_11221 ^ n_9110;
assign n_11233 = n_11222 ^ n_11220;
assign n_11234 = n_11226 ^ n_10596;
assign n_11235 = n_11228 ^ n_11225;
assign n_11236 = n_11229 ^ n_11226;
assign n_11237 = n_11229 ^ n_10596;
assign n_11238 = n_11232 ^ n_9154;
assign n_11239 = n_11230 ^ n_11232;
assign n_11240 = n_11233 & ~n_11231;
assign n_11241 = n_11233 ^ x13;
assign n_11242 = n_11235 ^ n_11227;
assign n_11243 = ~n_11236 & ~n_11234;
assign n_11244 = n_9959 & n_11236;
assign n_11245 = n_11237 ^ n_11226;
assign n_11246 = n_11230 ^ n_11238;
assign n_11247 = ~n_11238 & ~n_11239;
assign n_11248 = n_11240 ^ x13;
assign n_11249 = n_11223 & n_11241;
assign n_11250 = n_11241 ^ n_11223;
assign n_11251 = n_11242 ^ n_10616;
assign n_11252 = n_11243 ^ n_10596;
assign n_11253 = n_11244 ^ n_10596;
assign n_11254 = n_11246 ^ x12;
assign n_11255 = n_11247 ^ n_9154;
assign n_11256 = n_11248 ^ n_11246;
assign n_11257 = n_11252 ^ n_11242;
assign n_11258 = n_11252 ^ n_10616;
assign n_11259 = n_11253 ^ n_9196;
assign n_11260 = n_11253 ^ n_11255;
assign n_11261 = n_11255 ^ n_9196;
assign n_11262 = ~n_11256 & n_11254;
assign n_11263 = n_11256 ^ x12;
assign n_11264 = ~n_11257 & ~n_11251;
assign n_11265 = ~n_9980 & n_11257;
assign n_11266 = n_11258 ^ n_11242;
assign n_11267 = n_11259 & ~n_11260;
assign n_11268 = n_11253 ^ n_11261;
assign n_11269 = n_11262 ^ x12;
assign n_11270 = ~n_11249 & n_11263;
assign n_11271 = n_11264 ^ n_10616;
assign n_11272 = n_11265 ^ n_10616;
assign n_11273 = n_11267 ^ n_9196;
assign n_11274 = n_11269 ^ n_11268;
assign n_11275 = n_11269 ^ x11;
assign n_11276 = n_10641 ^ n_11271;
assign n_11277 = n_11271 ^ n_10294;
assign n_11278 = n_11272 ^ n_9236;
assign n_11279 = n_11272 ^ n_11273;
assign n_11280 = n_11273 ^ n_9236;
assign n_11281 = n_11274 ^ x11;
assign n_11282 = ~n_11274 & n_11275;
assign n_11283 = ~n_11277 & n_10641;
assign n_11284 = ~n_10001 & n_11277;
assign n_11285 = ~n_11278 & n_11279;
assign n_11286 = n_11272 ^ n_11280;
assign n_11287 = n_11281 & n_11270;
assign n_11288 = n_11270 ^ n_11281;
assign n_11289 = n_11282 ^ x11;
assign n_11290 = n_11283 ^ n_10635;
assign n_11291 = n_11284 ^ n_10635;
assign n_11292 = n_11285 ^ n_9236;
assign n_11293 = n_11286 ^ x10;
assign n_11294 = n_10788 & n_11288;
assign n_11295 = n_11288 ^ n_10788;
assign n_11296 = n_11289 ^ n_11286;
assign n_11297 = n_11290 ^ n_10651;
assign n_11298 = n_11292 ^ n_9277;
assign n_11299 = n_11292 ^ n_11291;
assign n_11300 = n_10814 ^ n_11294;
assign n_11301 = n_11295 ^ n_10780;
assign n_11302 = n_11296 & ~n_11293;
assign n_11303 = n_11296 ^ x10;
assign n_11304 = ~n_11297 & n_10660;
assign n_11305 = n_11297 ^ n_10346;
assign n_11306 = n_11298 ^ n_11291;
assign n_11307 = ~n_11298 & n_11299;
assign n_11308 = n_10248 & n_11301;
assign n_11309 = n_11302 ^ x10;
assign n_11310 = ~n_11303 & n_11287;
assign n_11311 = n_11287 ^ n_11303;
assign n_11312 = n_11304 ^ n_10346;
assign n_11313 = n_11305 ^ n_10651;
assign n_11314 = n_11306 ^ x9;
assign n_11315 = n_11307 ^ n_9277;
assign n_11316 = n_11308 ^ n_10780;
assign n_11317 = n_11309 ^ n_11306;
assign n_11318 = n_11311 ^ n_11294;
assign n_11319 = n_11300 ^ n_11311;
assign n_11320 = n_10681 ^ n_11312;
assign n_11321 = n_10397 ^ n_11312;
assign n_11322 = ~n_10022 & n_11313;
assign n_11323 = n_11315 ^ n_9317;
assign n_11324 = n_9711 & n_11316;
assign n_11325 = n_11316 ^ n_9711;
assign n_11326 = ~n_11317 & n_11314;
assign n_11327 = n_11317 ^ x9;
assign n_11328 = n_11318 & n_11300;
assign n_11329 = n_10278 & ~n_11318;
assign n_11330 = ~n_10687 & n_11320;
assign n_11331 = n_10681 ^ n_11321;
assign n_11332 = n_11322 ^ n_10651;
assign n_11333 = n_11324 ^ n_9734;
assign n_11334 = x167 & n_11325;
assign n_11335 = n_11325 ^ x167;
assign n_11336 = n_11326 ^ x9;
assign n_11337 = ~n_11327 & ~n_11310;
assign n_11338 = n_11310 ^ n_11327;
assign n_11339 = n_11328 ^ n_10814;
assign n_11340 = n_10814 ^ n_11329;
assign n_11341 = n_11330 ^ n_10397;
assign n_11342 = n_11331 ^ n_10672;
assign n_11343 = n_11332 ^ n_9317;
assign n_11344 = n_11332 ^ n_11315;
assign n_11345 = n_11332 ^ n_11323;
assign n_11346 = n_11334 ^ x166;
assign n_11347 = n_11336 ^ x8;
assign n_11348 = n_10862 ^ n_11338;
assign n_11349 = n_11339 ^ n_11338;
assign n_11350 = n_10862 ^ n_11339;
assign n_11351 = n_11340 ^ n_11324;
assign n_11352 = n_11341 ^ n_10701;
assign n_11353 = n_10437 ^ n_11341;
assign n_11354 = ~n_10045 & ~n_11342;
assign n_11355 = n_11343 & ~n_11344;
assign n_11356 = n_11336 ^ n_11345;
assign n_11357 = n_11349 & n_11348;
assign n_11358 = n_10318 & ~n_11349;
assign n_11359 = n_11350 ^ n_11338;
assign n_11360 = ~n_11351 & n_11333;
assign n_11361 = n_11351 ^ n_9734;
assign n_11362 = n_10707 & n_11352;
assign n_11363 = n_11353 ^ n_10701;
assign n_11364 = n_11354 ^ n_10672;
assign n_11365 = n_11355 ^ n_9317;
assign n_11366 = n_11356 & n_11347;
assign n_11367 = n_11356 ^ x8;
assign n_11368 = n_11357 ^ n_10862;
assign n_11369 = n_10862 ^ n_11358;
assign n_11370 = n_11360 ^ n_9734;
assign n_11371 = n_11361 ^ n_11334;
assign n_11372 = n_11362 ^ n_10437;
assign n_11373 = n_11363 ^ n_10693;
assign n_11374 = n_11364 ^ n_9359;
assign n_11375 = n_11365 ^ n_11364;
assign n_11376 = n_11366 ^ x8;
assign n_11377 = n_11367 & n_11337;
assign n_11378 = n_11337 ^ n_11367;
assign n_11379 = n_10900 ^ n_11368;
assign n_11380 = n_11369 ^ n_9770;
assign n_11381 = n_11369 ^ n_11370;
assign n_11382 = n_11370 ^ n_9770;
assign n_11383 = ~n_11371 & n_11346;
assign n_11384 = n_11371 ^ x166;
assign n_11385 = n_11372 ^ n_10719;
assign n_11386 = ~n_10066 & n_11373;
assign n_11387 = ~n_11375 & ~n_11374;
assign n_11388 = n_11375 ^ n_9359;
assign n_11389 = n_11376 ^ x23;
assign n_11390 = n_11368 ^ n_11378;
assign n_11391 = n_10900 ^ n_11378;
assign n_11392 = n_11379 ^ n_11378;
assign n_11393 = n_11380 & n_11381;
assign n_11394 = n_11369 ^ n_11382;
assign n_11395 = n_11383 ^ x166;
assign n_11396 = n_11335 & n_11384;
assign n_11397 = n_11384 ^ n_11335;
assign n_11398 = ~n_11385 & ~n_10727;
assign n_11399 = n_11385 ^ n_10475;
assign n_11400 = n_11386 ^ n_10693;
assign n_11401 = n_11387 ^ n_9359;
assign n_11402 = n_11388 ^ x23;
assign n_11403 = n_11388 ^ n_11376;
assign n_11404 = n_11388 ^ n_11389;
assign n_11405 = ~n_10360 & n_11390;
assign n_11406 = ~n_11390 & ~n_11391;
assign n_11407 = n_11393 ^ n_9770;
assign n_11408 = n_11394 ^ x165;
assign n_11409 = n_11395 ^ n_11394;
assign n_11410 = n_11398 ^ n_10475;
assign n_11411 = n_11399 ^ n_10719;
assign n_11412 = n_11400 ^ n_9398;
assign n_11413 = n_11400 ^ n_11401;
assign n_11414 = n_11401 ^ n_9398;
assign n_11415 = n_11402 & ~n_11403;
assign n_11416 = n_11404 & ~n_11377;
assign n_11417 = n_11377 ^ n_11404;
assign n_11418 = n_10900 ^ n_11405;
assign n_11419 = n_11406 ^ n_10900;
assign n_11420 = n_11407 ^ n_9796;
assign n_11421 = ~n_11409 & n_11408;
assign n_11422 = n_11409 ^ x165;
assign n_11423 = n_11410 ^ n_10740;
assign n_11424 = ~n_10085 & ~n_11411;
assign n_11425 = ~n_11412 & n_11413;
assign n_11426 = n_11400 ^ n_11414;
assign n_11427 = n_11415 ^ x23;
assign n_11428 = n_10939 ^ n_11417;
assign n_11429 = n_11418 ^ n_9796;
assign n_11430 = n_11418 ^ n_11407;
assign n_11431 = n_11419 ^ n_11417;
assign n_11432 = n_10939 ^ n_11419;
assign n_11433 = n_11418 ^ n_11420;
assign n_11434 = n_11421 ^ x165;
assign n_11435 = ~n_11396 & ~n_11422;
assign n_11436 = n_11422 ^ n_11396;
assign n_11437 = n_11423 & ~n_10747;
assign n_11438 = n_10505 ^ n_11423;
assign n_11439 = n_11424 ^ n_10719;
assign n_11440 = n_11425 ^ n_9398;
assign n_11441 = n_11426 ^ x22;
assign n_11442 = n_11427 ^ n_11426;
assign n_11443 = n_11429 & n_11430;
assign n_11444 = n_11431 & n_11428;
assign n_11445 = ~n_10401 & ~n_11431;
assign n_11446 = n_11432 ^ n_11417;
assign n_11447 = n_11433 ^ x164;
assign n_11448 = n_11434 ^ n_11433;
assign n_11449 = n_11437 ^ n_10505;
assign n_11450 = n_11438 ^ n_10740;
assign n_11451 = n_11439 ^ n_9435;
assign n_11452 = n_11439 ^ n_11440;
assign n_11453 = n_11440 ^ n_9435;
assign n_11454 = n_11442 & ~n_11441;
assign n_11455 = n_11442 ^ x22;
assign n_11456 = n_11443 ^ n_9796;
assign n_11457 = n_11444 ^ n_10939;
assign n_11458 = n_10939 ^ n_11445;
assign n_11459 = n_11448 & ~n_11447;
assign n_11460 = n_11448 ^ x164;
assign n_11461 = n_11449 ^ n_10761;
assign n_11462 = ~n_10105 & n_11450;
assign n_11463 = n_11451 & ~n_11452;
assign n_11464 = n_11439 ^ n_11453;
assign n_11465 = n_11454 ^ x22;
assign n_11466 = n_11455 & ~n_11416;
assign n_11467 = n_11416 ^ n_11455;
assign n_11468 = n_11456 ^ n_9818;
assign n_11469 = n_10980 ^ n_11457;
assign n_11470 = n_11458 ^ n_9818;
assign n_11471 = n_11458 ^ n_11456;
assign n_11472 = n_11459 ^ x164;
assign n_11473 = n_11435 & n_11460;
assign n_11474 = n_11460 ^ n_11435;
assign n_11475 = n_11461 & n_10768;
assign n_11476 = n_10526 ^ n_11461;
assign n_11477 = n_11462 ^ n_10740;
assign n_11478 = n_11463 ^ n_9435;
assign n_11479 = n_11464 ^ x21;
assign n_11480 = n_11465 ^ n_11464;
assign n_11481 = n_11467 ^ n_11457;
assign n_11482 = n_10980 ^ n_11467;
assign n_11483 = n_11458 ^ n_11468;
assign n_11484 = n_11469 ^ n_11467;
assign n_11485 = n_11470 & n_11471;
assign n_11486 = n_11475 ^ n_10526;
assign n_11487 = n_11476 ^ n_10761;
assign n_11488 = n_10839 ^ n_11476;
assign n_11489 = n_11477 ^ n_9466;
assign n_11490 = n_11478 ^ n_11477;
assign n_11491 = n_11478 ^ n_9466;
assign n_11492 = ~n_11480 & n_11479;
assign n_11493 = n_11480 ^ x21;
assign n_11494 = ~n_10440 & ~n_11481;
assign n_11495 = n_11481 & n_11482;
assign n_11496 = n_11472 ^ n_11483;
assign n_11497 = n_11483 ^ x163;
assign n_11498 = n_11484 ^ n_11335;
assign n_11499 = n_11485 ^ n_9818;
assign n_11500 = n_11486 ^ n_10782;
assign n_11501 = n_10126 & ~n_11487;
assign n_11502 = ~n_11489 & ~n_11490;
assign n_11503 = n_11491 ^ n_11477;
assign n_11504 = n_11492 ^ x21;
assign n_11505 = ~n_11493 & n_11466;
assign n_11506 = n_11466 ^ n_11493;
assign n_11507 = n_10980 ^ n_11494;
assign n_11508 = n_11495 ^ n_10980;
assign n_11509 = n_11496 ^ x163;
assign n_11510 = ~n_11496 & n_11497;
assign n_11511 = n_11499 ^ n_9832;
assign n_11512 = n_11500 & n_10791;
assign n_11513 = n_10545 ^ n_11500;
assign n_11514 = n_11501 ^ n_10761;
assign n_11515 = n_11502 ^ n_9466;
assign n_11516 = n_11503 ^ x20;
assign n_11517 = n_11504 ^ n_11503;
assign n_11518 = n_11024 ^ n_11506;
assign n_11519 = n_11507 ^ n_9832;
assign n_11520 = n_11507 ^ n_11499;
assign n_11521 = n_11508 ^ n_11506;
assign n_11522 = n_11024 ^ n_11508;
assign n_11523 = n_11473 & ~n_11509;
assign n_11524 = n_11509 ^ n_11473;
assign n_11525 = n_11510 ^ x163;
assign n_11526 = n_11507 ^ n_11511;
assign n_11527 = n_11512 ^ n_10545;
assign n_11528 = n_11513 ^ n_10782;
assign n_11529 = n_11513 ^ n_10865;
assign n_11530 = n_11514 ^ n_9496;
assign n_11531 = n_11515 ^ n_11514;
assign n_11532 = n_11515 ^ n_9496;
assign n_11533 = n_11517 & ~n_11516;
assign n_11534 = n_11517 ^ x20;
assign n_11535 = n_11519 & n_11520;
assign n_11536 = ~n_11521 & n_11518;
assign n_11537 = ~n_10478 & n_11521;
assign n_11538 = n_11522 ^ n_11506;
assign n_11539 = n_11525 ^ n_11526;
assign n_11540 = n_11526 ^ x162;
assign n_11541 = n_11527 ^ n_10808;
assign n_11542 = ~n_10147 & ~n_11528;
assign n_11543 = n_11530 & n_11531;
assign n_11544 = n_11532 ^ n_11514;
assign n_11545 = n_11533 ^ x20;
assign n_11546 = ~n_11505 & ~n_11534;
assign n_11547 = n_11534 ^ n_11505;
assign n_11548 = n_11535 ^ n_9832;
assign n_11549 = n_11536 ^ n_11024;
assign n_11550 = n_11024 ^ n_11537;
assign n_11551 = n_11397 ^ n_11538;
assign n_11552 = n_11539 ^ x162;
assign n_11553 = n_11539 & ~n_11540;
assign n_11554 = n_11541 & ~n_10818;
assign n_11555 = n_10565 ^ n_11541;
assign n_11556 = n_11542 ^ n_10782;
assign n_11557 = n_11543 ^ n_9496;
assign n_11558 = n_11544 ^ x19;
assign n_11559 = n_11545 ^ n_11544;
assign n_11560 = n_11064 ^ n_11547;
assign n_11561 = n_11548 ^ n_9850;
assign n_11562 = n_11549 ^ n_11547;
assign n_11563 = n_11064 ^ n_11549;
assign n_11564 = n_11550 ^ n_9850;
assign n_11565 = n_11550 ^ n_11548;
assign n_11566 = ~n_11523 & ~n_11552;
assign n_11567 = n_11552 ^ n_11523;
assign n_11568 = n_11553 ^ x162;
assign n_11569 = n_11554 ^ n_10565;
assign n_11570 = n_11555 ^ n_10808;
assign n_11571 = n_10943 ^ n_11555;
assign n_11572 = n_11556 ^ n_9521;
assign n_11573 = n_11557 ^ n_11556;
assign n_11574 = n_11557 ^ n_9521;
assign n_11575 = n_11559 & ~n_11558;
assign n_11576 = n_11559 ^ x19;
assign n_11577 = n_11550 ^ n_11561;
assign n_11578 = ~n_11562 & n_11560;
assign n_11579 = ~n_10508 & n_11562;
assign n_11580 = n_11563 ^ n_11547;
assign n_11581 = ~n_11564 & ~n_11565;
assign n_11582 = n_11569 ^ n_10840;
assign n_11583 = ~n_10168 & n_11570;
assign n_11584 = ~n_11572 & n_11573;
assign n_11585 = n_11574 ^ n_11556;
assign n_11586 = n_11575 ^ x19;
assign n_11587 = ~n_11546 & n_11576;
assign n_11588 = n_11576 ^ n_11546;
assign n_11589 = n_11568 ^ n_11577;
assign n_11590 = n_11577 ^ x161;
assign n_11591 = n_11578 ^ n_11064;
assign n_11592 = n_11579 ^ n_11064;
assign n_11593 = n_11436 ^ n_11580;
assign n_11594 = n_11581 ^ n_9850;
assign n_11595 = n_10589 ^ n_11582;
assign n_11596 = n_11582 & ~n_10853;
assign n_11597 = n_11583 ^ n_10808;
assign n_11598 = n_11584 ^ n_9521;
assign n_11599 = n_11585 ^ x18;
assign n_11600 = n_11586 ^ n_11585;
assign n_11601 = n_11107 ^ n_11588;
assign n_11602 = n_11589 ^ x161;
assign n_11603 = n_11589 & ~n_11590;
assign n_11604 = n_11591 ^ n_11588;
assign n_11605 = n_11107 ^ n_11591;
assign n_11606 = n_11592 ^ n_9863;
assign n_11607 = n_11594 ^ n_11592;
assign n_11608 = n_11594 ^ n_9863;
assign n_11609 = n_11595 ^ n_10840;
assign n_11610 = n_10985 ^ n_11595;
assign n_11611 = n_11596 ^ n_10589;
assign n_11612 = n_11597 ^ n_9536;
assign n_11613 = n_11598 ^ n_11597;
assign n_11614 = n_11598 ^ n_9536;
assign n_11615 = n_11600 & ~n_11599;
assign n_11616 = n_11600 ^ x18;
assign n_11617 = ~n_11566 & n_11602;
assign n_11618 = n_11602 ^ n_11566;
assign n_11619 = n_11603 ^ x161;
assign n_11620 = ~n_11604 & n_11601;
assign n_11621 = ~n_10531 & n_11604;
assign n_11622 = n_11605 ^ n_11588;
assign n_11623 = ~n_11606 & n_11607;
assign n_11624 = n_11608 ^ n_11592;
assign n_11625 = ~n_10189 & n_11609;
assign n_11626 = n_11611 ^ n_10892;
assign n_11627 = n_11611 ^ n_10878;
assign n_11628 = n_11612 & ~n_11613;
assign n_11629 = n_11614 ^ n_11597;
assign n_11630 = n_11615 ^ x18;
assign n_11631 = n_11616 & n_11587;
assign n_11632 = n_11587 ^ n_11616;
assign n_11633 = n_11620 ^ n_11107;
assign n_11634 = n_11621 ^ n_11107;
assign n_11635 = n_11474 ^ n_11622;
assign n_11636 = n_11623 ^ n_9863;
assign n_11637 = n_11619 ^ n_11624;
assign n_11638 = n_11624 ^ x160;
assign n_11639 = n_11625 ^ n_10840;
assign n_11640 = n_11626 ^ n_10878;
assign n_11641 = n_11626 ^ n_11029;
assign n_11642 = ~n_10892 & ~n_11627;
assign n_11643 = n_11628 ^ n_9536;
assign n_11644 = n_11629 ^ x17;
assign n_11645 = n_11630 ^ n_11629;
assign n_11646 = n_11147 ^ n_11632;
assign n_11647 = n_11633 ^ n_11632;
assign n_11648 = n_11147 ^ n_11633;
assign n_11649 = n_11634 ^ n_9878;
assign n_11650 = n_11636 ^ n_11634;
assign n_11651 = n_11636 ^ n_9878;
assign n_11652 = n_11637 ^ x160;
assign n_11653 = ~n_11637 & n_11638;
assign n_11654 = n_11639 ^ n_9561;
assign n_11655 = n_10212 & ~n_11640;
assign n_11656 = n_11642 ^ n_10613;
assign n_11657 = n_11643 ^ n_11639;
assign n_11658 = n_11643 ^ n_9561;
assign n_11659 = ~n_11645 & n_11644;
assign n_11660 = n_11645 ^ x17;
assign n_11661 = n_11647 & ~n_11646;
assign n_11662 = ~n_10548 & ~n_11647;
assign n_11663 = n_11648 ^ n_11632;
assign n_11664 = ~n_11649 & n_11650;
assign n_11665 = n_11651 ^ n_11634;
assign n_11666 = ~n_11617 & n_11652;
assign n_11667 = n_11652 ^ n_11617;
assign n_11668 = n_11653 ^ x160;
assign n_11669 = n_11655 ^ n_10878;
assign n_11670 = n_11656 ^ n_10634;
assign n_11671 = n_11656 ^ n_10918;
assign n_11672 = ~n_11654 & ~n_11657;
assign n_11673 = n_11658 ^ n_11639;
assign n_11674 = n_11659 ^ x17;
assign n_11675 = ~n_11631 & n_11660;
assign n_11676 = n_11660 ^ n_11631;
assign n_11677 = n_11661 ^ n_11147;
assign n_11678 = n_11662 ^ n_11147;
assign n_11679 = n_11524 ^ n_11663;
assign n_11680 = n_11664 ^ n_9878;
assign n_11681 = n_11665 ^ x175;
assign n_11682 = n_11668 ^ n_11665;
assign n_11683 = n_11669 ^ n_9580;
assign n_11684 = n_11670 ^ n_10918;
assign n_11685 = n_10932 & n_11671;
assign n_11686 = n_11672 ^ n_9561;
assign n_11687 = n_11673 ^ x16;
assign n_11688 = n_11674 ^ n_11673;
assign n_11689 = n_11186 ^ n_11676;
assign n_11690 = n_11677 ^ n_11676;
assign n_11691 = n_11186 ^ n_11677;
assign n_11692 = n_11678 ^ n_9898;
assign n_11693 = n_11680 ^ n_11678;
assign n_11694 = n_11680 ^ n_9898;
assign n_11695 = ~n_11682 & n_11681;
assign n_11696 = n_11682 ^ x175;
assign n_11697 = n_11684 ^ n_10904;
assign n_11698 = n_11684 ^ n_11069;
assign n_11699 = n_11685 ^ n_10634;
assign n_11700 = n_11686 ^ n_11669;
assign n_11701 = n_11688 & ~n_11687;
assign n_11702 = n_11688 ^ x16;
assign n_11703 = n_11690 & n_11689;
assign n_11704 = ~n_10562 & ~n_11690;
assign n_11705 = n_11691 ^ n_11676;
assign n_11706 = n_11692 & n_11693;
assign n_11707 = n_11694 ^ n_11678;
assign n_11708 = n_11695 ^ x175;
assign n_11709 = n_11666 & n_11696;
assign n_11710 = n_11696 ^ n_11666;
assign n_11711 = n_10232 & ~n_11697;
assign n_11712 = n_11699 ^ n_10957;
assign n_11713 = n_11700 ^ n_9580;
assign n_11714 = ~n_11700 & ~n_11683;
assign n_11715 = n_11701 ^ x16;
assign n_11716 = ~n_11675 & n_11702;
assign n_11717 = n_11702 ^ n_11675;
assign n_11718 = n_11703 ^ n_11186;
assign n_11719 = n_11704 ^ n_11186;
assign n_11720 = n_11567 ^ n_11705;
assign n_11721 = n_11706 ^ n_9898;
assign n_11722 = n_11707 ^ x174;
assign n_11723 = n_11708 ^ n_11707;
assign n_11724 = n_11711 ^ n_10904;
assign n_11725 = n_10656 ^ n_11712;
assign n_11726 = n_11712 & n_10972;
assign n_11727 = n_11713 ^ x31;
assign n_11728 = n_11714 ^ n_9580;
assign n_11729 = n_11715 ^ n_11713;
assign n_11730 = n_11715 ^ x31;
assign n_11731 = n_11717 ^ n_11219;
assign n_11732 = n_11717 ^ n_11718;
assign n_11733 = n_11718 ^ n_11219;
assign n_11734 = n_11719 ^ n_9918;
assign n_11735 = n_11721 ^ n_11719;
assign n_11736 = n_11721 ^ n_9918;
assign n_11737 = n_11723 & ~n_11722;
assign n_11738 = n_11723 ^ x174;
assign n_11739 = n_11724 ^ n_9600;
assign n_11740 = n_11725 ^ n_10957;
assign n_11741 = n_11725 ^ n_11112;
assign n_11742 = n_11726 ^ n_10656;
assign n_11743 = n_11728 ^ n_9600;
assign n_11744 = n_11728 ^ n_11724;
assign n_11745 = n_11727 & ~n_11729;
assign n_11746 = n_11730 ^ n_11713;
assign n_11747 = n_11732 & n_11731;
assign n_11748 = ~n_10578 & ~n_11732;
assign n_11749 = n_11733 ^ n_11717;
assign n_11750 = ~n_11734 & n_11735;
assign n_11751 = n_11736 ^ n_11719;
assign n_11752 = n_11737 ^ x174;
assign n_11753 = n_11709 & ~n_11738;
assign n_11754 = n_11738 ^ n_11709;
assign n_11755 = ~n_10256 & ~n_11740;
assign n_11756 = n_11001 ^ n_11742;
assign n_11757 = n_11743 ^ n_11724;
assign n_11758 = n_11739 & n_11744;
assign n_11759 = n_11745 ^ x31;
assign n_11760 = n_11716 & ~n_11746;
assign n_11761 = n_11746 ^ n_11716;
assign n_11762 = n_11747 ^ n_11219;
assign n_11763 = n_11748 ^ n_11219;
assign n_11764 = n_11749 ^ n_11618;
assign n_11765 = n_11750 ^ n_9918;
assign n_11766 = n_11751 ^ x173;
assign n_11767 = n_11752 ^ n_11751;
assign n_11768 = n_11755 ^ n_10957;
assign n_11769 = n_10678 ^ n_11756;
assign n_11770 = n_11756 & ~n_11016;
assign n_11771 = n_11757 ^ x30;
assign n_11772 = n_11758 ^ n_9600;
assign n_11773 = n_11759 ^ n_11757;
assign n_11774 = n_11245 ^ n_11761;
assign n_11775 = n_11762 ^ n_11761;
assign n_11776 = n_11763 ^ n_9938;
assign n_11777 = n_11765 ^ n_9938;
assign n_11778 = n_11765 ^ n_11763;
assign n_11779 = n_11767 & ~n_11766;
assign n_11780 = n_11767 ^ x173;
assign n_11781 = n_11768 ^ n_9620;
assign n_11782 = n_11769 ^ n_10987;
assign n_11783 = n_11152 ^ n_11769;
assign n_11784 = n_11770 ^ n_10678;
assign n_11785 = n_11772 ^ n_11768;
assign n_11786 = n_11773 ^ x30;
assign n_11787 = ~n_11773 & n_11771;
assign n_11788 = ~n_11775 & n_11774;
assign n_11789 = n_10596 & n_11775;
assign n_11790 = n_11245 ^ n_11775;
assign n_11791 = n_11777 ^ n_11763;
assign n_11792 = n_11776 & ~n_11778;
assign n_11793 = n_11779 ^ x173;
assign n_11794 = n_11753 & ~n_11780;
assign n_11795 = n_11780 ^ n_11753;
assign n_11796 = n_10282 & n_11782;
assign n_11797 = n_11784 ^ n_11042;
assign n_11798 = n_11785 ^ n_9620;
assign n_11799 = n_11785 & ~n_11781;
assign n_11800 = n_11786 & ~n_11760;
assign n_11801 = n_11760 ^ n_11786;
assign n_11802 = n_11787 ^ x30;
assign n_11803 = n_11788 ^ n_11245;
assign n_11804 = n_11789 ^ n_11245;
assign n_11805 = n_11790 ^ n_11667;
assign n_11806 = n_11791 ^ x172;
assign n_11807 = n_11792 ^ n_9938;
assign n_11808 = n_11793 ^ n_11791;
assign n_11809 = n_11793 ^ x172;
assign n_11810 = n_11796 ^ n_10987;
assign n_11811 = n_10698 ^ n_11797;
assign n_11812 = n_11797 & n_11056;
assign n_11813 = n_11798 ^ x29;
assign n_11814 = n_11799 ^ n_9620;
assign n_11815 = n_11266 ^ n_11801;
assign n_11816 = n_11802 ^ n_11798;
assign n_11817 = n_11803 ^ n_11801;
assign n_11818 = n_11803 ^ n_11266;
assign n_11819 = n_11804 ^ n_9959;
assign n_11820 = n_11807 ^ n_9959;
assign n_11821 = n_11807 ^ n_11804;
assign n_11822 = n_11806 & ~n_11808;
assign n_11823 = n_11809 ^ n_11791;
assign n_11824 = n_11810 ^ n_9641;
assign n_11825 = n_11811 ^ n_11042;
assign n_11826 = n_11191 ^ n_11811;
assign n_11827 = n_11812 ^ n_10698;
assign n_11828 = n_11814 ^ n_9641;
assign n_11829 = n_11814 ^ n_11810;
assign n_11830 = n_11816 ^ x29;
assign n_11831 = ~n_11816 & n_11813;
assign n_11832 = n_11815 & n_11817;
assign n_11833 = ~n_10616 & ~n_11817;
assign n_11834 = n_11818 ^ n_11801;
assign n_11835 = n_11820 ^ n_11804;
assign n_11836 = n_11819 & ~n_11821;
assign n_11837 = n_11822 ^ x172;
assign n_11838 = n_11794 & n_11823;
assign n_11839 = n_11823 ^ n_11794;
assign n_11840 = n_10316 & ~n_11825;
assign n_11841 = n_11085 ^ n_11827;
assign n_11842 = n_11828 ^ n_11810;
assign n_11843 = n_11824 & ~n_11829;
assign n_11844 = n_11800 ^ n_11830;
assign n_11845 = n_11830 & n_11800;
assign n_11846 = n_11831 ^ x29;
assign n_11847 = n_11832 ^ n_11266;
assign n_11848 = n_11833 ^ n_11266;
assign n_11849 = n_11834 ^ n_11710;
assign n_11850 = n_11835 ^ x171;
assign n_11851 = n_11836 ^ n_9959;
assign n_11852 = n_11837 ^ n_11835;
assign n_11853 = n_11840 ^ n_11042;
assign n_11854 = n_10717 ^ n_11841;
assign n_11855 = n_11841 & ~n_11099;
assign n_11856 = n_11842 ^ x28;
assign n_11857 = n_11843 ^ n_9641;
assign n_11858 = n_11276 ^ n_11844;
assign n_11859 = n_11846 ^ n_11842;
assign n_11860 = n_11847 ^ n_11844;
assign n_11861 = n_11847 ^ n_11276;
assign n_11862 = n_11848 ^ n_9980;
assign n_11863 = n_11851 ^ n_9980;
assign n_11864 = n_11851 ^ n_11848;
assign n_11865 = ~n_11852 & n_11850;
assign n_11866 = n_11852 ^ x171;
assign n_11867 = n_11853 ^ n_9662;
assign n_11868 = n_11854 ^ n_11071;
assign n_11869 = n_11224 ^ n_11854;
assign n_11870 = n_11855 ^ n_10717;
assign n_11871 = n_11857 ^ n_9662;
assign n_11872 = n_11857 ^ n_11853;
assign n_11873 = n_11859 ^ x28;
assign n_11874 = n_11859 & ~n_11856;
assign n_11875 = ~n_11858 & n_11860;
assign n_11876 = ~n_10635 & ~n_11860;
assign n_11877 = n_11861 ^ n_11844;
assign n_11878 = n_11863 ^ n_11848;
assign n_11879 = n_11862 & n_11864;
assign n_11880 = n_11865 ^ x171;
assign n_11881 = ~n_11838 & ~n_11866;
assign n_11882 = n_11866 ^ n_11838;
assign n_11883 = ~n_10356 & ~n_11868;
assign n_11884 = n_11870 ^ n_11125;
assign n_11885 = n_11871 ^ n_11853;
assign n_11886 = ~n_11867 & ~n_11872;
assign n_11887 = n_11845 ^ n_11873;
assign n_11888 = n_11873 & ~n_11845;
assign n_11889 = n_11874 ^ x28;
assign n_11890 = n_11875 ^ n_11276;
assign n_11891 = n_11876 ^ n_11276;
assign n_11892 = n_11877 ^ n_11754;
assign n_11893 = n_11878 ^ x170;
assign n_11894 = n_11879 ^ n_9980;
assign n_11895 = n_11880 ^ n_11878;
assign n_11896 = n_11883 ^ n_11071;
assign n_11897 = n_10738 ^ n_11884;
assign n_11898 = ~n_11884 & ~n_11139;
assign n_11899 = n_11885 ^ x27;
assign n_11900 = n_11886 ^ n_9662;
assign n_11901 = n_11887 ^ n_11305;
assign n_11902 = n_11889 ^ n_11885;
assign n_11903 = n_11890 ^ n_11305;
assign n_11904 = n_11890 ^ n_11887;
assign n_11905 = n_11891 ^ n_10001;
assign n_11906 = n_11894 ^ n_10001;
assign n_11907 = n_11894 ^ n_11891;
assign n_11908 = ~n_11895 & n_11893;
assign n_11909 = n_11895 ^ x170;
assign n_11910 = n_11896 ^ n_9685;
assign n_11911 = n_11897 ^ n_11125;
assign n_11912 = n_11250 ^ n_11897;
assign n_11913 = n_11898 ^ n_10738;
assign n_11914 = n_11900 ^ n_9685;
assign n_11915 = n_11900 ^ n_11896;
assign n_11916 = n_11902 ^ x27;
assign n_11917 = ~n_11902 & n_11899;
assign n_11918 = n_11903 ^ n_11887;
assign n_11919 = ~n_10651 & ~n_11904;
assign n_11920 = n_11904 & ~n_11901;
assign n_11921 = n_11906 ^ n_11891;
assign n_11922 = n_11905 & ~n_11907;
assign n_11923 = n_11908 ^ x170;
assign n_11924 = ~n_11881 & n_11909;
assign n_11925 = n_11909 ^ n_11881;
assign n_11926 = n_10394 & ~n_11911;
assign n_11927 = n_11913 ^ n_11154;
assign n_11928 = n_11914 ^ n_11896;
assign n_11929 = ~n_11910 & n_11915;
assign n_11930 = n_11916 ^ n_11888;
assign n_11931 = ~n_11888 & n_11916;
assign n_11932 = n_11917 ^ x27;
assign n_11933 = n_11795 ^ n_11918;
assign n_11934 = n_11919 ^ n_11305;
assign n_11935 = n_11920 ^ n_11305;
assign n_11936 = n_11921 ^ x169;
assign n_11937 = n_11922 ^ n_10001;
assign n_11938 = n_11923 ^ n_11921;
assign n_11939 = n_11926 ^ n_11125;
assign n_11940 = n_11927 ^ n_10759;
assign n_11941 = n_11928 ^ x26;
assign n_11942 = n_11929 ^ n_9685;
assign n_11943 = n_11930 ^ n_11331;
assign n_11944 = n_11932 ^ n_11928;
assign n_11945 = n_11934 ^ n_10022;
assign n_11946 = n_11935 ^ n_11930;
assign n_11947 = n_11937 ^ n_10022;
assign n_11948 = n_11937 ^ n_11934;
assign n_11949 = n_11938 & ~n_11936;
assign n_11950 = n_11938 ^ x169;
assign n_11951 = n_11939 ^ n_9705;
assign n_11952 = n_11940 ^ n_11154;
assign n_11953 = n_11940 ^ n_11249;
assign n_11954 = n_11942 ^ n_9705;
assign n_11955 = n_11939 ^ n_11942;
assign n_11956 = n_11935 ^ n_11943;
assign n_11957 = n_11944 ^ x26;
assign n_11958 = n_11944 & ~n_11941;
assign n_11959 = ~n_11943 & ~n_11946;
assign n_11960 = n_11947 ^ n_11934;
assign n_11961 = n_11945 & ~n_11948;
assign n_11962 = n_11949 ^ x169;
assign n_11963 = n_11924 & ~n_11950;
assign n_11964 = n_11950 ^ n_11924;
assign n_11965 = ~n_10435 & ~n_11952;
assign n_11966 = n_11953 ^ n_11263;
assign n_11967 = n_11939 ^ n_11954;
assign n_11968 = n_11951 & n_11955;
assign n_11969 = n_11956 ^ n_11321;
assign n_11970 = n_11839 ^ n_11956;
assign n_11971 = n_11931 ^ n_11957;
assign n_11972 = n_11957 & ~n_11931;
assign n_11973 = n_11958 ^ x26;
assign n_11974 = n_11959 ^ n_11331;
assign n_11975 = n_11960 ^ x168;
assign n_11976 = n_11961 ^ n_10022;
assign n_11977 = n_11962 ^ n_11960;
assign n_11978 = n_11965 ^ n_11154;
assign n_11979 = n_11967 ^ x25;
assign n_11980 = n_11968 ^ n_9705;
assign n_11981 = n_10681 & n_11969;
assign n_11982 = n_11971 ^ n_11363;
assign n_11983 = n_11973 ^ n_11967;
assign n_11984 = n_11974 ^ n_11363;
assign n_11985 = n_11974 ^ n_11971;
assign n_11986 = n_11977 & ~n_11975;
assign n_11987 = n_11977 ^ x168;
assign n_11988 = n_11978 ^ n_9730;
assign n_11989 = n_11980 ^ x24;
assign n_11990 = n_11981 ^ n_11321;
assign n_11991 = n_11983 ^ x25;
assign n_11992 = ~n_11983 & n_11979;
assign n_11993 = n_11984 ^ n_11971;
assign n_11994 = ~n_11982 & ~n_11985;
assign n_11995 = n_11986 ^ x168;
assign n_11996 = n_11963 & ~n_11987;
assign n_11997 = n_11987 ^ n_11963;
assign n_11998 = n_11989 ^ n_11988;
assign n_11999 = n_11976 ^ n_11990;
assign n_12000 = n_11990 ^ n_10045;
assign n_12001 = n_11991 ^ n_11972;
assign n_12002 = n_11972 & ~n_11991;
assign n_12003 = n_11992 ^ x25;
assign n_12004 = n_11993 ^ n_11353;
assign n_12005 = n_11882 ^ n_11993;
assign n_12006 = n_11994 ^ n_11363;
assign n_12007 = n_11995 ^ x183;
assign n_12008 = n_11999 ^ n_10045;
assign n_12009 = n_11999 & ~n_12000;
assign n_12010 = n_12001 ^ n_11399;
assign n_12011 = n_12003 ^ n_11998;
assign n_12012 = n_10701 & n_12004;
assign n_12013 = n_12006 ^ n_12001;
assign n_12014 = n_12006 ^ n_11399;
assign n_12015 = n_12007 ^ n_12008;
assign n_12016 = n_12008 ^ x183;
assign n_12017 = n_11995 ^ n_12008;
assign n_12018 = n_12009 ^ n_10045;
assign n_12019 = n_12011 ^ n_12002;
assign n_12020 = n_12012 ^ n_11353;
assign n_12021 = n_10719 & ~n_12013;
assign n_12022 = n_12013 & ~n_12010;
assign n_12023 = n_12014 ^ n_12001;
assign n_12024 = ~n_12015 & ~n_11996;
assign n_12025 = n_11996 ^ n_12015;
assign n_12026 = n_12016 & ~n_12017;
assign n_12027 = n_12018 ^ n_10066;
assign n_12028 = n_12019 ^ n_11438;
assign n_12029 = n_12020 ^ n_10066;
assign n_12030 = n_12018 ^ n_12020;
assign n_12031 = n_12021 ^ n_11399;
assign n_12032 = n_12022 ^ n_11399;
assign n_12033 = n_11925 ^ n_12023;
assign n_12034 = n_12026 ^ x183;
assign n_12035 = n_12027 ^ n_12020;
assign n_12036 = n_12029 & ~n_12030;
assign n_12037 = n_12031 ^ n_10085;
assign n_12038 = n_12032 ^ n_12019;
assign n_12039 = n_12032 ^ n_11438;
assign n_12040 = n_12034 ^ n_12035;
assign n_12041 = n_12035 ^ x182;
assign n_12042 = n_12036 ^ n_10066;
assign n_12043 = n_10740 & ~n_12038;
assign n_12044 = n_12038 & n_12028;
assign n_12045 = n_12039 ^ n_12019;
assign n_12046 = n_12040 ^ x182;
assign n_12047 = n_12040 & ~n_12041;
assign n_12048 = n_12042 ^ n_10085;
assign n_12049 = n_12042 ^ n_12031;
assign n_12050 = n_12043 ^ n_11438;
assign n_12051 = n_12044 ^ n_11438;
assign n_12052 = n_11964 ^ n_12045;
assign n_12053 = n_12024 & n_12046;
assign n_12054 = n_12046 ^ n_12024;
assign n_12055 = n_12047 ^ x182;
assign n_12056 = n_12048 ^ n_12031;
assign n_12057 = n_12037 & ~n_12049;
assign n_12058 = n_12050 ^ n_10105;
assign n_12059 = n_12051 ^ n_11476;
assign n_12060 = n_12055 ^ n_12056;
assign n_12061 = n_12056 ^ x181;
assign n_12062 = n_12057 ^ n_10085;
assign n_12063 = n_10839 ^ n_12059;
assign n_12064 = n_12059 & ~n_11488;
assign n_12065 = n_12060 ^ x181;
assign n_12066 = n_12060 & ~n_12061;
assign n_12067 = n_12062 ^ n_10105;
assign n_12068 = n_12062 ^ n_12050;
assign n_12069 = n_12063 ^ n_11476;
assign n_12070 = n_11997 ^ n_12063;
assign n_12071 = n_12064 ^ n_10839;
assign n_12072 = n_12053 & n_12065;
assign n_12073 = n_12065 ^ n_12053;
assign n_12074 = n_12066 ^ x181;
assign n_12075 = n_12067 ^ n_12050;
assign n_12076 = ~n_12058 & n_12068;
assign n_12077 = n_10761 & n_12069;
assign n_12078 = n_12071 ^ n_11513;
assign n_12079 = n_12074 ^ n_12075;
assign n_12080 = n_12075 ^ x180;
assign n_12081 = n_12076 ^ n_10105;
assign n_12082 = n_12077 ^ n_11476;
assign n_12083 = n_12078 ^ n_10865;
assign n_12084 = ~n_12078 & n_11529;
assign n_12085 = n_12079 ^ x180;
assign n_12086 = ~n_12079 & n_12080;
assign n_12087 = n_12081 ^ n_10126;
assign n_12088 = n_12082 ^ n_10126;
assign n_12089 = n_12081 ^ n_12082;
assign n_12090 = n_12083 ^ n_11513;
assign n_12091 = n_12025 ^ n_12083;
assign n_12092 = n_12084 ^ n_10865;
assign n_12093 = n_12072 & ~n_12085;
assign n_12094 = n_12085 ^ n_12072;
assign n_12095 = n_12086 ^ x180;
assign n_12096 = n_12087 ^ n_12082;
assign n_12097 = ~n_12088 & ~n_12089;
assign n_12098 = ~n_10782 & n_12090;
assign n_12099 = n_12092 ^ n_11555;
assign n_12100 = n_12095 ^ n_12096;
assign n_12101 = n_12096 ^ x179;
assign n_12102 = n_12097 ^ n_10126;
assign n_12103 = n_12098 ^ n_11513;
assign n_12104 = n_10943 ^ n_12099;
assign n_12105 = ~n_12099 & n_11571;
assign n_12106 = n_12100 ^ x179;
assign n_12107 = ~n_12100 & n_12101;
assign n_12108 = n_12102 ^ n_10147;
assign n_12109 = n_12103 ^ n_12102;
assign n_12110 = n_12104 ^ n_11555;
assign n_12111 = n_12054 ^ n_12104;
assign n_12112 = n_12105 ^ n_10943;
assign n_12113 = ~n_12093 & n_12106;
assign n_12114 = n_12106 ^ n_12093;
assign n_12115 = n_12107 ^ x179;
assign n_12116 = n_12103 ^ n_12108;
assign n_12117 = ~n_12108 & ~n_12109;
assign n_12118 = n_10808 & n_12110;
assign n_12119 = n_12112 ^ n_11595;
assign n_12120 = n_12115 ^ n_12116;
assign n_12121 = n_12116 ^ x178;
assign n_12122 = n_12117 ^ n_10147;
assign n_12123 = n_12118 ^ n_11555;
assign n_12124 = n_10985 ^ n_12119;
assign n_12125 = ~n_12119 & ~n_11610;
assign n_12126 = n_12120 ^ x178;
assign n_12127 = n_12120 & ~n_12121;
assign n_12128 = n_12122 ^ n_10168;
assign n_12129 = n_12123 ^ n_10168;
assign n_12130 = n_12122 ^ n_12123;
assign n_12131 = n_12124 ^ n_11595;
assign n_12132 = n_12073 ^ n_12124;
assign n_12133 = n_12125 ^ n_10985;
assign n_12134 = ~n_12113 & n_12126;
assign n_12135 = n_12126 ^ n_12113;
assign n_12136 = n_12127 ^ x178;
assign n_12137 = n_12128 ^ n_12123;
assign n_12138 = ~n_12129 & n_12130;
assign n_12139 = n_10840 & ~n_12131;
assign n_12140 = n_12133 ^ n_11641;
assign n_12141 = n_12133 ^ n_11626;
assign n_12142 = n_12136 ^ n_12137;
assign n_12143 = n_12137 ^ x177;
assign n_12144 = n_12138 ^ n_10168;
assign n_12145 = n_12139 ^ n_11595;
assign n_12146 = n_12140 ^ n_11626;
assign n_12147 = n_12094 ^ n_12140;
assign n_12148 = n_11641 & n_12141;
assign n_12149 = n_12142 ^ x177;
assign n_12150 = ~n_12142 & n_12143;
assign n_12151 = n_12144 ^ n_10189;
assign n_12152 = n_12145 ^ n_10189;
assign n_12153 = n_12144 ^ n_12145;
assign n_12154 = ~n_10878 & ~n_12146;
assign n_12155 = n_12148 ^ n_11029;
assign n_12156 = ~n_12134 & n_12149;
assign n_12157 = n_12149 ^ n_12134;
assign n_12158 = n_12150 ^ x177;
assign n_12159 = n_12151 ^ n_12145;
assign n_12160 = ~n_12152 & n_12153;
assign n_12161 = n_12154 ^ n_11626;
assign n_12162 = n_12155 ^ n_11069;
assign n_12163 = n_12155 ^ n_11684;
assign n_12164 = n_12158 ^ n_12159;
assign n_12165 = n_12159 ^ x176;
assign n_12166 = n_12160 ^ n_10189;
assign n_12167 = n_12161 ^ n_10212;
assign n_12168 = n_12162 ^ n_11684;
assign n_12169 = n_11698 & ~n_12163;
assign n_12170 = n_12164 ^ x176;
assign n_12171 = ~n_12164 & n_12165;
assign n_12172 = n_12161 ^ n_12166;
assign n_12173 = n_12168 ^ n_11670;
assign n_12174 = n_12114 ^ n_12168;
assign n_12175 = n_12169 ^ n_11069;
assign n_12176 = n_12156 & n_12170;
assign n_12177 = n_12170 ^ n_12156;
assign n_12178 = n_12171 ^ x176;
assign n_12179 = n_12172 ^ n_10212;
assign n_12180 = n_12172 & n_12167;
assign n_12181 = ~n_10918 & ~n_12173;
assign n_12182 = n_12175 ^ n_11112;
assign n_12183 = n_12175 ^ n_11725;
assign n_12184 = n_12178 ^ x191;
assign n_12185 = n_12179 ^ x191;
assign n_12186 = n_12178 ^ n_12179;
assign n_12187 = n_12180 ^ n_10212;
assign n_12188 = n_12181 ^ n_11670;
assign n_12189 = n_10957 & n_12182;
assign n_12190 = n_12182 ^ n_11725;
assign n_12191 = ~n_11741 & n_12183;
assign n_12192 = n_12184 ^ n_12179;
assign n_12193 = ~n_12185 & n_12186;
assign n_12194 = n_12187 ^ n_12188;
assign n_12195 = n_12188 ^ n_10232;
assign n_12196 = n_12189 ^ n_11725;
assign n_12197 = n_12135 ^ n_12190;
assign n_12198 = n_12191 ^ n_11112;
assign n_12199 = n_12176 & ~n_12192;
assign n_12200 = n_12192 ^ n_12176;
assign n_12201 = n_12193 ^ x191;
assign n_12202 = n_12194 ^ n_10232;
assign n_12203 = n_12194 & ~n_12195;
assign n_12204 = n_12196 ^ n_10256;
assign n_12205 = n_12198 ^ n_11769;
assign n_12206 = n_12201 ^ n_12202;
assign n_12207 = n_12202 ^ x190;
assign n_12208 = n_12203 ^ n_10232;
assign n_12209 = n_11152 ^ n_12205;
assign n_12210 = n_12205 & ~n_11783;
assign n_12211 = n_12206 ^ x190;
assign n_12212 = n_12206 & ~n_12207;
assign n_12213 = n_12208 ^ n_10256;
assign n_12214 = n_12208 ^ n_12196;
assign n_12215 = n_12209 ^ n_11769;
assign n_12216 = n_12157 ^ n_12209;
assign n_12217 = n_12210 ^ n_11152;
assign n_12218 = ~n_12199 & n_12211;
assign n_12219 = n_12211 ^ n_12199;
assign n_12220 = n_12212 ^ x190;
assign n_12221 = n_12213 ^ n_12196;
assign n_12222 = n_12204 & n_12214;
assign n_12223 = ~n_11001 & n_12215;
assign n_12224 = n_12217 ^ n_11811;
assign n_12225 = n_12220 ^ x189;
assign n_12226 = n_12220 ^ n_12221;
assign n_12227 = n_12222 ^ n_10256;
assign n_12228 = n_12223 ^ n_11769;
assign n_12229 = n_11191 ^ n_12224;
assign n_12230 = ~n_12224 & n_11826;
assign n_12231 = n_12226 ^ x189;
assign n_12232 = ~n_12226 & n_12225;
assign n_12233 = n_12227 ^ n_10282;
assign n_12234 = n_12228 ^ n_10282;
assign n_12235 = n_12227 ^ n_12228;
assign n_12236 = n_12229 ^ n_11811;
assign n_12237 = n_12177 ^ n_12229;
assign n_12238 = n_12230 ^ n_11191;
assign n_12239 = n_12218 & ~n_12231;
assign n_12240 = n_12231 ^ n_12218;
assign n_12241 = n_12232 ^ x189;
assign n_12242 = n_12233 ^ n_12228;
assign n_12243 = ~n_12234 & ~n_12235;
assign n_12244 = ~n_11042 & n_12236;
assign n_12245 = n_12238 ^ n_11854;
assign n_12246 = n_12241 ^ n_12242;
assign n_12247 = n_12242 ^ x188;
assign n_12248 = n_12243 ^ n_10282;
assign n_12249 = n_12244 ^ n_11811;
assign n_12250 = n_11224 ^ n_12245;
assign n_12251 = ~n_12245 & n_11869;
assign n_12252 = n_12246 ^ x188;
assign n_12253 = ~n_12246 & n_12247;
assign n_12254 = n_12248 ^ n_10316;
assign n_12255 = n_12249 ^ n_10316;
assign n_12256 = n_12248 ^ n_12249;
assign n_12257 = n_12250 ^ n_11854;
assign n_12258 = n_12200 ^ n_12250;
assign n_12259 = n_12251 ^ n_11224;
assign n_12260 = n_12239 ^ n_12252;
assign n_12261 = n_12252 & ~n_12239;
assign n_12262 = n_12253 ^ x188;
assign n_12263 = n_12254 ^ n_12249;
assign n_12264 = n_12255 & ~n_12256;
assign n_12265 = n_11085 & n_12257;
assign n_12266 = n_12259 ^ n_11897;
assign n_12267 = n_12260 ^ n_11295;
assign n_12268 = n_11295 & ~n_12260;
assign n_12269 = n_12262 ^ n_12263;
assign n_12270 = n_12263 ^ x187;
assign n_12271 = n_12264 ^ n_10316;
assign n_12272 = n_12265 ^ n_11854;
assign n_12273 = n_11250 ^ n_12266;
assign n_12274 = ~n_12266 & ~n_11912;
assign n_12275 = n_12267 ^ n_11288;
assign n_12276 = n_11319 ^ n_12268;
assign n_12277 = n_12269 ^ x187;
assign n_12278 = ~n_12269 & n_12270;
assign n_12279 = n_12271 ^ n_10356;
assign n_12280 = n_12272 ^ n_10356;
assign n_12281 = n_12271 ^ n_12272;
assign n_12282 = n_12273 ^ n_11897;
assign n_12283 = n_12219 ^ n_12273;
assign n_12284 = n_12274 ^ n_11250;
assign n_12285 = n_10788 & ~n_12275;
assign n_12286 = n_12261 ^ n_12277;
assign n_12287 = ~n_12277 & ~n_12261;
assign n_12288 = n_12278 ^ x187;
assign n_12289 = n_12279 ^ n_12272;
assign n_12290 = ~n_12280 & ~n_12281;
assign n_12291 = ~n_11125 & ~n_12282;
assign n_12292 = n_12284 ^ n_11966;
assign n_12293 = n_12285 ^ n_11288;
assign n_12294 = n_12286 ^ n_12268;
assign n_12295 = n_12276 ^ n_12286;
assign n_12296 = n_12288 ^ n_12289;
assign n_12297 = n_12289 ^ x186;
assign n_12298 = n_12290 ^ n_10356;
assign n_12299 = n_12291 ^ n_11897;
assign n_12300 = n_12292 ^ n_11940;
assign n_12301 = n_12240 ^ n_12292;
assign n_12302 = n_12293 ^ n_10248;
assign n_12303 = n_10248 & n_12293;
assign n_12304 = n_10814 & ~n_12294;
assign n_12305 = n_12294 & ~n_12276;
assign n_12306 = n_12296 ^ x186;
assign n_12307 = n_12296 & ~n_12297;
assign n_12308 = n_12298 ^ n_10394;
assign n_12309 = n_12299 ^ n_10394;
assign n_12310 = n_12298 ^ n_12299;
assign n_12311 = n_11154 & n_12300;
assign n_12312 = x327 & n_12302;
assign n_12313 = n_12302 ^ x327;
assign n_12314 = n_12303 ^ n_10278;
assign n_12315 = n_12304 ^ n_11319;
assign n_12316 = n_12305 ^ n_11319;
assign n_12317 = n_12306 ^ n_12287;
assign n_12318 = ~n_12287 & ~n_12306;
assign n_12319 = n_12307 ^ x186;
assign n_12320 = n_12308 ^ n_12299;
assign n_12321 = n_12309 & n_12310;
assign n_12322 = n_12311 ^ n_11940;
assign n_12323 = n_12312 ^ x326;
assign n_12324 = n_12315 ^ n_12314;
assign n_12325 = n_12315 ^ n_12303;
assign n_12326 = n_11359 ^ n_12316;
assign n_12327 = n_12316 ^ n_12317;
assign n_12328 = n_11359 ^ n_12317;
assign n_12329 = n_12319 ^ n_12320;
assign n_12330 = n_12320 ^ x185;
assign n_12331 = n_12321 ^ n_10394;
assign n_12332 = n_12322 ^ n_10435;
assign n_12333 = n_12324 ^ n_12312;
assign n_12334 = n_12324 ^ n_12323;
assign n_12335 = n_12314 & n_12325;
assign n_12336 = n_12326 ^ n_12317;
assign n_12337 = ~n_10862 & ~n_12327;
assign n_12338 = n_12327 & n_12328;
assign n_12339 = n_12329 ^ x185;
assign n_12340 = n_12329 & ~n_12330;
assign n_12341 = n_12331 ^ x184;
assign n_12342 = n_12323 & n_12333;
assign n_12343 = ~n_12313 & n_12334;
assign n_12344 = n_12334 ^ n_12313;
assign n_12345 = n_12335 ^ n_10278;
assign n_12346 = n_12337 ^ n_11359;
assign n_12347 = n_12338 ^ n_11359;
assign n_12348 = n_12339 ^ n_12318;
assign n_12349 = ~n_12318 & n_12339;
assign n_12350 = n_12340 ^ x185;
assign n_12351 = n_12341 ^ n_12332;
assign n_12352 = n_12342 ^ x326;
assign n_12353 = n_12345 ^ n_10318;
assign n_12354 = n_12346 ^ n_10318;
assign n_12355 = n_12345 ^ n_12346;
assign n_12356 = n_11392 ^ n_12347;
assign n_12357 = n_12347 ^ n_12348;
assign n_12358 = n_11392 ^ n_12348;
assign n_12359 = n_12350 ^ n_12349;
assign n_12360 = n_12353 ^ n_12346;
assign n_12361 = n_12354 & ~n_12355;
assign n_12362 = n_12356 ^ n_12348;
assign n_12363 = n_10900 & n_12357;
assign n_12364 = ~n_12357 & n_12358;
assign n_12365 = n_12359 ^ n_12351;
assign n_12366 = n_12352 ^ n_12360;
assign n_12367 = n_12360 ^ x325;
assign n_12368 = n_12361 ^ n_10318;
assign n_12369 = n_12363 ^ n_11392;
assign n_12370 = n_12364 ^ n_11392;
assign n_12371 = n_11446 ^ n_12365;
assign n_12372 = n_12366 ^ x325;
assign n_12373 = ~n_12366 & n_12367;
assign n_12374 = n_12368 ^ n_10360;
assign n_12375 = n_12369 ^ n_10360;
assign n_12376 = n_12368 ^ n_12369;
assign n_12377 = n_12370 ^ n_12365;
assign n_12378 = n_11446 ^ n_12370;
assign n_12379 = ~n_12343 & n_12372;
assign n_12380 = n_12372 ^ n_12343;
assign n_12381 = n_12373 ^ x325;
assign n_12382 = n_12374 ^ n_12369;
assign n_12383 = ~n_12375 & ~n_12376;
assign n_12384 = ~n_10939 & n_12377;
assign n_12385 = ~n_12377 & n_12371;
assign n_12386 = n_12378 ^ n_12365;
assign n_12387 = n_12381 ^ n_12382;
assign n_12388 = n_12382 ^ x324;
assign n_12389 = n_12383 ^ n_10360;
assign n_12390 = n_12384 ^ n_11446;
assign n_12391 = n_12385 ^ n_11446;
assign n_12392 = n_12387 ^ x324;
assign n_12393 = n_12387 & ~n_12388;
assign n_12394 = n_12389 ^ n_10401;
assign n_12395 = n_12390 ^ n_10401;
assign n_12396 = n_12389 ^ n_12390;
assign n_12397 = n_12391 ^ n_11335;
assign n_12398 = n_11498 ^ n_12391;
assign n_12399 = n_12379 & ~n_12392;
assign n_12400 = n_12392 ^ n_12379;
assign n_12401 = n_12393 ^ x324;
assign n_12402 = n_12394 ^ n_12390;
assign n_12403 = ~n_12395 & n_12396;
assign n_12404 = n_10980 & ~n_12397;
assign n_12405 = n_12397 & n_11498;
assign n_12406 = n_12401 ^ n_12402;
assign n_12407 = n_12402 ^ x323;
assign n_12408 = n_12403 ^ n_10401;
assign n_12409 = n_12404 ^ n_11484;
assign n_12410 = n_12405 ^ n_11484;
assign n_12411 = n_12406 ^ x323;
assign n_12412 = ~n_12406 & n_12407;
assign n_12413 = n_12408 ^ n_10440;
assign n_12414 = n_12409 ^ n_12408;
assign n_12415 = n_11538 ^ n_12410;
assign n_12416 = ~n_12399 & ~n_12411;
assign n_12417 = n_12411 ^ n_12399;
assign n_12418 = n_12412 ^ x323;
assign n_12419 = n_12409 ^ n_12413;
assign n_12420 = n_12413 & ~n_12414;
assign n_12421 = n_11397 ^ n_12415;
assign n_12422 = n_12415 & n_11551;
assign n_12423 = n_12418 ^ n_12419;
assign n_12424 = n_12419 ^ x322;
assign n_12425 = n_12420 ^ n_10440;
assign n_12426 = n_12421 ^ n_11538;
assign n_12427 = n_12422 ^ n_11397;
assign n_12428 = n_12423 ^ x322;
assign n_12429 = n_12423 & ~n_12424;
assign n_12430 = n_12425 ^ n_10478;
assign n_12431 = n_11024 & ~n_12426;
assign n_12432 = n_11580 ^ n_12427;
assign n_12433 = ~n_12416 & ~n_12428;
assign n_12434 = n_12428 ^ n_12416;
assign n_12435 = n_12429 ^ x322;
assign n_12436 = n_12431 ^ n_11538;
assign n_12437 = ~n_12432 & ~n_11593;
assign n_12438 = n_11436 ^ n_12432;
assign n_12439 = n_12435 ^ x321;
assign n_12440 = n_12430 ^ n_12436;
assign n_12441 = n_12436 ^ n_10478;
assign n_12442 = n_12425 ^ n_12436;
assign n_12443 = n_12437 ^ n_11436;
assign n_12444 = n_12438 ^ n_11580;
assign n_12445 = n_12435 ^ n_12440;
assign n_12446 = ~n_12441 & n_12442;
assign n_12447 = n_11622 ^ n_12443;
assign n_12448 = n_11064 & ~n_12444;
assign n_12449 = n_12445 ^ x321;
assign n_12450 = ~n_12445 & n_12439;
assign n_12451 = n_12446 ^ n_10478;
assign n_12452 = n_12447 & ~n_11635;
assign n_12453 = n_11474 ^ n_12447;
assign n_12454 = n_12448 ^ n_11580;
assign n_12455 = n_12449 ^ n_12433;
assign n_12456 = ~n_12433 & ~n_12449;
assign n_12457 = n_12450 ^ x321;
assign n_12458 = n_12451 ^ n_10508;
assign n_12459 = n_12452 ^ n_11474;
assign n_12460 = n_12453 ^ n_11622;
assign n_12461 = n_12454 ^ n_10508;
assign n_12462 = n_12451 ^ n_12454;
assign n_12463 = n_12458 ^ n_12454;
assign n_12464 = n_11663 ^ n_12459;
assign n_12465 = n_11107 & n_12460;
assign n_12466 = ~n_12461 & n_12462;
assign n_12467 = n_12457 ^ n_12463;
assign n_12468 = n_12463 ^ x320;
assign n_12469 = ~n_12464 & ~n_11679;
assign n_12470 = n_11524 ^ n_12464;
assign n_12471 = n_12465 ^ n_11622;
assign n_12472 = n_12466 ^ n_10508;
assign n_12473 = n_12467 ^ x320;
assign n_12474 = ~n_12467 & n_12468;
assign n_12475 = n_12469 ^ n_11524;
assign n_12476 = n_12470 ^ n_11663;
assign n_12477 = n_12313 ^ n_12470;
assign n_12478 = n_12471 ^ n_10531;
assign n_12479 = n_12472 ^ n_12471;
assign n_12480 = n_12472 ^ n_10531;
assign n_12481 = ~n_12456 & n_12473;
assign n_12482 = n_12473 ^ n_12456;
assign n_12483 = n_12474 ^ x320;
assign n_12484 = n_11705 ^ n_12475;
assign n_12485 = n_11147 & ~n_12476;
assign n_12486 = ~n_12478 & n_12479;
assign n_12487 = n_12480 ^ n_12471;
assign n_12488 = ~n_12484 & n_11720;
assign n_12489 = n_11567 ^ n_12484;
assign n_12490 = n_12485 ^ n_11663;
assign n_12491 = n_12486 ^ n_10531;
assign n_12492 = n_12483 ^ n_12487;
assign n_12493 = n_12487 ^ x335;
assign n_12494 = n_12488 ^ n_11567;
assign n_12495 = n_12489 ^ n_11705;
assign n_12496 = n_12344 ^ n_12489;
assign n_12497 = n_12490 ^ n_10548;
assign n_12498 = n_12491 ^ n_12490;
assign n_12499 = n_12491 ^ n_10548;
assign n_12500 = n_12492 ^ x335;
assign n_12501 = ~n_12492 & n_12493;
assign n_12502 = n_11749 ^ n_12494;
assign n_12503 = ~n_11186 & n_12495;
assign n_12504 = n_12497 & ~n_12498;
assign n_12505 = n_12499 ^ n_12490;
assign n_12506 = n_12500 & n_12481;
assign n_12507 = n_12481 ^ n_12500;
assign n_12508 = n_12501 ^ x335;
assign n_12509 = n_12502 & ~n_11764;
assign n_12510 = n_12502 ^ n_11618;
assign n_12511 = n_12503 ^ n_11705;
assign n_12512 = n_12504 ^ n_10548;
assign n_12513 = n_12505 ^ x334;
assign n_12514 = n_12508 ^ n_12505;
assign n_12515 = n_12509 ^ n_11618;
assign n_12516 = n_12510 ^ n_11749;
assign n_12517 = n_12380 ^ n_12510;
assign n_12518 = n_12511 ^ n_10562;
assign n_12519 = n_12512 ^ n_12511;
assign n_12520 = n_12512 ^ n_10562;
assign n_12521 = n_12514 & ~n_12513;
assign n_12522 = n_12514 ^ x334;
assign n_12523 = n_11790 ^ n_12515;
assign n_12524 = n_11219 & n_12516;
assign n_12525 = ~n_12518 & n_12519;
assign n_12526 = n_12520 ^ n_12511;
assign n_12527 = n_12521 ^ x334;
assign n_12528 = ~n_12522 & n_12506;
assign n_12529 = n_12506 ^ n_12522;
assign n_12530 = ~n_12523 & ~n_11805;
assign n_12531 = n_12523 ^ n_11667;
assign n_12532 = n_12524 ^ n_11749;
assign n_12533 = n_12525 ^ n_10562;
assign n_12534 = n_12526 ^ x333;
assign n_12535 = n_12527 ^ n_12526;
assign n_12536 = n_12530 ^ n_11667;
assign n_12537 = n_12400 ^ n_12531;
assign n_12538 = n_12531 ^ n_11775;
assign n_12539 = n_12532 ^ n_10578;
assign n_12540 = n_12533 ^ n_12532;
assign n_12541 = n_12533 ^ n_10578;
assign n_12542 = ~n_12535 & n_12534;
assign n_12543 = n_12535 ^ x333;
assign n_12544 = n_11834 ^ n_12536;
assign n_12545 = n_11245 & ~n_12538;
assign n_12546 = n_12539 & ~n_12540;
assign n_12547 = n_12541 ^ n_12532;
assign n_12548 = n_12542 ^ x333;
assign n_12549 = ~n_12528 & ~n_12543;
assign n_12550 = n_12543 ^ n_12528;
assign n_12551 = n_12544 & n_11849;
assign n_12552 = n_12544 ^ n_11710;
assign n_12553 = n_12545 ^ n_11775;
assign n_12554 = n_12546 ^ n_10578;
assign n_12555 = n_12547 ^ x332;
assign n_12556 = n_12548 ^ n_12547;
assign n_12557 = n_12551 ^ n_11710;
assign n_12558 = n_12552 ^ n_11834;
assign n_12559 = n_12417 ^ n_12552;
assign n_12560 = n_12553 ^ n_10596;
assign n_12561 = n_12553 ^ n_12554;
assign n_12562 = n_12554 ^ n_10596;
assign n_12563 = n_12556 & ~n_12555;
assign n_12564 = n_12556 ^ x332;
assign n_12565 = n_12557 ^ n_11754;
assign n_12566 = n_11877 ^ n_12557;
assign n_12567 = ~n_11266 & ~n_12558;
assign n_12568 = n_12560 & n_12561;
assign n_12569 = n_12553 ^ n_12562;
assign n_12570 = n_12563 ^ x332;
assign n_12571 = ~n_12549 & ~n_12564;
assign n_12572 = n_12564 ^ n_12549;
assign n_12573 = n_11877 ^ n_12565;
assign n_12574 = ~n_11276 & ~n_12565;
assign n_12575 = ~n_11892 & ~n_12566;
assign n_12576 = n_12567 ^ n_11834;
assign n_12577 = n_12568 ^ n_10596;
assign n_12578 = n_12569 ^ x331;
assign n_12579 = n_12570 ^ n_12569;
assign n_12580 = n_12434 ^ n_12573;
assign n_12581 = n_11877 ^ n_12574;
assign n_12582 = n_12575 ^ n_11754;
assign n_12583 = n_12576 ^ n_10616;
assign n_12584 = n_12576 ^ n_12577;
assign n_12585 = n_12577 ^ n_10616;
assign n_12586 = n_12579 & ~n_12578;
assign n_12587 = n_12579 ^ x331;
assign n_12588 = n_12581 ^ n_10635;
assign n_12589 = n_11918 ^ n_12582;
assign n_12590 = ~n_12583 & ~n_12584;
assign n_12591 = n_12576 ^ n_12585;
assign n_12592 = n_12586 ^ x331;
assign n_12593 = n_12587 & ~n_12571;
assign n_12594 = n_12571 ^ n_12587;
assign n_12595 = n_11795 ^ n_12589;
assign n_12596 = n_12589 & ~n_11933;
assign n_12597 = n_12590 ^ n_10616;
assign n_12598 = n_12591 ^ x330;
assign n_12599 = n_12592 ^ n_12591;
assign n_12600 = n_12595 ^ n_11918;
assign n_12601 = n_12455 ^ n_12595;
assign n_12602 = n_12596 ^ n_11795;
assign n_12603 = n_12581 ^ n_12597;
assign n_12604 = n_12597 ^ n_10635;
assign n_12605 = n_12599 & ~n_12598;
assign n_12606 = n_12599 ^ x330;
assign n_12607 = ~n_11305 & n_12600;
assign n_12608 = n_12602 ^ n_11970;
assign n_12609 = n_12602 ^ n_11956;
assign n_12610 = ~n_12588 & n_12603;
assign n_12611 = n_12581 ^ n_12604;
assign n_12612 = n_12605 ^ x330;
assign n_12613 = ~n_12593 & ~n_12606;
assign n_12614 = n_12606 ^ n_12593;
assign n_12615 = n_12607 ^ n_11918;
assign n_12616 = n_12608 ^ n_11956;
assign n_12617 = n_12482 ^ n_12608;
assign n_12618 = n_11970 & n_12609;
assign n_12619 = n_12610 ^ n_10635;
assign n_12620 = n_12611 ^ x329;
assign n_12621 = n_12612 ^ n_12611;
assign n_12622 = n_12615 ^ n_10651;
assign n_12623 = n_11331 & ~n_12616;
assign n_12624 = n_12618 ^ n_11839;
assign n_12625 = n_12615 ^ n_12619;
assign n_12626 = n_12619 ^ n_10651;
assign n_12627 = ~n_12621 & n_12620;
assign n_12628 = n_12621 ^ x329;
assign n_12629 = n_12623 ^ n_11956;
assign n_12630 = n_12624 ^ n_11882;
assign n_12631 = n_12624 ^ n_11993;
assign n_12632 = ~n_12622 & n_12625;
assign n_12633 = n_12615 ^ n_12626;
assign n_12634 = n_12627 ^ x329;
assign n_12635 = n_12613 & n_12628;
assign n_12636 = n_12628 ^ n_12613;
assign n_12637 = n_12629 ^ n_10681;
assign n_12638 = ~n_11363 & ~n_12630;
assign n_12639 = n_12630 ^ n_11993;
assign n_12640 = n_12005 & n_12631;
assign n_12641 = n_12632 ^ n_10651;
assign n_12642 = n_12633 ^ x328;
assign n_12643 = n_12634 ^ n_12633;
assign n_12644 = n_12638 ^ n_11993;
assign n_12645 = n_12507 ^ n_12639;
assign n_12646 = n_12640 ^ n_11882;
assign n_12647 = n_12641 ^ n_12629;
assign n_12648 = ~n_12643 & n_12642;
assign n_12649 = n_12643 ^ x328;
assign n_12650 = n_12644 ^ n_10701;
assign n_12651 = n_12646 ^ n_11925;
assign n_12652 = n_12646 ^ n_12023;
assign n_12653 = n_12647 & n_12637;
assign n_12654 = n_12647 ^ n_10681;
assign n_12655 = n_12648 ^ x328;
assign n_12656 = n_12635 & n_12649;
assign n_12657 = n_12649 ^ n_12635;
assign n_12658 = ~n_11399 & n_12651;
assign n_12659 = n_12651 ^ n_12023;
assign n_12660 = ~n_12033 & n_12652;
assign n_12661 = n_12653 ^ n_10681;
assign n_12662 = n_12654 ^ x343;
assign n_12663 = n_12654 ^ n_12655;
assign n_12664 = n_12655 ^ x343;
assign n_12665 = n_12658 ^ n_12023;
assign n_12666 = n_12529 ^ n_12659;
assign n_12667 = n_12660 ^ n_11925;
assign n_12668 = n_12661 ^ n_12644;
assign n_12669 = ~n_12662 & n_12663;
assign n_12670 = n_12654 ^ n_12664;
assign n_12671 = n_12665 ^ n_10719;
assign n_12672 = n_12045 ^ n_12667;
assign n_12673 = n_12668 & ~n_12650;
assign n_12674 = n_12668 ^ n_10701;
assign n_12675 = n_12669 ^ x343;
assign n_12676 = n_12656 & ~n_12670;
assign n_12677 = n_12670 ^ n_12656;
assign n_12678 = n_11964 ^ n_12672;
assign n_12679 = ~n_12672 & n_12052;
assign n_12680 = n_12673 ^ n_10701;
assign n_12681 = n_12674 ^ x342;
assign n_12682 = n_12675 ^ n_12674;
assign n_12683 = n_12678 ^ n_12045;
assign n_12684 = n_12550 ^ n_12678;
assign n_12685 = n_12679 ^ n_11964;
assign n_12686 = n_12680 ^ n_10719;
assign n_12687 = n_12680 ^ n_12665;
assign n_12688 = n_12682 & ~n_12681;
assign n_12689 = n_12682 ^ x342;
assign n_12690 = n_11438 & n_12683;
assign n_12691 = n_12685 ^ n_11997;
assign n_12692 = n_12685 ^ n_12063;
assign n_12693 = n_12686 ^ n_12665;
assign n_12694 = n_12671 & ~n_12687;
assign n_12695 = n_12688 ^ x342;
assign n_12696 = n_12676 & ~n_12689;
assign n_12697 = n_12689 ^ n_12676;
assign n_12698 = n_12690 ^ n_12045;
assign n_12699 = ~n_11476 & n_12691;
assign n_12700 = n_12691 ^ n_12063;
assign n_12701 = n_12070 & ~n_12692;
assign n_12702 = n_12693 ^ x341;
assign n_12703 = n_12694 ^ n_10719;
assign n_12704 = n_12695 ^ n_12693;
assign n_12705 = n_12695 ^ x341;
assign n_12706 = n_12698 ^ n_10740;
assign n_12707 = n_12699 ^ n_12063;
assign n_12708 = n_12572 ^ n_12700;
assign n_12709 = n_12701 ^ n_11997;
assign n_12710 = n_12703 ^ n_10740;
assign n_12711 = n_12703 ^ n_12698;
assign n_12712 = n_12702 & ~n_12704;
assign n_12713 = n_12705 ^ n_12693;
assign n_12714 = n_12707 ^ n_10761;
assign n_12715 = n_12709 ^ n_12083;
assign n_12716 = n_12710 ^ n_12698;
assign n_12717 = ~n_12706 & n_12711;
assign n_12718 = n_12712 ^ x341;
assign n_12719 = ~n_12696 & ~n_12713;
assign n_12720 = n_12713 ^ n_12696;
assign n_12721 = n_12025 ^ n_12715;
assign n_12722 = n_12715 & ~n_12091;
assign n_12723 = n_12716 ^ x340;
assign n_12724 = n_12717 ^ n_10740;
assign n_12725 = n_12718 ^ n_12716;
assign n_12726 = n_12721 ^ n_12083;
assign n_12727 = n_12594 ^ n_12721;
assign n_12728 = n_12722 ^ n_12025;
assign n_12729 = n_12724 ^ n_10761;
assign n_12730 = n_12724 ^ n_12707;
assign n_12731 = n_12725 & ~n_12723;
assign n_12732 = n_12725 ^ x340;
assign n_12733 = n_11513 & n_12726;
assign n_12734 = n_12728 ^ n_12104;
assign n_12735 = n_12729 ^ n_12707;
assign n_12736 = ~n_12714 & n_12730;
assign n_12737 = n_12731 ^ x340;
assign n_12738 = ~n_12732 & ~n_12719;
assign n_12739 = n_12719 ^ n_12732;
assign n_12740 = n_12733 ^ n_12083;
assign n_12741 = n_12054 ^ n_12734;
assign n_12742 = n_12734 & ~n_12111;
assign n_12743 = n_12735 ^ x339;
assign n_12744 = n_12736 ^ n_10761;
assign n_12745 = n_12737 ^ n_12735;
assign n_12746 = n_12740 ^ n_10782;
assign n_12747 = n_12741 ^ n_12104;
assign n_12748 = n_12614 ^ n_12741;
assign n_12749 = n_12742 ^ n_12054;
assign n_12750 = n_12744 ^ n_10782;
assign n_12751 = n_12744 ^ n_12740;
assign n_12752 = n_12745 & ~n_12743;
assign n_12753 = n_12745 ^ x339;
assign n_12754 = n_11555 & n_12747;
assign n_12755 = n_12749 ^ n_12124;
assign n_12756 = n_12750 ^ n_12740;
assign n_12757 = ~n_12746 & ~n_12751;
assign n_12758 = n_12752 ^ x339;
assign n_12759 = ~n_12753 & n_12738;
assign n_12760 = n_12738 ^ n_12753;
assign n_12761 = n_12754 ^ n_12104;
assign n_12762 = n_12073 ^ n_12755;
assign n_12763 = ~n_12755 & n_12132;
assign n_12764 = n_12756 ^ x338;
assign n_12765 = n_12757 ^ n_10782;
assign n_12766 = n_12758 ^ n_12756;
assign n_12767 = n_12761 ^ n_10808;
assign n_12768 = n_12762 ^ n_12124;
assign n_12769 = n_12636 ^ n_12762;
assign n_12770 = n_12763 ^ n_12073;
assign n_12771 = n_12765 ^ n_10808;
assign n_12772 = n_12765 ^ n_12761;
assign n_12773 = n_12766 & ~n_12764;
assign n_12774 = n_12766 ^ x338;
assign n_12775 = n_11595 & n_12768;
assign n_12776 = n_12770 ^ n_12094;
assign n_12777 = n_12770 ^ n_12140;
assign n_12778 = n_12771 ^ n_12761;
assign n_12779 = n_12767 & n_12772;
assign n_12780 = n_12773 ^ x338;
assign n_12781 = n_12759 & ~n_12774;
assign n_12782 = n_12774 ^ n_12759;
assign n_12783 = n_12775 ^ n_12124;
assign n_12784 = n_11626 & ~n_12776;
assign n_12785 = n_12776 ^ n_12140;
assign n_12786 = ~n_12147 & ~n_12777;
assign n_12787 = n_12778 ^ x337;
assign n_12788 = n_12779 ^ n_10808;
assign n_12789 = n_12780 ^ n_12778;
assign n_12790 = n_12783 ^ n_10840;
assign n_12791 = n_12784 ^ n_12140;
assign n_12792 = n_12785 ^ n_12657;
assign n_12793 = n_12786 ^ n_12094;
assign n_12794 = n_12788 ^ n_10840;
assign n_12795 = n_12788 ^ n_12783;
assign n_12796 = n_12789 & ~n_12787;
assign n_12797 = n_12789 ^ x337;
assign n_12798 = n_12791 ^ n_10878;
assign n_12799 = n_12793 ^ n_12114;
assign n_12800 = n_12793 ^ n_12168;
assign n_12801 = n_12794 ^ n_12783;
assign n_12802 = ~n_12790 & n_12795;
assign n_12803 = n_12796 ^ x337;
assign n_12804 = n_12797 & ~n_12781;
assign n_12805 = n_12781 ^ n_12797;
assign n_12806 = n_12799 ^ n_12168;
assign n_12807 = ~n_12174 & ~n_12800;
assign n_12808 = n_12801 ^ x336;
assign n_12809 = n_12802 ^ n_10840;
assign n_12810 = n_12803 ^ n_12801;
assign n_12811 = n_12806 ^ n_12162;
assign n_12812 = n_12806 ^ n_12677;
assign n_12813 = n_12807 ^ n_12114;
assign n_12814 = n_12798 ^ n_12809;
assign n_12815 = n_12809 ^ n_10878;
assign n_12816 = n_12791 ^ n_12809;
assign n_12817 = n_12810 & ~n_12808;
assign n_12818 = n_12810 ^ x336;
assign n_12819 = n_11684 & ~n_12811;
assign n_12820 = n_12190 ^ n_12813;
assign n_12821 = ~n_12815 & n_12816;
assign n_12822 = n_12817 ^ x336;
assign n_12823 = ~n_12818 & ~n_12804;
assign n_12824 = n_12804 ^ n_12818;
assign n_12825 = n_12819 ^ n_12162;
assign n_12826 = n_12135 ^ n_12820;
assign n_12827 = ~n_12820 & ~n_12197;
assign n_12828 = n_12821 ^ n_10878;
assign n_12829 = n_12822 ^ x351;
assign n_12830 = n_12814 ^ n_12822;
assign n_12831 = ~n_12267 & n_12824;
assign n_12832 = n_12824 ^ n_12267;
assign n_12833 = n_12825 ^ n_10918;
assign n_12834 = n_12826 ^ n_12182;
assign n_12835 = n_12826 ^ n_12697;
assign n_12836 = n_12827 ^ n_12135;
assign n_12837 = n_12828 ^ n_12825;
assign n_12838 = n_12814 ^ n_12829;
assign n_12839 = n_12829 & ~n_12830;
assign n_12840 = n_12295 ^ n_12831;
assign n_12841 = n_12832 ^ n_12260;
assign n_12842 = ~n_11725 & n_12834;
assign n_12843 = n_12836 ^ n_12209;
assign n_12844 = n_12837 ^ n_10918;
assign n_12845 = n_12837 & ~n_12833;
assign n_12846 = n_12838 & n_12823;
assign n_12847 = n_12823 ^ n_12838;
assign n_12848 = n_12839 ^ x351;
assign n_12849 = n_11295 & n_12841;
assign n_12850 = n_12842 ^ n_12182;
assign n_12851 = n_12157 ^ n_12843;
assign n_12852 = n_12843 & n_12216;
assign n_12853 = n_12844 ^ x350;
assign n_12854 = n_12845 ^ n_10918;
assign n_12855 = n_12847 ^ n_12831;
assign n_12856 = n_12840 ^ n_12847;
assign n_12857 = n_12848 ^ n_12844;
assign n_12858 = n_12849 ^ n_12260;
assign n_12859 = n_12850 ^ n_10957;
assign n_12860 = n_12851 ^ n_12209;
assign n_12861 = n_12720 ^ n_12851;
assign n_12862 = n_12852 ^ n_12157;
assign n_12863 = n_12854 ^ n_10957;
assign n_12864 = n_12854 ^ n_12850;
assign n_12865 = ~n_12855 & n_12840;
assign n_12866 = ~n_11319 & n_12855;
assign n_12867 = ~n_12857 & n_12853;
assign n_12868 = n_12857 ^ x350;
assign n_12869 = n_10788 & ~n_12858;
assign n_12870 = n_12858 ^ n_10788;
assign n_12871 = ~n_11769 & ~n_12860;
assign n_12872 = n_12862 ^ n_12229;
assign n_12873 = n_12863 ^ n_12850;
assign n_12874 = n_12859 & n_12864;
assign n_12875 = n_12865 ^ n_12295;
assign n_12876 = n_12866 ^ n_12295;
assign n_12877 = n_12867 ^ x350;
assign n_12878 = ~n_12868 & ~n_12846;
assign n_12879 = n_12846 ^ n_12868;
assign n_12880 = n_12869 ^ n_10814;
assign n_12881 = x487 & ~n_12870;
assign n_12882 = n_12870 ^ x487;
assign n_12883 = n_12871 ^ n_12209;
assign n_12884 = n_12177 ^ n_12872;
assign n_12885 = n_12872 & n_12237;
assign n_12886 = n_12873 ^ x349;
assign n_12887 = n_12874 ^ n_10957;
assign n_12888 = n_12336 ^ n_12875;
assign n_12889 = n_12876 ^ n_12869;
assign n_12890 = n_12877 ^ n_12873;
assign n_12891 = n_12879 ^ n_12875;
assign n_12892 = n_12876 ^ n_12880;
assign n_12893 = n_12881 ^ x486;
assign n_12894 = n_12883 ^ n_11001;
assign n_12895 = n_12884 ^ n_12229;
assign n_12896 = n_12739 ^ n_12884;
assign n_12897 = n_12885 ^ n_12177;
assign n_12898 = n_12887 ^ n_11001;
assign n_12899 = n_12887 ^ n_12883;
assign n_12900 = n_12888 ^ n_12879;
assign n_12901 = n_12880 & ~n_12889;
assign n_12902 = n_12890 & ~n_12886;
assign n_12903 = n_12890 ^ x349;
assign n_12904 = n_12891 & ~n_12888;
assign n_12905 = n_11359 & ~n_12891;
assign n_12906 = n_12892 ^ n_12881;
assign n_12907 = n_12892 ^ n_12893;
assign n_12908 = n_11811 & ~n_12895;
assign n_12909 = n_12897 ^ n_12250;
assign n_12910 = n_12898 ^ n_12883;
assign n_12911 = n_12894 & n_12899;
assign n_12912 = n_12901 ^ n_10814;
assign n_12913 = n_12902 ^ x349;
assign n_12914 = ~n_12903 & ~n_12878;
assign n_12915 = n_12878 ^ n_12903;
assign n_12916 = n_12904 ^ n_12336;
assign n_12917 = n_12905 ^ n_12336;
assign n_12918 = n_12893 & ~n_12906;
assign n_12919 = n_12907 & ~n_12882;
assign n_12920 = n_12882 ^ n_12907;
assign n_12921 = n_12908 ^ n_12229;
assign n_12922 = n_12200 ^ n_12909;
assign n_12923 = ~n_12909 & ~n_12258;
assign n_12924 = n_12910 ^ x348;
assign n_12925 = n_12911 ^ n_11001;
assign n_12926 = n_12912 ^ n_10862;
assign n_12927 = n_12913 ^ n_12910;
assign n_12928 = n_12362 ^ n_12915;
assign n_12929 = n_12916 ^ n_12915;
assign n_12930 = n_12362 ^ n_12916;
assign n_12931 = n_12917 ^ n_10862;
assign n_12932 = n_12912 ^ n_12917;
assign n_12933 = n_12918 ^ x486;
assign n_12934 = n_12921 ^ n_11042;
assign n_12935 = n_12922 ^ n_12250;
assign n_12936 = n_12760 ^ n_12922;
assign n_12937 = n_12923 ^ n_12200;
assign n_12938 = n_12925 ^ n_11042;
assign n_12939 = n_12925 ^ n_12921;
assign n_12940 = n_12926 ^ n_12917;
assign n_12941 = ~n_12927 & n_12924;
assign n_12942 = n_12927 ^ x348;
assign n_12943 = n_12929 & n_12928;
assign n_12944 = n_11392 & ~n_12929;
assign n_12945 = n_12930 ^ n_12915;
assign n_12946 = n_12931 & n_12932;
assign n_12947 = n_11854 & ~n_12935;
assign n_12948 = n_12937 ^ n_12273;
assign n_12949 = n_12938 ^ n_12921;
assign n_12950 = ~n_12934 & n_12939;
assign n_12951 = n_12933 ^ n_12940;
assign n_12952 = n_12940 ^ x485;
assign n_12953 = n_12941 ^ x348;
assign n_12954 = n_12942 & n_12914;
assign n_12955 = n_12914 ^ n_12942;
assign n_12956 = n_12943 ^ n_12362;
assign n_12957 = n_12944 ^ n_12362;
assign n_12958 = n_12946 ^ n_10862;
assign n_12959 = n_12947 ^ n_12250;
assign n_12960 = n_12219 ^ n_12948;
assign n_12961 = ~n_12948 & ~n_12283;
assign n_12962 = n_12949 ^ x347;
assign n_12963 = n_12950 ^ n_11042;
assign n_12964 = n_12951 ^ x485;
assign n_12965 = ~n_12951 & n_12952;
assign n_12966 = n_12953 ^ n_12949;
assign n_12967 = n_12386 ^ n_12955;
assign n_12968 = n_12956 ^ n_12955;
assign n_12969 = n_12386 ^ n_12956;
assign n_12970 = n_12958 ^ n_10900;
assign n_12971 = n_12957 ^ n_12958;
assign n_12972 = n_12959 ^ n_11085;
assign n_12973 = n_12960 ^ n_12273;
assign n_12974 = n_12782 ^ n_12960;
assign n_12975 = n_12961 ^ n_12219;
assign n_12976 = n_12963 ^ n_11085;
assign n_12977 = n_12963 ^ n_12959;
assign n_12978 = n_12919 & n_12964;
assign n_12979 = n_12964 ^ n_12919;
assign n_12980 = n_12965 ^ x485;
assign n_12981 = n_12966 ^ x347;
assign n_12982 = ~n_12966 & n_12962;
assign n_12983 = ~n_12968 & n_12967;
assign n_12984 = n_11446 & n_12968;
assign n_12985 = n_12969 ^ n_12955;
assign n_12986 = n_12957 ^ n_12970;
assign n_12987 = ~n_12970 & n_12971;
assign n_12988 = n_11897 & ~n_12973;
assign n_12989 = n_12975 ^ n_12301;
assign n_12990 = n_12976 ^ n_12959;
assign n_12991 = n_12972 & n_12977;
assign n_12992 = n_12981 ^ n_12954;
assign n_12993 = n_12954 & n_12981;
assign n_12994 = n_12982 ^ x347;
assign n_12995 = n_12983 ^ n_12386;
assign n_12996 = n_12984 ^ n_12386;
assign n_12997 = n_12980 ^ n_12986;
assign n_12998 = n_12986 ^ x484;
assign n_12999 = n_12987 ^ n_10900;
assign n_13000 = n_12988 ^ n_12273;
assign n_13001 = n_12989 ^ n_12292;
assign n_13002 = n_12805 ^ n_12989;
assign n_13003 = n_12990 ^ x346;
assign n_13004 = n_12991 ^ n_11085;
assign n_13005 = n_12398 ^ n_12992;
assign n_13006 = n_12994 ^ n_12990;
assign n_13007 = n_12992 ^ n_12995;
assign n_13008 = n_12398 ^ n_12995;
assign n_13009 = n_12996 ^ n_10939;
assign n_13010 = n_12997 ^ x484;
assign n_13011 = n_12997 & ~n_12998;
assign n_13012 = n_12999 ^ n_12996;
assign n_13013 = n_12999 ^ n_10939;
assign n_13014 = n_13000 ^ n_11125;
assign n_13015 = ~n_11940 & n_13001;
assign n_13016 = n_13004 ^ n_11125;
assign n_13017 = n_13000 ^ n_13004;
assign n_13018 = n_13006 ^ x346;
assign n_13019 = n_13006 & ~n_13003;
assign n_13020 = ~n_13007 & n_13005;
assign n_13021 = ~n_11484 & n_13007;
assign n_13022 = n_13008 ^ n_12992;
assign n_13023 = n_12978 & ~n_13010;
assign n_13024 = n_13010 ^ n_12978;
assign n_13025 = n_13011 ^ x484;
assign n_13026 = ~n_13009 & ~n_13012;
assign n_13027 = n_13013 ^ n_12996;
assign n_13028 = n_13015 ^ n_12292;
assign n_13029 = n_13000 ^ n_13016;
assign n_13030 = n_13014 & n_13017;
assign n_13031 = n_13018 ^ n_12993;
assign n_13032 = n_12993 & ~n_13018;
assign n_13033 = n_13019 ^ x346;
assign n_13034 = n_13020 ^ n_12398;
assign n_13035 = n_13021 ^ n_12398;
assign n_13036 = n_13026 ^ n_10939;
assign n_13037 = n_13025 ^ n_13027;
assign n_13038 = n_13027 ^ x483;
assign n_13039 = n_13028 ^ n_11154;
assign n_13040 = n_13029 ^ x345;
assign n_13041 = n_13030 ^ n_11125;
assign n_13042 = n_13031 ^ n_12421;
assign n_13043 = n_13033 ^ n_13029;
assign n_13044 = n_13034 ^ n_13031;
assign n_13045 = n_13034 ^ n_12421;
assign n_13046 = n_13035 ^ n_10980;
assign n_13047 = n_13036 ^ n_13035;
assign n_13048 = n_13036 ^ n_10980;
assign n_13049 = n_13037 ^ x483;
assign n_13050 = n_13037 & ~n_13038;
assign n_13051 = n_13041 ^ x344;
assign n_13052 = n_13043 ^ x345;
assign n_13053 = ~n_13043 & n_13040;
assign n_13054 = n_13044 & n_13042;
assign n_13055 = n_11538 & ~n_13044;
assign n_13056 = n_13045 ^ n_13031;
assign n_13057 = n_13046 & n_13047;
assign n_13058 = n_13048 ^ n_13035;
assign n_13059 = n_13023 & ~n_13049;
assign n_13060 = n_13049 ^ n_13023;
assign n_13061 = n_13050 ^ x483;
assign n_13062 = n_13051 ^ n_13039;
assign n_13063 = n_13052 ^ n_13032;
assign n_13064 = n_13032 & n_13052;
assign n_13065 = n_13053 ^ x345;
assign n_13066 = n_13054 ^ n_12421;
assign n_13067 = n_13055 ^ n_12421;
assign n_13068 = n_13057 ^ n_10980;
assign n_13069 = n_13058 ^ x482;
assign n_13070 = n_13061 ^ n_13058;
assign n_13071 = n_13063 ^ n_12438;
assign n_13072 = n_13065 ^ n_13062;
assign n_13073 = n_13066 ^ n_13063;
assign n_13074 = n_13066 ^ n_12438;
assign n_13075 = n_13067 ^ n_11024;
assign n_13076 = n_13068 ^ n_13067;
assign n_13077 = n_13068 ^ n_11024;
assign n_13078 = n_13070 & ~n_13069;
assign n_13079 = n_13070 ^ x482;
assign n_13080 = n_13072 ^ n_13064;
assign n_13081 = n_13073 & ~n_13071;
assign n_13082 = n_11580 & ~n_13073;
assign n_13083 = n_13074 ^ n_13063;
assign n_13084 = ~n_13075 & n_13076;
assign n_13085 = n_13077 ^ n_13067;
assign n_13086 = n_13078 ^ x482;
assign n_13087 = n_13059 & ~n_13079;
assign n_13088 = n_13079 ^ n_13059;
assign n_13089 = n_13080 ^ n_12453;
assign n_13090 = n_13081 ^ n_12438;
assign n_13091 = n_13082 ^ n_12438;
assign n_13092 = n_13084 ^ n_11024;
assign n_13093 = n_13085 ^ x481;
assign n_13094 = n_13086 ^ n_13085;
assign n_13095 = n_13090 ^ n_13080;
assign n_13096 = n_13090 ^ n_12453;
assign n_13097 = n_13091 ^ n_11064;
assign n_13098 = n_13092 ^ n_13091;
assign n_13099 = n_13092 ^ n_11064;
assign n_13100 = n_13094 & ~n_13093;
assign n_13101 = n_13094 ^ x481;
assign n_13102 = n_13095 & n_13089;
assign n_13103 = n_11622 & ~n_13095;
assign n_13104 = n_13096 ^ n_13080;
assign n_13105 = ~n_13097 & n_13098;
assign n_13106 = n_13099 ^ n_13091;
assign n_13107 = n_13100 ^ x481;
assign n_13108 = n_13087 & ~n_13101;
assign n_13109 = n_13101 ^ n_13087;
assign n_13110 = n_13102 ^ n_12453;
assign n_13111 = n_13103 ^ n_12453;
assign n_13112 = n_13105 ^ n_11064;
assign n_13113 = n_13106 ^ x480;
assign n_13114 = n_13107 ^ n_13106;
assign n_13115 = n_13110 ^ n_12313;
assign n_13116 = n_12477 ^ n_13110;
assign n_13117 = n_13111 ^ n_11107;
assign n_13118 = n_13112 ^ n_13111;
assign n_13119 = n_13112 ^ n_11107;
assign n_13120 = n_13114 & ~n_13113;
assign n_13121 = n_13114 ^ x480;
assign n_13122 = n_13115 & ~n_12477;
assign n_13123 = ~n_11663 & ~n_13115;
assign n_13124 = n_13117 & ~n_13118;
assign n_13125 = n_13119 ^ n_13111;
assign n_13126 = n_13120 ^ x480;
assign n_13127 = ~n_13108 & n_13121;
assign n_13128 = n_13121 ^ n_13108;
assign n_13129 = n_13122 ^ n_12470;
assign n_13130 = n_13123 ^ n_12470;
assign n_13131 = n_13124 ^ n_11107;
assign n_13132 = n_13125 ^ x495;
assign n_13133 = n_13126 ^ n_13125;
assign n_13134 = n_13129 ^ n_12489;
assign n_13135 = n_13131 ^ n_11147;
assign n_13136 = n_13130 ^ n_13131;
assign n_13137 = ~n_13133 & n_13132;
assign n_13138 = n_13133 ^ x495;
assign n_13139 = ~n_13134 & n_12496;
assign n_13140 = n_12344 ^ n_13134;
assign n_13141 = n_13130 ^ n_13135;
assign n_13142 = n_13135 & ~n_13136;
assign n_13143 = n_13137 ^ x495;
assign n_13144 = ~n_13127 & n_13138;
assign n_13145 = n_13138 ^ n_13127;
assign n_13146 = n_13139 ^ n_12344;
assign n_13147 = n_13140 ^ n_12489;
assign n_13148 = n_13141 ^ x494;
assign n_13149 = n_13142 ^ n_11147;
assign n_13150 = n_13143 ^ n_13141;
assign n_13151 = n_13146 ^ n_12510;
assign n_13152 = n_11705 & n_13147;
assign n_13153 = n_13149 ^ n_11186;
assign n_13154 = ~n_13150 & n_13148;
assign n_13155 = n_13150 ^ x494;
assign n_13156 = n_13151 & n_12517;
assign n_13157 = n_12380 ^ n_13151;
assign n_13158 = n_13152 ^ n_12489;
assign n_13159 = n_13154 ^ x494;
assign n_13160 = ~n_13144 & ~n_13155;
assign n_13161 = n_13155 ^ n_13144;
assign n_13162 = n_13156 ^ n_12380;
assign n_13163 = n_13157 ^ n_12510;
assign n_13164 = n_13158 ^ n_11186;
assign n_13165 = n_13149 ^ n_13158;
assign n_13166 = n_13153 ^ n_13158;
assign n_13167 = n_13162 ^ n_12531;
assign n_13168 = n_13162 ^ n_12400;
assign n_13169 = ~n_11749 & ~n_13163;
assign n_13170 = ~n_13164 & ~n_13165;
assign n_13171 = n_13159 ^ n_13166;
assign n_13172 = n_13166 ^ x493;
assign n_13173 = n_12537 & ~n_13167;
assign n_13174 = n_11790 & n_13168;
assign n_13175 = n_13168 ^ n_12531;
assign n_13176 = n_13169 ^ n_12510;
assign n_13177 = n_13170 ^ n_11186;
assign n_13178 = n_13171 ^ x493;
assign n_13179 = n_13171 & ~n_13172;
assign n_13180 = n_13173 ^ n_12400;
assign n_13181 = n_13174 ^ n_12531;
assign n_13182 = n_13176 ^ n_11219;
assign n_13183 = n_13177 ^ n_13176;
assign n_13184 = n_13177 ^ n_11219;
assign n_13185 = n_13160 & n_13178;
assign n_13186 = n_13178 ^ n_13160;
assign n_13187 = n_13179 ^ x493;
assign n_13188 = n_13180 ^ n_12552;
assign n_13189 = n_13181 ^ n_11245;
assign n_13190 = ~n_13182 & ~n_13183;
assign n_13191 = n_13184 ^ n_13176;
assign n_13192 = ~n_13188 & n_12559;
assign n_13193 = n_12417 ^ n_13188;
assign n_13194 = n_13190 ^ n_11219;
assign n_13195 = n_13187 ^ n_13191;
assign n_13196 = n_13191 ^ x492;
assign n_13197 = n_13192 ^ n_12417;
assign n_13198 = n_13193 ^ n_12552;
assign n_13199 = n_13194 ^ n_13181;
assign n_13200 = n_13194 ^ n_11245;
assign n_13201 = n_13195 ^ x492;
assign n_13202 = ~n_13195 & n_13196;
assign n_13203 = n_12573 ^ n_13197;
assign n_13204 = n_11834 & n_13198;
assign n_13205 = ~n_13189 & n_13199;
assign n_13206 = n_13200 ^ n_13181;
assign n_13207 = ~n_13185 & n_13201;
assign n_13208 = n_13201 ^ n_13185;
assign n_13209 = n_13202 ^ x492;
assign n_13210 = ~n_13203 & ~n_12580;
assign n_13211 = n_12434 ^ n_13203;
assign n_13212 = n_13204 ^ n_12552;
assign n_13213 = n_13205 ^ n_11245;
assign n_13214 = n_13206 ^ x491;
assign n_13215 = n_13209 ^ n_13206;
assign n_13216 = n_13210 ^ n_12434;
assign n_13217 = n_13211 ^ n_12565;
assign n_13218 = n_12882 ^ n_13211;
assign n_13219 = n_13212 ^ n_11266;
assign n_13220 = n_13213 ^ n_13212;
assign n_13221 = n_13213 ^ n_11266;
assign n_13222 = n_13215 & ~n_13214;
assign n_13223 = n_13215 ^ x491;
assign n_13224 = n_13216 ^ n_12595;
assign n_13225 = n_11877 & ~n_13217;
assign n_13226 = n_13219 & n_13220;
assign n_13227 = n_13221 ^ n_13212;
assign n_13228 = n_13222 ^ x491;
assign n_13229 = n_13207 & ~n_13223;
assign n_13230 = n_13223 ^ n_13207;
assign n_13231 = n_12455 ^ n_13224;
assign n_13232 = ~n_13224 & ~n_12601;
assign n_13233 = n_13225 ^ n_12565;
assign n_13234 = n_13226 ^ n_11266;
assign n_13235 = n_13227 ^ x490;
assign n_13236 = n_13228 ^ n_13227;
assign n_13237 = n_13231 ^ n_12595;
assign n_13238 = n_12920 ^ n_13231;
assign n_13239 = n_13232 ^ n_12455;
assign n_13240 = n_13233 ^ n_11276;
assign n_13241 = n_13234 ^ n_13233;
assign n_13242 = n_13234 ^ n_11276;
assign n_13243 = ~n_13236 & n_13235;
assign n_13244 = n_13236 ^ x490;
assign n_13245 = n_11918 & ~n_13237;
assign n_13246 = n_13239 ^ n_12617;
assign n_13247 = n_13239 ^ n_12608;
assign n_13248 = n_13240 & ~n_13241;
assign n_13249 = n_13242 ^ n_13233;
assign n_13250 = n_13243 ^ x490;
assign n_13251 = ~n_13229 & ~n_13244;
assign n_13252 = n_13244 ^ n_13229;
assign n_13253 = n_13245 ^ n_12595;
assign n_13254 = n_13246 ^ n_12608;
assign n_13255 = n_12979 ^ n_13246;
assign n_13256 = n_12617 & ~n_13247;
assign n_13257 = n_13248 ^ n_11276;
assign n_13258 = n_13249 ^ x489;
assign n_13259 = n_13250 ^ n_13249;
assign n_13260 = n_13253 ^ n_11305;
assign n_13261 = n_11956 & n_13254;
assign n_13262 = n_13256 ^ n_12482;
assign n_13263 = n_13257 ^ n_13253;
assign n_13264 = n_13257 ^ n_11305;
assign n_13265 = n_13259 & ~n_13258;
assign n_13266 = n_13259 ^ x489;
assign n_13267 = n_13261 ^ n_12608;
assign n_13268 = n_13262 ^ n_12507;
assign n_13269 = n_13262 ^ n_12639;
assign n_13270 = ~n_13260 & n_13263;
assign n_13271 = n_13264 ^ n_13253;
assign n_13272 = n_13265 ^ x489;
assign n_13273 = n_13251 & n_13266;
assign n_13274 = n_13266 ^ n_13251;
assign n_13275 = n_13267 ^ n_11331;
assign n_13276 = n_13268 ^ n_12639;
assign n_13277 = n_12645 & n_13269;
assign n_13278 = n_13270 ^ n_11305;
assign n_13279 = n_13271 ^ x488;
assign n_13280 = n_13272 ^ n_13271;
assign n_13281 = n_13276 ^ n_12630;
assign n_13282 = n_13024 ^ n_13276;
assign n_13283 = n_13277 ^ n_12507;
assign n_13284 = n_13278 ^ n_13275;
assign n_13285 = n_13278 ^ n_13267;
assign n_13286 = ~n_13280 & n_13279;
assign n_13287 = n_13280 ^ x488;
assign n_13288 = ~n_11993 & n_13281;
assign n_13289 = n_13283 ^ n_12529;
assign n_13290 = n_13283 ^ n_12659;
assign n_13291 = n_13284 ^ x503;
assign n_13292 = ~n_13275 & ~n_13285;
assign n_13293 = n_13286 ^ x488;
assign n_13294 = n_13273 & ~n_13287;
assign n_13295 = n_13287 ^ n_13273;
assign n_13296 = n_13288 ^ n_12630;
assign n_13297 = n_13289 ^ n_12659;
assign n_13298 = ~n_12666 & ~n_13290;
assign n_13299 = n_13292 ^ n_11331;
assign n_13300 = n_13293 ^ n_13284;
assign n_13301 = n_13293 ^ x503;
assign n_13302 = n_13296 ^ n_11363;
assign n_13303 = n_13297 ^ n_12651;
assign n_13304 = n_13060 ^ n_13297;
assign n_13305 = n_13298 ^ n_12529;
assign n_13306 = n_13299 ^ n_13296;
assign n_13307 = n_13291 & ~n_13300;
assign n_13308 = n_13301 ^ n_13284;
assign n_13309 = n_12023 & ~n_13303;
assign n_13310 = n_13305 ^ n_12678;
assign n_13311 = n_13306 ^ n_11363;
assign n_13312 = n_13306 & n_13302;
assign n_13313 = n_13307 ^ x503;
assign n_13314 = n_13294 & ~n_13308;
assign n_13315 = n_13308 ^ n_13294;
assign n_13316 = n_13309 ^ n_12651;
assign n_13317 = n_12550 ^ n_13310;
assign n_13318 = ~n_13310 & n_12684;
assign n_13319 = n_13311 ^ x502;
assign n_13320 = n_13312 ^ n_11363;
assign n_13321 = n_13313 ^ n_13311;
assign n_13322 = n_13316 ^ n_11399;
assign n_13323 = n_13317 ^ n_12678;
assign n_13324 = n_13088 ^ n_13317;
assign n_13325 = n_13318 ^ n_12550;
assign n_13326 = n_13320 ^ n_11399;
assign n_13327 = n_13320 ^ n_13316;
assign n_13328 = n_13321 ^ x502;
assign n_13329 = ~n_13321 & n_13319;
assign n_13330 = ~n_12045 & n_13323;
assign n_13331 = n_12700 ^ n_13325;
assign n_13332 = n_13326 ^ n_13316;
assign n_13333 = ~n_13322 & n_13327;
assign n_13334 = n_13328 & ~n_13314;
assign n_13335 = n_13314 ^ n_13328;
assign n_13336 = n_13329 ^ x502;
assign n_13337 = n_13330 ^ n_12678;
assign n_13338 = n_12572 ^ n_13331;
assign n_13339 = ~n_13331 & ~n_12708;
assign n_13340 = n_13332 ^ x501;
assign n_13341 = n_13333 ^ n_11399;
assign n_13342 = n_13336 ^ n_13332;
assign n_13343 = n_13337 ^ n_11438;
assign n_13344 = n_13338 ^ n_12691;
assign n_13345 = n_13109 ^ n_13338;
assign n_13346 = n_13339 ^ n_12572;
assign n_13347 = n_13341 ^ n_11438;
assign n_13348 = n_13341 ^ n_13337;
assign n_13349 = n_13342 ^ x501;
assign n_13350 = ~n_13342 & n_13340;
assign n_13351 = ~n_12063 & n_13344;
assign n_13352 = n_13346 ^ n_12721;
assign n_13353 = n_13347 ^ n_13337;
assign n_13354 = ~n_13343 & ~n_13348;
assign n_13355 = n_13334 ^ n_13349;
assign n_13356 = n_13349 & n_13334;
assign n_13357 = n_13350 ^ x501;
assign n_13358 = n_13351 ^ n_12691;
assign n_13359 = n_12594 ^ n_13352;
assign n_13360 = ~n_13352 & n_12727;
assign n_13361 = n_13353 ^ x500;
assign n_13362 = n_13354 ^ n_11438;
assign n_13363 = n_13355 ^ n_12832;
assign n_13364 = ~n_12832 & n_13355;
assign n_13365 = n_13357 ^ n_13353;
assign n_13366 = n_13358 ^ n_11476;
assign n_13367 = n_13359 ^ n_12721;
assign n_13368 = n_13128 ^ n_13359;
assign n_13369 = n_13360 ^ n_12594;
assign n_13370 = n_13362 ^ n_11476;
assign n_13371 = n_13362 ^ n_13358;
assign n_13372 = n_13363 ^ n_12824;
assign n_13373 = n_12856 ^ n_13364;
assign n_13374 = n_13365 ^ x500;
assign n_13375 = ~n_13365 & n_13361;
assign n_13376 = n_12083 & n_13367;
assign n_13377 = n_13369 ^ n_12741;
assign n_13378 = n_13370 ^ n_13358;
assign n_13379 = ~n_13366 & ~n_13371;
assign n_13380 = ~n_12267 & ~n_13372;
assign n_13381 = n_13374 ^ n_13356;
assign n_13382 = n_13356 & n_13374;
assign n_13383 = n_13375 ^ x500;
assign n_13384 = n_13376 ^ n_12721;
assign n_13385 = n_12614 ^ n_13377;
assign n_13386 = ~n_13377 & n_12748;
assign n_13387 = n_13378 ^ x499;
assign n_13388 = n_13379 ^ n_11476;
assign n_13389 = n_13380 ^ n_12824;
assign n_13390 = n_13381 ^ n_13364;
assign n_13391 = n_13373 ^ n_13381;
assign n_13392 = n_13383 ^ n_13378;
assign n_13393 = n_13384 ^ n_11513;
assign n_13394 = n_13385 ^ n_12741;
assign n_13395 = n_13145 ^ n_13385;
assign n_13396 = n_13386 ^ n_12614;
assign n_13397 = n_13388 ^ n_11513;
assign n_13398 = n_13388 ^ n_13384;
assign n_13399 = n_13389 ^ n_11295;
assign n_13400 = n_11295 & n_13389;
assign n_13401 = n_12295 & n_13390;
assign n_13402 = ~n_13390 & n_13373;
assign n_13403 = n_13392 ^ x499;
assign n_13404 = n_13392 & ~n_13387;
assign n_13405 = n_12104 & n_13394;
assign n_13406 = n_13396 ^ n_12762;
assign n_13407 = n_13397 ^ n_13384;
assign n_13408 = n_13393 & n_13398;
assign n_13409 = x135 & n_13399;
assign n_13410 = n_13399 ^ x135;
assign n_13411 = n_13400 ^ n_11319;
assign n_13412 = n_13401 ^ n_12856;
assign n_13413 = n_13402 ^ n_12856;
assign n_13414 = n_13382 ^ n_13403;
assign n_13415 = ~n_13403 & n_13382;
assign n_13416 = n_13404 ^ x499;
assign n_13417 = n_13405 ^ n_12741;
assign n_13418 = n_12636 ^ n_13406;
assign n_13419 = n_13406 & ~n_12769;
assign n_13420 = n_13407 ^ x498;
assign n_13421 = n_13408 ^ n_11513;
assign n_13422 = n_13409 ^ x134;
assign n_13423 = n_13412 ^ n_13411;
assign n_13424 = n_13412 ^ n_13400;
assign n_13425 = n_12900 ^ n_13413;
assign n_13426 = n_13413 ^ n_13414;
assign n_13427 = n_12900 ^ n_13414;
assign n_13428 = n_13416 ^ n_13407;
assign n_13429 = n_13417 ^ n_11555;
assign n_13430 = n_13418 ^ n_12762;
assign n_13431 = n_13161 ^ n_13418;
assign n_13432 = n_13419 ^ n_12636;
assign n_13433 = n_13421 ^ n_11555;
assign n_13434 = n_13421 ^ n_13417;
assign n_13435 = n_13423 ^ n_13409;
assign n_13436 = n_13423 ^ n_13422;
assign n_13437 = ~n_13411 & ~n_13424;
assign n_13438 = n_13425 ^ n_13414;
assign n_13439 = ~n_12336 & ~n_13426;
assign n_13440 = n_13426 & ~n_13427;
assign n_13441 = n_13428 ^ x498;
assign n_13442 = n_13428 & ~n_13420;
assign n_13443 = ~n_12124 & n_13430;
assign n_13444 = n_13432 ^ n_12792;
assign n_13445 = n_13432 ^ n_12785;
assign n_13446 = n_13433 ^ n_13417;
assign n_13447 = n_13429 & ~n_13434;
assign n_13448 = n_13422 & n_13435;
assign n_13449 = n_13437 ^ n_11319;
assign n_13450 = n_13439 ^ n_12900;
assign n_13451 = n_13440 ^ n_12900;
assign n_13452 = n_13441 ^ n_13415;
assign n_13453 = ~n_13415 & n_13441;
assign n_13454 = n_13442 ^ x498;
assign n_13455 = n_13443 ^ n_12762;
assign n_13456 = n_13444 ^ n_12785;
assign n_13457 = n_13186 ^ n_13444;
assign n_13458 = n_12792 & ~n_13445;
assign n_13459 = n_13446 ^ x497;
assign n_13460 = n_13447 ^ n_11555;
assign n_13461 = n_13448 ^ x134;
assign n_13462 = n_13449 ^ n_11359;
assign n_13463 = n_13450 ^ n_11359;
assign n_13464 = n_13449 ^ n_13450;
assign n_13465 = n_12945 ^ n_13451;
assign n_13466 = n_13452 ^ n_13451;
assign n_13467 = n_12945 ^ n_13452;
assign n_13468 = n_13454 ^ n_13446;
assign n_13469 = n_13455 ^ n_11595;
assign n_13470 = ~n_12140 & n_13456;
assign n_13471 = n_13458 ^ n_12657;
assign n_13472 = n_13460 ^ n_11595;
assign n_13473 = n_13460 ^ n_13455;
assign n_13474 = n_13462 ^ n_13450;
assign n_13475 = n_13463 & n_13464;
assign n_13476 = n_13465 ^ n_13452;
assign n_13477 = n_12362 & n_13466;
assign n_13478 = ~n_13466 & ~n_13467;
assign n_13479 = n_13468 ^ x497;
assign n_13480 = ~n_13468 & n_13459;
assign n_13481 = n_13470 ^ n_12785;
assign n_13482 = n_13471 ^ n_12677;
assign n_13483 = n_13471 ^ n_12806;
assign n_13484 = n_13472 ^ n_13455;
assign n_13485 = ~n_13469 & n_13473;
assign n_13486 = n_13461 ^ n_13474;
assign n_13487 = n_13474 ^ x133;
assign n_13488 = n_13475 ^ n_11359;
assign n_13489 = n_13477 ^ n_12945;
assign n_13490 = n_13478 ^ n_12945;
assign n_13491 = n_13479 ^ n_13453;
assign n_13492 = ~n_13453 & n_13479;
assign n_13493 = n_13480 ^ x497;
assign n_13494 = n_13481 ^ n_11626;
assign n_13495 = n_13482 ^ n_12806;
assign n_13496 = n_12812 & n_13483;
assign n_13497 = n_13484 ^ x496;
assign n_13498 = n_13485 ^ n_11595;
assign n_13499 = n_13486 ^ x133;
assign n_13500 = n_13486 & ~n_13487;
assign n_13501 = n_13488 ^ n_11392;
assign n_13502 = n_13489 ^ n_11392;
assign n_13503 = n_13488 ^ n_13489;
assign n_13504 = n_12985 ^ n_13490;
assign n_13505 = n_13490 ^ n_13491;
assign n_13506 = n_12985 ^ n_13491;
assign n_13507 = n_13493 ^ n_13484;
assign n_13508 = n_13495 ^ n_12799;
assign n_13509 = n_13208 ^ n_13495;
assign n_13510 = n_13496 ^ n_12677;
assign n_13511 = n_13498 ^ n_13494;
assign n_13512 = n_13498 ^ n_13481;
assign n_13513 = n_13500 ^ x133;
assign n_13514 = n_13501 ^ n_13489;
assign n_13515 = ~n_13502 & n_13503;
assign n_13516 = n_13504 ^ n_13491;
assign n_13517 = n_12386 & n_13505;
assign n_13518 = ~n_13505 & ~n_13506;
assign n_13519 = n_13507 ^ x496;
assign n_13520 = n_13507 & ~n_13497;
assign n_13521 = n_12168 & ~n_13508;
assign n_13522 = n_13510 ^ n_12697;
assign n_13523 = n_13510 ^ n_12826;
assign n_13524 = n_13511 ^ x511;
assign n_13525 = n_13494 & ~n_13512;
assign n_13526 = n_13513 ^ n_13514;
assign n_13527 = n_13514 ^ x132;
assign n_13528 = n_13515 ^ n_11392;
assign n_13529 = n_13517 ^ n_12985;
assign n_13530 = n_13518 ^ n_12985;
assign n_13531 = n_13492 ^ n_13519;
assign n_13532 = n_13519 & ~n_13492;
assign n_13533 = n_13520 ^ x496;
assign n_13534 = n_13521 ^ n_12799;
assign n_13535 = ~n_12190 & n_13522;
assign n_13536 = n_13522 ^ n_12826;
assign n_13537 = ~n_12835 & n_13523;
assign n_13538 = n_13525 ^ n_11626;
assign n_13539 = n_13526 ^ x132;
assign n_13540 = n_13526 & ~n_13527;
assign n_13541 = n_13528 ^ n_11446;
assign n_13542 = n_13529 ^ n_11446;
assign n_13543 = n_13528 ^ n_13529;
assign n_13544 = n_13530 ^ n_13022;
assign n_13545 = n_13530 ^ n_13531;
assign n_13546 = n_13531 ^ n_13022;
assign n_13547 = n_13533 ^ x511;
assign n_13548 = n_13533 ^ n_13511;
assign n_13549 = n_13534 ^ n_11684;
assign n_13550 = n_13535 ^ n_12826;
assign n_13551 = n_13230 ^ n_13536;
assign n_13552 = n_13537 ^ n_12697;
assign n_13553 = n_13538 ^ n_13534;
assign n_13554 = n_13540 ^ x132;
assign n_13555 = n_13541 ^ n_13529;
assign n_13556 = n_13542 & ~n_13543;
assign n_13557 = n_13544 ^ n_13531;
assign n_13558 = n_12398 & n_13545;
assign n_13559 = ~n_13545 & n_13546;
assign n_13560 = n_13547 ^ n_13511;
assign n_13561 = n_13524 & ~n_13548;
assign n_13562 = n_13550 ^ n_11725;
assign n_13563 = n_13552 ^ n_12851;
assign n_13564 = n_13553 ^ n_11684;
assign n_13565 = n_13553 & ~n_13549;
assign n_13566 = n_13554 ^ n_13555;
assign n_13567 = n_13555 ^ x131;
assign n_13568 = n_13556 ^ n_11446;
assign n_13569 = n_13558 ^ n_13022;
assign n_13570 = n_13559 ^ n_13022;
assign n_13571 = n_13532 ^ n_13560;
assign n_13572 = n_13560 & ~n_13532;
assign n_13573 = n_13561 ^ x511;
assign n_13574 = n_12720 ^ n_13563;
assign n_13575 = n_13563 & ~n_12861;
assign n_13576 = n_13564 ^ x510;
assign n_13577 = n_13565 ^ n_11684;
assign n_13578 = n_13566 ^ x131;
assign n_13579 = ~n_13566 & n_13567;
assign n_13580 = n_13568 ^ n_11484;
assign n_13581 = n_13569 ^ n_11484;
assign n_13582 = n_13568 ^ n_13569;
assign n_13583 = n_13570 ^ n_13056;
assign n_13584 = n_13570 ^ n_13571;
assign n_13585 = n_13571 ^ n_13056;
assign n_13586 = n_13573 ^ n_13564;
assign n_13587 = n_13574 ^ n_12851;
assign n_13588 = n_13252 ^ n_13574;
assign n_13589 = n_13575 ^ n_12720;
assign n_13590 = n_13577 ^ n_11725;
assign n_13591 = n_13577 ^ n_13550;
assign n_13592 = ~n_13539 & n_13578;
assign n_13593 = n_13578 ^ n_13539;
assign n_13594 = n_13579 ^ x131;
assign n_13595 = n_13580 ^ n_13569;
assign n_13596 = ~n_13581 & ~n_13582;
assign n_13597 = n_13583 ^ n_13571;
assign n_13598 = ~n_12421 & ~n_13584;
assign n_13599 = n_13584 & ~n_13585;
assign n_13600 = n_13586 ^ x510;
assign n_13601 = n_13586 & ~n_13576;
assign n_13602 = ~n_12209 & n_13587;
assign n_13603 = n_13589 ^ n_12884;
assign n_13604 = n_13590 ^ n_13550;
assign n_13605 = ~n_13562 & ~n_13591;
assign n_13606 = n_13594 ^ n_13595;
assign n_13607 = n_13595 ^ x130;
assign n_13608 = n_13596 ^ n_11484;
assign n_13609 = n_13598 ^ n_13056;
assign n_13610 = n_13599 ^ n_13056;
assign n_13611 = n_13572 ^ n_13600;
assign n_13612 = ~n_13600 & n_13572;
assign n_13613 = n_13601 ^ x510;
assign n_13614 = n_13602 ^ n_12851;
assign n_13615 = n_12739 ^ n_13603;
assign n_13616 = ~n_13603 & ~n_12896;
assign n_13617 = n_13604 ^ x509;
assign n_13618 = n_13605 ^ n_11725;
assign n_13619 = n_13606 ^ x130;
assign n_13620 = n_13606 & ~n_13607;
assign n_13621 = n_13608 ^ n_11538;
assign n_13622 = n_13609 ^ n_11538;
assign n_13623 = n_13608 ^ n_13609;
assign n_13624 = n_13610 ^ n_13083;
assign n_13625 = n_13610 ^ n_13611;
assign n_13626 = n_13611 ^ n_13083;
assign n_13627 = n_13613 ^ n_13604;
assign n_13628 = n_13614 ^ n_11769;
assign n_13629 = n_13615 ^ n_12884;
assign n_13630 = n_13274 ^ n_13615;
assign n_13631 = n_13616 ^ n_12739;
assign n_13632 = n_13618 ^ n_11769;
assign n_13633 = n_13618 ^ n_13614;
assign n_13634 = ~n_13619 & n_13592;
assign n_13635 = n_13592 ^ n_13619;
assign n_13636 = n_13620 ^ x130;
assign n_13637 = n_13621 ^ n_13609;
assign n_13638 = n_13622 & n_13623;
assign n_13639 = n_13624 ^ n_13611;
assign n_13640 = ~n_12438 & ~n_13625;
assign n_13641 = n_13625 & ~n_13626;
assign n_13642 = n_13627 ^ x509;
assign n_13643 = n_13627 & ~n_13617;
assign n_13644 = n_12229 & ~n_13629;
assign n_13645 = n_13631 ^ n_12922;
assign n_13646 = n_13632 ^ n_13614;
assign n_13647 = ~n_13628 & n_13633;
assign n_13648 = n_13636 ^ n_13637;
assign n_13649 = n_13637 ^ x129;
assign n_13650 = n_13638 ^ n_11538;
assign n_13651 = n_13640 ^ n_13083;
assign n_13652 = n_13641 ^ n_13083;
assign n_13653 = n_13612 ^ n_13642;
assign n_13654 = ~n_13642 & n_13612;
assign n_13655 = n_13643 ^ x509;
assign n_13656 = n_13644 ^ n_12884;
assign n_13657 = n_12760 ^ n_13645;
assign n_13658 = n_13645 & n_12936;
assign n_13659 = n_13646 ^ x508;
assign n_13660 = n_13647 ^ n_11769;
assign n_13661 = n_13648 ^ x129;
assign n_13662 = n_13648 & ~n_13649;
assign n_13663 = n_13650 ^ n_11580;
assign n_13664 = n_13651 ^ n_11580;
assign n_13665 = n_13650 ^ n_13651;
assign n_13666 = n_13652 ^ n_13104;
assign n_13667 = n_13652 ^ n_13653;
assign n_13668 = n_13653 ^ n_13104;
assign n_13669 = n_13655 ^ n_13646;
assign n_13670 = n_13656 ^ n_11811;
assign n_13671 = n_13657 ^ n_12922;
assign n_13672 = n_13295 ^ n_13657;
assign n_13673 = n_13658 ^ n_12760;
assign n_13674 = n_13660 ^ n_11811;
assign n_13675 = n_13660 ^ n_13656;
assign n_13676 = ~n_13634 & n_13661;
assign n_13677 = n_13661 ^ n_13634;
assign n_13678 = n_13662 ^ x129;
assign n_13679 = n_13663 ^ n_13651;
assign n_13680 = n_13664 & ~n_13665;
assign n_13681 = n_13666 ^ n_13653;
assign n_13682 = n_12453 & ~n_13667;
assign n_13683 = n_13667 & n_13668;
assign n_13684 = n_13669 ^ x508;
assign n_13685 = ~n_13669 & n_13659;
assign n_13686 = n_12250 & ~n_13671;
assign n_13687 = n_13673 ^ n_12960;
assign n_13688 = n_13674 ^ n_13656;
assign n_13689 = ~n_13670 & ~n_13675;
assign n_13690 = n_13678 ^ n_13679;
assign n_13691 = n_13679 ^ x128;
assign n_13692 = n_13680 ^ n_11580;
assign n_13693 = n_13682 ^ n_13104;
assign n_13694 = n_13683 ^ n_13104;
assign n_13695 = n_13684 ^ n_13654;
assign n_13696 = ~n_13654 & ~n_13684;
assign n_13697 = n_13685 ^ x508;
assign n_13698 = n_13686 ^ n_12922;
assign n_13699 = n_12782 ^ n_13687;
assign n_13700 = n_13687 & ~n_12974;
assign n_13701 = n_13688 ^ x507;
assign n_13702 = n_13689 ^ n_11811;
assign n_13703 = n_13690 ^ x128;
assign n_13704 = ~n_13690 & n_13691;
assign n_13705 = n_13692 ^ n_11622;
assign n_13706 = n_13693 ^ n_11622;
assign n_13707 = n_13692 ^ n_13693;
assign n_13708 = n_13694 ^ n_13116;
assign n_13709 = n_13694 ^ n_13695;
assign n_13710 = n_13695 ^ n_13116;
assign n_13711 = n_13697 ^ n_13688;
assign n_13712 = n_13698 ^ n_11854;
assign n_13713 = n_13699 ^ n_12960;
assign n_13714 = n_13315 ^ n_13699;
assign n_13715 = n_13700 ^ n_12782;
assign n_13716 = n_13702 ^ n_11854;
assign n_13717 = n_13702 ^ n_13698;
assign n_13718 = n_13676 & ~n_13703;
assign n_13719 = n_13703 ^ n_13676;
assign n_13720 = n_13704 ^ x128;
assign n_13721 = n_13705 ^ n_13693;
assign n_13722 = ~n_13706 & n_13707;
assign n_13723 = n_13708 ^ n_13695;
assign n_13724 = n_12470 & n_13709;
assign n_13725 = ~n_13709 & n_13710;
assign n_13726 = n_13711 ^ x507;
assign n_13727 = ~n_13711 & n_13701;
assign n_13728 = ~n_12273 & n_13713;
assign n_13729 = n_13715 ^ n_13002;
assign n_13730 = n_13716 ^ n_13698;
assign n_13731 = ~n_13712 & n_13717;
assign n_13732 = n_13720 ^ n_13721;
assign n_13733 = n_13721 ^ x143;
assign n_13734 = n_13722 ^ n_11622;
assign n_13735 = n_13724 ^ n_13116;
assign n_13736 = n_13725 ^ n_13116;
assign n_13737 = n_13726 ^ n_13696;
assign n_13738 = n_13696 & ~n_13726;
assign n_13739 = n_13727 ^ x507;
assign n_13740 = n_13728 ^ n_12960;
assign n_13741 = n_13729 ^ n_12989;
assign n_13742 = n_13335 ^ n_13729;
assign n_13743 = n_13730 ^ x506;
assign n_13744 = n_13731 ^ n_11854;
assign n_13745 = n_13732 ^ x143;
assign n_13746 = n_13732 & ~n_13733;
assign n_13747 = n_13734 ^ n_11663;
assign n_13748 = n_13735 ^ n_11663;
assign n_13749 = n_13734 ^ n_13735;
assign n_13750 = n_13736 ^ n_13140;
assign n_13751 = n_13736 ^ n_13737;
assign n_13752 = n_13737 ^ n_13140;
assign n_13753 = n_13739 ^ n_13730;
assign n_13754 = n_13740 ^ n_11897;
assign n_13755 = ~n_12292 & ~n_13741;
assign n_13756 = n_13744 ^ n_11897;
assign n_13757 = n_13744 ^ n_13740;
assign n_13758 = n_13718 & n_13745;
assign n_13759 = n_13745 ^ n_13718;
assign n_13760 = n_13746 ^ x143;
assign n_13761 = n_13747 ^ n_13735;
assign n_13762 = n_13748 & n_13749;
assign n_13763 = n_13750 ^ n_13737;
assign n_13764 = n_12489 & ~n_13751;
assign n_13765 = n_13751 & n_13752;
assign n_13766 = n_13753 ^ x506;
assign n_13767 = n_13753 & ~n_13743;
assign n_13768 = n_13755 ^ n_12989;
assign n_13769 = n_13756 ^ n_13740;
assign n_13770 = n_13754 & ~n_13757;
assign n_13771 = n_13760 ^ n_13761;
assign n_13772 = n_13761 ^ x142;
assign n_13773 = n_13762 ^ n_11663;
assign n_13774 = n_13764 ^ n_13140;
assign n_13775 = n_13765 ^ n_13140;
assign n_13776 = n_13766 ^ n_13738;
assign n_13777 = ~n_13738 & ~n_13766;
assign n_13778 = n_13767 ^ x506;
assign n_13779 = n_13768 ^ n_11940;
assign n_13780 = n_13769 ^ x505;
assign n_13781 = n_13770 ^ n_11897;
assign n_13782 = n_13771 ^ x142;
assign n_13783 = ~n_13771 & n_13772;
assign n_13784 = n_13773 ^ n_11705;
assign n_13785 = n_13774 ^ n_11705;
assign n_13786 = n_13773 ^ n_13774;
assign n_13787 = n_13775 ^ n_13157;
assign n_13788 = n_13775 ^ n_13776;
assign n_13789 = n_13776 ^ n_13157;
assign n_13790 = n_13778 ^ n_13769;
assign n_13791 = n_13781 ^ x504;
assign n_13792 = n_13758 & ~n_13782;
assign n_13793 = n_13782 ^ n_13758;
assign n_13794 = n_13783 ^ x142;
assign n_13795 = n_13784 ^ n_13774;
assign n_13796 = n_13785 & n_13786;
assign n_13797 = n_13787 ^ n_13776;
assign n_13798 = ~n_12510 & n_13788;
assign n_13799 = ~n_13788 & n_13789;
assign n_13800 = n_13790 ^ x505;
assign n_13801 = ~n_13790 & n_13780;
assign n_13802 = n_13791 ^ n_13779;
assign n_13803 = n_13794 ^ n_13795;
assign n_13804 = n_13795 ^ x141;
assign n_13805 = n_13796 ^ n_11705;
assign n_13806 = n_13798 ^ n_13157;
assign n_13807 = n_13799 ^ n_13157;
assign n_13808 = n_13777 ^ n_13800;
assign n_13809 = ~n_13800 & ~n_13777;
assign n_13810 = n_13801 ^ x505;
assign n_13811 = n_13803 ^ x141;
assign n_13812 = n_13803 & ~n_13804;
assign n_13813 = n_13805 ^ n_11749;
assign n_13814 = n_13806 ^ n_11749;
assign n_13815 = n_13805 ^ n_13806;
assign n_13816 = n_13807 ^ n_13175;
assign n_13817 = n_13175 ^ n_13808;
assign n_13818 = n_13807 ^ n_13808;
assign n_13819 = n_13810 ^ n_13809;
assign n_13820 = ~n_13792 & ~n_13811;
assign n_13821 = n_13811 ^ n_13792;
assign n_13822 = n_13812 ^ x141;
assign n_13823 = n_13813 ^ n_13806;
assign n_13824 = ~n_13814 & ~n_13815;
assign n_13825 = n_13816 ^ n_13808;
assign n_13826 = n_13817 & n_13818;
assign n_13827 = n_13819 ^ n_13802;
assign n_13828 = n_13822 ^ n_13823;
assign n_13829 = n_13823 ^ x140;
assign n_13830 = n_13824 ^ n_11749;
assign n_13831 = n_13825 ^ n_13168;
assign n_13832 = n_13826 ^ n_13175;
assign n_13833 = n_13827 ^ n_13193;
assign n_13834 = n_13828 ^ x140;
assign n_13835 = n_13828 & ~n_13829;
assign n_13836 = n_13830 ^ n_11790;
assign n_13837 = ~n_12531 & n_13831;
assign n_13838 = n_13832 ^ n_13827;
assign n_13839 = n_13832 ^ n_13193;
assign n_13840 = ~n_13820 & n_13834;
assign n_13841 = n_13835 ^ x140;
assign n_13842 = n_13837 ^ n_13168;
assign n_13843 = ~n_12552 & ~n_13838;
assign n_13844 = n_13838 & ~n_13833;
assign n_13845 = n_13839 ^ n_13827;
assign n_13846 = n_13836 ^ n_13842;
assign n_13847 = n_13842 ^ n_11790;
assign n_13848 = n_13830 ^ n_13842;
assign n_13849 = n_13843 ^ n_13193;
assign n_13850 = n_13844 ^ n_13193;
assign n_13851 = n_13841 ^ n_13846;
assign n_13852 = n_13846 ^ x139;
assign n_13853 = n_13847 & n_13848;
assign n_13854 = n_13849 ^ n_11834;
assign n_13855 = n_13850 ^ n_12882;
assign n_13856 = n_13218 ^ n_13850;
assign n_13857 = n_13851 ^ x139;
assign n_13858 = n_13851 & ~n_13852;
assign n_13859 = n_13853 ^ n_11790;
assign n_13860 = ~n_12573 & ~n_13855;
assign n_13861 = n_13855 & n_13218;
assign n_13862 = n_13840 & n_13857;
assign n_13863 = n_13857 ^ n_13840;
assign n_13864 = n_13858 ^ x139;
assign n_13865 = n_13859 ^ n_11834;
assign n_13866 = n_13859 ^ n_13849;
assign n_13867 = n_13860 ^ n_13211;
assign n_13868 = n_13861 ^ n_13211;
assign n_13869 = ~n_13363 & ~n_13863;
assign n_13870 = n_13863 ^ n_13363;
assign n_13871 = n_13865 ^ n_13849;
assign n_13872 = ~n_13854 & n_13866;
assign n_13873 = n_13868 ^ n_13231;
assign n_13874 = n_13391 ^ n_13869;
assign n_13875 = n_13870 ^ n_13355;
assign n_13876 = n_13864 ^ n_13871;
assign n_13877 = n_13871 ^ x138;
assign n_13878 = n_13872 ^ n_11834;
assign n_13879 = n_12920 ^ n_13873;
assign n_13880 = n_13873 & n_13238;
assign n_13881 = ~n_12832 & n_13875;
assign n_13882 = n_13876 ^ x138;
assign n_13883 = n_13876 & ~n_13877;
assign n_13884 = n_13878 ^ n_11877;
assign n_13885 = n_13867 ^ n_13878;
assign n_13886 = n_13879 ^ n_13231;
assign n_13887 = n_13880 ^ n_12920;
assign n_13888 = n_13881 ^ n_13355;
assign n_13889 = n_13862 & n_13882;
assign n_13890 = n_13882 ^ n_13862;
assign n_13891 = n_13883 ^ x138;
assign n_13892 = n_13867 ^ n_13884;
assign n_13893 = n_13884 & ~n_13885;
assign n_13894 = n_12595 & ~n_13886;
assign n_13895 = n_13887 ^ n_12979;
assign n_13896 = n_13887 ^ n_13246;
assign n_13897 = ~n_12267 & n_13888;
assign n_13898 = n_13888 ^ n_12267;
assign n_13899 = n_13890 ^ n_13869;
assign n_13900 = n_13874 ^ n_13890;
assign n_13901 = n_13891 ^ n_13892;
assign n_13902 = n_13892 ^ x137;
assign n_13903 = n_13893 ^ n_11877;
assign n_13904 = n_13894 ^ n_13231;
assign n_13905 = ~n_12608 & ~n_13895;
assign n_13906 = n_13895 ^ n_13246;
assign n_13907 = ~n_13255 & ~n_13896;
assign n_13908 = n_13897 ^ n_12295;
assign n_13909 = x295 & ~n_13898;
assign n_13910 = n_13898 ^ x295;
assign n_13911 = n_13899 & n_13874;
assign n_13912 = n_12856 & ~n_13899;
assign n_13913 = n_13901 ^ x137;
assign n_13914 = ~n_13901 & n_13902;
assign n_13915 = n_13903 ^ n_11918;
assign n_13916 = n_13904 ^ n_11918;
assign n_13917 = n_13903 ^ n_13904;
assign n_13918 = n_13905 ^ n_13246;
assign n_13919 = n_13907 ^ n_12979;
assign n_13920 = n_13909 ^ x294;
assign n_13921 = n_13911 ^ n_13391;
assign n_13922 = n_13912 ^ n_13391;
assign n_13923 = n_13889 & ~n_13913;
assign n_13924 = n_13913 ^ n_13889;
assign n_13925 = n_13914 ^ x137;
assign n_13926 = n_13915 ^ n_13904;
assign n_13927 = ~n_13916 & n_13917;
assign n_13928 = n_13918 ^ n_11956;
assign n_13929 = n_13919 ^ n_13024;
assign n_13930 = n_13919 ^ n_13276;
assign n_13931 = n_13438 ^ n_13921;
assign n_13932 = n_13922 ^ n_13897;
assign n_13933 = n_13922 ^ n_13908;
assign n_13934 = n_13921 ^ n_13924;
assign n_13935 = n_13438 ^ n_13924;
assign n_13936 = n_13925 ^ n_13926;
assign n_13937 = n_13926 ^ x136;
assign n_13938 = n_13927 ^ n_11918;
assign n_13939 = n_13929 ^ n_13276;
assign n_13940 = n_13282 & n_13930;
assign n_13941 = n_13931 ^ n_13924;
assign n_13942 = n_13908 & ~n_13932;
assign n_13943 = n_13933 ^ n_13909;
assign n_13944 = n_13933 ^ n_13920;
assign n_13945 = n_12900 & n_13934;
assign n_13946 = ~n_13934 & ~n_13935;
assign n_13947 = n_13936 ^ x136;
assign n_13948 = n_13936 & ~n_13937;
assign n_13949 = n_13918 ^ n_13938;
assign n_13950 = n_13939 ^ n_13268;
assign n_13951 = n_13940 ^ n_13024;
assign n_13952 = n_13942 ^ n_12295;
assign n_13953 = n_13920 & ~n_13943;
assign n_13954 = n_13945 ^ n_13438;
assign n_13955 = n_13946 ^ n_13438;
assign n_13956 = n_13923 ^ n_13947;
assign n_13957 = n_13947 & n_13923;
assign n_13958 = n_13948 ^ x136;
assign n_13959 = n_13949 ^ n_11956;
assign n_13960 = n_13949 & ~n_13928;
assign n_13961 = n_12639 & ~n_13950;
assign n_13962 = n_13951 ^ n_13297;
assign n_13963 = n_13952 ^ n_12336;
assign n_13964 = n_13953 ^ x294;
assign n_13965 = n_13954 ^ n_12336;
assign n_13966 = n_13952 ^ n_13954;
assign n_13967 = n_13476 ^ n_13955;
assign n_13968 = n_13956 ^ n_13955;
assign n_13969 = n_13476 ^ n_13956;
assign n_13970 = n_13958 ^ x151;
assign n_13971 = n_13959 ^ x151;
assign n_13972 = n_13958 ^ n_13959;
assign n_13973 = n_13960 ^ n_11956;
assign n_13974 = n_13961 ^ n_13268;
assign n_13975 = n_13060 ^ n_13962;
assign n_13976 = ~n_13962 & n_13304;
assign n_13977 = n_13963 ^ n_13954;
assign n_13978 = n_13965 & n_13966;
assign n_13979 = n_13967 ^ n_13956;
assign n_13980 = ~n_12945 & n_13968;
assign n_13981 = ~n_13968 & n_13969;
assign n_13982 = n_13970 ^ n_13959;
assign n_13983 = ~n_13971 & n_13972;
assign n_13984 = n_13973 ^ n_11993;
assign n_13985 = n_13974 ^ n_11993;
assign n_13986 = n_13973 ^ n_13974;
assign n_13987 = n_13975 ^ n_13289;
assign n_13988 = n_13976 ^ n_13060;
assign n_13989 = n_13964 ^ n_13977;
assign n_13990 = n_13977 ^ x293;
assign n_13991 = n_13978 ^ n_12336;
assign n_13992 = n_13980 ^ n_13476;
assign n_13993 = n_13981 ^ n_13476;
assign n_13994 = n_13982 ^ n_13957;
assign n_13995 = n_13957 & n_13982;
assign n_13996 = n_13983 ^ x151;
assign n_13997 = n_13984 ^ n_13974;
assign n_13998 = n_13985 & n_13986;
assign n_13999 = n_12659 & n_13987;
assign n_14000 = n_13988 ^ n_13088;
assign n_14001 = n_13988 ^ n_13317;
assign n_14002 = n_13989 ^ x293;
assign n_14003 = ~n_13989 & n_13990;
assign n_14004 = n_13991 ^ n_12362;
assign n_14005 = n_13992 ^ n_12362;
assign n_14006 = n_13991 ^ n_13992;
assign n_14007 = n_13516 ^ n_13993;
assign n_14008 = n_13993 ^ n_13994;
assign n_14009 = n_13516 ^ n_13994;
assign n_14010 = n_13996 ^ n_13997;
assign n_14011 = n_13997 ^ x150;
assign n_14012 = n_13998 ^ n_11993;
assign n_14013 = n_13999 ^ n_13289;
assign n_14014 = ~n_12678 & n_14000;
assign n_14015 = n_14000 ^ n_13317;
assign n_14016 = n_13324 & ~n_14001;
assign n_14017 = ~n_14002 & ~n_13944;
assign n_14018 = n_13944 ^ n_14002;
assign n_14019 = n_14003 ^ x293;
assign n_14020 = n_14004 ^ n_13992;
assign n_14021 = ~n_14005 & ~n_14006;
assign n_14022 = n_14007 ^ n_13994;
assign n_14023 = n_12985 & n_14008;
assign n_14024 = ~n_14008 & ~n_14009;
assign n_14025 = n_14010 ^ x150;
assign n_14026 = ~n_14010 & n_14011;
assign n_14027 = n_14012 ^ n_14013;
assign n_14028 = n_14013 ^ n_12023;
assign n_14029 = n_14014 ^ n_13317;
assign n_14030 = n_14016 ^ n_13088;
assign n_14031 = n_14019 ^ n_14020;
assign n_14032 = n_14020 ^ x292;
assign n_14033 = n_14021 ^ n_12362;
assign n_14034 = n_14023 ^ n_13516;
assign n_14035 = n_14024 ^ n_13516;
assign n_14036 = n_13995 ^ n_14025;
assign n_14037 = ~n_14025 & n_13995;
assign n_14038 = n_14026 ^ x150;
assign n_14039 = n_14027 ^ n_12023;
assign n_14040 = ~n_14027 & ~n_14028;
assign n_14041 = n_14029 ^ n_12045;
assign n_14042 = n_14030 ^ n_13338;
assign n_14043 = n_14031 ^ x292;
assign n_14044 = ~n_14031 & n_14032;
assign n_14045 = n_14033 ^ n_12386;
assign n_14046 = n_14034 ^ n_12386;
assign n_14047 = n_14033 ^ n_14034;
assign n_14048 = n_13557 ^ n_14035;
assign n_14049 = n_14035 ^ n_14036;
assign n_14050 = n_13557 ^ n_14036;
assign n_14051 = n_14038 ^ n_14039;
assign n_14052 = n_14039 ^ x149;
assign n_14053 = n_14040 ^ n_12023;
assign n_14054 = n_13109 ^ n_14042;
assign n_14055 = n_14042 & ~n_13345;
assign n_14056 = ~n_14017 & n_14043;
assign n_14057 = n_14043 ^ n_14017;
assign n_14058 = n_14044 ^ x292;
assign n_14059 = n_14045 ^ n_14034;
assign n_14060 = n_14046 & ~n_14047;
assign n_14061 = n_14048 ^ n_14036;
assign n_14062 = n_13022 & n_14049;
assign n_14063 = ~n_14049 & n_14050;
assign n_14064 = n_14051 ^ x149;
assign n_14065 = ~n_14051 & n_14052;
assign n_14066 = n_14053 ^ n_12045;
assign n_14067 = n_14053 ^ n_14029;
assign n_14068 = n_14054 ^ n_13338;
assign n_14069 = n_13410 ^ n_14054;
assign n_14070 = n_14055 ^ n_13109;
assign n_14071 = n_14058 ^ n_14059;
assign n_14072 = n_14059 ^ x291;
assign n_14073 = n_14060 ^ n_12386;
assign n_14074 = n_13910 ^ n_14061;
assign n_14075 = n_14062 ^ n_13557;
assign n_14076 = n_14063 ^ n_13557;
assign n_14077 = n_14037 ^ n_14064;
assign n_14078 = n_14064 & ~n_14037;
assign n_14079 = n_14065 ^ x149;
assign n_14080 = n_14066 ^ n_14029;
assign n_14081 = n_14041 & n_14067;
assign n_14082 = ~n_12700 & n_14068;
assign n_14083 = n_14070 ^ n_13359;
assign n_14084 = n_14071 ^ x291;
assign n_14085 = ~n_14071 & n_14072;
assign n_14086 = n_14073 ^ n_12398;
assign n_14087 = n_14075 ^ n_12398;
assign n_14088 = n_14073 ^ n_14075;
assign n_14089 = n_13597 ^ n_14076;
assign n_14090 = n_14076 ^ n_14077;
assign n_14091 = n_13597 ^ n_14077;
assign n_14092 = n_14079 ^ n_14080;
assign n_14093 = n_14080 ^ x148;
assign n_14094 = n_14081 ^ n_12045;
assign n_14095 = n_14082 ^ n_13338;
assign n_14096 = n_13128 ^ n_14083;
assign n_14097 = n_14083 & n_13368;
assign n_14098 = n_14056 & n_14084;
assign n_14099 = n_14084 ^ n_14056;
assign n_14100 = n_14085 ^ x291;
assign n_14101 = n_14086 ^ n_14075;
assign n_14102 = n_14087 & ~n_14088;
assign n_14103 = n_14089 ^ n_14077;
assign n_14104 = n_13056 & ~n_14090;
assign n_14105 = n_14090 & n_14091;
assign n_14106 = n_14092 ^ x148;
assign n_14107 = ~n_14092 & n_14093;
assign n_14108 = n_14094 ^ n_12063;
assign n_14109 = n_14095 ^ n_12063;
assign n_14110 = n_14094 ^ n_14095;
assign n_14111 = n_14096 ^ n_13359;
assign n_14112 = n_13436 ^ n_14096;
assign n_14113 = n_14097 ^ n_13128;
assign n_14114 = n_14100 ^ n_14101;
assign n_14115 = n_14101 ^ x290;
assign n_14116 = n_14102 ^ n_12398;
assign n_14117 = n_14103 ^ n_13944;
assign n_14118 = n_14104 ^ n_13597;
assign n_14119 = n_14105 ^ n_13597;
assign n_14120 = n_14078 ^ n_14106;
assign n_14121 = n_14106 & n_14078;
assign n_14122 = n_14107 ^ x148;
assign n_14123 = n_14108 ^ n_14095;
assign n_14124 = ~n_14109 & n_14110;
assign n_14125 = n_12721 & ~n_14111;
assign n_14126 = n_14113 ^ n_13385;
assign n_14127 = n_14114 ^ x290;
assign n_14128 = ~n_14114 & n_14115;
assign n_14129 = n_14116 ^ n_12421;
assign n_14130 = n_14118 ^ n_12421;
assign n_14131 = n_14116 ^ n_14118;
assign n_14132 = n_13639 ^ n_14119;
assign n_14133 = n_14119 ^ n_14120;
assign n_14134 = n_13639 ^ n_14120;
assign n_14135 = n_14122 ^ n_14123;
assign n_14136 = n_14123 ^ x147;
assign n_14137 = n_14124 ^ n_12063;
assign n_14138 = n_14125 ^ n_13359;
assign n_14139 = n_13145 ^ n_14126;
assign n_14140 = ~n_14126 & ~n_13395;
assign n_14141 = ~n_14098 & ~n_14127;
assign n_14142 = n_14127 ^ n_14098;
assign n_14143 = n_14128 ^ x290;
assign n_14144 = n_14129 ^ n_14118;
assign n_14145 = n_14130 & n_14131;
assign n_14146 = n_14132 ^ n_14120;
assign n_14147 = n_13083 & ~n_14133;
assign n_14148 = n_14133 & ~n_14134;
assign n_14149 = n_14135 ^ x147;
assign n_14150 = ~n_14135 & n_14136;
assign n_14151 = n_14137 ^ n_12083;
assign n_14152 = n_14138 ^ n_12083;
assign n_14153 = n_14137 ^ n_14138;
assign n_14154 = n_14139 ^ n_13385;
assign n_14155 = n_13499 ^ n_14139;
assign n_14156 = n_14140 ^ n_13145;
assign n_14157 = n_14143 ^ n_14144;
assign n_14158 = n_14144 ^ x289;
assign n_14159 = n_14145 ^ n_12421;
assign n_14160 = n_14018 ^ n_14146;
assign n_14161 = n_14147 ^ n_13639;
assign n_14162 = n_14148 ^ n_13639;
assign n_14163 = n_14149 ^ n_14121;
assign n_14164 = ~n_14121 & ~n_14149;
assign n_14165 = n_14150 ^ x147;
assign n_14166 = n_14151 ^ n_14138;
assign n_14167 = n_14152 & n_14153;
assign n_14168 = n_12741 & ~n_14154;
assign n_14169 = n_14156 ^ n_13418;
assign n_14170 = n_14157 ^ x289;
assign n_14171 = ~n_14157 & n_14158;
assign n_14172 = n_14159 ^ n_12438;
assign n_14173 = n_14161 ^ n_12438;
assign n_14174 = n_14159 ^ n_14161;
assign n_14175 = n_13681 ^ n_14162;
assign n_14176 = n_14162 ^ n_14163;
assign n_14177 = n_13681 ^ n_14163;
assign n_14178 = n_14165 ^ n_14166;
assign n_14179 = n_14166 ^ x146;
assign n_14180 = n_14167 ^ n_12083;
assign n_14181 = n_14168 ^ n_13385;
assign n_14182 = n_13161 ^ n_14169;
assign n_14183 = ~n_14169 & n_13431;
assign n_14184 = n_14141 & ~n_14170;
assign n_14185 = n_14170 ^ n_14141;
assign n_14186 = n_14171 ^ x289;
assign n_14187 = n_14172 ^ n_14161;
assign n_14188 = n_14173 & ~n_14174;
assign n_14189 = n_14175 ^ n_14163;
assign n_14190 = ~n_13104 & n_14176;
assign n_14191 = ~n_14176 & ~n_14177;
assign n_14192 = n_14178 ^ x146;
assign n_14193 = n_14178 & ~n_14179;
assign n_14194 = n_14180 ^ n_12104;
assign n_14195 = n_14181 ^ n_12104;
assign n_14196 = n_14180 ^ n_14181;
assign n_14197 = n_14182 ^ n_13418;
assign n_14198 = n_14182 ^ n_13539;
assign n_14199 = n_14183 ^ n_13161;
assign n_14200 = n_14186 ^ n_14187;
assign n_14201 = n_14187 ^ x288;
assign n_14202 = n_14188 ^ n_12438;
assign n_14203 = n_14057 ^ n_14189;
assign n_14204 = n_14190 ^ n_13681;
assign n_14205 = n_14191 ^ n_13681;
assign n_14206 = n_14164 ^ n_14192;
assign n_14207 = ~n_14192 & ~n_14164;
assign n_14208 = n_14193 ^ x146;
assign n_14209 = n_14194 ^ n_14181;
assign n_14210 = n_14195 & ~n_14196;
assign n_14211 = ~n_12762 & n_14197;
assign n_14212 = n_14199 ^ n_13457;
assign n_14213 = n_14199 ^ n_13444;
assign n_14214 = n_14200 ^ x288;
assign n_14215 = n_14200 & ~n_14201;
assign n_14216 = n_14202 ^ n_12453;
assign n_14217 = n_14204 ^ n_12453;
assign n_14218 = n_14202 ^ n_14204;
assign n_14219 = n_13723 ^ n_14205;
assign n_14220 = n_14205 ^ n_14206;
assign n_14221 = n_13723 ^ n_14206;
assign n_14222 = n_14208 ^ n_14209;
assign n_14223 = n_14209 ^ x145;
assign n_14224 = n_14210 ^ n_12104;
assign n_14225 = n_14211 ^ n_13418;
assign n_14226 = n_14212 ^ n_13444;
assign n_14227 = n_14212 ^ n_13593;
assign n_14228 = ~n_13457 & n_14213;
assign n_14229 = n_14214 & n_14184;
assign n_14230 = n_14184 ^ n_14214;
assign n_14231 = n_14215 ^ x288;
assign n_14232 = n_14216 ^ n_14204;
assign n_14233 = n_14217 & n_14218;
assign n_14234 = n_14219 ^ n_14206;
assign n_14235 = ~n_13116 & n_14220;
assign n_14236 = ~n_14220 & ~n_14221;
assign n_14237 = n_14222 ^ x145;
assign n_14238 = ~n_14222 & n_14223;
assign n_14239 = n_14224 ^ n_12124;
assign n_14240 = n_14225 ^ n_12124;
assign n_14241 = n_14224 ^ n_14225;
assign n_14242 = n_12785 & n_14226;
assign n_14243 = n_14228 ^ n_13186;
assign n_14244 = n_14231 ^ n_14232;
assign n_14245 = n_14232 ^ x303;
assign n_14246 = n_14233 ^ n_12453;
assign n_14247 = n_14099 ^ n_14234;
assign n_14248 = n_14235 ^ n_13723;
assign n_14249 = n_14236 ^ n_13723;
assign n_14250 = n_14237 ^ n_14207;
assign n_14251 = ~n_14207 & ~n_14237;
assign n_14252 = n_14238 ^ x145;
assign n_14253 = n_14239 ^ n_14225;
assign n_14254 = n_14240 & n_14241;
assign n_14255 = n_14242 ^ n_13444;
assign n_14256 = n_14243 ^ n_13208;
assign n_14257 = n_14243 ^ n_13495;
assign n_14258 = n_14244 ^ x303;
assign n_14259 = n_14244 & ~n_14245;
assign n_14260 = n_14246 ^ n_12470;
assign n_14261 = n_14248 ^ n_12470;
assign n_14262 = n_14246 ^ n_14248;
assign n_14263 = n_13763 ^ n_14249;
assign n_14264 = n_14249 ^ n_14250;
assign n_14265 = n_13763 ^ n_14250;
assign n_14266 = n_14252 ^ n_14253;
assign n_14267 = n_14253 ^ x144;
assign n_14268 = n_14254 ^ n_12124;
assign n_14269 = n_14255 ^ n_12140;
assign n_14270 = n_14256 ^ n_13495;
assign n_14271 = ~n_13509 & n_14257;
assign n_14272 = n_14229 & n_14258;
assign n_14273 = n_14258 ^ n_14229;
assign n_14274 = n_14259 ^ x303;
assign n_14275 = n_14260 ^ n_14248;
assign n_14276 = ~n_14261 & n_14262;
assign n_14277 = n_14263 ^ n_14250;
assign n_14278 = n_13140 & n_14264;
assign n_14279 = ~n_14264 & n_14265;
assign n_14280 = n_14266 ^ x144;
assign n_14281 = ~n_14266 & n_14267;
assign n_14282 = n_14268 ^ n_14255;
assign n_14283 = n_14268 ^ n_14269;
assign n_14284 = n_14270 ^ n_13482;
assign n_14285 = n_14270 ^ n_13635;
assign n_14286 = n_14271 ^ n_13208;
assign n_14287 = n_14274 ^ n_14275;
assign n_14288 = n_14275 ^ x302;
assign n_14289 = n_14276 ^ n_12470;
assign n_14290 = n_14142 ^ n_14277;
assign n_14291 = n_14278 ^ n_13763;
assign n_14292 = n_14279 ^ n_13763;
assign n_14293 = n_14251 ^ n_14280;
assign n_14294 = ~n_14280 & n_14251;
assign n_14295 = n_14281 ^ x144;
assign n_14296 = ~n_14269 & n_14282;
assign n_14297 = n_14283 ^ x159;
assign n_14298 = ~n_12806 & ~n_14284;
assign n_14299 = n_14286 ^ n_13230;
assign n_14300 = n_14286 ^ n_13536;
assign n_14301 = n_14287 ^ x302;
assign n_14302 = n_14287 & ~n_14288;
assign n_14303 = n_14289 ^ n_12489;
assign n_14304 = n_14291 ^ n_12489;
assign n_14305 = n_14289 ^ n_14291;
assign n_14306 = n_13797 ^ n_14292;
assign n_14307 = n_14292 ^ n_14293;
assign n_14308 = n_13797 ^ n_14293;
assign n_14309 = n_14295 ^ x159;
assign n_14310 = n_14295 ^ n_14283;
assign n_14311 = n_14296 ^ n_12140;
assign n_14312 = n_14298 ^ n_13482;
assign n_14313 = n_14299 ^ n_13536;
assign n_14314 = ~n_13551 & n_14300;
assign n_14315 = ~n_14272 & ~n_14301;
assign n_14316 = n_14301 ^ n_14272;
assign n_14317 = n_14302 ^ x302;
assign n_14318 = n_14303 ^ n_14291;
assign n_14319 = ~n_14304 & n_14305;
assign n_14320 = n_14306 ^ n_14293;
assign n_14321 = n_13157 & ~n_14307;
assign n_14322 = n_14307 & n_14308;
assign n_14323 = n_14309 ^ n_14283;
assign n_14324 = n_14297 & ~n_14310;
assign n_14325 = n_14311 ^ n_14312;
assign n_14326 = n_14312 ^ n_12168;
assign n_14327 = n_14313 ^ n_13522;
assign n_14328 = n_13677 ^ n_14313;
assign n_14329 = n_14314 ^ n_13230;
assign n_14330 = n_14317 ^ n_14318;
assign n_14331 = n_14318 ^ x301;
assign n_14332 = n_14319 ^ n_12489;
assign n_14333 = n_14185 ^ n_14320;
assign n_14334 = n_14321 ^ n_13797;
assign n_14335 = n_14322 ^ n_13797;
assign n_14336 = n_14294 ^ n_14323;
assign n_14337 = ~n_14323 & n_14294;
assign n_14338 = n_14324 ^ x159;
assign n_14339 = n_14325 ^ n_12168;
assign n_14340 = ~n_14325 & ~n_14326;
assign n_14341 = n_12826 & n_14327;
assign n_14342 = n_14329 ^ n_13574;
assign n_14343 = n_14330 ^ x301;
assign n_14344 = n_14330 & ~n_14331;
assign n_14345 = n_14332 ^ n_12510;
assign n_14346 = n_14334 ^ n_12510;
assign n_14347 = n_14332 ^ n_14334;
assign n_14348 = n_14335 ^ n_13825;
assign n_14349 = n_14335 ^ n_14336;
assign n_14350 = n_14336 ^ n_13825;
assign n_14351 = n_14338 ^ n_14339;
assign n_14352 = n_14339 ^ x158;
assign n_14353 = n_14340 ^ n_12168;
assign n_14354 = n_14341 ^ n_13522;
assign n_14355 = n_13252 ^ n_14342;
assign n_14356 = n_14342 & ~n_13588;
assign n_14357 = n_14343 & ~n_14315;
assign n_14358 = n_14315 ^ n_14343;
assign n_14359 = n_14344 ^ x301;
assign n_14360 = n_14345 ^ n_14334;
assign n_14361 = ~n_14346 & ~n_14347;
assign n_14362 = n_14348 ^ n_14336;
assign n_14363 = ~n_13175 & n_14349;
assign n_14364 = ~n_14349 & n_14350;
assign n_14365 = n_14351 ^ x158;
assign n_14366 = ~n_14351 & n_14352;
assign n_14367 = n_14353 ^ n_12190;
assign n_14368 = n_14354 ^ n_12190;
assign n_14369 = n_14353 ^ n_14354;
assign n_14370 = n_14355 ^ n_13574;
assign n_14371 = n_13719 ^ n_14355;
assign n_14372 = n_14356 ^ n_13252;
assign n_14373 = n_14359 ^ n_14360;
assign n_14374 = n_14360 ^ x300;
assign n_14375 = n_14361 ^ n_12510;
assign n_14376 = n_14230 ^ n_14362;
assign n_14377 = n_14363 ^ n_13825;
assign n_14378 = n_14364 ^ n_13825;
assign n_14379 = n_14337 ^ n_14365;
assign n_14380 = ~n_14365 & n_14337;
assign n_14381 = n_14366 ^ x158;
assign n_14382 = n_14367 ^ n_14354;
assign n_14383 = ~n_14368 & ~n_14369;
assign n_14384 = n_12851 & n_14370;
assign n_14385 = n_14372 ^ n_13615;
assign n_14386 = n_14373 ^ x300;
assign n_14387 = n_14373 & ~n_14374;
assign n_14388 = n_14375 ^ n_12531;
assign n_14389 = n_14377 ^ n_12531;
assign n_14390 = n_14375 ^ n_14377;
assign n_14391 = n_13845 ^ n_14378;
assign n_14392 = n_14378 ^ n_14379;
assign n_14393 = n_13845 ^ n_14379;
assign n_14394 = n_14381 ^ n_14382;
assign n_14395 = n_14382 ^ x157;
assign n_14396 = n_14383 ^ n_12190;
assign n_14397 = n_14384 ^ n_13574;
assign n_14398 = n_13274 ^ n_14385;
assign n_14399 = n_14385 & ~n_13630;
assign n_14400 = n_14357 & n_14386;
assign n_14401 = n_14386 ^ n_14357;
assign n_14402 = n_14387 ^ x300;
assign n_14403 = n_14388 ^ n_14377;
assign n_14404 = ~n_14389 & n_14390;
assign n_14405 = n_14391 ^ n_14379;
assign n_14406 = ~n_13193 & n_14392;
assign n_14407 = ~n_14392 & n_14393;
assign n_14408 = n_14394 ^ x157;
assign n_14409 = n_14394 & ~n_14395;
assign n_14410 = n_14396 ^ n_12209;
assign n_14411 = n_14397 ^ n_12209;
assign n_14412 = n_14396 ^ n_14397;
assign n_14413 = n_14398 ^ n_13615;
assign n_14414 = n_13759 ^ n_14398;
assign n_14415 = n_14399 ^ n_13274;
assign n_14416 = n_14402 ^ n_14403;
assign n_14417 = n_14403 ^ x299;
assign n_14418 = n_14404 ^ n_12531;
assign n_14419 = n_14273 ^ n_14405;
assign n_14420 = n_14406 ^ n_13845;
assign n_14421 = n_14407 ^ n_13845;
assign n_14422 = n_14408 ^ n_14380;
assign n_14423 = n_14380 & n_14408;
assign n_14424 = n_14409 ^ x157;
assign n_14425 = n_14410 ^ n_14397;
assign n_14426 = ~n_14411 & n_14412;
assign n_14427 = ~n_12884 & n_14413;
assign n_14428 = n_14415 ^ n_13657;
assign n_14429 = n_14416 ^ x299;
assign n_14430 = ~n_14416 & n_14417;
assign n_14431 = n_14418 ^ n_12552;
assign n_14432 = n_14420 ^ n_12552;
assign n_14433 = n_14418 ^ n_14420;
assign n_14434 = n_13856 ^ n_14421;
assign n_14435 = n_14421 ^ n_14422;
assign n_14436 = n_13856 ^ n_14422;
assign n_14437 = n_14424 ^ n_14425;
assign n_14438 = n_14425 ^ x156;
assign n_14439 = n_14426 ^ n_12209;
assign n_14440 = n_14427 ^ n_13615;
assign n_14441 = n_13295 ^ n_14428;
assign n_14442 = n_14428 & n_13672;
assign n_14443 = ~n_14400 & n_14429;
assign n_14444 = n_14429 ^ n_14400;
assign n_14445 = n_14430 ^ x299;
assign n_14446 = n_14431 ^ n_14420;
assign n_14447 = ~n_14432 & n_14433;
assign n_14448 = n_14434 ^ n_14422;
assign n_14449 = n_13211 & ~n_14435;
assign n_14450 = n_14435 & n_14436;
assign n_14451 = n_14437 ^ x156;
assign n_14452 = ~n_14437 & n_14438;
assign n_14453 = n_14439 ^ n_12229;
assign n_14454 = n_14440 ^ n_12229;
assign n_14455 = n_14439 ^ n_14440;
assign n_14456 = n_14441 ^ n_13657;
assign n_14457 = n_14441 ^ n_13793;
assign n_14458 = n_14442 ^ n_13295;
assign n_14459 = n_14445 ^ n_14446;
assign n_14460 = n_14446 ^ x298;
assign n_14461 = n_14447 ^ n_12552;
assign n_14462 = n_14448 ^ n_14316;
assign n_14463 = n_14449 ^ n_13856;
assign n_14464 = n_14450 ^ n_13856;
assign n_14465 = n_14451 ^ n_14423;
assign n_14466 = ~n_14423 & n_14451;
assign n_14467 = n_14452 ^ x156;
assign n_14468 = n_14453 ^ n_14440;
assign n_14469 = n_14454 & n_14455;
assign n_14470 = ~n_12922 & ~n_14456;
assign n_14471 = n_14458 ^ n_13699;
assign n_14472 = n_14459 ^ x298;
assign n_14473 = ~n_14459 & n_14460;
assign n_14474 = n_14461 ^ n_12573;
assign n_14475 = n_14463 ^ n_14461;
assign n_14476 = n_14464 ^ n_13879;
assign n_14477 = n_14464 ^ n_14465;
assign n_14478 = n_14465 ^ n_13879;
assign n_14479 = n_14467 ^ n_14468;
assign n_14480 = n_14468 ^ x155;
assign n_14481 = n_14469 ^ n_12229;
assign n_14482 = n_14470 ^ n_13657;
assign n_14483 = n_13315 ^ n_14471;
assign n_14484 = ~n_14471 & n_13714;
assign n_14485 = n_14443 & n_14472;
assign n_14486 = n_14472 ^ n_14443;
assign n_14487 = n_14473 ^ x298;
assign n_14488 = n_14463 ^ n_14474;
assign n_14489 = n_14474 & ~n_14475;
assign n_14490 = n_14476 ^ n_14465;
assign n_14491 = ~n_13231 & n_14477;
assign n_14492 = ~n_14477 & ~n_14478;
assign n_14493 = n_14479 ^ x155;
assign n_14494 = n_14479 & ~n_14480;
assign n_14495 = n_14481 ^ n_12250;
assign n_14496 = n_14482 ^ n_12250;
assign n_14497 = n_14481 ^ n_14482;
assign n_14498 = n_14483 ^ n_13699;
assign n_14499 = n_13821 ^ n_14483;
assign n_14500 = n_14484 ^ n_13315;
assign n_14501 = n_14487 ^ n_14488;
assign n_14502 = n_14488 ^ x297;
assign n_14503 = n_14489 ^ n_12573;
assign n_14504 = n_14490 ^ n_14358;
assign n_14505 = n_14491 ^ n_13879;
assign n_14506 = n_14492 ^ n_13879;
assign n_14507 = n_14493 ^ n_14466;
assign n_14508 = n_14466 & ~n_14493;
assign n_14509 = n_14494 ^ x155;
assign n_14510 = n_14495 ^ n_14482;
assign n_14511 = n_14496 & ~n_14497;
assign n_14512 = n_12960 & n_14498;
assign n_14513 = n_14500 ^ n_13742;
assign n_14514 = n_14501 ^ x297;
assign n_14515 = n_14501 & ~n_14502;
assign n_14516 = n_14503 ^ n_12595;
assign n_14517 = n_14505 ^ n_12595;
assign n_14518 = n_14503 ^ n_14505;
assign n_14519 = n_14506 ^ n_13906;
assign n_14520 = n_13906 ^ n_14507;
assign n_14521 = n_14506 ^ n_14507;
assign n_14522 = n_14509 ^ n_14510;
assign n_14523 = n_14510 ^ x154;
assign n_14524 = n_14511 ^ n_12250;
assign n_14525 = n_14512 ^ n_13699;
assign n_14526 = n_14513 ^ n_13729;
assign n_14527 = n_14513 ^ n_13820;
assign n_14528 = ~n_14485 & n_14514;
assign n_14529 = n_14514 ^ n_14485;
assign n_14530 = n_14515 ^ x297;
assign n_14531 = n_14516 ^ n_14505;
assign n_14532 = n_14517 & n_14518;
assign n_14533 = n_14519 ^ n_14507;
assign n_14534 = ~n_14520 & n_14521;
assign n_14535 = n_14522 ^ x154;
assign n_14536 = ~n_14522 & n_14523;
assign n_14537 = n_14524 ^ n_12273;
assign n_14538 = n_14525 ^ n_12273;
assign n_14539 = n_14525 ^ n_14524;
assign n_14540 = ~n_12989 & ~n_14526;
assign n_14541 = n_14527 ^ n_13834;
assign n_14542 = n_14530 ^ n_14531;
assign n_14543 = n_14531 ^ x296;
assign n_14544 = n_14532 ^ n_12595;
assign n_14545 = n_14533 ^ n_13895;
assign n_14546 = n_14401 ^ n_14533;
assign n_14547 = n_14534 ^ n_13906;
assign n_14548 = n_14535 ^ n_14508;
assign n_14549 = ~n_14508 & ~n_14535;
assign n_14550 = n_14536 ^ x154;
assign n_14551 = n_14525 ^ n_14537;
assign n_14552 = ~n_14538 & ~n_14539;
assign n_14553 = n_14540 ^ n_13729;
assign n_14554 = n_14542 ^ x296;
assign n_14555 = n_14542 & ~n_14543;
assign n_14556 = ~n_13246 & n_14545;
assign n_14557 = n_14547 ^ n_13939;
assign n_14558 = n_14548 ^ n_13939;
assign n_14559 = n_14547 ^ n_14548;
assign n_14560 = n_14550 ^ n_14551;
assign n_14561 = n_14551 ^ x153;
assign n_14562 = n_14552 ^ n_12273;
assign n_14563 = n_14553 ^ n_12292;
assign n_14564 = n_14528 & n_14554;
assign n_14565 = n_14554 ^ n_14528;
assign n_14566 = n_14555 ^ x296;
assign n_14567 = n_14556 ^ n_13895;
assign n_14568 = n_14557 ^ n_14548;
assign n_14569 = ~n_14558 & n_14559;
assign n_14570 = n_14560 ^ x153;
assign n_14571 = n_14560 & ~n_14561;
assign n_14572 = n_14562 ^ x152;
assign n_14573 = n_14566 ^ x311;
assign n_14574 = n_14544 ^ n_14567;
assign n_14575 = n_14567 ^ n_12608;
assign n_14576 = n_14568 ^ n_13929;
assign n_14577 = n_14444 ^ n_14568;
assign n_14578 = n_14569 ^ n_13939;
assign n_14579 = n_14570 ^ n_14549;
assign n_14580 = n_14549 & n_14570;
assign n_14581 = n_14571 ^ x153;
assign n_14582 = n_14572 ^ n_14563;
assign n_14583 = n_14574 ^ n_12608;
assign n_14584 = n_14574 & n_14575;
assign n_14585 = ~n_13276 & n_14576;
assign n_14586 = n_14578 ^ n_13975;
assign n_14587 = n_14578 ^ n_14579;
assign n_14588 = n_14579 ^ n_13975;
assign n_14589 = n_14581 ^ n_14582;
assign n_14590 = n_14583 ^ x311;
assign n_14591 = n_14566 ^ n_14583;
assign n_14592 = n_14573 ^ n_14583;
assign n_14593 = n_14584 ^ n_12608;
assign n_14594 = n_14585 ^ n_13929;
assign n_14595 = n_14586 ^ n_14579;
assign n_14596 = ~n_13297 & ~n_14587;
assign n_14597 = n_14587 & n_14588;
assign n_14598 = n_14589 ^ n_14580;
assign n_14599 = n_14590 & ~n_14591;
assign n_14600 = n_14564 & ~n_14592;
assign n_14601 = n_14592 ^ n_14564;
assign n_14602 = n_14593 ^ n_12639;
assign n_14603 = n_14594 ^ n_12639;
assign n_14604 = n_14593 ^ n_14594;
assign n_14605 = n_14486 ^ n_14595;
assign n_14606 = n_14596 ^ n_13975;
assign n_14607 = n_14597 ^ n_13975;
assign n_14608 = n_14015 ^ n_14598;
assign n_14609 = n_14599 ^ x311;
assign n_14610 = n_14602 ^ n_14594;
assign n_14611 = ~n_14603 & ~n_14604;
assign n_14612 = n_14606 ^ n_12659;
assign n_14613 = n_14607 ^ n_14015;
assign n_14614 = n_14607 ^ n_14598;
assign n_14615 = n_14609 ^ n_14610;
assign n_14616 = n_14610 ^ x310;
assign n_14617 = n_14611 ^ n_12639;
assign n_14618 = n_14613 ^ n_14598;
assign n_14619 = ~n_14608 & n_14614;
assign n_14620 = n_14615 ^ x310;
assign n_14621 = ~n_14615 & n_14616;
assign n_14622 = n_14617 ^ n_12659;
assign n_14623 = n_14617 ^ n_14606;
assign n_14624 = n_14618 ^ n_14000;
assign n_14625 = n_14529 ^ n_14618;
assign n_14626 = n_14619 ^ n_14015;
assign n_14627 = ~n_14600 & n_14620;
assign n_14628 = n_14620 ^ n_14600;
assign n_14629 = n_14621 ^ x310;
assign n_14630 = n_14622 ^ n_14606;
assign n_14631 = ~n_14612 & n_14623;
assign n_14632 = ~n_13317 & n_14624;
assign n_14633 = n_14626 ^ n_14054;
assign n_14634 = n_14629 ^ n_14630;
assign n_14635 = n_14630 ^ x309;
assign n_14636 = n_14631 ^ n_12659;
assign n_14637 = n_14632 ^ n_14000;
assign n_14638 = n_13410 ^ n_14633;
assign n_14639 = n_14633 & n_14069;
assign n_14640 = n_14634 ^ x309;
assign n_14641 = n_14634 & ~n_14635;
assign n_14642 = n_14636 ^ n_12678;
assign n_14643 = n_14637 ^ n_12678;
assign n_14644 = n_14636 ^ n_14637;
assign n_14645 = n_14638 ^ n_14054;
assign n_14646 = n_14565 ^ n_14638;
assign n_14647 = n_14639 ^ n_13410;
assign n_14648 = n_14627 & ~n_14640;
assign n_14649 = n_14640 ^ n_14627;
assign n_14650 = n_14641 ^ x309;
assign n_14651 = n_14642 ^ n_14637;
assign n_14652 = ~n_14643 & ~n_14644;
assign n_14653 = n_13338 & ~n_14645;
assign n_14654 = n_14647 ^ n_14096;
assign n_14655 = n_14650 ^ n_14651;
assign n_14656 = n_14651 ^ x308;
assign n_14657 = n_14652 ^ n_12678;
assign n_14658 = n_14653 ^ n_14054;
assign n_14659 = n_13436 ^ n_14654;
assign n_14660 = n_14654 & n_14112;
assign n_14661 = n_14655 ^ x308;
assign n_14662 = n_14655 & ~n_14656;
assign n_14663 = n_14657 ^ n_12700;
assign n_14664 = n_14658 ^ n_12700;
assign n_14665 = n_14657 ^ n_14658;
assign n_14666 = n_14659 ^ n_14096;
assign n_14667 = n_14601 ^ n_14659;
assign n_14668 = n_14660 ^ n_13436;
assign n_14669 = n_14648 & ~n_14661;
assign n_14670 = n_14661 ^ n_14648;
assign n_14671 = n_14662 ^ x308;
assign n_14672 = n_14663 ^ n_14658;
assign n_14673 = ~n_14664 & n_14665;
assign n_14674 = n_13359 & ~n_14666;
assign n_14675 = n_14668 ^ n_14139;
assign n_14676 = n_14671 ^ n_14672;
assign n_14677 = n_14672 ^ x307;
assign n_14678 = n_14673 ^ n_12700;
assign n_14679 = n_14674 ^ n_14096;
assign n_14680 = n_13499 ^ n_14675;
assign n_14681 = ~n_14675 & n_14155;
assign n_14682 = n_14676 ^ x307;
assign n_14683 = ~n_14676 & n_14677;
assign n_14684 = n_14678 ^ n_14679;
assign n_14685 = n_14679 ^ n_12721;
assign n_14686 = n_14680 ^ n_14139;
assign n_14687 = n_14628 ^ n_14680;
assign n_14688 = n_14681 ^ n_13499;
assign n_14689 = n_14669 & n_14682;
assign n_14690 = n_14682 ^ n_14669;
assign n_14691 = n_14683 ^ x307;
assign n_14692 = n_14684 ^ n_12721;
assign n_14693 = ~n_14684 & ~n_14685;
assign n_14694 = n_13385 & n_14686;
assign n_14695 = n_14688 ^ n_14198;
assign n_14696 = n_14688 ^ n_14182;
assign n_14697 = n_14691 ^ n_14692;
assign n_14698 = n_14692 ^ x306;
assign n_14699 = n_14693 ^ n_12721;
assign n_14700 = n_14694 ^ n_14139;
assign n_14701 = n_14695 ^ n_14182;
assign n_14702 = n_14649 ^ n_14695;
assign n_14703 = ~n_14198 & ~n_14696;
assign n_14704 = n_14697 ^ x306;
assign n_14705 = ~n_14697 & n_14698;
assign n_14706 = n_14699 ^ n_12741;
assign n_14707 = n_14700 ^ n_12741;
assign n_14708 = n_14699 ^ n_14700;
assign n_14709 = ~n_13418 & ~n_14701;
assign n_14710 = n_14703 ^ n_13539;
assign n_14711 = ~n_14689 & ~n_14704;
assign n_14712 = n_14704 ^ n_14689;
assign n_14713 = n_14705 ^ x306;
assign n_14714 = n_14706 ^ n_14700;
assign n_14715 = ~n_14707 & n_14708;
assign n_14716 = n_14709 ^ n_14182;
assign n_14717 = n_14710 ^ n_14227;
assign n_14718 = n_14710 ^ n_14212;
assign n_14719 = n_14713 ^ n_14714;
assign n_14720 = n_14714 ^ x305;
assign n_14721 = n_14715 ^ n_12741;
assign n_14722 = n_14717 ^ n_14212;
assign n_14723 = n_14670 ^ n_14717;
assign n_14724 = ~n_14227 & ~n_14718;
assign n_14725 = n_14719 ^ x305;
assign n_14726 = n_14719 & ~n_14720;
assign n_14727 = n_14721 ^ n_12762;
assign n_14728 = n_14716 ^ n_14721;
assign n_14729 = n_13444 & ~n_14722;
assign n_14730 = n_14724 ^ n_13593;
assign n_14731 = n_14711 & n_14725;
assign n_14732 = n_14725 ^ n_14711;
assign n_14733 = n_14726 ^ x305;
assign n_14734 = n_14716 ^ n_14727;
assign n_14735 = ~n_14727 & n_14728;
assign n_14736 = n_14729 ^ n_14212;
assign n_14737 = n_14730 ^ n_13635;
assign n_14738 = n_14730 ^ n_14270;
assign n_14739 = n_14733 ^ n_14734;
assign n_14740 = n_14734 ^ x304;
assign n_14741 = n_14735 ^ n_12762;
assign n_14742 = n_14736 ^ n_12785;
assign n_14743 = n_14737 ^ n_14270;
assign n_14744 = ~n_14285 & n_14738;
assign n_14745 = n_14739 ^ x304;
assign n_14746 = ~n_14739 & n_14740;
assign n_14747 = n_14741 ^ n_14736;
assign n_14748 = n_14741 ^ n_14742;
assign n_14749 = n_14743 ^ n_14256;
assign n_14750 = n_14690 ^ n_14743;
assign n_14751 = n_14744 ^ n_13635;
assign n_14752 = n_14731 & ~n_14745;
assign n_14753 = n_14745 ^ n_14731;
assign n_14754 = n_14746 ^ x304;
assign n_14755 = n_14742 & n_14747;
assign n_14756 = n_13495 & n_14749;
assign n_14757 = n_14751 ^ n_14313;
assign n_14758 = n_14754 ^ x319;
assign n_14759 = n_14748 ^ n_14754;
assign n_14760 = n_14755 ^ n_12785;
assign n_14761 = n_14756 ^ n_14256;
assign n_14762 = n_13677 ^ n_14757;
assign n_14763 = n_14757 & n_14328;
assign n_14764 = n_14748 ^ n_14758;
assign n_14765 = n_14758 & n_14759;
assign n_14766 = n_14760 ^ n_14761;
assign n_14767 = n_14761 ^ n_12806;
assign n_14768 = n_14762 ^ n_14299;
assign n_14769 = n_14712 ^ n_14762;
assign n_14770 = n_14763 ^ n_13677;
assign n_14771 = n_14752 & n_14764;
assign n_14772 = n_14764 ^ n_14752;
assign n_14773 = n_14765 ^ x319;
assign n_14774 = n_14766 ^ n_12806;
assign n_14775 = ~n_14766 & ~n_14767;
assign n_14776 = n_13536 & ~n_14768;
assign n_14777 = n_14770 ^ n_14355;
assign n_14778 = n_14773 ^ n_14774;
assign n_14779 = n_14774 ^ x318;
assign n_14780 = n_14775 ^ n_12806;
assign n_14781 = n_14776 ^ n_14299;
assign n_14782 = n_13719 ^ n_14777;
assign n_14783 = ~n_14777 & n_14371;
assign n_14784 = n_14778 ^ x318;
assign n_14785 = n_14778 & ~n_14779;
assign n_14786 = n_14780 ^ n_14781;
assign n_14787 = n_14781 ^ n_12826;
assign n_14788 = n_14782 ^ n_14355;
assign n_14789 = n_14732 ^ n_14782;
assign n_14790 = n_14783 ^ n_13719;
assign n_14791 = ~n_14771 & ~n_14784;
assign n_14792 = n_14784 ^ n_14771;
assign n_14793 = n_14785 ^ x318;
assign n_14794 = n_14786 ^ n_12826;
assign n_14795 = n_14786 & n_14787;
assign n_14796 = n_13574 & n_14788;
assign n_14797 = n_14790 ^ n_14398;
assign n_14798 = n_14793 ^ n_14794;
assign n_14799 = n_14794 ^ x317;
assign n_14800 = n_14795 ^ n_12826;
assign n_14801 = n_14796 ^ n_14355;
assign n_14802 = n_13759 ^ n_14797;
assign n_14803 = ~n_14797 & ~n_14414;
assign n_14804 = n_14798 ^ x317;
assign n_14805 = n_14798 & ~n_14799;
assign n_14806 = n_14800 ^ n_12851;
assign n_14807 = n_14801 ^ n_12851;
assign n_14808 = n_14800 ^ n_14801;
assign n_14809 = n_14802 ^ n_14398;
assign n_14810 = n_14753 ^ n_14802;
assign n_14811 = n_14803 ^ n_13759;
assign n_14812 = ~n_14804 & n_14791;
assign n_14813 = n_14791 ^ n_14804;
assign n_14814 = n_14805 ^ x317;
assign n_14815 = n_14806 ^ n_14801;
assign n_14816 = n_14807 & ~n_14808;
assign n_14817 = n_13615 & ~n_14809;
assign n_14818 = n_14811 ^ n_14441;
assign n_14819 = n_14814 ^ n_14815;
assign n_14820 = n_14815 ^ x316;
assign n_14821 = n_14816 ^ n_12851;
assign n_14822 = n_14817 ^ n_14398;
assign n_14823 = n_14818 ^ n_13793;
assign n_14824 = ~n_14818 & ~n_14457;
assign n_14825 = n_14819 ^ x316;
assign n_14826 = ~n_14819 & n_14820;
assign n_14827 = n_14821 ^ n_12884;
assign n_14828 = n_14822 ^ n_12884;
assign n_14829 = n_14821 ^ n_14822;
assign n_14830 = n_14823 ^ n_14441;
assign n_14831 = n_14772 ^ n_14823;
assign n_14832 = n_14824 ^ n_13793;
assign n_14833 = n_14825 ^ n_14812;
assign n_14834 = n_14812 & n_14825;
assign n_14835 = n_14826 ^ x316;
assign n_14836 = n_14827 ^ n_14822;
assign n_14837 = ~n_14828 & ~n_14829;
assign n_14838 = n_13657 & ~n_14830;
assign n_14839 = n_14832 ^ n_14483;
assign n_14840 = n_14833 ^ n_13870;
assign n_14841 = n_13870 & n_14833;
assign n_14842 = n_14835 ^ n_14836;
assign n_14843 = n_14836 ^ x315;
assign n_14844 = n_14837 ^ n_12884;
assign n_14845 = n_14838 ^ n_14441;
assign n_14846 = n_14839 ^ n_13821;
assign n_14847 = ~n_14839 & n_14499;
assign n_14848 = n_14840 ^ n_13863;
assign n_14849 = n_14840 ^ x423;
assign n_14850 = n_13900 ^ n_14841;
assign n_14851 = n_14842 ^ x315;
assign n_14852 = n_14842 & ~n_14843;
assign n_14853 = n_14844 ^ n_12922;
assign n_14854 = n_14845 ^ n_12922;
assign n_14855 = n_14844 ^ n_14845;
assign n_14856 = n_14846 ^ n_14483;
assign n_14857 = n_14792 ^ n_14846;
assign n_14858 = n_14847 ^ n_13821;
assign n_14859 = ~n_13363 & ~n_14848;
assign n_14860 = n_14834 ^ n_14851;
assign n_14861 = ~n_14851 & n_14834;
assign n_14862 = n_14852 ^ x315;
assign n_14863 = n_14853 ^ n_14845;
assign n_14864 = n_14854 & ~n_14855;
assign n_14865 = n_13699 & n_14856;
assign n_14866 = n_14858 ^ n_14541;
assign n_14867 = n_14859 ^ n_13863;
assign n_14868 = n_14860 ^ n_14841;
assign n_14869 = n_14850 ^ n_14860;
assign n_14870 = n_14862 ^ n_14863;
assign n_14871 = n_14863 ^ x314;
assign n_14872 = n_14864 ^ n_12922;
assign n_14873 = n_14865 ^ n_14483;
assign n_14874 = n_14866 ^ n_14513;
assign n_14875 = n_14867 ^ n_12832;
assign n_14876 = ~n_12832 & ~n_14867;
assign n_14877 = n_13391 & ~n_14868;
assign n_14878 = n_14868 & ~n_14850;
assign n_14879 = n_14870 ^ x314;
assign n_14880 = n_14870 & ~n_14871;
assign n_14881 = n_14872 ^ n_12960;
assign n_14882 = n_14873 ^ n_12960;
assign n_14883 = n_14873 ^ n_14872;
assign n_14884 = n_13729 & n_14874;
assign n_14885 = x455 & n_14875;
assign n_14886 = n_14875 ^ x455;
assign n_14887 = n_14876 ^ n_12856;
assign n_14888 = n_14877 ^ n_13900;
assign n_14889 = n_14878 ^ n_13900;
assign n_14890 = n_14879 ^ n_14861;
assign n_14891 = ~n_14861 & n_14879;
assign n_14892 = n_14880 ^ x314;
assign n_14893 = n_14873 ^ n_14881;
assign n_14894 = n_14882 & n_14883;
assign n_14895 = n_14884 ^ n_14513;
assign n_14896 = n_14885 ^ x454;
assign n_14897 = n_14888 ^ n_14887;
assign n_14898 = n_14888 ^ n_14876;
assign n_14899 = n_13941 ^ n_14889;
assign n_14900 = n_14889 ^ n_14890;
assign n_14901 = n_13941 ^ n_14890;
assign n_14902 = n_14892 ^ n_14893;
assign n_14903 = n_14893 ^ x313;
assign n_14904 = n_14894 ^ n_12960;
assign n_14905 = n_14895 ^ n_12989;
assign n_14906 = n_14897 ^ n_14885;
assign n_14907 = n_14897 ^ n_14896;
assign n_14908 = n_14887 & n_14898;
assign n_14909 = n_14899 ^ n_14890;
assign n_14910 = ~n_13438 & ~n_14900;
assign n_14911 = n_14900 & ~n_14901;
assign n_14912 = n_14902 ^ x313;
assign n_14913 = n_14902 & ~n_14903;
assign n_14914 = n_14904 ^ x312;
assign n_14915 = n_14896 & n_14906;
assign n_14916 = n_14908 ^ n_12856;
assign n_14917 = n_14910 ^ n_13941;
assign n_14918 = n_14911 ^ n_13941;
assign n_14919 = n_14891 ^ n_14912;
assign n_14920 = ~n_14912 & ~n_14891;
assign n_14921 = n_14913 ^ x313;
assign n_14922 = n_14914 ^ n_14905;
assign n_14923 = n_14915 ^ x454;
assign n_14924 = n_14916 ^ n_12900;
assign n_14925 = n_14917 ^ n_12900;
assign n_14926 = n_14916 ^ n_14917;
assign n_14927 = n_13979 ^ n_14918;
assign n_14928 = n_14918 ^ n_14919;
assign n_14929 = n_13979 ^ n_14919;
assign n_14930 = n_14921 ^ n_14922;
assign n_14931 = n_14924 ^ n_14917;
assign n_14932 = ~n_14925 & n_14926;
assign n_14933 = n_14927 ^ n_14919;
assign n_14934 = ~n_13476 & ~n_14928;
assign n_14935 = n_14928 & ~n_14929;
assign n_14936 = n_14930 ^ n_14920;
assign n_14937 = n_14923 ^ n_14931;
assign n_14938 = n_14931 ^ x453;
assign n_14939 = n_14932 ^ n_12900;
assign n_14940 = n_14934 ^ n_13979;
assign n_14941 = n_14935 ^ n_13979;
assign n_14942 = n_14022 ^ n_14936;
assign n_14943 = n_14937 ^ x453;
assign n_14944 = n_14937 & ~n_14938;
assign n_14945 = n_14939 ^ n_12945;
assign n_14946 = n_14940 ^ n_12945;
assign n_14947 = n_14939 ^ n_14940;
assign n_14948 = n_14941 ^ n_14936;
assign n_14949 = n_14022 ^ n_14941;
assign n_14950 = n_14943 & n_14907;
assign n_14951 = n_14907 ^ n_14943;
assign n_14952 = n_14944 ^ x453;
assign n_14953 = n_14945 ^ n_14940;
assign n_14954 = n_14946 & n_14947;
assign n_14955 = n_13516 & ~n_14948;
assign n_14956 = n_14948 & n_14942;
assign n_14957 = n_14949 ^ n_14936;
assign n_14958 = n_14952 ^ n_14953;
assign n_14959 = n_14953 ^ x452;
assign n_14960 = n_14954 ^ n_12945;
assign n_14961 = n_14955 ^ n_14022;
assign n_14962 = n_14956 ^ n_14022;
assign n_14963 = n_14958 ^ x452;
assign n_14964 = ~n_14958 & n_14959;
assign n_14965 = n_14960 ^ n_12985;
assign n_14966 = n_14961 ^ n_12985;
assign n_14967 = n_14960 ^ n_14961;
assign n_14968 = n_14061 ^ n_14962;
assign n_14969 = n_14963 & ~n_14950;
assign n_14970 = n_14950 ^ n_14963;
assign n_14971 = n_14964 ^ x452;
assign n_14972 = n_14965 ^ n_14961;
assign n_14973 = n_14966 & n_14967;
assign n_14974 = n_13910 ^ n_14968;
assign n_14975 = ~n_14968 & ~n_14074;
assign n_14976 = n_14971 ^ n_14972;
assign n_14977 = n_14972 ^ x451;
assign n_14978 = n_14973 ^ n_12985;
assign n_14979 = n_14974 ^ n_14061;
assign n_14980 = n_14975 ^ n_13910;
assign n_14981 = n_14976 ^ x451;
assign n_14982 = n_14976 & ~n_14977;
assign n_14983 = n_14978 ^ n_13022;
assign n_14984 = n_13557 & ~n_14979;
assign n_14985 = n_14980 ^ n_13944;
assign n_14986 = n_14103 ^ n_14980;
assign n_14987 = ~n_14969 & n_14981;
assign n_14988 = n_14981 ^ n_14969;
assign n_14989 = n_14982 ^ x451;
assign n_14990 = n_14984 ^ n_14061;
assign n_14991 = ~n_13597 & n_14985;
assign n_14992 = ~n_14985 & ~n_14117;
assign n_14993 = n_14986 ^ n_13944;
assign n_14994 = n_14983 ^ n_14990;
assign n_14995 = n_14990 ^ n_13022;
assign n_14996 = n_14978 ^ n_14990;
assign n_14997 = n_14991 ^ n_14103;
assign n_14998 = n_14992 ^ n_14103;
assign n_14999 = n_14989 ^ n_14994;
assign n_15000 = n_14994 ^ x450;
assign n_15001 = n_14995 & ~n_14996;
assign n_15002 = n_14146 ^ n_14998;
assign n_15003 = n_14999 ^ x450;
assign n_15004 = ~n_14999 & n_15000;
assign n_15005 = n_15001 ^ n_13022;
assign n_15006 = n_14018 ^ n_15002;
assign n_15007 = ~n_15002 & ~n_14160;
assign n_15008 = n_15003 & ~n_14987;
assign n_15009 = n_14987 ^ n_15003;
assign n_15010 = n_15004 ^ x450;
assign n_15011 = n_15005 ^ n_13056;
assign n_15012 = n_14997 ^ n_15005;
assign n_15013 = n_15006 ^ n_14146;
assign n_15014 = n_15007 ^ n_14018;
assign n_15015 = n_14997 ^ n_15011;
assign n_15016 = n_15011 & ~n_15012;
assign n_15017 = ~n_13639 & ~n_15013;
assign n_15018 = n_14189 ^ n_15014;
assign n_15019 = n_15010 ^ n_15015;
assign n_15020 = n_15015 ^ x449;
assign n_15021 = n_15016 ^ n_13056;
assign n_15022 = n_15017 ^ n_14146;
assign n_15023 = n_15018 & ~n_14203;
assign n_15024 = n_14057 ^ n_15018;
assign n_15025 = n_15019 ^ x449;
assign n_15026 = ~n_15019 & n_15020;
assign n_15027 = n_15021 ^ n_13083;
assign n_15028 = n_15022 ^ n_13083;
assign n_15029 = n_15021 ^ n_15022;
assign n_15030 = n_15023 ^ n_14057;
assign n_15031 = n_15024 ^ n_14189;
assign n_15032 = ~n_15025 & ~n_15008;
assign n_15033 = n_15008 ^ n_15025;
assign n_15034 = n_15026 ^ x449;
assign n_15035 = n_15027 ^ n_15022;
assign n_15036 = n_15028 & ~n_15029;
assign n_15037 = n_14234 ^ n_15030;
assign n_15038 = n_13681 & n_15031;
assign n_15039 = n_15034 ^ n_15035;
assign n_15040 = n_15035 ^ x448;
assign n_15041 = n_15036 ^ n_13083;
assign n_15042 = ~n_15037 & ~n_14247;
assign n_15043 = n_14099 ^ n_15037;
assign n_15044 = n_15038 ^ n_14189;
assign n_15045 = n_15039 ^ x448;
assign n_15046 = ~n_15039 & n_15040;
assign n_15047 = n_15041 ^ n_13104;
assign n_15048 = n_15042 ^ n_14099;
assign n_15049 = n_15043 ^ n_14234;
assign n_15050 = n_14886 ^ n_15043;
assign n_15051 = n_15044 ^ n_13104;
assign n_15052 = n_15041 ^ n_15044;
assign n_15053 = n_15032 ^ n_15045;
assign n_15054 = ~n_15045 & n_15032;
assign n_15055 = n_15046 ^ x448;
assign n_15056 = n_15047 ^ n_15044;
assign n_15057 = n_14277 ^ n_15048;
assign n_15058 = ~n_13723 & ~n_15049;
assign n_15059 = ~n_15051 & ~n_15052;
assign n_15060 = n_15055 ^ n_15056;
assign n_15061 = n_15056 ^ x463;
assign n_15062 = n_15057 & n_14290;
assign n_15063 = n_14142 ^ n_15057;
assign n_15064 = n_15058 ^ n_14234;
assign n_15065 = n_15059 ^ n_13104;
assign n_15066 = n_15060 ^ x463;
assign n_15067 = n_15060 & ~n_15061;
assign n_15068 = n_15062 ^ n_14142;
assign n_15069 = n_15063 ^ n_14277;
assign n_15070 = n_14907 ^ n_15063;
assign n_15071 = n_15064 ^ n_13116;
assign n_15072 = n_15065 ^ n_15064;
assign n_15073 = n_15065 ^ n_13116;
assign n_15074 = n_15054 & n_15066;
assign n_15075 = n_15066 ^ n_15054;
assign n_15076 = n_15067 ^ x463;
assign n_15077 = n_14320 ^ n_15068;
assign n_15078 = ~n_13763 & ~n_15069;
assign n_15079 = n_15071 & ~n_15072;
assign n_15080 = n_15073 ^ n_15064;
assign n_15081 = ~n_15077 & ~n_14333;
assign n_15082 = n_14185 ^ n_15077;
assign n_15083 = n_15078 ^ n_14277;
assign n_15084 = n_15079 ^ n_13116;
assign n_15085 = n_15076 ^ n_15080;
assign n_15086 = n_15080 ^ x462;
assign n_15087 = n_15081 ^ n_14185;
assign n_15088 = n_15082 ^ n_14320;
assign n_15089 = n_14951 ^ n_15082;
assign n_15090 = n_15083 ^ n_13140;
assign n_15091 = n_15084 ^ n_15083;
assign n_15092 = n_15084 ^ n_13140;
assign n_15093 = n_15085 ^ x462;
assign n_15094 = n_15085 & ~n_15086;
assign n_15095 = n_14362 ^ n_15087;
assign n_15096 = n_13797 & ~n_15088;
assign n_15097 = ~n_15090 & ~n_15091;
assign n_15098 = n_15092 ^ n_15083;
assign n_15099 = n_15074 & n_15093;
assign n_15100 = n_15093 ^ n_15074;
assign n_15101 = n_15094 ^ x462;
assign n_15102 = ~n_15095 & ~n_14376;
assign n_15103 = n_14230 ^ n_15095;
assign n_15104 = n_15096 ^ n_14320;
assign n_15105 = n_15097 ^ n_13140;
assign n_15106 = n_15098 ^ x461;
assign n_15107 = n_15101 ^ n_15098;
assign n_15108 = n_15102 ^ n_14230;
assign n_15109 = n_15103 ^ n_14362;
assign n_15110 = n_14970 ^ n_15103;
assign n_15111 = n_15104 ^ n_13157;
assign n_15112 = n_15105 ^ n_15104;
assign n_15113 = n_15105 ^ n_13157;
assign n_15114 = ~n_15107 & n_15106;
assign n_15115 = n_15107 ^ x461;
assign n_15116 = n_14405 ^ n_15108;
assign n_15117 = n_13825 & ~n_15109;
assign n_15118 = ~n_15111 & n_15112;
assign n_15119 = n_15113 ^ n_15104;
assign n_15120 = n_15114 ^ x461;
assign n_15121 = n_15099 & ~n_15115;
assign n_15122 = n_15115 ^ n_15099;
assign n_15123 = n_15116 & ~n_14419;
assign n_15124 = n_14273 ^ n_15116;
assign n_15125 = n_15117 ^ n_14362;
assign n_15126 = n_15118 ^ n_13157;
assign n_15127 = n_15119 ^ x460;
assign n_15128 = n_15120 ^ n_15119;
assign n_15129 = n_15123 ^ n_14273;
assign n_15130 = n_15124 ^ n_14405;
assign n_15131 = n_14988 ^ n_15124;
assign n_15132 = n_15125 ^ n_13175;
assign n_15133 = n_15126 ^ n_15125;
assign n_15134 = n_15126 ^ n_13175;
assign n_15135 = n_15128 & ~n_15127;
assign n_15136 = n_15128 ^ x460;
assign n_15137 = n_14448 ^ n_15129;
assign n_15138 = n_13845 & n_15130;
assign n_15139 = ~n_15132 & ~n_15133;
assign n_15140 = n_15134 ^ n_15125;
assign n_15141 = n_15135 ^ x460;
assign n_15142 = ~n_15121 & ~n_15136;
assign n_15143 = n_15136 ^ n_15121;
assign n_15144 = n_15137 & n_14462;
assign n_15145 = n_15137 ^ n_14316;
assign n_15146 = n_15138 ^ n_14405;
assign n_15147 = n_15139 ^ n_13175;
assign n_15148 = n_15140 ^ x459;
assign n_15149 = n_15141 ^ n_15140;
assign n_15150 = n_15144 ^ n_14316;
assign n_15151 = n_15145 ^ n_14448;
assign n_15152 = n_15009 ^ n_15145;
assign n_15153 = n_15146 ^ n_13193;
assign n_15154 = n_15147 ^ n_15146;
assign n_15155 = n_15147 ^ n_13193;
assign n_15156 = n_15149 & ~n_15148;
assign n_15157 = n_15149 ^ x459;
assign n_15158 = n_14490 ^ n_15150;
assign n_15159 = ~n_13856 & ~n_15151;
assign n_15160 = ~n_15153 & n_15154;
assign n_15161 = n_15155 ^ n_15146;
assign n_15162 = n_15156 ^ x459;
assign n_15163 = n_15142 & ~n_15157;
assign n_15164 = n_15157 ^ n_15142;
assign n_15165 = ~n_15158 & n_14504;
assign n_15166 = n_15158 ^ n_14358;
assign n_15167 = n_15159 ^ n_14448;
assign n_15168 = n_15160 ^ n_13193;
assign n_15169 = n_15161 ^ x458;
assign n_15170 = n_15162 ^ n_15161;
assign n_15171 = n_15165 ^ n_14358;
assign n_15172 = n_15166 ^ n_14490;
assign n_15173 = n_15033 ^ n_15166;
assign n_15174 = n_15167 ^ n_13211;
assign n_15175 = n_15168 ^ n_15167;
assign n_15176 = n_15168 ^ n_13211;
assign n_15177 = ~n_15170 & n_15169;
assign n_15178 = n_15170 ^ x458;
assign n_15179 = n_14401 ^ n_15171;
assign n_15180 = n_15171 ^ n_14533;
assign n_15181 = n_13879 & n_15172;
assign n_15182 = n_15174 & n_15175;
assign n_15183 = n_15176 ^ n_15167;
assign n_15184 = n_15177 ^ x458;
assign n_15185 = n_15163 & n_15178;
assign n_15186 = n_15178 ^ n_15163;
assign n_15187 = n_15179 ^ n_14533;
assign n_15188 = n_13906 & ~n_15179;
assign n_15189 = n_14546 & n_15180;
assign n_15190 = n_15181 ^ n_14490;
assign n_15191 = n_15182 ^ n_13211;
assign n_15192 = n_15183 ^ x457;
assign n_15193 = n_15184 ^ n_15183;
assign n_15194 = n_15053 ^ n_15187;
assign n_15195 = n_15188 ^ n_14533;
assign n_15196 = n_15189 ^ n_14401;
assign n_15197 = n_15190 ^ n_13231;
assign n_15198 = n_15190 ^ n_15191;
assign n_15199 = n_15191 ^ n_13231;
assign n_15200 = n_15193 & ~n_15192;
assign n_15201 = n_15193 ^ x457;
assign n_15202 = n_15195 ^ n_13246;
assign n_15203 = n_15196 ^ n_14444;
assign n_15204 = n_15196 ^ n_14568;
assign n_15205 = ~n_15197 & ~n_15198;
assign n_15206 = n_15190 ^ n_15199;
assign n_15207 = n_15200 ^ x457;
assign n_15208 = ~n_15201 & n_15185;
assign n_15209 = n_15185 ^ n_15201;
assign n_15210 = n_13939 & n_15203;
assign n_15211 = n_15203 ^ n_14568;
assign n_15212 = n_14577 & ~n_15204;
assign n_15213 = n_15205 ^ n_13231;
assign n_15214 = n_15206 ^ x456;
assign n_15215 = n_15207 ^ n_15206;
assign n_15216 = n_15210 ^ n_14568;
assign n_15217 = n_15075 ^ n_15211;
assign n_15218 = n_15212 ^ n_14444;
assign n_15219 = n_15213 ^ n_15195;
assign n_15220 = n_15215 & ~n_15214;
assign n_15221 = n_15215 ^ x456;
assign n_15222 = n_15216 ^ n_13276;
assign n_15223 = n_14595 ^ n_15218;
assign n_15224 = n_15219 ^ n_13246;
assign n_15225 = ~n_15219 & n_15202;
assign n_15226 = n_15220 ^ x456;
assign n_15227 = n_15208 & ~n_15221;
assign n_15228 = n_15221 ^ n_15208;
assign n_15229 = n_14486 ^ n_15223;
assign n_15230 = n_15223 & n_14605;
assign n_15231 = n_15224 ^ x471;
assign n_15232 = n_15225 ^ n_13246;
assign n_15233 = n_15224 ^ n_15226;
assign n_15234 = n_15226 ^ x471;
assign n_15235 = n_15229 ^ n_14595;
assign n_15236 = n_15100 ^ n_15229;
assign n_15237 = n_15230 ^ n_14486;
assign n_15238 = n_15232 ^ n_15216;
assign n_15239 = ~n_15231 & n_15233;
assign n_15240 = n_15224 ^ n_15234;
assign n_15241 = ~n_13975 & ~n_15235;
assign n_15242 = n_15237 ^ n_14618;
assign n_15243 = n_15238 ^ n_13276;
assign n_15244 = ~n_15238 & n_15222;
assign n_15245 = n_15239 ^ x471;
assign n_15246 = ~n_15227 & n_15240;
assign n_15247 = n_15240 ^ n_15227;
assign n_15248 = n_15241 ^ n_14595;
assign n_15249 = n_14529 ^ n_15242;
assign n_15250 = ~n_15242 & n_14625;
assign n_15251 = n_15243 ^ x470;
assign n_15252 = n_15244 ^ n_13276;
assign n_15253 = n_15245 ^ n_15243;
assign n_15254 = n_15248 ^ n_13297;
assign n_15255 = n_15249 ^ n_14618;
assign n_15256 = n_15122 ^ n_15249;
assign n_15257 = n_15250 ^ n_14529;
assign n_15258 = n_15252 ^ n_13297;
assign n_15259 = n_15252 ^ n_15248;
assign n_15260 = n_15253 & ~n_15251;
assign n_15261 = n_15253 ^ x470;
assign n_15262 = ~n_14015 & n_15255;
assign n_15263 = n_15257 ^ n_14638;
assign n_15264 = n_15258 ^ n_15248;
assign n_15265 = ~n_15254 & n_15259;
assign n_15266 = n_15260 ^ x470;
assign n_15267 = n_15246 & n_15261;
assign n_15268 = n_15261 ^ n_15246;
assign n_15269 = n_15262 ^ n_14618;
assign n_15270 = n_14565 ^ n_15263;
assign n_15271 = n_15263 & n_14646;
assign n_15272 = n_15264 ^ x469;
assign n_15273 = n_15265 ^ n_13297;
assign n_15274 = n_15266 ^ n_15264;
assign n_15275 = n_15269 ^ n_13317;
assign n_15276 = n_15270 ^ n_14638;
assign n_15277 = n_15143 ^ n_15270;
assign n_15278 = n_15271 ^ n_14565;
assign n_15279 = n_15273 ^ n_13317;
assign n_15280 = n_15273 ^ n_15269;
assign n_15281 = ~n_15274 & n_15272;
assign n_15282 = n_15274 ^ x469;
assign n_15283 = n_14054 & ~n_15276;
assign n_15284 = n_15278 ^ n_14659;
assign n_15285 = n_15279 ^ n_15269;
assign n_15286 = ~n_15275 & n_15280;
assign n_15287 = n_15281 ^ x469;
assign n_15288 = n_15267 & ~n_15282;
assign n_15289 = n_15282 ^ n_15267;
assign n_15290 = n_15283 ^ n_14638;
assign n_15291 = n_14601 ^ n_15284;
assign n_15292 = n_15284 & n_14667;
assign n_15293 = n_15285 ^ x468;
assign n_15294 = n_15286 ^ n_13317;
assign n_15295 = n_15287 ^ n_15285;
assign n_15296 = n_15290 ^ n_13338;
assign n_15297 = n_15291 ^ n_14659;
assign n_15298 = n_15164 ^ n_15291;
assign n_15299 = n_15292 ^ n_14601;
assign n_15300 = n_15294 ^ n_13338;
assign n_15301 = n_15294 ^ n_15290;
assign n_15302 = ~n_15295 & n_15293;
assign n_15303 = n_15295 ^ x468;
assign n_15304 = ~n_14096 & ~n_15297;
assign n_15305 = n_15299 ^ n_14680;
assign n_15306 = n_15300 ^ n_15290;
assign n_15307 = ~n_15296 & ~n_15301;
assign n_15308 = n_15302 ^ x468;
assign n_15309 = ~n_15288 & n_15303;
assign n_15310 = n_15303 ^ n_15288;
assign n_15311 = n_15304 ^ n_14659;
assign n_15312 = n_14628 ^ n_15305;
assign n_15313 = n_15305 & n_14687;
assign n_15314 = n_15306 ^ x467;
assign n_15315 = n_15307 ^ n_13338;
assign n_15316 = n_15308 ^ n_15306;
assign n_15317 = n_15311 ^ n_13359;
assign n_15318 = n_15312 ^ n_14680;
assign n_15319 = n_15186 ^ n_15312;
assign n_15320 = n_15313 ^ n_14628;
assign n_15321 = n_15315 ^ n_13359;
assign n_15322 = n_15315 ^ n_15311;
assign n_15323 = ~n_15316 & n_15314;
assign n_15324 = n_15316 ^ x467;
assign n_15325 = ~n_14139 & ~n_15318;
assign n_15326 = n_15320 ^ n_14695;
assign n_15327 = n_15321 ^ n_15311;
assign n_15328 = n_15317 & ~n_15322;
assign n_15329 = n_15323 ^ x467;
assign n_15330 = ~n_15309 & ~n_15324;
assign n_15331 = n_15324 ^ n_15309;
assign n_15332 = n_15325 ^ n_14680;
assign n_15333 = n_14649 ^ n_15326;
assign n_15334 = n_15326 & ~n_14702;
assign n_15335 = n_15327 ^ x466;
assign n_15336 = n_15328 ^ n_13359;
assign n_15337 = n_15329 ^ n_15327;
assign n_15338 = n_15332 ^ n_13385;
assign n_15339 = n_15333 ^ n_14695;
assign n_15340 = n_15209 ^ n_15333;
assign n_15341 = n_15334 ^ n_14649;
assign n_15342 = n_15336 ^ n_13385;
assign n_15343 = n_15336 ^ n_15332;
assign n_15344 = ~n_15337 & n_15335;
assign n_15345 = n_15337 ^ x466;
assign n_15346 = ~n_14182 & n_15339;
assign n_15347 = n_15341 ^ n_14717;
assign n_15348 = n_15342 ^ n_15332;
assign n_15349 = ~n_15338 & n_15343;
assign n_15350 = n_15344 ^ x466;
assign n_15351 = n_15330 & ~n_15345;
assign n_15352 = n_15345 ^ n_15330;
assign n_15353 = n_15346 ^ n_14695;
assign n_15354 = n_14670 ^ n_15347;
assign n_15355 = ~n_15347 & n_14723;
assign n_15356 = n_15348 ^ x465;
assign n_15357 = n_15349 ^ n_13385;
assign n_15358 = n_15350 ^ n_15348;
assign n_15359 = n_15353 ^ n_13418;
assign n_15360 = n_15354 ^ n_14717;
assign n_15361 = n_15354 ^ n_15228;
assign n_15362 = n_15355 ^ n_14670;
assign n_15363 = n_15357 ^ n_13418;
assign n_15364 = n_15357 ^ n_15353;
assign n_15365 = n_15358 & ~n_15356;
assign n_15366 = n_15358 ^ x465;
assign n_15367 = n_14212 & n_15360;
assign n_15368 = n_15362 ^ n_14690;
assign n_15369 = n_15362 ^ n_14743;
assign n_15370 = n_15363 ^ n_15353;
assign n_15371 = ~n_15359 & ~n_15364;
assign n_15372 = n_15365 ^ x465;
assign n_15373 = ~n_15351 & ~n_15366;
assign n_15374 = n_15366 ^ n_15351;
assign n_15375 = n_15367 ^ n_14717;
assign n_15376 = n_15368 ^ n_14743;
assign n_15377 = n_14750 & n_15369;
assign n_15378 = n_15370 ^ x464;
assign n_15379 = n_15371 ^ n_13418;
assign n_15380 = n_15372 ^ n_15370;
assign n_15381 = n_15375 ^ n_13444;
assign n_15382 = n_15376 ^ n_14737;
assign n_15383 = n_15376 ^ n_15247;
assign n_15384 = n_15377 ^ n_14690;
assign n_15385 = n_15375 ^ n_15379;
assign n_15386 = n_15380 ^ x464;
assign n_15387 = n_15380 & ~n_15378;
assign n_15388 = n_14270 & ~n_15382;
assign n_15389 = n_15384 ^ n_14762;
assign n_15390 = n_15385 ^ n_13444;
assign n_15391 = ~n_15385 & ~n_15381;
assign n_15392 = ~n_15386 & n_15373;
assign n_15393 = n_15373 ^ n_15386;
assign n_15394 = n_15387 ^ x464;
assign n_15395 = n_15388 ^ n_14737;
assign n_15396 = n_14712 ^ n_15389;
assign n_15397 = n_15389 & n_14769;
assign n_15398 = n_15390 ^ x479;
assign n_15399 = n_15391 ^ n_13444;
assign n_15400 = n_14840 & ~n_15393;
assign n_15401 = n_15393 ^ n_14840;
assign n_15402 = n_15394 ^ x479;
assign n_15403 = n_15394 ^ n_15390;
assign n_15404 = n_15395 ^ n_13495;
assign n_15405 = n_15396 ^ n_14762;
assign n_15406 = n_15268 ^ n_15396;
assign n_15407 = n_15397 ^ n_14712;
assign n_15408 = n_15399 ^ n_15395;
assign n_15409 = n_14869 ^ n_15400;
assign n_15410 = n_15401 ^ n_14833;
assign n_15411 = n_15402 ^ n_15390;
assign n_15412 = n_15398 & ~n_15403;
assign n_15413 = n_14313 & ~n_15405;
assign n_15414 = n_15407 ^ n_14782;
assign n_15415 = n_15408 ^ n_13495;
assign n_15416 = ~n_15408 & n_15404;
assign n_15417 = n_13870 & ~n_15410;
assign n_15418 = n_15392 ^ n_15411;
assign n_15419 = ~n_15411 & ~n_15392;
assign n_15420 = n_15412 ^ x479;
assign n_15421 = n_15413 ^ n_14762;
assign n_15422 = n_14732 ^ n_15414;
assign n_15423 = n_15414 & ~n_14789;
assign n_15424 = n_15415 ^ x478;
assign n_15425 = n_15416 ^ n_13495;
assign n_15426 = n_15417 ^ n_14833;
assign n_15427 = n_15418 ^ n_15400;
assign n_15428 = n_15409 ^ n_15418;
assign n_15429 = n_15420 ^ n_15415;
assign n_15430 = n_15421 ^ n_13536;
assign n_15431 = n_15422 ^ n_14782;
assign n_15432 = n_15289 ^ n_15422;
assign n_15433 = n_15423 ^ n_14732;
assign n_15434 = n_15425 ^ n_13536;
assign n_15435 = n_15425 ^ n_15421;
assign n_15436 = n_15426 ^ n_13363;
assign n_15437 = ~n_13363 & n_15426;
assign n_15438 = n_15427 & n_15409;
assign n_15439 = ~n_13900 & ~n_15427;
assign n_15440 = n_15429 ^ x478;
assign n_15441 = ~n_15429 & n_15424;
assign n_15442 = n_14355 & n_15431;
assign n_15443 = n_15433 ^ n_14802;
assign n_15444 = n_15434 ^ n_15421;
assign n_15445 = ~n_15430 & n_15435;
assign n_15446 = x103 & ~n_15436;
assign n_15447 = n_15436 ^ x103;
assign n_15448 = n_15437 ^ n_13391;
assign n_15449 = n_15438 ^ n_14869;
assign n_15450 = n_15439 ^ n_14869;
assign n_15451 = n_15440 ^ n_15419;
assign n_15452 = n_15419 & ~n_15440;
assign n_15453 = n_15441 ^ x478;
assign n_15454 = n_15442 ^ n_14782;
assign n_15455 = n_14753 ^ n_15443;
assign n_15456 = ~n_15443 & ~n_14810;
assign n_15457 = n_15444 ^ x477;
assign n_15458 = n_15445 ^ n_13536;
assign n_15459 = n_15446 ^ x102;
assign n_15460 = n_14909 ^ n_15449;
assign n_15461 = n_15450 ^ n_15448;
assign n_15462 = n_15450 ^ n_15437;
assign n_15463 = n_15449 ^ n_15451;
assign n_15464 = n_14909 ^ n_15451;
assign n_15465 = n_15453 ^ n_15444;
assign n_15466 = n_15454 ^ n_13574;
assign n_15467 = n_15455 ^ n_14802;
assign n_15468 = n_15310 ^ n_15455;
assign n_15469 = n_15456 ^ n_14753;
assign n_15470 = n_15458 ^ n_13574;
assign n_15471 = n_15458 ^ n_15454;
assign n_15472 = n_15460 ^ n_15451;
assign n_15473 = n_15461 ^ n_15446;
assign n_15474 = n_15461 ^ n_15459;
assign n_15475 = n_15448 & ~n_15462;
assign n_15476 = ~n_13941 & n_15463;
assign n_15477 = ~n_15463 & n_15464;
assign n_15478 = n_15465 ^ x477;
assign n_15479 = n_15465 & ~n_15457;
assign n_15480 = n_14398 & ~n_15467;
assign n_15481 = n_15469 ^ n_14823;
assign n_15482 = n_15470 ^ n_15454;
assign n_15483 = n_15466 & ~n_15471;
assign n_15484 = n_15459 & ~n_15473;
assign n_15485 = n_15447 & ~n_15474;
assign n_15486 = n_15474 ^ n_15447;
assign n_15487 = n_15475 ^ n_13391;
assign n_15488 = n_15476 ^ n_14909;
assign n_15489 = n_15477 ^ n_14909;
assign n_15490 = n_15478 ^ n_15452;
assign n_15491 = ~n_15452 & ~n_15478;
assign n_15492 = n_15479 ^ x477;
assign n_15493 = n_15480 ^ n_14802;
assign n_15494 = n_14772 ^ n_15481;
assign n_15495 = ~n_15481 & ~n_14831;
assign n_15496 = n_15482 ^ x476;
assign n_15497 = n_15483 ^ n_13574;
assign n_15498 = n_15484 ^ x102;
assign n_15499 = n_15487 ^ n_13438;
assign n_15500 = n_15488 ^ n_13438;
assign n_15501 = n_15487 ^ n_15488;
assign n_15502 = n_14933 ^ n_15489;
assign n_15503 = n_15489 ^ n_15490;
assign n_15504 = n_14933 ^ n_15490;
assign n_15505 = n_15492 ^ n_15482;
assign n_15506 = n_15493 ^ n_13615;
assign n_15507 = n_15494 ^ n_14823;
assign n_15508 = n_15331 ^ n_15494;
assign n_15509 = n_15495 ^ n_14772;
assign n_15510 = n_15497 ^ n_13615;
assign n_15511 = n_15497 ^ n_15493;
assign n_15512 = n_15499 ^ n_15488;
assign n_15513 = ~n_15500 & ~n_15501;
assign n_15514 = n_15502 ^ n_15490;
assign n_15515 = ~n_13979 & n_15503;
assign n_15516 = ~n_15503 & n_15504;
assign n_15517 = n_15505 ^ x476;
assign n_15518 = ~n_15505 & n_15496;
assign n_15519 = ~n_14441 & ~n_15507;
assign n_15520 = n_15509 ^ n_14846;
assign n_15521 = n_15510 ^ n_15493;
assign n_15522 = ~n_15506 & n_15511;
assign n_15523 = n_15498 ^ n_15512;
assign n_15524 = n_15512 ^ x101;
assign n_15525 = n_15513 ^ n_13438;
assign n_15526 = n_15515 ^ n_14933;
assign n_15527 = n_15516 ^ n_14933;
assign n_15528 = n_15517 ^ n_15491;
assign n_15529 = n_15491 & n_15517;
assign n_15530 = n_15518 ^ x476;
assign n_15531 = n_15519 ^ n_14823;
assign n_15532 = n_14792 ^ n_15520;
assign n_15533 = n_15520 & n_14857;
assign n_15534 = n_15521 ^ x475;
assign n_15535 = n_15522 ^ n_13615;
assign n_15536 = n_15523 ^ x101;
assign n_15537 = n_15523 & ~n_15524;
assign n_15538 = n_15525 ^ n_13476;
assign n_15539 = n_15526 ^ n_13476;
assign n_15540 = n_15525 ^ n_15526;
assign n_15541 = n_14957 ^ n_15527;
assign n_15542 = n_15527 ^ n_15528;
assign n_15543 = n_14957 ^ n_15528;
assign n_15544 = n_15530 ^ n_15521;
assign n_15545 = n_15531 ^ n_13657;
assign n_15546 = n_15532 ^ n_14846;
assign n_15547 = n_15352 ^ n_15532;
assign n_15548 = n_15533 ^ n_14792;
assign n_15549 = n_15535 ^ n_13657;
assign n_15550 = n_15535 ^ n_15531;
assign n_15551 = n_15485 & n_15536;
assign n_15552 = n_15536 ^ n_15485;
assign n_15553 = n_15537 ^ x101;
assign n_15554 = n_15538 ^ n_15526;
assign n_15555 = ~n_15539 & n_15540;
assign n_15556 = n_15541 ^ n_15528;
assign n_15557 = n_14022 & n_15542;
assign n_15558 = ~n_15542 & ~n_15543;
assign n_15559 = n_15544 ^ x475;
assign n_15560 = n_15544 & ~n_15534;
assign n_15561 = n_14483 & ~n_15546;
assign n_15562 = n_15548 ^ n_14866;
assign n_15563 = n_15549 ^ n_15531;
assign n_15564 = n_15545 & ~n_15550;
assign n_15565 = n_15553 ^ n_15554;
assign n_15566 = n_15554 ^ x100;
assign n_15567 = n_15555 ^ n_13476;
assign n_15568 = n_15557 ^ n_14957;
assign n_15569 = n_15558 ^ n_14957;
assign n_15570 = n_15559 ^ n_15529;
assign n_15571 = n_15529 & ~n_15559;
assign n_15572 = n_15560 ^ x475;
assign n_15573 = n_15561 ^ n_14846;
assign n_15574 = n_15562 ^ n_14813;
assign n_15575 = n_15563 ^ x474;
assign n_15576 = n_15564 ^ n_13657;
assign n_15577 = n_15565 ^ x100;
assign n_15578 = ~n_15565 & n_15566;
assign n_15579 = n_15567 ^ n_15568;
assign n_15580 = n_15568 ^ n_13516;
assign n_15581 = n_15569 ^ n_14974;
assign n_15582 = n_15569 ^ n_15570;
assign n_15583 = n_15570 ^ n_14974;
assign n_15584 = n_15572 ^ n_15563;
assign n_15585 = n_15573 ^ n_13699;
assign n_15586 = n_15574 ^ n_14866;
assign n_15587 = n_15576 ^ n_13699;
assign n_15588 = n_15576 ^ n_15573;
assign n_15589 = ~n_15551 & n_15577;
assign n_15590 = n_15577 ^ n_15551;
assign n_15591 = n_15578 ^ x100;
assign n_15592 = n_15579 ^ n_13516;
assign n_15593 = ~n_15579 & ~n_15580;
assign n_15594 = n_15581 ^ n_15570;
assign n_15595 = n_14061 & n_15582;
assign n_15596 = ~n_15582 & n_15583;
assign n_15597 = n_15584 ^ x474;
assign n_15598 = ~n_15584 & n_15575;
assign n_15599 = ~n_14513 & ~n_15586;
assign n_15600 = n_15587 ^ n_15573;
assign n_15601 = n_15585 & ~n_15588;
assign n_15602 = n_15591 ^ n_15592;
assign n_15603 = n_15592 ^ x99;
assign n_15604 = n_15593 ^ n_13516;
assign n_15605 = n_15595 ^ n_14974;
assign n_15606 = n_15596 ^ n_14974;
assign n_15607 = n_15597 ^ n_15571;
assign n_15608 = n_15571 & n_15597;
assign n_15609 = n_15598 ^ x474;
assign n_15610 = n_15599 ^ n_14866;
assign n_15611 = n_15600 ^ x473;
assign n_15612 = n_15601 ^ n_13699;
assign n_15613 = n_15602 ^ x99;
assign n_15614 = ~n_15602 & n_15603;
assign n_15615 = n_15604 ^ n_15605;
assign n_15616 = n_15605 ^ n_13557;
assign n_15617 = n_14993 ^ n_15606;
assign n_15618 = n_15606 ^ n_15607;
assign n_15619 = n_14993 ^ n_15607;
assign n_15620 = n_15609 ^ n_15600;
assign n_15621 = n_15610 ^ n_13729;
assign n_15622 = n_15612 ^ x472;
assign n_15623 = n_15589 & n_15613;
assign n_15624 = n_15613 ^ n_15589;
assign n_15625 = n_15614 ^ x99;
assign n_15626 = n_15615 ^ n_13557;
assign n_15627 = n_15615 & ~n_15616;
assign n_15628 = n_15617 ^ n_15607;
assign n_15629 = n_14103 & ~n_15618;
assign n_15630 = n_15618 & n_15619;
assign n_15631 = n_15620 ^ x473;
assign n_15632 = ~n_15620 & n_15611;
assign n_15633 = n_15622 ^ n_15621;
assign n_15634 = n_15625 ^ n_15626;
assign n_15635 = n_15626 ^ x98;
assign n_15636 = n_15627 ^ n_13557;
assign n_15637 = n_15629 ^ n_14993;
assign n_15638 = n_15630 ^ n_14993;
assign n_15639 = n_15631 ^ n_15608;
assign n_15640 = ~n_15608 & ~n_15631;
assign n_15641 = n_15632 ^ x473;
assign n_15642 = n_15634 ^ x98;
assign n_15643 = n_15634 & ~n_15635;
assign n_15644 = n_15636 ^ n_13597;
assign n_15645 = n_15637 ^ n_13597;
assign n_15646 = n_15636 ^ n_15637;
assign n_15647 = n_15638 ^ n_15006;
assign n_15648 = n_15638 ^ n_15639;
assign n_15649 = n_15639 ^ n_15006;
assign n_15650 = n_15641 ^ n_15640;
assign n_15651 = ~n_15642 & n_15623;
assign n_15652 = n_15623 ^ n_15642;
assign n_15653 = n_15643 ^ x98;
assign n_15654 = n_15644 ^ n_15637;
assign n_15655 = ~n_15645 & ~n_15646;
assign n_15656 = n_15647 ^ n_15639;
assign n_15657 = n_14146 & ~n_15648;
assign n_15658 = n_15648 & n_15649;
assign n_15659 = n_15650 ^ n_15633;
assign n_15660 = n_15653 ^ n_15654;
assign n_15661 = n_15654 ^ x97;
assign n_15662 = n_15655 ^ n_13597;
assign n_15663 = n_15657 ^ n_15006;
assign n_15664 = n_15658 ^ n_15006;
assign n_15665 = n_15659 ^ n_15024;
assign n_15666 = n_15660 ^ x97;
assign n_15667 = n_15660 & ~n_15661;
assign n_15668 = n_15662 ^ n_13639;
assign n_15669 = n_15663 ^ n_13639;
assign n_15670 = n_15662 ^ n_15663;
assign n_15671 = n_15664 ^ n_15659;
assign n_15672 = n_15664 ^ n_15024;
assign n_15673 = n_15651 & ~n_15666;
assign n_15674 = n_15666 ^ n_15651;
assign n_15675 = n_15667 ^ x97;
assign n_15676 = n_15668 ^ n_15663;
assign n_15677 = n_15669 & ~n_15670;
assign n_15678 = ~n_15671 & ~n_15665;
assign n_15679 = n_14189 & n_15671;
assign n_15680 = n_15672 ^ n_15659;
assign n_15681 = n_15675 ^ n_15676;
assign n_15682 = n_15676 ^ x96;
assign n_15683 = n_15677 ^ n_13639;
assign n_15684 = n_15678 ^ n_15024;
assign n_15685 = n_15679 ^ n_15024;
assign n_15686 = n_15681 ^ x96;
assign n_15687 = n_15681 & ~n_15682;
assign n_15688 = n_15683 ^ n_13681;
assign n_15689 = n_15684 ^ n_15043;
assign n_15690 = n_15685 ^ n_13681;
assign n_15691 = n_15683 ^ n_15685;
assign n_15692 = ~n_15673 & n_15686;
assign n_15693 = n_15686 ^ n_15673;
assign n_15694 = n_15687 ^ x96;
assign n_15695 = n_15688 ^ n_15685;
assign n_15696 = ~n_15689 & n_15050;
assign n_15697 = n_14886 ^ n_15689;
assign n_15698 = n_15690 & n_15691;
assign n_15699 = n_15694 ^ n_15695;
assign n_15700 = n_15695 ^ x111;
assign n_15701 = n_15696 ^ n_14886;
assign n_15702 = n_15697 ^ n_15043;
assign n_15703 = n_15698 ^ n_13681;
assign n_15704 = n_15699 ^ x111;
assign n_15705 = n_15699 & ~n_15700;
assign n_15706 = n_15701 ^ n_15063;
assign n_15707 = ~n_14234 & n_15702;
assign n_15708 = n_15703 ^ n_13723;
assign n_15709 = n_15692 & n_15704;
assign n_15710 = n_15704 ^ n_15692;
assign n_15711 = n_15705 ^ x111;
assign n_15712 = ~n_15706 & n_15070;
assign n_15713 = n_15706 ^ n_14907;
assign n_15714 = n_15707 ^ n_15043;
assign n_15715 = n_15712 ^ n_14907;
assign n_15716 = n_15713 ^ n_15063;
assign n_15717 = n_15708 ^ n_15714;
assign n_15718 = n_15714 ^ n_13723;
assign n_15719 = n_15703 ^ n_15714;
assign n_15720 = n_15715 ^ n_15082;
assign n_15721 = ~n_14277 & n_15716;
assign n_15722 = n_15711 ^ n_15717;
assign n_15723 = n_15717 ^ x110;
assign n_15724 = ~n_15718 & ~n_15719;
assign n_15725 = ~n_15720 & ~n_15089;
assign n_15726 = n_14951 ^ n_15720;
assign n_15727 = n_15721 ^ n_15063;
assign n_15728 = n_15722 ^ x110;
assign n_15729 = n_15722 & ~n_15723;
assign n_15730 = n_15724 ^ n_13723;
assign n_15731 = n_15725 ^ n_14951;
assign n_15732 = n_15726 ^ n_15082;
assign n_15733 = n_15709 ^ n_15728;
assign n_15734 = ~n_15728 & ~n_15709;
assign n_15735 = n_15729 ^ x110;
assign n_15736 = n_15730 ^ n_13763;
assign n_15737 = n_15727 ^ n_15730;
assign n_15738 = n_15731 ^ n_15103;
assign n_15739 = ~n_14320 & ~n_15732;
assign n_15740 = n_15727 ^ n_15736;
assign n_15741 = n_15736 & n_15737;
assign n_15742 = ~n_15738 & n_15110;
assign n_15743 = n_14970 ^ n_15738;
assign n_15744 = n_15739 ^ n_15082;
assign n_15745 = n_15735 ^ n_15740;
assign n_15746 = n_15740 ^ x109;
assign n_15747 = n_15741 ^ n_13763;
assign n_15748 = n_15742 ^ n_14970;
assign n_15749 = n_15743 ^ n_15103;
assign n_15750 = n_15744 ^ n_13797;
assign n_15751 = n_15745 ^ x109;
assign n_15752 = ~n_15745 & n_15746;
assign n_15753 = n_15747 ^ n_15744;
assign n_15754 = n_15747 ^ n_13797;
assign n_15755 = n_15748 ^ n_15124;
assign n_15756 = n_14362 & n_15749;
assign n_15757 = ~n_15751 & ~n_15734;
assign n_15758 = n_15734 ^ n_15751;
assign n_15759 = n_15752 ^ x109;
assign n_15760 = n_15750 & n_15753;
assign n_15761 = n_15754 ^ n_15744;
assign n_15762 = n_15755 & n_15131;
assign n_15763 = n_14988 ^ n_15755;
assign n_15764 = n_15756 ^ n_15103;
assign n_15765 = n_15759 ^ x108;
assign n_15766 = n_15760 ^ n_13797;
assign n_15767 = n_15759 ^ n_15761;
assign n_15768 = n_15762 ^ n_14988;
assign n_15769 = n_15763 ^ n_15124;
assign n_15770 = n_15764 ^ n_13825;
assign n_15771 = n_15766 ^ n_15764;
assign n_15772 = n_15766 ^ n_13825;
assign n_15773 = n_15767 & n_15765;
assign n_15774 = n_15767 ^ x108;
assign n_15775 = n_15768 ^ n_15145;
assign n_15776 = n_14405 & ~n_15769;
assign n_15777 = ~n_15770 & n_15771;
assign n_15778 = n_15772 ^ n_15764;
assign n_15779 = n_15773 ^ x108;
assign n_15780 = n_15757 & n_15774;
assign n_15781 = n_15774 ^ n_15757;
assign n_15782 = n_15775 & n_15152;
assign n_15783 = n_15009 ^ n_15775;
assign n_15784 = n_15776 ^ n_15124;
assign n_15785 = n_15777 ^ n_13825;
assign n_15786 = n_15778 ^ x107;
assign n_15787 = n_15779 ^ n_15778;
assign n_15788 = n_15782 ^ n_15009;
assign n_15789 = n_15447 ^ n_15783;
assign n_15790 = n_15783 ^ n_15145;
assign n_15791 = n_15784 ^ n_13845;
assign n_15792 = n_15785 ^ n_15784;
assign n_15793 = n_15785 ^ n_13845;
assign n_15794 = n_15787 & ~n_15786;
assign n_15795 = n_15787 ^ x107;
assign n_15796 = n_15788 ^ n_15166;
assign n_15797 = n_14448 & ~n_15790;
assign n_15798 = n_15791 & ~n_15792;
assign n_15799 = n_15793 ^ n_15784;
assign n_15800 = n_15794 ^ x107;
assign n_15801 = ~n_15780 & ~n_15795;
assign n_15802 = n_15795 ^ n_15780;
assign n_15803 = n_15796 & ~n_15173;
assign n_15804 = n_15033 ^ n_15796;
assign n_15805 = n_15797 ^ n_15145;
assign n_15806 = n_15798 ^ n_13845;
assign n_15807 = n_15799 ^ x106;
assign n_15808 = n_15800 ^ n_15799;
assign n_15809 = n_15803 ^ n_15033;
assign n_15810 = n_15804 ^ n_15166;
assign n_15811 = n_15486 ^ n_15804;
assign n_15812 = n_15805 ^ n_13856;
assign n_15813 = n_15806 ^ n_15805;
assign n_15814 = n_15806 ^ n_13856;
assign n_15815 = ~n_15808 & n_15807;
assign n_15816 = n_15808 ^ x106;
assign n_15817 = n_15187 ^ n_15809;
assign n_15818 = n_14490 & n_15810;
assign n_15819 = n_15812 & n_15813;
assign n_15820 = n_15814 ^ n_15805;
assign n_15821 = n_15815 ^ x106;
assign n_15822 = n_15801 & n_15816;
assign n_15823 = n_15816 ^ n_15801;
assign n_15824 = n_15053 ^ n_15817;
assign n_15825 = n_15817 & n_15194;
assign n_15826 = n_15818 ^ n_15166;
assign n_15827 = n_15819 ^ n_13856;
assign n_15828 = n_15820 ^ x105;
assign n_15829 = n_15821 ^ n_15820;
assign n_15830 = n_15824 ^ n_15179;
assign n_15831 = n_15552 ^ n_15824;
assign n_15832 = n_15825 ^ n_15053;
assign n_15833 = n_15826 ^ n_13879;
assign n_15834 = n_15827 ^ n_15826;
assign n_15835 = n_15827 ^ n_13879;
assign n_15836 = ~n_15829 & n_15828;
assign n_15837 = n_15829 ^ x105;
assign n_15838 = ~n_14533 & n_15830;
assign n_15839 = n_15211 ^ n_15832;
assign n_15840 = n_15833 & n_15834;
assign n_15841 = n_15835 ^ n_15826;
assign n_15842 = n_15836 ^ x105;
assign n_15843 = n_15822 & n_15837;
assign n_15844 = n_15837 ^ n_15822;
assign n_15845 = n_15838 ^ n_15179;
assign n_15846 = n_15839 & n_15217;
assign n_15847 = n_15075 ^ n_15839;
assign n_15848 = n_15840 ^ n_13879;
assign n_15849 = n_15841 ^ x104;
assign n_15850 = n_15842 ^ n_15841;
assign n_15851 = n_15845 ^ n_13906;
assign n_15852 = n_15846 ^ n_15075;
assign n_15853 = n_15590 ^ n_15847;
assign n_15854 = n_15847 ^ n_15203;
assign n_15855 = n_15848 ^ n_15845;
assign n_15856 = n_15842 ^ n_15849;
assign n_15857 = ~n_15849 & n_15850;
assign n_15858 = n_15852 ^ n_15229;
assign n_15859 = ~n_14568 & n_15854;
assign n_15860 = n_15855 & ~n_15851;
assign n_15861 = n_15855 ^ n_13906;
assign n_15862 = n_15843 & ~n_15856;
assign n_15863 = n_15856 ^ n_15843;
assign n_15864 = n_15857 ^ x104;
assign n_15865 = ~n_15858 & n_15236;
assign n_15866 = n_15100 ^ n_15858;
assign n_15867 = n_15859 ^ n_15203;
assign n_15868 = n_15860 ^ n_13906;
assign n_15869 = n_15861 ^ x119;
assign n_15870 = n_15864 ^ n_15861;
assign n_15871 = n_15864 ^ x119;
assign n_15872 = n_15865 ^ n_15100;
assign n_15873 = n_15866 ^ n_15229;
assign n_15874 = n_15624 ^ n_15866;
assign n_15875 = n_15867 ^ n_13939;
assign n_15876 = n_15868 ^ n_15867;
assign n_15877 = n_15868 ^ n_13939;
assign n_15878 = ~n_15869 & n_15870;
assign n_15879 = n_15871 ^ n_15861;
assign n_15880 = n_15872 ^ n_15249;
assign n_15881 = n_14595 & n_15873;
assign n_15882 = n_15875 & ~n_15876;
assign n_15883 = n_15877 ^ n_15867;
assign n_15884 = n_15878 ^ x119;
assign n_15885 = ~n_15862 & n_15879;
assign n_15886 = n_15879 ^ n_15862;
assign n_15887 = n_15122 ^ n_15880;
assign n_15888 = n_15880 & n_15256;
assign n_15889 = n_15881 ^ n_15229;
assign n_15890 = n_15882 ^ n_13939;
assign n_15891 = n_15883 ^ x118;
assign n_15892 = n_15884 ^ n_15883;
assign n_15893 = n_15652 ^ n_15887;
assign n_15894 = n_15887 ^ n_15249;
assign n_15895 = n_15888 ^ n_15122;
assign n_15896 = n_15889 ^ n_13975;
assign n_15897 = n_15890 ^ n_15889;
assign n_15898 = ~n_15892 & n_15891;
assign n_15899 = n_15892 ^ x118;
assign n_15900 = n_14618 & ~n_15894;
assign n_15901 = n_15895 ^ n_15270;
assign n_15902 = n_15897 & n_15896;
assign n_15903 = n_15897 ^ n_13975;
assign n_15904 = n_15898 ^ x118;
assign n_15905 = ~n_15885 & n_15899;
assign n_15906 = n_15900 ^ n_15249;
assign n_15907 = ~n_15901 & n_15277;
assign n_15908 = n_15143 ^ n_15901;
assign n_15909 = n_15902 ^ n_13975;
assign n_15910 = n_15903 ^ x117;
assign n_15911 = n_15904 ^ n_15903;
assign n_15912 = n_15904 ^ x117;
assign n_15913 = n_15906 ^ n_14015;
assign n_15914 = n_15907 ^ n_15143;
assign n_15915 = n_15908 ^ n_15270;
assign n_15916 = n_15674 ^ n_15908;
assign n_15917 = n_15909 ^ n_15906;
assign n_15918 = n_15909 ^ n_14015;
assign n_15919 = n_15910 & ~n_15911;
assign n_15920 = n_15912 ^ n_15903;
assign n_15921 = n_15914 ^ n_15291;
assign n_15922 = ~n_14638 & n_15915;
assign n_15923 = ~n_15913 & n_15917;
assign n_15924 = n_15918 ^ n_15906;
assign n_15925 = n_15919 ^ x117;
assign n_15926 = ~n_15920 & ~n_15905;
assign n_15927 = n_15905 ^ n_15920;
assign n_15928 = n_15921 & n_15298;
assign n_15929 = n_15164 ^ n_15921;
assign n_15930 = n_15922 ^ n_15270;
assign n_15931 = n_15923 ^ n_14015;
assign n_15932 = n_15924 ^ x116;
assign n_15933 = n_15925 ^ n_15924;
assign n_15934 = ~n_15401 & ~n_15927;
assign n_15935 = n_15927 ^ n_15401;
assign n_15936 = n_15928 ^ n_15164;
assign n_15937 = n_15929 ^ n_15291;
assign n_15938 = n_15693 ^ n_15929;
assign n_15939 = n_15930 ^ n_14054;
assign n_15940 = n_15931 ^ n_15930;
assign n_15941 = n_15931 ^ n_14054;
assign n_15942 = ~n_15933 & n_15932;
assign n_15943 = n_15933 ^ x116;
assign n_15944 = n_15428 ^ n_15934;
assign n_15945 = n_15935 ^ n_15393;
assign n_15946 = n_15936 ^ n_15312;
assign n_15947 = n_14659 & ~n_15937;
assign n_15948 = n_15939 & n_15940;
assign n_15949 = n_15941 ^ n_15930;
assign n_15950 = n_15942 ^ x116;
assign n_15951 = n_15943 & ~n_15926;
assign n_15952 = n_15926 ^ n_15943;
assign n_15953 = n_14840 & ~n_15945;
assign n_15954 = n_15946 & n_15319;
assign n_15955 = n_15186 ^ n_15946;
assign n_15956 = n_15947 ^ n_15291;
assign n_15957 = n_15948 ^ n_14054;
assign n_15958 = n_15949 ^ x115;
assign n_15959 = n_15950 ^ n_15949;
assign n_15960 = n_15934 ^ n_15952;
assign n_15961 = n_15428 ^ n_15952;
assign n_15962 = n_15944 ^ n_15952;
assign n_15963 = n_15953 ^ n_15393;
assign n_15964 = n_15954 ^ n_15186;
assign n_15965 = n_15955 ^ n_15312;
assign n_15966 = n_15710 ^ n_15955;
assign n_15967 = n_15956 ^ n_14096;
assign n_15968 = n_15957 ^ n_15956;
assign n_15969 = n_15957 ^ n_14096;
assign n_15970 = n_15959 & ~n_15958;
assign n_15971 = n_15959 ^ x115;
assign n_15972 = n_14869 & ~n_15960;
assign n_15973 = n_15960 & n_15961;
assign n_15974 = n_13870 & ~n_15963;
assign n_15975 = n_15963 ^ n_13870;
assign n_15976 = n_15964 ^ n_15333;
assign n_15977 = ~n_14680 & ~n_15965;
assign n_15978 = n_15967 & n_15968;
assign n_15979 = n_15969 ^ n_15956;
assign n_15980 = n_15970 ^ x115;
assign n_15981 = n_15971 & ~n_15951;
assign n_15982 = n_15951 ^ n_15971;
assign n_15983 = n_15972 ^ n_15428;
assign n_15984 = n_15973 ^ n_15428;
assign n_15985 = n_15974 ^ n_13900;
assign n_15986 = x263 & ~n_15975;
assign n_15987 = n_15975 ^ x263;
assign n_15988 = n_15209 ^ n_15976;
assign n_15989 = ~n_15976 & ~n_15340;
assign n_15990 = n_15977 ^ n_15312;
assign n_15991 = n_15978 ^ n_14096;
assign n_15992 = n_15979 ^ x114;
assign n_15993 = n_15980 ^ n_15979;
assign n_15994 = n_15472 ^ n_15982;
assign n_15995 = n_15983 ^ n_15974;
assign n_15996 = n_15984 ^ n_15982;
assign n_15997 = n_15472 ^ n_15984;
assign n_15998 = n_15983 ^ n_15985;
assign n_15999 = n_15986 ^ x262;
assign n_16000 = n_15988 ^ n_15333;
assign n_16001 = n_15733 ^ n_15988;
assign n_16002 = n_15989 ^ n_15209;
assign n_16003 = n_15990 ^ n_14139;
assign n_16004 = n_15991 ^ n_15990;
assign n_16005 = n_15991 ^ n_14139;
assign n_16006 = ~n_15993 & n_15992;
assign n_16007 = n_15993 ^ x114;
assign n_16008 = ~n_15985 & n_15995;
assign n_16009 = n_15996 & n_15994;
assign n_16010 = n_14909 & ~n_15996;
assign n_16011 = n_15997 ^ n_15982;
assign n_16012 = n_15998 ^ n_15986;
assign n_16013 = n_15998 ^ n_15999;
assign n_16014 = n_14695 & ~n_16000;
assign n_16015 = n_16002 ^ n_15228;
assign n_16016 = n_16002 ^ n_15354;
assign n_16017 = ~n_16003 & n_16004;
assign n_16018 = n_16005 ^ n_15990;
assign n_16019 = n_16006 ^ x114;
assign n_16020 = ~n_15981 & n_16007;
assign n_16021 = n_16007 ^ n_15981;
assign n_16022 = n_16008 ^ n_13900;
assign n_16023 = n_16009 ^ n_15472;
assign n_16024 = n_16010 ^ n_15472;
assign n_16025 = n_15999 & ~n_16012;
assign n_16026 = ~n_15987 & n_16013;
assign n_16027 = n_16013 ^ n_15987;
assign n_16028 = n_16014 ^ n_15333;
assign n_16029 = ~n_14717 & n_16015;
assign n_16030 = n_16015 ^ n_15354;
assign n_16031 = n_15361 & ~n_16016;
assign n_16032 = n_16017 ^ n_14139;
assign n_16033 = n_16018 ^ x113;
assign n_16034 = n_16019 ^ n_16018;
assign n_16035 = n_15514 ^ n_16021;
assign n_16036 = n_16022 ^ n_13941;
assign n_16037 = n_16023 ^ n_16021;
assign n_16038 = n_15514 ^ n_16023;
assign n_16039 = n_16024 ^ n_13941;
assign n_16040 = n_16022 ^ n_16024;
assign n_16041 = n_16025 ^ x262;
assign n_16042 = n_16028 ^ n_14182;
assign n_16043 = n_16029 ^ n_15354;
assign n_16044 = n_15758 ^ n_16030;
assign n_16045 = n_16031 ^ n_15228;
assign n_16046 = n_16032 ^ n_16028;
assign n_16047 = n_16032 ^ n_14182;
assign n_16048 = ~n_16034 & n_16033;
assign n_16049 = n_16034 ^ x113;
assign n_16050 = n_16036 ^ n_16024;
assign n_16051 = n_16037 & ~n_16035;
assign n_16052 = n_14933 & ~n_16037;
assign n_16053 = n_16038 ^ n_16021;
assign n_16054 = ~n_16039 & n_16040;
assign n_16055 = n_16043 ^ n_14212;
assign n_16056 = n_16045 ^ n_15247;
assign n_16057 = n_16045 ^ n_15376;
assign n_16058 = ~n_16042 & n_16046;
assign n_16059 = n_16047 ^ n_16028;
assign n_16060 = n_16048 ^ x113;
assign n_16061 = ~n_16049 & ~n_16020;
assign n_16062 = n_16020 ^ n_16049;
assign n_16063 = n_16041 ^ n_16050;
assign n_16064 = n_16050 ^ x261;
assign n_16065 = n_16051 ^ n_15514;
assign n_16066 = n_16052 ^ n_15514;
assign n_16067 = n_16054 ^ n_13941;
assign n_16068 = n_16056 ^ n_15376;
assign n_16069 = ~n_15383 & ~n_16057;
assign n_16070 = n_16058 ^ n_14182;
assign n_16071 = n_16059 ^ x112;
assign n_16072 = n_16060 ^ n_16059;
assign n_16073 = n_15556 ^ n_16062;
assign n_16074 = n_16063 ^ x261;
assign n_16075 = ~n_16063 & n_16064;
assign n_16076 = n_16065 ^ n_16062;
assign n_16077 = n_15556 ^ n_16065;
assign n_16078 = n_16066 ^ n_13979;
assign n_16079 = n_16067 ^ n_16066;
assign n_16080 = n_16067 ^ n_13979;
assign n_16081 = n_16068 ^ n_15368;
assign n_16082 = n_15781 ^ n_16068;
assign n_16083 = n_16069 ^ n_15247;
assign n_16084 = n_16070 ^ n_16043;
assign n_16085 = ~n_16072 & n_16071;
assign n_16086 = n_16072 ^ x112;
assign n_16087 = ~n_16074 & ~n_16026;
assign n_16088 = n_16026 ^ n_16074;
assign n_16089 = n_16075 ^ x261;
assign n_16090 = n_16076 & n_16073;
assign n_16091 = ~n_14957 & ~n_16076;
assign n_16092 = n_16077 ^ n_16062;
assign n_16093 = ~n_16078 & n_16079;
assign n_16094 = n_16080 ^ n_16066;
assign n_16095 = n_14743 & ~n_16081;
assign n_16096 = n_16083 ^ n_15396;
assign n_16097 = n_16084 ^ n_14212;
assign n_16098 = ~n_16084 & ~n_16055;
assign n_16099 = n_16085 ^ x112;
assign n_16100 = n_16061 & ~n_16086;
assign n_16101 = n_16086 ^ n_16061;
assign n_16102 = n_16090 ^ n_15556;
assign n_16103 = n_16091 ^ n_15556;
assign n_16104 = n_16093 ^ n_13979;
assign n_16105 = n_16089 ^ n_16094;
assign n_16106 = n_16094 ^ x260;
assign n_16107 = n_16095 ^ n_15368;
assign n_16108 = n_15268 ^ n_16096;
assign n_16109 = ~n_16096 & ~n_15406;
assign n_16110 = n_16097 ^ x127;
assign n_16111 = n_16098 ^ n_14212;
assign n_16112 = n_16099 ^ n_16097;
assign n_16113 = n_16099 ^ x127;
assign n_16114 = n_15594 ^ n_16101;
assign n_16115 = n_16102 ^ n_16101;
assign n_16116 = n_15594 ^ n_16102;
assign n_16117 = n_16103 ^ n_14022;
assign n_16118 = n_16104 ^ n_16103;
assign n_16119 = n_16104 ^ n_14022;
assign n_16120 = n_16105 ^ x260;
assign n_16121 = ~n_16105 & n_16106;
assign n_16122 = n_16107 ^ n_14270;
assign n_16123 = n_16108 ^ n_15396;
assign n_16124 = n_15802 ^ n_16108;
assign n_16125 = n_16109 ^ n_15268;
assign n_16126 = n_16111 ^ n_16107;
assign n_16127 = n_16110 & ~n_16112;
assign n_16128 = n_16113 ^ n_16097;
assign n_16129 = n_16115 & ~n_16114;
assign n_16130 = ~n_14974 & ~n_16115;
assign n_16131 = n_16116 ^ n_16101;
assign n_16132 = ~n_16117 & ~n_16118;
assign n_16133 = n_16119 ^ n_16103;
assign n_16134 = n_16087 & ~n_16120;
assign n_16135 = n_16120 ^ n_16087;
assign n_16136 = n_16121 ^ x260;
assign n_16137 = ~n_14762 & ~n_16123;
assign n_16138 = n_16125 ^ n_15422;
assign n_16139 = n_16126 ^ n_14270;
assign n_16140 = n_16126 & ~n_16122;
assign n_16141 = n_16127 ^ x127;
assign n_16142 = ~n_16100 & n_16128;
assign n_16143 = n_16128 ^ n_16100;
assign n_16144 = n_16129 ^ n_15594;
assign n_16145 = n_16130 ^ n_15594;
assign n_16146 = n_16132 ^ n_14022;
assign n_16147 = n_16133 ^ x259;
assign n_16148 = n_16136 ^ n_16133;
assign n_16149 = n_16137 ^ n_15396;
assign n_16150 = n_15289 ^ n_16138;
assign n_16151 = n_16138 & n_15432;
assign n_16152 = n_16139 ^ x126;
assign n_16153 = n_16140 ^ n_14270;
assign n_16154 = n_16141 ^ n_16139;
assign n_16155 = n_15628 ^ n_16143;
assign n_16156 = n_16144 ^ n_16143;
assign n_16157 = n_15628 ^ n_16144;
assign n_16158 = n_16145 ^ n_14061;
assign n_16159 = n_16146 ^ n_16145;
assign n_16160 = n_16146 ^ n_14061;
assign n_16161 = ~n_16148 & n_16147;
assign n_16162 = n_16148 ^ x259;
assign n_16163 = n_16149 ^ n_14313;
assign n_16164 = n_16150 ^ n_15422;
assign n_16165 = n_15823 ^ n_16150;
assign n_16166 = n_16151 ^ n_15289;
assign n_16167 = n_16153 ^ n_14313;
assign n_16168 = n_16153 ^ n_16149;
assign n_16169 = n_16154 & ~n_16152;
assign n_16170 = n_16154 ^ x126;
assign n_16171 = ~n_16156 & n_16155;
assign n_16172 = n_14993 & n_16156;
assign n_16173 = n_16157 ^ n_16143;
assign n_16174 = ~n_16158 & n_16159;
assign n_16175 = n_16160 ^ n_16145;
assign n_16176 = n_16161 ^ x259;
assign n_16177 = n_16162 & ~n_16134;
assign n_16178 = n_16134 ^ n_16162;
assign n_16179 = n_14782 & ~n_16164;
assign n_16180 = n_16166 ^ n_15455;
assign n_16181 = n_16167 ^ n_16149;
assign n_16182 = n_16163 & ~n_16168;
assign n_16183 = n_16169 ^ x126;
assign n_16184 = n_16142 & ~n_16170;
assign n_16185 = n_16170 ^ n_16142;
assign n_16186 = n_16171 ^ n_15628;
assign n_16187 = n_16172 ^ n_15628;
assign n_16188 = n_16174 ^ n_14061;
assign n_16189 = n_16175 ^ x258;
assign n_16190 = n_16176 ^ n_16175;
assign n_16191 = n_16179 ^ n_15422;
assign n_16192 = n_15310 ^ n_16180;
assign n_16193 = ~n_16180 & ~n_15468;
assign n_16194 = n_16181 ^ x125;
assign n_16195 = n_16182 ^ n_14313;
assign n_16196 = n_16183 ^ n_16181;
assign n_16197 = n_15656 ^ n_16185;
assign n_16198 = n_16186 ^ n_16185;
assign n_16199 = n_15656 ^ n_16186;
assign n_16200 = n_16187 ^ n_14103;
assign n_16201 = n_16188 ^ n_16187;
assign n_16202 = n_16188 ^ n_14103;
assign n_16203 = n_16190 & ~n_16189;
assign n_16204 = n_16190 ^ x258;
assign n_16205 = n_16191 ^ n_14355;
assign n_16206 = n_16192 ^ n_15455;
assign n_16207 = n_15844 ^ n_16192;
assign n_16208 = n_16193 ^ n_15310;
assign n_16209 = n_16195 ^ n_14355;
assign n_16210 = n_16195 ^ n_16191;
assign n_16211 = ~n_16196 & n_16194;
assign n_16212 = n_16196 ^ x125;
assign n_16213 = ~n_16198 & ~n_16197;
assign n_16214 = ~n_15006 & n_16198;
assign n_16215 = n_16199 ^ n_16185;
assign n_16216 = ~n_16200 & n_16201;
assign n_16217 = n_16202 ^ n_16187;
assign n_16218 = n_16203 ^ x258;
assign n_16219 = ~n_16177 & n_16204;
assign n_16220 = n_16204 ^ n_16177;
assign n_16221 = ~n_14802 & ~n_16206;
assign n_16222 = n_16208 ^ n_15494;
assign n_16223 = n_16209 ^ n_16191;
assign n_16224 = n_16205 & ~n_16210;
assign n_16225 = n_16211 ^ x125;
assign n_16226 = ~n_16212 & ~n_16184;
assign n_16227 = n_16184 ^ n_16212;
assign n_16228 = n_16213 ^ n_15656;
assign n_16229 = n_16214 ^ n_15656;
assign n_16230 = n_16216 ^ n_14103;
assign n_16231 = n_16217 ^ x257;
assign n_16232 = n_16218 ^ n_16217;
assign n_16233 = n_16221 ^ n_15455;
assign n_16234 = n_15331 ^ n_16222;
assign n_16235 = ~n_16222 & n_15508;
assign n_16236 = n_16223 ^ x124;
assign n_16237 = n_16224 ^ n_14355;
assign n_16238 = n_16225 ^ n_16223;
assign n_16239 = n_15680 ^ n_16227;
assign n_16240 = n_16228 ^ n_16227;
assign n_16241 = n_15680 ^ n_16228;
assign n_16242 = n_16229 ^ n_14146;
assign n_16243 = n_16230 ^ n_16229;
assign n_16244 = n_16230 ^ n_14146;
assign n_16245 = n_16232 & ~n_16231;
assign n_16246 = n_16232 ^ x257;
assign n_16247 = n_16233 ^ n_14398;
assign n_16248 = n_16234 ^ n_15494;
assign n_16249 = n_15863 ^ n_16234;
assign n_16250 = n_16235 ^ n_15331;
assign n_16251 = n_16237 ^ n_14398;
assign n_16252 = n_16237 ^ n_16233;
assign n_16253 = ~n_16238 & n_16236;
assign n_16254 = n_16238 ^ x124;
assign n_16255 = n_16240 & ~n_16239;
assign n_16256 = n_15024 & ~n_16240;
assign n_16257 = n_16241 ^ n_16227;
assign n_16258 = n_16242 & ~n_16243;
assign n_16259 = n_16244 ^ n_16229;
assign n_16260 = n_16245 ^ x257;
assign n_16261 = n_16219 & n_16246;
assign n_16262 = n_16246 ^ n_16219;
assign n_16263 = n_14823 & n_16248;
assign n_16264 = n_16250 ^ n_15532;
assign n_16265 = n_16251 ^ n_16233;
assign n_16266 = n_16247 & ~n_16252;
assign n_16267 = n_16253 ^ x124;
assign n_16268 = ~n_16226 & n_16254;
assign n_16269 = n_16254 ^ n_16226;
assign n_16270 = n_16255 ^ n_15680;
assign n_16271 = n_16256 ^ n_15680;
assign n_16272 = n_16258 ^ n_14146;
assign n_16273 = n_16259 ^ x256;
assign n_16274 = n_16260 ^ n_16259;
assign n_16275 = n_16263 ^ n_15494;
assign n_16276 = n_15352 ^ n_16264;
assign n_16277 = ~n_16264 & ~n_15547;
assign n_16278 = n_16265 ^ x123;
assign n_16279 = n_16266 ^ n_14398;
assign n_16280 = n_16267 ^ n_16265;
assign n_16281 = n_16269 ^ n_15697;
assign n_16282 = n_16270 ^ n_16269;
assign n_16283 = n_16270 ^ n_15697;
assign n_16284 = n_16271 ^ n_14189;
assign n_16285 = n_16272 ^ n_16271;
assign n_16286 = n_16272 ^ n_14189;
assign n_16287 = ~n_16274 & n_16273;
assign n_16288 = n_16274 ^ x256;
assign n_16289 = n_16275 ^ n_14441;
assign n_16290 = n_16276 ^ n_15532;
assign n_16291 = n_15886 ^ n_16276;
assign n_16292 = n_16277 ^ n_15352;
assign n_16293 = n_16279 ^ n_14441;
assign n_16294 = n_16279 ^ n_16275;
assign n_16295 = ~n_16280 & n_16278;
assign n_16296 = n_16280 ^ x123;
assign n_16297 = n_16282 & ~n_16281;
assign n_16298 = n_15043 & ~n_16282;
assign n_16299 = n_16283 ^ n_16269;
assign n_16300 = n_16284 & ~n_16285;
assign n_16301 = n_16286 ^ n_16271;
assign n_16302 = n_16287 ^ x256;
assign n_16303 = n_16261 & ~n_16288;
assign n_16304 = n_16288 ^ n_16261;
assign n_16305 = n_14846 & ~n_16290;
assign n_16306 = n_16292 ^ n_15574;
assign n_16307 = n_16293 ^ n_16275;
assign n_16308 = n_16289 & n_16294;
assign n_16309 = n_16295 ^ x123;
assign n_16310 = ~n_16268 & ~n_16296;
assign n_16311 = n_16296 ^ n_16268;
assign n_16312 = n_16297 ^ n_15697;
assign n_16313 = n_16298 ^ n_15697;
assign n_16314 = n_16300 ^ n_14189;
assign n_16315 = n_16301 ^ x271;
assign n_16316 = n_16302 ^ n_16301;
assign n_16317 = n_16305 ^ n_15532;
assign n_16318 = n_16306 ^ n_15374;
assign n_16319 = n_16307 ^ x122;
assign n_16320 = n_16308 ^ n_14441;
assign n_16321 = n_16309 ^ n_16307;
assign n_16322 = n_16311 ^ n_15713;
assign n_16323 = n_16311 ^ n_16312;
assign n_16324 = n_16312 ^ n_15713;
assign n_16325 = n_16314 ^ n_14234;
assign n_16326 = n_16313 ^ n_16314;
assign n_16327 = ~n_16316 & n_16315;
assign n_16328 = n_16316 ^ x271;
assign n_16329 = n_16317 ^ n_14483;
assign n_16330 = n_16318 ^ n_15574;
assign n_16331 = n_16318 ^ n_15885;
assign n_16332 = n_16320 ^ n_14483;
assign n_16333 = n_16320 ^ n_16317;
assign n_16334 = ~n_16321 & n_16319;
assign n_16335 = n_16321 ^ x122;
assign n_16336 = n_16323 & ~n_16322;
assign n_16337 = n_15063 & ~n_16323;
assign n_16338 = n_16324 ^ n_16311;
assign n_16339 = n_16313 ^ n_16325;
assign n_16340 = ~n_16325 & ~n_16326;
assign n_16341 = n_16327 ^ x271;
assign n_16342 = n_16328 & ~n_16303;
assign n_16343 = n_16303 ^ n_16328;
assign n_16344 = ~n_14866 & n_16330;
assign n_16345 = n_16331 ^ n_15899;
assign n_16346 = n_16332 ^ n_16317;
assign n_16347 = ~n_16329 & ~n_16333;
assign n_16348 = n_16334 ^ x122;
assign n_16349 = n_16310 & ~n_16335;
assign n_16350 = n_16335 ^ n_16310;
assign n_16351 = n_16336 ^ n_15713;
assign n_16352 = n_16337 ^ n_15713;
assign n_16353 = n_16339 ^ x270;
assign n_16354 = n_16340 ^ n_14234;
assign n_16355 = n_16341 ^ n_16339;
assign n_16356 = n_16344 ^ n_15574;
assign n_16357 = n_16346 ^ x121;
assign n_16358 = n_16347 ^ n_14483;
assign n_16359 = n_16348 ^ n_16346;
assign n_16360 = n_16350 ^ n_15726;
assign n_16361 = n_16350 ^ n_16351;
assign n_16362 = n_16351 ^ n_15726;
assign n_16363 = n_16352 ^ n_14277;
assign n_16364 = n_16354 ^ n_16352;
assign n_16365 = n_16354 ^ n_14277;
assign n_16366 = n_16355 & ~n_16353;
assign n_16367 = n_16355 ^ x270;
assign n_16368 = n_16356 ^ n_14513;
assign n_16369 = n_16358 ^ x120;
assign n_16370 = ~n_16359 & n_16357;
assign n_16371 = n_16359 ^ x121;
assign n_16372 = ~n_16361 & ~n_16360;
assign n_16373 = n_15082 & n_16361;
assign n_16374 = n_16362 ^ n_16350;
assign n_16375 = ~n_16363 & n_16364;
assign n_16376 = n_16365 ^ n_16352;
assign n_16377 = n_16366 ^ x270;
assign n_16378 = n_16342 & ~n_16367;
assign n_16379 = n_16367 ^ n_16342;
assign n_16380 = n_16369 ^ n_16368;
assign n_16381 = n_16370 ^ x121;
assign n_16382 = n_16349 & ~n_16371;
assign n_16383 = n_16371 ^ n_16349;
assign n_16384 = n_16372 ^ n_15726;
assign n_16385 = n_16373 ^ n_15726;
assign n_16386 = n_16375 ^ n_14277;
assign n_16387 = n_16376 ^ x269;
assign n_16388 = n_16377 ^ n_16376;
assign n_16389 = n_16381 ^ n_16382;
assign n_16390 = n_16383 ^ n_15743;
assign n_16391 = n_16383 ^ n_16384;
assign n_16392 = n_16384 ^ n_15743;
assign n_16393 = n_16385 ^ n_14320;
assign n_16394 = n_16386 ^ n_16385;
assign n_16395 = n_16386 ^ n_14320;
assign n_16396 = ~n_16388 & n_16387;
assign n_16397 = n_16388 ^ x269;
assign n_16398 = n_16389 ^ n_16380;
assign n_16399 = n_16391 & ~n_16390;
assign n_16400 = ~n_15103 & ~n_16391;
assign n_16401 = n_16392 ^ n_16383;
assign n_16402 = n_16393 & ~n_16394;
assign n_16403 = n_16395 ^ n_16385;
assign n_16404 = n_16396 ^ x269;
assign n_16405 = ~n_16378 & ~n_16397;
assign n_16406 = n_16397 ^ n_16378;
assign n_16407 = n_16398 ^ n_15763;
assign n_16408 = n_16399 ^ n_15743;
assign n_16409 = n_16400 ^ n_15743;
assign n_16410 = n_16402 ^ n_14320;
assign n_16411 = n_16403 ^ x268;
assign n_16412 = n_16404 ^ n_16403;
assign n_16413 = n_16398 ^ n_16408;
assign n_16414 = n_16408 ^ n_15763;
assign n_16415 = n_16409 ^ n_14362;
assign n_16416 = n_16410 ^ n_16409;
assign n_16417 = n_16410 ^ n_14362;
assign n_16418 = n_16412 & ~n_16411;
assign n_16419 = n_16412 ^ x268;
assign n_16420 = ~n_16413 & n_16407;
assign n_16421 = n_15124 & n_16413;
assign n_16422 = n_16414 ^ n_16398;
assign n_16423 = ~n_16415 & ~n_16416;
assign n_16424 = n_16417 ^ n_16409;
assign n_16425 = n_16418 ^ x268;
assign n_16426 = ~n_16405 & ~n_16419;
assign n_16427 = n_16419 ^ n_16405;
assign n_16428 = n_16420 ^ n_15763;
assign n_16429 = n_16421 ^ n_15763;
assign n_16430 = n_16423 ^ n_14362;
assign n_16431 = n_16424 ^ x267;
assign n_16432 = n_16425 ^ n_16424;
assign n_16433 = n_16425 ^ x267;
assign n_16434 = n_16428 ^ n_15783;
assign n_16435 = n_15789 ^ n_16428;
assign n_16436 = n_16429 ^ n_14405;
assign n_16437 = n_16430 ^ n_16429;
assign n_16438 = n_16430 ^ n_14405;
assign n_16439 = n_16431 & ~n_16432;
assign n_16440 = n_16433 ^ n_16424;
assign n_16441 = n_15789 & n_16434;
assign n_16442 = n_16435 ^ n_15783;
assign n_16443 = ~n_16436 & n_16437;
assign n_16444 = n_16438 ^ n_16429;
assign n_16445 = n_16439 ^ x267;
assign n_16446 = ~n_16426 & ~n_16440;
assign n_16447 = n_16440 ^ n_16426;
assign n_16448 = n_16441 ^ n_15447;
assign n_16449 = ~n_15145 & ~n_16442;
assign n_16450 = n_16443 ^ n_14405;
assign n_16451 = n_16444 ^ x266;
assign n_16452 = n_16445 ^ n_16444;
assign n_16453 = n_15935 & ~n_16447;
assign n_16454 = n_16447 ^ n_15935;
assign n_16455 = n_16448 ^ n_15804;
assign n_16456 = n_16449 ^ n_15783;
assign n_16457 = n_16450 ^ n_14448;
assign n_16458 = n_16452 & ~n_16451;
assign n_16459 = n_16452 ^ x266;
assign n_16460 = n_15962 ^ n_16453;
assign n_16461 = n_16454 ^ n_15927;
assign n_16462 = ~n_16455 & n_15811;
assign n_16463 = n_16455 ^ n_15486;
assign n_16464 = n_16456 ^ n_16450;
assign n_16465 = n_16456 ^ n_16457;
assign n_16466 = n_16458 ^ x266;
assign n_16467 = ~n_16446 & ~n_16459;
assign n_16468 = n_16459 ^ n_16446;
assign n_16469 = ~n_15401 & n_16461;
assign n_16470 = n_16462 ^ n_15486;
assign n_16471 = n_16463 ^ n_15804;
assign n_16472 = n_16457 & ~n_16464;
assign n_16473 = n_16465 ^ x265;
assign n_16474 = n_16466 ^ n_16465;
assign n_16475 = n_16468 ^ n_16453;
assign n_16476 = n_16468 ^ n_16460;
assign n_16477 = n_16469 ^ n_15927;
assign n_16478 = n_16470 ^ n_15824;
assign n_16479 = n_15166 & n_16471;
assign n_16480 = n_16472 ^ n_14448;
assign n_16481 = ~n_16474 & n_16473;
assign n_16482 = n_16474 ^ x265;
assign n_16483 = n_16460 & ~n_16475;
assign n_16484 = ~n_15428 & n_16475;
assign n_16485 = n_14840 & ~n_16477;
assign n_16486 = n_16477 ^ n_14840;
assign n_16487 = n_16477 ^ n_14849;
assign n_16488 = n_16478 & n_15831;
assign n_16489 = n_16478 ^ n_15552;
assign n_16490 = n_16479 ^ n_15804;
assign n_16491 = n_16480 ^ n_14490;
assign n_16492 = n_16481 ^ x265;
assign n_16493 = n_16482 & n_16467;
assign n_16494 = n_16467 ^ n_16482;
assign n_16495 = n_16483 ^ n_15962;
assign n_16496 = n_16484 ^ n_15962;
assign n_16497 = n_16485 ^ n_14869;
assign n_16498 = x423 & ~n_16486;
assign n_16499 = n_16488 ^ n_15552;
assign n_16500 = n_16489 ^ n_15824;
assign n_16501 = n_16490 ^ n_14490;
assign n_16502 = n_16490 ^ n_16480;
assign n_16503 = n_16490 ^ n_16491;
assign n_16504 = n_16492 ^ x264;
assign n_16505 = n_16011 ^ n_16494;
assign n_16506 = n_16495 ^ n_16494;
assign n_16507 = n_16495 ^ n_16011;
assign n_16508 = n_16496 ^ n_16485;
assign n_16509 = n_16496 ^ n_16497;
assign n_16510 = n_16498 ^ x422;
assign n_16511 = n_16499 ^ n_15847;
assign n_16512 = n_15590 ^ n_16499;
assign n_16513 = n_15187 & ~n_16500;
assign n_16514 = n_16501 & ~n_16502;
assign n_16515 = n_16492 ^ n_16503;
assign n_16516 = ~n_16505 & ~n_16506;
assign n_16517 = n_15472 & n_16506;
assign n_16518 = n_16507 ^ n_16494;
assign n_16519 = n_16497 & ~n_16508;
assign n_16520 = n_16509 ^ n_16498;
assign n_16521 = ~n_15853 & n_16511;
assign n_16522 = ~n_15211 & n_16512;
assign n_16523 = n_16512 ^ n_15847;
assign n_16524 = n_16513 ^ n_15824;
assign n_16525 = n_16514 ^ n_14490;
assign n_16526 = ~n_16515 & n_16504;
assign n_16527 = n_16515 ^ x264;
assign n_16528 = n_16516 ^ n_16011;
assign n_16529 = n_16517 ^ n_16011;
assign n_16530 = n_16519 ^ n_14869;
assign n_16531 = ~n_16520 & n_16510;
assign n_16532 = n_16520 ^ x422;
assign n_16533 = n_16521 ^ n_15590;
assign n_16534 = n_16522 ^ n_15847;
assign n_16535 = n_16524 ^ n_14533;
assign n_16536 = n_16525 ^ n_16524;
assign n_16537 = n_16526 ^ x264;
assign n_16538 = n_16527 & n_16493;
assign n_16539 = n_16493 ^ n_16527;
assign n_16540 = n_16053 ^ n_16528;
assign n_16541 = n_16529 ^ n_14909;
assign n_16542 = n_16530 ^ n_16529;
assign n_16543 = n_16530 ^ n_14909;
assign n_16544 = n_16531 ^ x422;
assign n_16545 = ~n_16487 & n_16532;
assign n_16546 = n_16532 ^ n_16487;
assign n_16547 = n_16533 ^ n_15866;
assign n_16548 = n_16534 ^ n_14568;
assign n_16549 = n_16536 & n_16535;
assign n_16550 = n_16536 ^ n_14533;
assign n_16551 = n_16537 ^ x279;
assign n_16552 = n_16539 ^ n_16528;
assign n_16553 = n_16539 ^ n_16540;
assign n_16554 = ~n_16541 & n_16542;
assign n_16555 = n_16543 ^ n_16529;
assign n_16556 = n_16544 ^ x421;
assign n_16557 = ~n_16547 & ~n_15874;
assign n_16558 = n_15624 ^ n_16547;
assign n_16559 = n_16549 ^ n_14533;
assign n_16560 = n_16550 ^ x279;
assign n_16561 = n_16550 ^ n_16537;
assign n_16562 = n_16550 ^ n_16551;
assign n_16563 = n_16540 & n_16552;
assign n_16564 = n_15514 & ~n_16552;
assign n_16565 = n_16554 ^ n_14909;
assign n_16566 = n_16544 ^ n_16555;
assign n_16567 = n_16557 ^ n_15624;
assign n_16568 = n_16558 ^ n_15866;
assign n_16569 = n_16534 ^ n_16559;
assign n_16570 = n_16559 ^ n_14568;
assign n_16571 = n_16560 & ~n_16561;
assign n_16572 = n_16562 & n_16538;
assign n_16573 = n_16538 ^ n_16562;
assign n_16574 = n_16563 ^ n_16053;
assign n_16575 = n_16564 ^ n_16053;
assign n_16576 = n_16565 ^ n_14933;
assign n_16577 = n_16566 & n_16556;
assign n_16578 = n_16566 ^ x421;
assign n_16579 = n_16567 ^ n_15887;
assign n_16580 = n_16567 ^ n_15652;
assign n_16581 = ~n_15229 & ~n_16568;
assign n_16582 = ~n_16548 & n_16569;
assign n_16583 = n_16534 ^ n_16570;
assign n_16584 = n_16571 ^ x279;
assign n_16585 = n_16092 ^ n_16573;
assign n_16586 = n_16574 ^ n_16573;
assign n_16587 = n_16574 ^ n_16092;
assign n_16588 = n_16575 ^ n_14933;
assign n_16589 = n_16565 ^ n_16575;
assign n_16590 = n_16576 ^ n_16575;
assign n_16591 = n_16577 ^ x421;
assign n_16592 = ~n_16545 & n_16578;
assign n_16593 = n_16578 ^ n_16545;
assign n_16594 = n_15893 & n_16579;
assign n_16595 = n_15249 & ~n_16580;
assign n_16596 = n_16580 ^ n_15887;
assign n_16597 = n_16581 ^ n_15866;
assign n_16598 = n_16582 ^ n_14568;
assign n_16599 = n_16583 ^ x278;
assign n_16600 = n_16584 ^ n_16583;
assign n_16601 = n_16585 & n_16586;
assign n_16602 = ~n_15556 & ~n_16586;
assign n_16603 = n_16587 ^ n_16573;
assign n_16604 = ~n_16588 & n_16589;
assign n_16605 = n_16591 ^ n_16590;
assign n_16606 = n_16591 ^ x420;
assign n_16607 = n_16594 ^ n_15652;
assign n_16608 = n_16595 ^ n_15887;
assign n_16609 = n_16597 ^ n_14595;
assign n_16610 = n_16598 ^ n_16597;
assign n_16611 = n_16598 ^ n_14595;
assign n_16612 = ~n_16600 & n_16599;
assign n_16613 = n_16600 ^ x278;
assign n_16614 = n_16601 ^ n_16092;
assign n_16615 = n_16602 ^ n_16092;
assign n_16616 = n_16604 ^ n_14933;
assign n_16617 = n_16605 ^ x420;
assign n_16618 = n_16605 & n_16606;
assign n_16619 = n_16607 ^ n_15908;
assign n_16620 = n_16608 ^ n_14618;
assign n_16621 = ~n_16609 & ~n_16610;
assign n_16622 = n_16611 ^ n_16597;
assign n_16623 = n_16612 ^ x278;
assign n_16624 = ~n_16613 & ~n_16572;
assign n_16625 = n_16572 ^ n_16613;
assign n_16626 = n_16131 ^ n_16614;
assign n_16627 = n_16615 ^ n_14957;
assign n_16628 = n_16616 ^ n_16615;
assign n_16629 = n_16616 ^ n_14957;
assign n_16630 = ~n_16592 & ~n_16617;
assign n_16631 = n_16617 ^ n_16592;
assign n_16632 = n_16618 ^ x420;
assign n_16633 = n_16619 & ~n_15916;
assign n_16634 = n_15674 ^ n_16619;
assign n_16635 = n_16621 ^ n_14595;
assign n_16636 = n_16622 ^ x277;
assign n_16637 = n_16623 ^ n_16622;
assign n_16638 = n_16625 ^ n_16131;
assign n_16639 = n_16625 ^ n_16614;
assign n_16640 = n_16625 ^ n_16626;
assign n_16641 = ~n_16627 & ~n_16628;
assign n_16642 = n_16629 ^ n_16615;
assign n_16643 = n_16632 ^ x419;
assign n_16644 = n_16633 ^ n_15674;
assign n_16645 = n_16634 ^ n_15908;
assign n_16646 = n_16634 ^ n_15987;
assign n_16647 = n_16635 ^ n_16608;
assign n_16648 = n_16635 ^ n_14618;
assign n_16649 = ~n_16637 & n_16636;
assign n_16650 = n_16637 ^ x277;
assign n_16651 = ~n_16638 & n_16639;
assign n_16652 = ~n_15594 & ~n_16639;
assign n_16653 = n_16487 ^ n_16640;
assign n_16654 = n_16641 ^ n_14957;
assign n_16655 = n_16632 ^ n_16642;
assign n_16656 = n_16644 ^ n_15929;
assign n_16657 = n_15270 & n_16645;
assign n_16658 = ~n_16620 & n_16647;
assign n_16659 = n_16648 ^ n_16608;
assign n_16660 = n_16649 ^ x277;
assign n_16661 = n_16650 & ~n_16624;
assign n_16662 = n_16624 ^ n_16650;
assign n_16663 = n_16651 ^ n_16131;
assign n_16664 = n_16652 ^ n_16131;
assign n_16665 = n_16654 ^ n_14974;
assign n_16666 = n_16655 & n_16643;
assign n_16667 = n_16655 ^ x419;
assign n_16668 = n_16656 & n_15938;
assign n_16669 = n_15693 ^ n_16656;
assign n_16670 = n_16657 ^ n_15908;
assign n_16671 = n_16658 ^ n_14618;
assign n_16672 = n_16659 ^ x276;
assign n_16673 = n_16660 ^ n_16659;
assign n_16674 = n_16173 ^ n_16662;
assign n_16675 = n_16663 ^ n_16662;
assign n_16676 = n_16663 ^ n_16173;
assign n_16677 = n_16664 ^ n_16654;
assign n_16678 = n_16664 ^ n_16665;
assign n_16679 = n_16666 ^ x419;
assign n_16680 = n_16630 & ~n_16667;
assign n_16681 = n_16667 ^ n_16630;
assign n_16682 = n_16668 ^ n_15693;
assign n_16683 = n_16669 ^ n_15929;
assign n_16684 = n_16027 ^ n_16669;
assign n_16685 = n_16670 ^ n_14638;
assign n_16686 = n_16671 ^ n_16670;
assign n_16687 = n_16671 ^ n_14638;
assign n_16688 = n_16673 & ~n_16672;
assign n_16689 = n_16673 ^ x276;
assign n_16690 = n_16674 & n_16675;
assign n_16691 = ~n_15628 & ~n_16675;
assign n_16692 = n_16676 ^ n_16662;
assign n_16693 = n_16665 & n_16677;
assign n_16694 = n_16678 ^ x418;
assign n_16695 = n_16679 ^ n_16678;
assign n_16696 = n_16682 ^ n_15955;
assign n_16697 = ~n_15291 & ~n_16683;
assign n_16698 = ~n_16685 & ~n_16686;
assign n_16699 = n_16687 ^ n_16670;
assign n_16700 = n_16688 ^ x276;
assign n_16701 = n_16689 & ~n_16661;
assign n_16702 = n_16661 ^ n_16689;
assign n_16703 = n_16690 ^ n_16173;
assign n_16704 = n_16691 ^ n_16173;
assign n_16705 = n_16546 ^ n_16692;
assign n_16706 = n_16693 ^ n_14974;
assign n_16707 = ~n_16695 & n_16694;
assign n_16708 = n_16695 ^ x418;
assign n_16709 = n_16696 & n_15966;
assign n_16710 = n_15710 ^ n_16696;
assign n_16711 = n_16697 ^ n_15929;
assign n_16712 = n_16698 ^ n_14638;
assign n_16713 = n_16699 ^ x275;
assign n_16714 = n_16700 ^ n_16699;
assign n_16715 = n_16215 ^ n_16702;
assign n_16716 = n_16703 ^ n_16702;
assign n_16717 = n_16703 ^ n_16215;
assign n_16718 = n_16706 ^ n_14993;
assign n_16719 = n_16704 ^ n_16706;
assign n_16720 = n_16707 ^ x418;
assign n_16721 = n_16680 & n_16708;
assign n_16722 = n_16708 ^ n_16680;
assign n_16723 = n_16709 ^ n_15710;
assign n_16724 = n_16710 ^ n_15955;
assign n_16725 = n_16088 ^ n_16710;
assign n_16726 = n_16711 ^ n_14659;
assign n_16727 = n_16712 ^ n_16711;
assign n_16728 = n_16714 & ~n_16713;
assign n_16729 = n_16714 ^ x275;
assign n_16730 = n_16715 & n_16716;
assign n_16731 = n_15656 & ~n_16716;
assign n_16732 = n_16717 ^ n_16702;
assign n_16733 = n_16704 ^ n_16718;
assign n_16734 = ~n_16718 & ~n_16719;
assign n_16735 = n_16720 ^ x417;
assign n_16736 = n_16723 ^ n_15988;
assign n_16737 = n_15312 & ~n_16724;
assign n_16738 = n_16727 & n_16726;
assign n_16739 = n_16727 ^ n_14659;
assign n_16740 = n_16728 ^ x275;
assign n_16741 = n_16729 & n_16701;
assign n_16742 = n_16701 ^ n_16729;
assign n_16743 = n_16730 ^ n_16215;
assign n_16744 = n_16731 ^ n_16215;
assign n_16745 = n_16593 ^ n_16732;
assign n_16746 = n_16720 ^ n_16733;
assign n_16747 = n_16734 ^ n_14993;
assign n_16748 = n_15733 ^ n_16736;
assign n_16749 = ~n_16736 & ~n_16001;
assign n_16750 = n_16737 ^ n_15955;
assign n_16751 = n_16738 ^ n_14659;
assign n_16752 = n_16739 ^ x274;
assign n_16753 = n_16740 ^ n_16739;
assign n_16754 = n_16257 ^ n_16742;
assign n_16755 = n_16743 ^ n_16742;
assign n_16756 = n_16743 ^ n_16257;
assign n_16757 = n_16744 ^ n_15006;
assign n_16758 = ~n_16746 & n_16735;
assign n_16759 = n_16746 ^ x417;
assign n_16760 = n_16747 ^ n_16744;
assign n_16761 = n_16747 ^ n_15006;
assign n_16762 = n_16748 ^ n_15988;
assign n_16763 = n_16135 ^ n_16748;
assign n_16764 = n_16749 ^ n_15733;
assign n_16765 = n_16750 ^ n_14680;
assign n_16766 = n_16751 ^ n_16750;
assign n_16767 = n_16751 ^ n_14680;
assign n_16768 = n_16753 & ~n_16752;
assign n_16769 = n_16753 ^ x274;
assign n_16770 = n_16754 & n_16755;
assign n_16771 = n_15680 & ~n_16755;
assign n_16772 = n_16756 ^ n_16742;
assign n_16773 = n_16758 ^ x417;
assign n_16774 = n_16721 & n_16759;
assign n_16775 = n_16759 ^ n_16721;
assign n_16776 = ~n_16757 & ~n_16760;
assign n_16777 = n_16761 ^ n_16744;
assign n_16778 = n_15333 & ~n_16762;
assign n_16779 = n_16030 ^ n_16764;
assign n_16780 = n_16765 & n_16766;
assign n_16781 = n_16767 ^ n_16750;
assign n_16782 = n_16768 ^ x274;
assign n_16783 = ~n_16769 & ~n_16741;
assign n_16784 = n_16741 ^ n_16769;
assign n_16785 = n_16770 ^ n_16257;
assign n_16786 = n_16771 ^ n_16257;
assign n_16787 = n_16631 ^ n_16772;
assign n_16788 = n_16773 ^ x416;
assign n_16789 = n_16776 ^ n_15006;
assign n_16790 = n_16773 ^ n_16777;
assign n_16791 = n_16778 ^ n_15988;
assign n_16792 = n_15758 ^ n_16779;
assign n_16793 = n_16779 & n_16044;
assign n_16794 = n_16780 ^ n_14680;
assign n_16795 = n_16781 ^ x273;
assign n_16796 = n_16782 ^ n_16781;
assign n_16797 = n_16299 ^ n_16784;
assign n_16798 = n_16785 ^ n_16784;
assign n_16799 = n_16785 ^ n_16299;
assign n_16800 = n_16786 ^ n_15024;
assign n_16801 = n_16789 ^ n_16786;
assign n_16802 = n_16789 ^ n_15024;
assign n_16803 = n_16790 & n_16788;
assign n_16804 = n_16790 ^ x416;
assign n_16805 = n_16791 ^ n_14695;
assign n_16806 = n_16792 ^ n_16015;
assign n_16807 = n_16792 ^ n_16178;
assign n_16808 = n_16793 ^ n_15758;
assign n_16809 = n_16794 ^ n_16791;
assign n_16810 = n_16794 ^ n_14695;
assign n_16811 = ~n_16796 & n_16795;
assign n_16812 = n_16796 ^ x273;
assign n_16813 = ~n_16797 & n_16798;
assign n_16814 = n_15697 & ~n_16798;
assign n_16815 = n_16799 ^ n_16784;
assign n_16816 = ~n_16800 & ~n_16801;
assign n_16817 = n_16802 ^ n_16786;
assign n_16818 = n_16803 ^ x416;
assign n_16819 = n_16774 & ~n_16804;
assign n_16820 = n_16804 ^ n_16774;
assign n_16821 = ~n_15354 & n_16806;
assign n_16822 = n_15781 ^ n_16808;
assign n_16823 = n_16808 ^ n_16068;
assign n_16824 = ~n_16805 & ~n_16809;
assign n_16825 = n_16810 ^ n_16791;
assign n_16826 = n_16811 ^ x273;
assign n_16827 = ~n_16812 & ~n_16783;
assign n_16828 = n_16783 ^ n_16812;
assign n_16829 = n_16813 ^ n_16299;
assign n_16830 = n_16814 ^ n_16299;
assign n_16831 = n_16681 ^ n_16815;
assign n_16832 = n_16816 ^ n_15024;
assign n_16833 = n_16817 ^ x431;
assign n_16834 = n_16818 ^ n_16817;
assign n_16835 = n_16821 ^ n_16015;
assign n_16836 = n_16822 ^ n_16068;
assign n_16837 = ~n_16082 & n_16823;
assign n_16838 = n_16824 ^ n_14695;
assign n_16839 = n_16825 ^ x272;
assign n_16840 = n_16826 ^ n_16825;
assign n_16841 = n_16338 ^ n_16828;
assign n_16842 = n_16829 ^ n_16828;
assign n_16843 = n_16829 ^ n_16338;
assign n_16844 = n_16830 ^ n_15043;
assign n_16845 = n_16832 ^ n_16830;
assign n_16846 = n_16832 ^ n_15043;
assign n_16847 = ~n_16834 & n_16833;
assign n_16848 = n_16834 ^ x431;
assign n_16849 = n_16835 ^ n_14717;
assign n_16850 = n_16836 ^ n_16056;
assign n_16851 = n_16836 ^ n_16220;
assign n_16852 = n_16837 ^ n_15781;
assign n_16853 = n_16838 ^ n_16835;
assign n_16854 = ~n_16840 & n_16839;
assign n_16855 = n_16840 ^ x272;
assign n_16856 = n_16841 & ~n_16842;
assign n_16857 = n_15713 & n_16842;
assign n_16858 = n_16843 ^ n_16828;
assign n_16859 = ~n_16844 & n_16845;
assign n_16860 = n_16846 ^ n_16830;
assign n_16861 = n_16847 ^ x431;
assign n_16862 = ~n_16819 & ~n_16848;
assign n_16863 = n_16848 ^ n_16819;
assign n_16864 = ~n_15376 & ~n_16850;
assign n_16865 = n_16852 ^ n_16108;
assign n_16866 = n_16853 ^ n_14717;
assign n_16867 = ~n_16853 & ~n_16849;
assign n_16868 = n_16854 ^ x272;
assign n_16869 = n_16855 & ~n_16827;
assign n_16870 = n_16827 ^ n_16855;
assign n_16871 = n_16856 ^ n_16338;
assign n_16872 = n_16857 ^ n_16338;
assign n_16873 = n_16722 ^ n_16858;
assign n_16874 = n_16859 ^ n_15043;
assign n_16875 = n_16860 ^ x430;
assign n_16876 = n_16861 ^ n_16860;
assign n_16877 = n_16864 ^ n_16056;
assign n_16878 = n_15802 ^ n_16865;
assign n_16879 = ~n_16865 & ~n_16124;
assign n_16880 = n_16866 ^ x287;
assign n_16881 = n_16867 ^ n_14717;
assign n_16882 = n_16868 ^ n_16866;
assign n_16883 = n_16868 ^ x287;
assign n_16884 = n_16374 ^ n_16870;
assign n_16885 = n_16871 ^ n_16870;
assign n_16886 = n_16871 ^ n_16374;
assign n_16887 = n_16872 ^ n_15063;
assign n_16888 = n_16874 ^ n_16872;
assign n_16889 = n_16874 ^ n_15063;
assign n_16890 = n_16876 & ~n_16875;
assign n_16891 = n_16876 ^ x430;
assign n_16892 = n_16877 ^ n_14743;
assign n_16893 = n_16878 ^ n_16108;
assign n_16894 = n_16262 ^ n_16878;
assign n_16895 = n_16879 ^ n_15802;
assign n_16896 = n_16881 ^ n_14743;
assign n_16897 = n_16881 ^ n_16877;
assign n_16898 = ~n_16880 & n_16882;
assign n_16899 = n_16883 ^ n_16866;
assign n_16900 = n_16884 & ~n_16885;
assign n_16901 = ~n_15726 & n_16885;
assign n_16902 = n_16886 ^ n_16870;
assign n_16903 = ~n_16887 & n_16888;
assign n_16904 = n_16889 ^ n_16872;
assign n_16905 = n_16890 ^ x430;
assign n_16906 = ~n_16862 & ~n_16891;
assign n_16907 = n_16891 ^ n_16862;
assign n_16908 = n_15396 & ~n_16893;
assign n_16909 = n_16895 ^ n_16150;
assign n_16910 = n_16896 ^ n_16877;
assign n_16911 = ~n_16892 & ~n_16897;
assign n_16912 = n_16898 ^ x287;
assign n_16913 = n_16899 & ~n_16869;
assign n_16914 = n_16869 ^ n_16899;
assign n_16915 = n_16900 ^ n_16374;
assign n_16916 = n_16901 ^ n_16374;
assign n_16917 = n_16775 ^ n_16902;
assign n_16918 = n_16903 ^ n_15063;
assign n_16919 = n_16904 ^ x429;
assign n_16920 = n_16905 ^ n_16904;
assign n_16921 = n_16908 ^ n_16108;
assign n_16922 = n_15823 ^ n_16909;
assign n_16923 = n_16909 & ~n_16165;
assign n_16924 = n_16910 ^ x286;
assign n_16925 = n_16911 ^ n_14743;
assign n_16926 = n_16912 ^ n_16910;
assign n_16927 = n_16401 ^ n_16914;
assign n_16928 = n_16914 ^ n_16915;
assign n_16929 = n_16401 ^ n_16915;
assign n_16930 = n_16916 ^ n_15082;
assign n_16931 = n_16918 ^ n_16916;
assign n_16932 = n_16918 ^ n_15082;
assign n_16933 = n_16920 & ~n_16919;
assign n_16934 = n_16920 ^ x429;
assign n_16935 = n_16921 ^ n_14762;
assign n_16936 = n_16922 ^ n_16150;
assign n_16937 = n_16304 ^ n_16922;
assign n_16938 = n_16923 ^ n_15823;
assign n_16939 = n_16925 ^ n_14762;
assign n_16940 = n_16925 ^ n_16921;
assign n_16941 = n_16926 ^ x286;
assign n_16942 = ~n_16926 & n_16924;
assign n_16943 = n_16928 & n_16927;
assign n_16944 = ~n_15743 & ~n_16928;
assign n_16945 = n_16929 ^ n_16914;
assign n_16946 = ~n_16930 & n_16931;
assign n_16947 = n_16932 ^ n_16916;
assign n_16948 = n_16933 ^ x429;
assign n_16949 = ~n_16934 & n_16906;
assign n_16950 = n_16906 ^ n_16934;
assign n_16951 = n_15422 & n_16936;
assign n_16952 = n_16938 ^ n_16192;
assign n_16953 = n_16939 ^ n_16921;
assign n_16954 = n_16935 & n_16940;
assign n_16955 = n_16941 & ~n_16913;
assign n_16956 = n_16913 ^ n_16941;
assign n_16957 = n_16942 ^ x286;
assign n_16958 = n_16943 ^ n_16401;
assign n_16959 = n_16944 ^ n_16401;
assign n_16960 = n_16820 ^ n_16945;
assign n_16961 = n_16946 ^ n_15082;
assign n_16962 = n_16947 ^ x428;
assign n_16963 = n_16948 ^ n_16947;
assign n_16964 = n_16951 ^ n_16150;
assign n_16965 = n_15844 ^ n_16952;
assign n_16966 = n_16952 & ~n_16207;
assign n_16967 = n_16953 ^ x285;
assign n_16968 = n_16954 ^ n_14762;
assign n_16969 = n_16422 ^ n_16956;
assign n_16970 = n_16957 ^ n_16953;
assign n_16971 = n_16956 ^ n_16958;
assign n_16972 = n_16422 ^ n_16958;
assign n_16973 = n_16959 ^ n_15103;
assign n_16974 = n_16961 ^ n_16959;
assign n_16975 = n_16961 ^ n_15103;
assign n_16976 = n_16963 & ~n_16962;
assign n_16977 = n_16963 ^ x428;
assign n_16978 = n_16964 ^ n_14782;
assign n_16979 = n_16965 ^ n_16192;
assign n_16980 = n_16343 ^ n_16965;
assign n_16981 = n_16966 ^ n_15844;
assign n_16982 = n_16968 ^ n_14782;
assign n_16983 = n_16968 ^ n_16964;
assign n_16984 = n_16970 ^ x285;
assign n_16985 = ~n_16970 & n_16967;
assign n_16986 = n_16971 & n_16969;
assign n_16987 = ~n_15763 & ~n_16971;
assign n_16988 = n_16972 ^ n_16956;
assign n_16989 = ~n_16973 & ~n_16974;
assign n_16990 = n_16975 ^ n_16959;
assign n_16991 = n_16976 ^ x428;
assign n_16992 = ~n_16949 & n_16977;
assign n_16993 = n_16977 ^ n_16949;
assign n_16994 = n_15455 & n_16979;
assign n_16995 = n_16981 ^ n_16234;
assign n_16996 = n_16982 ^ n_16964;
assign n_16997 = ~n_16978 & ~n_16983;
assign n_16998 = n_16955 ^ n_16984;
assign n_16999 = ~n_16984 & ~n_16955;
assign n_17000 = n_16985 ^ x285;
assign n_17001 = n_16986 ^ n_16422;
assign n_17002 = n_16987 ^ n_16422;
assign n_17003 = n_16863 ^ n_16988;
assign n_17004 = n_16989 ^ n_15103;
assign n_17005 = n_16990 ^ x427;
assign n_17006 = n_16991 ^ n_16990;
assign n_17007 = n_16994 ^ n_16192;
assign n_17008 = n_15863 ^ n_16995;
assign n_17009 = n_16995 & n_16249;
assign n_17010 = n_16996 ^ x284;
assign n_17011 = n_16997 ^ n_14782;
assign n_17012 = n_16998 ^ n_16435;
assign n_17013 = n_17000 ^ n_16996;
assign n_17014 = n_16998 ^ n_17001;
assign n_17015 = n_17001 ^ n_16435;
assign n_17016 = n_17002 ^ n_15124;
assign n_17017 = n_17004 ^ n_17002;
assign n_17018 = n_17004 ^ n_15124;
assign n_17019 = n_17006 & ~n_17005;
assign n_17020 = n_17006 ^ x427;
assign n_17021 = n_17007 ^ n_14802;
assign n_17022 = n_17008 ^ n_16234;
assign n_17023 = n_16379 ^ n_17008;
assign n_17024 = n_17009 ^ n_15863;
assign n_17025 = n_17000 ^ n_17010;
assign n_17026 = n_17011 ^ n_17007;
assign n_17027 = n_17010 & ~n_17013;
assign n_17028 = ~n_17014 & n_17012;
assign n_17029 = n_15783 & n_17014;
assign n_17030 = n_17015 ^ n_16998;
assign n_17031 = ~n_17016 & ~n_17017;
assign n_17032 = n_17018 ^ n_17002;
assign n_17033 = n_17019 ^ x427;
assign n_17034 = ~n_16992 & ~n_17020;
assign n_17035 = n_17020 ^ n_16992;
assign n_17036 = n_17011 ^ n_17021;
assign n_17037 = ~n_15494 & ~n_17022;
assign n_17038 = n_17024 ^ n_16276;
assign n_17039 = n_17025 ^ n_16999;
assign n_17040 = ~n_16999 & n_17025;
assign n_17041 = n_17021 & n_17026;
assign n_17042 = n_17027 ^ x284;
assign n_17043 = n_17028 ^ n_16435;
assign n_17044 = n_17029 ^ n_16435;
assign n_17045 = n_16907 ^ n_17030;
assign n_17046 = n_17031 ^ n_15124;
assign n_17047 = n_17032 ^ x426;
assign n_17048 = n_17033 ^ n_17032;
assign n_17049 = n_17036 ^ x283;
assign n_17050 = n_17037 ^ n_16234;
assign n_17051 = n_15886 ^ n_17038;
assign n_17052 = n_17038 & n_16291;
assign n_17053 = n_17041 ^ n_14802;
assign n_17054 = n_17042 ^ n_17036;
assign n_17055 = n_17043 ^ n_16463;
assign n_17056 = n_17039 ^ n_17043;
assign n_17057 = n_17044 ^ n_15145;
assign n_17058 = n_17046 ^ n_17044;
assign n_17059 = n_17046 ^ n_15145;
assign n_17060 = ~n_17048 & n_17047;
assign n_17061 = n_17048 ^ x426;
assign n_17062 = n_17050 ^ n_14823;
assign n_17063 = n_17051 ^ n_16276;
assign n_17064 = n_16406 ^ n_17051;
assign n_17065 = n_17052 ^ n_15886;
assign n_17066 = n_17053 ^ n_14823;
assign n_17067 = n_17053 ^ n_17050;
assign n_17068 = n_17054 ^ x283;
assign n_17069 = ~n_17054 & n_17049;
assign n_17070 = n_17039 ^ n_17055;
assign n_17071 = ~n_17055 & ~n_17056;
assign n_17072 = n_15804 & n_17056;
assign n_17073 = n_17057 & n_17058;
assign n_17074 = n_17059 ^ n_17044;
assign n_17075 = n_17060 ^ x426;
assign n_17076 = ~n_17061 & ~n_17034;
assign n_17077 = n_17034 ^ n_17061;
assign n_17078 = ~n_15532 & ~n_17063;
assign n_17079 = n_17065 ^ n_16345;
assign n_17080 = n_17066 ^ n_17050;
assign n_17081 = ~n_17062 & ~n_17067;
assign n_17082 = n_17040 ^ n_17068;
assign n_17083 = n_17068 & n_17040;
assign n_17084 = n_17069 ^ x283;
assign n_17085 = n_16950 ^ n_17070;
assign n_17086 = n_17071 ^ n_16463;
assign n_17087 = n_17072 ^ n_16463;
assign n_17088 = n_17073 ^ n_15145;
assign n_17089 = n_17074 ^ x425;
assign n_17090 = n_17075 ^ n_17074;
assign n_17091 = n_17078 ^ n_16276;
assign n_17092 = n_17079 ^ n_16318;
assign n_17093 = n_17080 ^ x282;
assign n_17094 = n_17081 ^ n_14823;
assign n_17095 = n_17082 ^ n_16489;
assign n_17096 = n_17084 ^ n_17080;
assign n_17097 = n_17086 ^ n_17082;
assign n_17098 = n_17087 ^ n_15166;
assign n_17099 = n_17088 ^ n_17087;
assign n_17100 = n_17088 ^ n_15166;
assign n_17101 = ~n_17090 & n_17089;
assign n_17102 = n_17090 ^ x425;
assign n_17103 = n_17091 ^ n_14846;
assign n_17104 = n_15574 & ~n_17092;
assign n_17105 = n_17094 ^ n_14846;
assign n_17106 = n_17094 ^ n_17091;
assign n_17107 = n_17095 ^ n_17086;
assign n_17108 = n_17096 ^ x282;
assign n_17109 = ~n_17096 & n_17093;
assign n_17110 = ~n_15824 & n_17097;
assign n_17111 = ~n_17097 & n_17095;
assign n_17112 = n_17098 & n_17099;
assign n_17113 = n_17100 ^ n_17087;
assign n_17114 = n_17101 ^ x425;
assign n_17115 = ~n_17102 & n_17076;
assign n_17116 = n_17076 ^ n_17102;
assign n_17117 = n_17104 ^ n_16318;
assign n_17118 = n_17105 ^ n_17091;
assign n_17119 = n_17103 & ~n_17106;
assign n_17120 = n_17107 ^ n_16993;
assign n_17121 = n_17108 ^ n_17083;
assign n_17122 = n_17083 & n_17108;
assign n_17123 = n_17109 ^ x282;
assign n_17124 = n_17110 ^ n_16489;
assign n_17125 = n_17111 ^ n_16489;
assign n_17126 = n_17112 ^ n_15166;
assign n_17127 = n_17113 ^ x424;
assign n_17128 = n_17114 ^ n_17113;
assign n_17129 = n_17117 ^ n_14866;
assign n_17130 = n_17118 ^ x281;
assign n_17131 = n_17119 ^ n_14846;
assign n_17132 = n_16523 ^ n_17121;
assign n_17133 = n_17123 ^ n_17118;
assign n_17134 = n_17125 ^ n_17121;
assign n_17135 = n_17124 ^ n_17126;
assign n_17136 = n_17126 ^ n_15187;
assign n_17137 = n_17128 & ~n_17127;
assign n_17138 = n_17128 ^ x424;
assign n_17139 = n_17131 ^ x280;
assign n_17140 = n_17133 ^ x281;
assign n_17141 = ~n_17133 & n_17130;
assign n_17142 = n_16523 ^ n_17134;
assign n_17143 = ~n_17134 & n_17132;
assign n_17144 = n_17135 ^ n_15187;
assign n_17145 = ~n_17135 & n_17136;
assign n_17146 = n_17137 ^ x424;
assign n_17147 = n_17138 & n_17115;
assign n_17148 = n_17115 ^ n_17138;
assign n_17149 = n_17139 ^ n_17129;
assign n_17150 = n_17122 ^ n_17140;
assign n_17151 = ~n_17140 & ~n_17122;
assign n_17152 = n_17141 ^ x281;
assign n_17153 = n_17142 ^ n_16512;
assign n_17154 = n_17035 ^ n_17142;
assign n_17155 = n_17143 ^ n_16523;
assign n_17156 = n_17144 ^ x439;
assign n_17157 = n_17145 ^ n_15187;
assign n_17158 = n_17146 ^ n_17144;
assign n_17159 = n_17146 ^ x439;
assign n_17160 = n_17150 ^ n_16558;
assign n_17161 = n_17152 ^ n_17151;
assign n_17162 = n_15847 & n_17153;
assign n_17163 = n_17155 ^ n_17150;
assign n_17164 = n_17155 ^ n_16558;
assign n_17165 = n_17156 & ~n_17158;
assign n_17166 = n_17159 ^ n_17144;
assign n_17167 = n_17161 ^ n_17149;
assign n_17168 = n_17162 ^ n_16512;
assign n_17169 = ~n_15866 & ~n_17163;
assign n_17170 = n_17163 & ~n_17160;
assign n_17171 = n_17164 ^ n_17150;
assign n_17172 = n_17165 ^ x439;
assign n_17173 = n_17147 & ~n_17166;
assign n_17174 = n_17166 ^ n_17147;
assign n_17175 = n_16596 ^ n_17167;
assign n_17176 = n_17157 ^ n_17168;
assign n_17177 = n_17168 ^ n_15211;
assign n_17178 = n_17169 ^ n_16558;
assign n_17179 = n_17170 ^ n_16558;
assign n_17180 = n_17077 ^ n_17171;
assign n_17181 = n_17176 ^ n_15211;
assign n_17182 = ~n_17176 & ~n_17177;
assign n_17183 = n_17178 ^ n_15229;
assign n_17184 = n_17179 ^ n_16596;
assign n_17185 = n_17179 ^ n_17167;
assign n_17186 = n_17172 ^ n_17181;
assign n_17187 = n_17181 ^ x438;
assign n_17188 = n_17182 ^ n_15211;
assign n_17189 = n_17184 ^ n_17167;
assign n_17190 = n_17175 & ~n_17185;
assign n_17191 = n_17186 ^ x438;
assign n_17192 = n_17186 & ~n_17187;
assign n_17193 = n_17188 ^ n_15229;
assign n_17194 = n_17188 ^ n_17178;
assign n_17195 = n_17189 ^ n_16580;
assign n_17196 = n_17116 ^ n_17189;
assign n_17197 = n_17190 ^ n_16596;
assign n_17198 = n_17173 & n_17191;
assign n_17199 = n_17191 ^ n_17173;
assign n_17200 = n_17192 ^ x438;
assign n_17201 = n_17193 ^ n_17178;
assign n_17202 = ~n_17183 & n_17194;
assign n_17203 = ~n_15887 & ~n_17195;
assign n_17204 = n_17197 ^ n_16646;
assign n_17205 = n_17197 ^ n_16634;
assign n_17206 = n_17200 ^ n_17201;
assign n_17207 = n_17201 ^ x437;
assign n_17208 = n_17202 ^ n_15229;
assign n_17209 = n_17203 ^ n_16580;
assign n_17210 = n_17204 ^ n_16634;
assign n_17211 = n_17148 ^ n_17204;
assign n_17212 = n_16646 & ~n_17205;
assign n_17213 = n_17206 ^ x437;
assign n_17214 = ~n_17206 & n_17207;
assign n_17215 = n_17208 ^ n_15249;
assign n_17216 = n_17209 ^ n_15249;
assign n_17217 = n_17208 ^ n_17209;
assign n_17218 = n_15908 & n_17210;
assign n_17219 = n_17212 ^ n_15987;
assign n_17220 = n_17213 & ~n_17198;
assign n_17221 = n_17198 ^ n_17213;
assign n_17222 = n_17214 ^ x437;
assign n_17223 = n_17215 ^ n_17209;
assign n_17224 = ~n_17216 & ~n_17217;
assign n_17225 = n_17218 ^ n_16634;
assign n_17226 = n_17219 ^ n_16669;
assign n_17227 = n_17222 ^ n_17223;
assign n_17228 = n_17223 ^ x436;
assign n_17229 = n_17224 ^ n_15249;
assign n_17230 = n_16027 ^ n_17226;
assign n_17231 = n_17226 & n_16684;
assign n_17232 = n_17227 ^ x436;
assign n_17233 = ~n_17227 & n_17228;
assign n_17234 = n_17229 ^ n_15270;
assign n_17235 = n_17225 ^ n_17229;
assign n_17236 = n_17230 ^ n_16669;
assign n_17237 = n_17174 ^ n_17230;
assign n_17238 = n_17231 ^ n_16027;
assign n_17239 = n_17220 & n_17232;
assign n_17240 = n_17232 ^ n_17220;
assign n_17241 = n_17233 ^ x436;
assign n_17242 = n_17225 ^ n_17234;
assign n_17243 = n_17234 & ~n_17235;
assign n_17244 = n_15929 & ~n_17236;
assign n_17245 = n_17238 ^ n_16710;
assign n_17246 = n_17241 ^ n_17242;
assign n_17247 = n_17242 ^ x435;
assign n_17248 = n_17243 ^ n_15270;
assign n_17249 = n_17244 ^ n_16669;
assign n_17250 = n_16088 ^ n_17245;
assign n_17251 = n_17245 & ~n_16725;
assign n_17252 = n_17246 ^ x435;
assign n_17253 = ~n_17246 & n_17247;
assign n_17254 = n_17248 ^ n_15291;
assign n_17255 = n_17249 ^ n_15291;
assign n_17256 = n_17248 ^ n_17249;
assign n_17257 = n_17250 ^ n_16710;
assign n_17258 = n_17199 ^ n_17250;
assign n_17259 = n_17251 ^ n_16088;
assign n_17260 = n_17239 & n_17252;
assign n_17261 = n_17252 ^ n_17239;
assign n_17262 = n_17253 ^ x435;
assign n_17263 = n_17254 ^ n_17249;
assign n_17264 = n_17255 & n_17256;
assign n_17265 = ~n_15955 & n_17257;
assign n_17266 = n_17259 ^ n_16748;
assign n_17267 = n_17262 ^ x434;
assign n_17268 = n_17262 ^ n_17263;
assign n_17269 = n_17264 ^ n_15291;
assign n_17270 = n_17265 ^ n_16710;
assign n_17271 = n_16135 ^ n_17266;
assign n_17272 = n_17266 & n_16763;
assign n_17273 = ~n_17268 & n_17267;
assign n_17274 = n_17268 ^ x434;
assign n_17275 = n_17269 ^ n_15312;
assign n_17276 = n_17270 ^ n_15312;
assign n_17277 = n_17269 ^ n_17270;
assign n_17278 = n_17271 ^ n_16748;
assign n_17279 = n_17221 ^ n_17271;
assign n_17280 = n_17272 ^ n_16135;
assign n_17281 = n_17273 ^ x434;
assign n_17282 = ~n_17260 & ~n_17274;
assign n_17283 = n_17274 ^ n_17260;
assign n_17284 = n_17275 ^ n_17270;
assign n_17285 = n_17276 & n_17277;
assign n_17286 = ~n_15988 & ~n_17278;
assign n_17287 = n_17280 ^ n_16807;
assign n_17288 = n_17280 ^ n_16792;
assign n_17289 = n_17281 ^ n_17284;
assign n_17290 = n_17284 ^ x433;
assign n_17291 = n_17285 ^ n_15312;
assign n_17292 = n_17286 ^ n_16748;
assign n_17293 = n_17287 ^ n_16792;
assign n_17294 = n_17240 ^ n_17287;
assign n_17295 = ~n_16807 & ~n_17288;
assign n_17296 = n_17289 ^ x433;
assign n_17297 = n_17289 & ~n_17290;
assign n_17298 = n_17291 ^ n_15333;
assign n_17299 = n_17292 ^ n_15333;
assign n_17300 = n_17291 ^ n_17292;
assign n_17301 = ~n_16030 & ~n_17293;
assign n_17302 = n_17295 ^ n_16178;
assign n_17303 = n_17282 & n_17296;
assign n_17304 = n_17296 ^ n_17282;
assign n_17305 = n_17297 ^ x433;
assign n_17306 = n_17298 ^ n_17292;
assign n_17307 = n_17299 & ~n_17300;
assign n_17308 = n_17301 ^ n_16792;
assign n_17309 = n_17302 ^ n_16220;
assign n_17310 = n_17302 ^ n_16836;
assign n_17311 = n_17305 ^ n_17306;
assign n_17312 = n_17306 ^ x432;
assign n_17313 = n_17307 ^ n_15333;
assign n_17314 = n_17308 ^ n_15354;
assign n_17315 = n_17309 ^ n_16836;
assign n_17316 = n_16851 & n_17310;
assign n_17317 = n_17311 ^ x432;
assign n_17318 = ~n_17311 & n_17312;
assign n_17319 = n_17313 ^ n_17308;
assign n_17320 = n_17315 ^ n_16822;
assign n_17321 = n_17261 ^ n_17315;
assign n_17322 = n_17316 ^ n_16220;
assign n_17323 = n_17303 & ~n_17317;
assign n_17324 = n_17317 ^ n_17303;
assign n_17325 = n_17318 ^ x432;
assign n_17326 = n_17319 ^ n_15354;
assign n_17327 = ~n_17319 & ~n_17314;
assign n_17328 = n_16068 & ~n_17320;
assign n_17329 = n_17322 ^ n_16878;
assign n_17330 = n_17325 ^ x447;
assign n_17331 = n_17326 ^ x447;
assign n_17332 = n_17325 ^ n_17326;
assign n_17333 = n_17327 ^ n_15354;
assign n_17334 = n_17328 ^ n_16822;
assign n_17335 = n_16262 ^ n_17329;
assign n_17336 = ~n_17329 & ~n_16894;
assign n_17337 = n_17330 ^ n_17326;
assign n_17338 = ~n_17331 & n_17332;
assign n_17339 = n_17333 ^ n_15376;
assign n_17340 = n_17334 ^ n_15376;
assign n_17341 = n_17333 ^ n_17334;
assign n_17342 = n_17335 ^ n_16878;
assign n_17343 = n_17283 ^ n_17335;
assign n_17344 = n_17336 ^ n_16262;
assign n_17345 = n_17337 & n_17323;
assign n_17346 = n_17323 ^ n_17337;
assign n_17347 = n_17338 ^ x447;
assign n_17348 = n_17339 ^ n_17334;
assign n_17349 = ~n_17340 & n_17341;
assign n_17350 = ~n_16108 & ~n_17342;
assign n_17351 = n_17344 ^ n_16922;
assign n_17352 = n_17347 ^ n_17348;
assign n_17353 = n_17348 ^ x446;
assign n_17354 = n_17349 ^ n_15376;
assign n_17355 = n_17350 ^ n_16878;
assign n_17356 = n_16304 ^ n_17351;
assign n_17357 = ~n_17351 & ~n_16937;
assign n_17358 = n_17352 ^ x446;
assign n_17359 = ~n_17352 & n_17353;
assign n_17360 = n_17354 ^ n_15396;
assign n_17361 = n_17355 ^ n_15396;
assign n_17362 = n_17354 ^ n_17355;
assign n_17363 = n_17356 ^ n_16922;
assign n_17364 = n_17304 ^ n_17356;
assign n_17365 = n_17357 ^ n_16304;
assign n_17366 = ~n_17345 & n_17358;
assign n_17367 = n_17358 ^ n_17345;
assign n_17368 = n_17359 ^ x446;
assign n_17369 = n_17360 ^ n_17355;
assign n_17370 = n_17361 & n_17362;
assign n_17371 = ~n_16150 & ~n_17363;
assign n_17372 = n_17365 ^ n_16965;
assign n_17373 = n_17368 ^ n_17369;
assign n_17374 = n_17369 ^ x445;
assign n_17375 = n_17370 ^ n_15396;
assign n_17376 = n_17371 ^ n_16922;
assign n_17377 = n_16343 ^ n_17372;
assign n_17378 = n_17372 & n_16980;
assign n_17379 = n_17373 ^ x445;
assign n_17380 = n_17373 & ~n_17374;
assign n_17381 = n_17375 ^ n_15422;
assign n_17382 = n_17376 ^ n_15422;
assign n_17383 = n_17375 ^ n_17376;
assign n_17384 = n_17377 ^ n_16965;
assign n_17385 = n_17324 ^ n_17377;
assign n_17386 = n_17378 ^ n_16343;
assign n_17387 = n_17366 & ~n_17379;
assign n_17388 = n_17379 ^ n_17366;
assign n_17389 = n_17380 ^ x445;
assign n_17390 = n_17381 ^ n_17376;
assign n_17391 = ~n_17382 & n_17383;
assign n_17392 = ~n_16192 & ~n_17384;
assign n_17393 = n_17386 ^ n_16379;
assign n_17394 = n_17386 ^ n_17008;
assign n_17395 = n_17389 ^ n_17390;
assign n_17396 = n_17390 ^ x444;
assign n_17397 = n_17391 ^ n_15422;
assign n_17398 = n_17392 ^ n_16965;
assign n_17399 = ~n_16234 & n_17393;
assign n_17400 = n_17393 ^ n_17008;
assign n_17401 = ~n_17023 & n_17394;
assign n_17402 = n_17395 ^ x444;
assign n_17403 = n_17395 & ~n_17396;
assign n_17404 = n_17397 ^ n_15455;
assign n_17405 = n_17398 ^ n_15455;
assign n_17406 = n_17397 ^ n_17398;
assign n_17407 = n_17399 ^ n_17008;
assign n_17408 = n_17400 ^ n_17346;
assign n_17409 = n_17401 ^ n_16379;
assign n_17410 = n_17387 ^ n_17402;
assign n_17411 = n_17402 & ~n_17387;
assign n_17412 = n_17403 ^ x444;
assign n_17413 = n_17404 ^ n_17398;
assign n_17414 = ~n_17405 & n_17406;
assign n_17415 = n_17407 ^ n_15494;
assign n_17416 = n_17409 ^ n_17051;
assign n_17417 = n_17410 ^ n_16454;
assign n_17418 = ~n_16454 & n_17410;
assign n_17419 = n_17412 ^ n_17413;
assign n_17420 = n_17413 ^ x443;
assign n_17421 = n_17414 ^ n_15455;
assign n_17422 = n_17416 ^ n_16406;
assign n_17423 = ~n_17416 & n_17064;
assign n_17424 = n_17417 ^ n_16447;
assign n_17425 = n_16476 ^ n_17418;
assign n_17426 = n_17419 ^ x443;
assign n_17427 = n_17419 & ~n_17420;
assign n_17428 = n_17421 ^ n_15494;
assign n_17429 = n_17421 ^ n_17407;
assign n_17430 = n_17422 ^ n_17051;
assign n_17431 = n_17367 ^ n_17422;
assign n_17432 = n_17423 ^ n_16406;
assign n_17433 = n_15935 & n_17424;
assign n_17434 = n_17411 ^ n_17426;
assign n_17435 = ~n_17426 & ~n_17411;
assign n_17436 = n_17427 ^ x443;
assign n_17437 = n_17428 ^ n_17407;
assign n_17438 = ~n_17415 & ~n_17429;
assign n_17439 = n_16276 & n_17430;
assign n_17440 = n_17432 ^ n_16427;
assign n_17441 = n_17433 ^ n_16447;
assign n_17442 = n_17434 ^ n_17418;
assign n_17443 = n_17425 ^ n_17434;
assign n_17444 = n_17436 ^ n_17437;
assign n_17445 = n_17437 ^ x442;
assign n_17446 = n_17438 ^ n_15494;
assign n_17447 = n_17439 ^ n_17051;
assign n_17448 = n_16318 & ~n_17440;
assign n_17449 = n_17440 ^ n_17079;
assign n_17450 = n_17441 ^ n_15401;
assign n_17451 = ~n_15401 & ~n_17441;
assign n_17452 = n_15962 & n_17442;
assign n_17453 = ~n_17442 & n_17425;
assign n_17454 = n_17444 ^ x442;
assign n_17455 = n_17444 & ~n_17445;
assign n_17456 = n_17446 ^ n_15532;
assign n_17457 = n_17447 ^ n_15532;
assign n_17458 = n_17447 ^ n_17446;
assign n_17459 = n_17448 ^ n_17079;
assign n_17460 = x71 & n_17450;
assign n_17461 = n_17450 ^ x71;
assign n_17462 = n_17451 ^ n_15428;
assign n_17463 = n_17452 ^ n_16476;
assign n_17464 = n_17453 ^ n_16476;
assign n_17465 = n_17454 ^ n_17435;
assign n_17466 = ~n_17435 & n_17454;
assign n_17467 = n_17455 ^ x442;
assign n_17468 = n_17447 ^ n_17456;
assign n_17469 = n_17457 & ~n_17458;
assign n_17470 = n_17459 ^ n_15574;
assign n_17471 = n_17460 ^ x70;
assign n_17472 = n_17463 ^ n_17462;
assign n_17473 = n_17463 ^ n_17451;
assign n_17474 = n_16518 ^ n_17464;
assign n_17475 = n_17464 ^ n_17465;
assign n_17476 = n_16518 ^ n_17465;
assign n_17477 = n_17467 ^ n_17468;
assign n_17478 = n_17468 ^ x441;
assign n_17479 = n_17469 ^ n_15532;
assign n_17480 = n_17472 ^ n_17460;
assign n_17481 = n_17472 ^ n_17471;
assign n_17482 = ~n_17462 & ~n_17473;
assign n_17483 = n_17474 ^ n_17465;
assign n_17484 = ~n_16011 & n_17475;
assign n_17485 = ~n_17475 & ~n_17476;
assign n_17486 = n_17477 ^ x441;
assign n_17487 = n_17477 & ~n_17478;
assign n_17488 = n_17479 ^ x440;
assign n_17489 = n_17471 & n_17480;
assign n_17490 = n_17482 ^ n_15428;
assign n_17491 = n_17484 ^ n_16518;
assign n_17492 = n_17485 ^ n_16518;
assign n_17493 = n_17486 ^ n_17466;
assign n_17494 = ~n_17466 & ~n_17486;
assign n_17495 = n_17487 ^ x441;
assign n_17496 = n_17488 ^ n_17470;
assign n_17497 = n_17489 ^ x70;
assign n_17498 = n_17490 ^ n_15472;
assign n_17499 = n_17491 ^ n_15472;
assign n_17500 = n_17490 ^ n_17491;
assign n_17501 = n_16553 ^ n_17492;
assign n_17502 = n_17492 ^ n_17493;
assign n_17503 = n_16553 ^ n_17493;
assign n_17504 = n_17495 ^ n_17496;
assign n_17505 = n_17498 ^ n_17491;
assign n_17506 = ~n_17499 & ~n_17500;
assign n_17507 = n_17501 ^ n_17493;
assign n_17508 = ~n_16053 & ~n_17502;
assign n_17509 = n_17502 & n_17503;
assign n_17510 = n_17504 ^ n_17494;
assign n_17511 = n_17497 ^ n_17505;
assign n_17512 = n_17505 ^ x69;
assign n_17513 = n_17506 ^ n_15472;
assign n_17514 = n_17508 ^ n_16553;
assign n_17515 = n_17509 ^ n_16553;
assign n_17516 = n_16603 ^ n_17510;
assign n_17517 = n_17511 ^ x69;
assign n_17518 = ~n_17511 & n_17512;
assign n_17519 = n_17513 ^ n_15514;
assign n_17520 = n_17514 ^ n_15514;
assign n_17521 = n_17513 ^ n_17514;
assign n_17522 = n_17515 ^ n_17510;
assign n_17523 = n_16603 ^ n_17515;
assign n_17524 = n_17518 ^ x69;
assign n_17525 = n_17519 ^ n_17514;
assign n_17526 = n_17520 & ~n_17521;
assign n_17527 = n_16092 & ~n_17522;
assign n_17528 = n_17522 & n_17516;
assign n_17529 = n_17523 ^ n_17510;
assign n_17530 = n_17524 ^ n_17525;
assign n_17531 = n_17525 ^ x68;
assign n_17532 = n_17526 ^ n_15514;
assign n_17533 = n_17527 ^ n_16603;
assign n_17534 = n_17528 ^ n_16603;
assign n_17535 = n_17530 ^ x68;
assign n_17536 = ~n_17530 & n_17531;
assign n_17537 = n_17532 ^ n_15556;
assign n_17538 = n_17533 ^ n_15556;
assign n_17539 = n_17532 ^ n_17533;
assign n_17540 = n_17534 ^ n_16653;
assign n_17541 = n_17534 ^ n_16640;
assign n_17542 = n_17536 ^ x68;
assign n_17543 = n_17537 ^ n_17533;
assign n_17544 = n_17538 & n_17539;
assign n_17545 = n_17540 ^ n_16640;
assign n_17546 = ~n_16653 & ~n_17541;
assign n_17547 = n_17542 ^ n_17543;
assign n_17548 = n_17543 ^ x67;
assign n_17549 = n_17544 ^ n_15556;
assign n_17550 = n_16131 & ~n_17545;
assign n_17551 = n_17546 ^ n_16487;
assign n_17552 = n_17547 ^ x67;
assign n_17553 = ~n_17547 & n_17548;
assign n_17554 = n_17549 ^ n_15594;
assign n_17555 = n_17550 ^ n_16640;
assign n_17556 = n_16692 ^ n_17551;
assign n_17557 = ~n_17535 & ~n_17552;
assign n_17558 = n_17552 ^ n_17535;
assign n_17559 = n_17553 ^ x67;
assign n_17560 = n_17554 ^ n_17555;
assign n_17561 = n_17555 ^ n_15594;
assign n_17562 = n_17549 ^ n_17555;
assign n_17563 = n_16546 ^ n_17556;
assign n_17564 = ~n_17556 & ~n_16705;
assign n_17565 = n_17559 ^ n_17560;
assign n_17566 = n_17560 ^ x66;
assign n_17567 = n_17561 & ~n_17562;
assign n_17568 = n_17563 ^ n_16692;
assign n_17569 = n_17564 ^ n_16546;
assign n_17570 = n_17565 ^ x66;
assign n_17571 = n_17565 & ~n_17566;
assign n_17572 = n_17567 ^ n_15594;
assign n_17573 = ~n_16173 & ~n_17568;
assign n_17574 = n_16732 ^ n_17569;
assign n_17575 = n_17557 & n_17570;
assign n_17576 = n_17570 ^ n_17557;
assign n_17577 = n_17571 ^ x66;
assign n_17578 = n_17572 ^ n_15628;
assign n_17579 = n_17573 ^ n_16692;
assign n_17580 = ~n_17574 & ~n_16745;
assign n_17581 = n_16593 ^ n_17574;
assign n_17582 = n_17578 ^ n_17579;
assign n_17583 = n_17579 ^ n_15628;
assign n_17584 = n_17572 ^ n_17579;
assign n_17585 = n_17580 ^ n_16593;
assign n_17586 = n_17581 ^ n_16732;
assign n_17587 = n_17577 ^ n_17582;
assign n_17588 = n_17582 ^ x65;
assign n_17589 = ~n_17583 & n_17584;
assign n_17590 = n_16772 ^ n_17585;
assign n_17591 = n_16215 & ~n_17586;
assign n_17592 = n_17587 ^ x65;
assign n_17593 = ~n_17587 & n_17588;
assign n_17594 = n_17589 ^ n_15628;
assign n_17595 = ~n_17590 & n_16787;
assign n_17596 = n_16631 ^ n_17590;
assign n_17597 = n_17591 ^ n_16732;
assign n_17598 = n_17592 ^ n_17575;
assign n_17599 = n_17575 & ~n_17592;
assign n_17600 = n_17593 ^ x65;
assign n_17601 = n_17594 ^ n_15656;
assign n_17602 = n_17595 ^ n_16631;
assign n_17603 = n_17596 ^ n_16772;
assign n_17604 = n_17597 ^ n_15656;
assign n_17605 = n_17594 ^ n_17597;
assign n_17606 = n_17601 ^ n_17597;
assign n_17607 = n_16815 ^ n_17602;
assign n_17608 = ~n_16257 & n_17603;
assign n_17609 = ~n_17604 & ~n_17605;
assign n_17610 = n_17600 ^ n_17606;
assign n_17611 = n_17606 ^ x64;
assign n_17612 = ~n_17607 & ~n_16831;
assign n_17613 = n_16681 ^ n_17607;
assign n_17614 = n_17608 ^ n_16772;
assign n_17615 = n_17609 ^ n_15656;
assign n_17616 = n_17610 ^ x64;
assign n_17617 = ~n_17610 & n_17611;
assign n_17618 = n_17612 ^ n_16681;
assign n_17619 = n_17613 ^ n_16815;
assign n_17620 = n_17461 ^ n_17613;
assign n_17621 = n_17614 ^ n_15680;
assign n_17622 = n_17615 ^ n_17614;
assign n_17623 = n_17615 ^ n_15680;
assign n_17624 = n_17599 & ~n_17616;
assign n_17625 = n_17616 ^ n_17599;
assign n_17626 = n_17617 ^ x64;
assign n_17627 = n_17618 ^ n_16858;
assign n_17628 = n_17618 ^ n_16722;
assign n_17629 = ~n_16299 & ~n_17619;
assign n_17630 = n_17621 & ~n_17622;
assign n_17631 = n_17623 ^ n_17614;
assign n_17632 = ~n_16873 & ~n_17627;
assign n_17633 = n_17628 ^ n_16858;
assign n_17634 = ~n_16338 & ~n_17628;
assign n_17635 = n_17629 ^ n_16815;
assign n_17636 = n_17630 ^ n_15680;
assign n_17637 = n_17626 ^ n_17631;
assign n_17638 = n_17631 ^ x79;
assign n_17639 = n_17632 ^ n_16722;
assign n_17640 = n_17481 ^ n_17633;
assign n_17641 = n_17634 ^ n_16858;
assign n_17642 = n_17635 ^ n_15697;
assign n_17643 = n_17636 ^ n_17635;
assign n_17644 = n_17636 ^ n_15697;
assign n_17645 = n_17637 ^ x79;
assign n_17646 = ~n_17637 & n_17638;
assign n_17647 = n_16902 ^ n_17639;
assign n_17648 = n_17641 ^ n_15713;
assign n_17649 = n_17642 & ~n_17643;
assign n_17650 = n_17644 ^ n_17635;
assign n_17651 = n_17624 & ~n_17645;
assign n_17652 = n_17645 ^ n_17624;
assign n_17653 = n_17646 ^ x79;
assign n_17654 = n_17647 & ~n_16917;
assign n_17655 = n_16775 ^ n_17647;
assign n_17656 = n_17649 ^ n_15697;
assign n_17657 = n_17650 ^ x78;
assign n_17658 = n_17653 ^ n_17650;
assign n_17659 = n_17654 ^ n_16775;
assign n_17660 = n_17655 ^ n_16902;
assign n_17661 = n_17517 ^ n_17655;
assign n_17662 = n_17656 ^ n_17641;
assign n_17663 = n_17656 ^ n_15713;
assign n_17664 = ~n_17658 & n_17657;
assign n_17665 = n_17658 ^ x78;
assign n_17666 = n_17659 ^ n_16820;
assign n_17667 = n_17659 ^ n_16945;
assign n_17668 = ~n_16374 & n_17660;
assign n_17669 = ~n_17648 & n_17662;
assign n_17670 = n_17663 ^ n_17641;
assign n_17671 = n_17664 ^ x78;
assign n_17672 = n_17651 & ~n_17665;
assign n_17673 = n_17665 ^ n_17651;
assign n_17674 = n_17666 ^ n_16945;
assign n_17675 = n_16401 & ~n_17666;
assign n_17676 = n_16960 & n_17667;
assign n_17677 = n_17668 ^ n_16902;
assign n_17678 = n_17669 ^ n_15713;
assign n_17679 = n_17670 ^ x77;
assign n_17680 = n_17671 ^ n_17670;
assign n_17681 = n_17674 ^ n_17535;
assign n_17682 = n_17675 ^ n_16945;
assign n_17683 = n_17676 ^ n_16820;
assign n_17684 = n_17677 ^ n_15726;
assign n_17685 = n_17678 ^ n_17677;
assign n_17686 = n_17678 ^ n_15726;
assign n_17687 = n_17680 & ~n_17679;
assign n_17688 = n_17680 ^ x77;
assign n_17689 = n_17682 ^ n_15743;
assign n_17690 = n_16988 ^ n_17683;
assign n_17691 = n_17684 & n_17685;
assign n_17692 = n_17686 ^ n_17677;
assign n_17693 = n_17687 ^ x77;
assign n_17694 = ~n_17672 & ~n_17688;
assign n_17695 = n_17688 ^ n_17672;
assign n_17696 = n_17690 & ~n_17003;
assign n_17697 = n_16863 ^ n_17690;
assign n_17698 = n_17691 ^ n_15726;
assign n_17699 = n_17692 ^ x76;
assign n_17700 = n_17693 ^ n_17692;
assign n_17701 = n_17696 ^ n_16863;
assign n_17702 = n_17697 ^ n_16988;
assign n_17703 = n_17558 ^ n_17697;
assign n_17704 = n_17698 ^ n_17682;
assign n_17705 = n_17698 ^ n_15743;
assign n_17706 = ~n_17700 & n_17699;
assign n_17707 = n_17700 ^ x76;
assign n_17708 = n_17030 ^ n_17701;
assign n_17709 = ~n_16422 & n_17702;
assign n_17710 = n_17689 & ~n_17704;
assign n_17711 = n_17705 ^ n_17682;
assign n_17712 = n_17706 ^ x76;
assign n_17713 = n_17707 & n_17694;
assign n_17714 = n_17694 ^ n_17707;
assign n_17715 = ~n_17708 & ~n_17045;
assign n_17716 = n_16907 ^ n_17708;
assign n_17717 = n_17709 ^ n_16988;
assign n_17718 = n_17710 ^ n_15743;
assign n_17719 = n_17711 ^ x75;
assign n_17720 = n_17712 ^ n_17711;
assign n_17721 = n_17715 ^ n_16907;
assign n_17722 = n_17716 ^ n_17030;
assign n_17723 = n_17576 ^ n_17716;
assign n_17724 = n_17717 ^ n_15763;
assign n_17725 = n_17718 ^ n_17717;
assign n_17726 = n_17718 ^ n_15763;
assign n_17727 = n_17720 & ~n_17719;
assign n_17728 = n_17720 ^ x75;
assign n_17729 = n_17070 ^ n_17721;
assign n_17730 = ~n_16435 & ~n_17722;
assign n_17731 = ~n_17724 & n_17725;
assign n_17732 = n_17726 ^ n_17717;
assign n_17733 = n_17727 ^ x75;
assign n_17734 = n_17713 & ~n_17728;
assign n_17735 = n_17728 ^ n_17713;
assign n_17736 = ~n_17729 & ~n_17085;
assign n_17737 = n_16950 ^ n_17729;
assign n_17738 = n_17730 ^ n_17030;
assign n_17739 = n_17731 ^ n_15763;
assign n_17740 = n_17732 ^ x74;
assign n_17741 = n_17733 ^ n_17732;
assign n_17742 = n_17736 ^ n_16950;
assign n_17743 = n_17737 ^ n_17070;
assign n_17744 = n_17598 ^ n_17737;
assign n_17745 = n_17738 ^ n_15783;
assign n_17746 = n_17739 ^ n_17738;
assign n_17747 = n_17739 ^ n_15783;
assign n_17748 = ~n_17741 & n_17740;
assign n_17749 = n_17741 ^ x74;
assign n_17750 = n_17742 ^ n_17107;
assign n_17751 = n_17742 ^ n_17120;
assign n_17752 = n_16463 & ~n_17743;
assign n_17753 = ~n_17745 & ~n_17746;
assign n_17754 = n_17747 ^ n_17738;
assign n_17755 = n_17748 ^ x74;
assign n_17756 = ~n_17749 & ~n_17734;
assign n_17757 = n_17734 ^ n_17749;
assign n_17758 = n_17120 & n_17750;
assign n_17759 = n_17751 ^ n_17107;
assign n_17760 = n_17625 ^ n_17751;
assign n_17761 = n_17752 ^ n_17070;
assign n_17762 = n_17753 ^ n_15783;
assign n_17763 = n_17754 ^ x73;
assign n_17764 = n_17755 ^ n_17754;
assign n_17765 = n_17758 ^ n_16993;
assign n_17766 = n_16489 & ~n_17759;
assign n_17767 = n_17761 ^ n_15804;
assign n_17768 = n_17762 ^ n_17761;
assign n_17769 = n_17762 ^ n_15804;
assign n_17770 = ~n_17764 & n_17763;
assign n_17771 = n_17764 ^ x73;
assign n_17772 = n_17765 ^ n_17142;
assign n_17773 = n_17035 ^ n_17765;
assign n_17774 = n_17766 ^ n_17107;
assign n_17775 = n_17767 & ~n_17768;
assign n_17776 = n_17769 ^ n_17761;
assign n_17777 = n_17770 ^ x73;
assign n_17778 = ~n_17756 & n_17771;
assign n_17779 = n_17771 ^ n_17756;
assign n_17780 = n_17154 & ~n_17772;
assign n_17781 = n_17773 ^ n_17142;
assign n_17782 = n_17774 ^ n_15824;
assign n_17783 = n_17775 ^ n_15804;
assign n_17784 = n_17776 ^ x72;
assign n_17785 = n_17777 ^ n_17776;
assign n_17786 = n_17780 ^ n_17035;
assign n_17787 = n_17781 ^ n_17134;
assign n_17788 = n_17781 ^ n_17652;
assign n_17789 = n_17783 ^ n_17774;
assign n_17790 = n_17783 ^ n_17782;
assign n_17791 = ~n_17785 & n_17784;
assign n_17792 = n_17785 ^ x72;
assign n_17793 = n_17171 ^ n_17786;
assign n_17794 = n_16523 & n_17787;
assign n_17795 = ~n_17782 & ~n_17789;
assign n_17796 = n_17791 ^ x72;
assign n_17797 = ~n_17778 & ~n_17792;
assign n_17798 = n_17792 ^ n_17778;
assign n_17799 = n_17793 & n_17180;
assign n_17800 = n_17077 ^ n_17793;
assign n_17801 = n_17794 ^ n_17134;
assign n_17802 = n_17795 ^ n_15824;
assign n_17803 = n_17796 ^ x87;
assign n_17804 = n_17790 ^ n_17796;
assign n_17805 = n_17799 ^ n_17077;
assign n_17806 = n_17800 ^ n_17171;
assign n_17807 = n_17673 ^ n_17800;
assign n_17808 = n_17801 ^ n_15847;
assign n_17809 = n_17802 ^ n_17801;
assign n_17810 = n_17790 ^ n_17803;
assign n_17811 = n_17803 & n_17804;
assign n_17812 = n_17805 ^ n_17189;
assign n_17813 = n_16558 & ~n_17806;
assign n_17814 = n_17809 & n_17808;
assign n_17815 = n_17809 ^ n_15847;
assign n_17816 = n_17810 & n_17797;
assign n_17817 = n_17797 ^ n_17810;
assign n_17818 = n_17811 ^ x87;
assign n_17819 = n_17812 & n_17196;
assign n_17820 = n_17116 ^ n_17812;
assign n_17821 = n_17813 ^ n_17171;
assign n_17822 = n_17814 ^ n_15847;
assign n_17823 = n_17815 ^ x86;
assign n_17824 = n_17818 ^ n_17815;
assign n_17825 = n_17819 ^ n_17116;
assign n_17826 = n_17820 ^ n_17189;
assign n_17827 = n_17695 ^ n_17820;
assign n_17828 = n_17821 ^ n_15866;
assign n_17829 = n_17822 ^ n_17821;
assign n_17830 = n_17822 ^ n_15866;
assign n_17831 = n_17824 & ~n_17823;
assign n_17832 = n_17824 ^ x86;
assign n_17833 = n_17825 ^ n_17204;
assign n_17834 = n_16596 & ~n_17826;
assign n_17835 = n_17828 & n_17829;
assign n_17836 = n_17830 ^ n_17821;
assign n_17837 = n_17831 ^ x86;
assign n_17838 = n_17816 & n_17832;
assign n_17839 = n_17832 ^ n_17816;
assign n_17840 = ~n_17833 & ~n_17211;
assign n_17841 = n_17148 ^ n_17833;
assign n_17842 = n_17834 ^ n_17189;
assign n_17843 = n_17835 ^ n_15866;
assign n_17844 = n_17836 ^ x85;
assign n_17845 = n_17837 ^ n_17836;
assign n_17846 = n_17840 ^ n_17148;
assign n_17847 = n_17841 ^ n_17204;
assign n_17848 = n_17714 ^ n_17841;
assign n_17849 = n_17842 ^ n_15887;
assign n_17850 = n_17843 ^ n_17842;
assign n_17851 = n_17843 ^ n_15887;
assign n_17852 = ~n_17845 & n_17844;
assign n_17853 = n_17845 ^ x85;
assign n_17854 = n_17846 ^ n_17230;
assign n_17855 = n_16634 & ~n_17847;
assign n_17856 = ~n_17849 & n_17850;
assign n_17857 = n_17851 ^ n_17842;
assign n_17858 = n_17852 ^ x85;
assign n_17859 = n_17838 & ~n_17853;
assign n_17860 = n_17853 ^ n_17838;
assign n_17861 = n_17854 & n_17237;
assign n_17862 = n_17174 ^ n_17854;
assign n_17863 = n_17855 ^ n_17204;
assign n_17864 = n_17856 ^ n_15887;
assign n_17865 = n_17857 ^ x84;
assign n_17866 = n_17858 ^ n_17857;
assign n_17867 = n_17861 ^ n_17174;
assign n_17868 = n_17862 ^ n_17230;
assign n_17869 = n_17735 ^ n_17862;
assign n_17870 = n_17863 ^ n_15908;
assign n_17871 = n_17864 ^ n_17863;
assign n_17872 = n_17864 ^ n_15908;
assign n_17873 = ~n_17866 & n_17865;
assign n_17874 = n_17866 ^ x84;
assign n_17875 = n_17867 ^ n_17250;
assign n_17876 = ~n_16669 & ~n_17868;
assign n_17877 = n_17870 & n_17871;
assign n_17878 = n_17872 ^ n_17863;
assign n_17879 = n_17873 ^ x84;
assign n_17880 = n_17859 & ~n_17874;
assign n_17881 = n_17874 ^ n_17859;
assign n_17882 = ~n_17875 & ~n_17258;
assign n_17883 = n_17199 ^ n_17875;
assign n_17884 = n_17876 ^ n_17230;
assign n_17885 = n_17877 ^ n_15908;
assign n_17886 = n_17878 ^ x83;
assign n_17887 = n_17879 ^ n_17878;
assign n_17888 = n_17882 ^ n_17199;
assign n_17889 = n_17883 ^ n_17250;
assign n_17890 = n_17883 ^ n_17757;
assign n_17891 = n_17884 ^ n_15929;
assign n_17892 = n_17885 ^ n_17884;
assign n_17893 = n_17885 ^ n_15929;
assign n_17894 = n_17887 & ~n_17886;
assign n_17895 = n_17887 ^ x83;
assign n_17896 = n_17888 ^ n_17271;
assign n_17897 = n_16710 & ~n_17889;
assign n_17898 = n_17891 & ~n_17892;
assign n_17899 = n_17893 ^ n_17884;
assign n_17900 = n_17894 ^ x83;
assign n_17901 = ~n_17880 & ~n_17895;
assign n_17902 = n_17895 ^ n_17880;
assign n_17903 = ~n_17896 & n_17279;
assign n_17904 = n_17221 ^ n_17896;
assign n_17905 = n_17897 ^ n_17250;
assign n_17906 = n_17898 ^ n_15929;
assign n_17907 = n_17899 ^ x82;
assign n_17908 = n_17900 ^ n_17899;
assign n_17909 = n_17903 ^ n_17221;
assign n_17910 = n_17904 ^ n_17271;
assign n_17911 = n_17779 ^ n_17904;
assign n_17912 = n_17905 ^ n_15955;
assign n_17913 = n_17906 ^ n_17905;
assign n_17914 = n_17906 ^ n_15955;
assign n_17915 = ~n_17908 & n_17907;
assign n_17916 = n_17908 ^ x82;
assign n_17917 = n_17909 ^ n_17240;
assign n_17918 = n_17909 ^ n_17287;
assign n_17919 = n_16748 & n_17910;
assign n_17920 = ~n_17912 & ~n_17913;
assign n_17921 = n_17914 ^ n_17905;
assign n_17922 = n_17915 ^ x82;
assign n_17923 = ~n_17901 & ~n_17916;
assign n_17924 = n_17916 ^ n_17901;
assign n_17925 = n_16792 & ~n_17917;
assign n_17926 = n_17917 ^ n_17287;
assign n_17927 = ~n_17294 & ~n_17918;
assign n_17928 = n_17919 ^ n_17271;
assign n_17929 = n_17920 ^ n_15955;
assign n_17930 = n_17921 ^ x81;
assign n_17931 = n_17922 ^ n_17921;
assign n_17932 = n_17925 ^ n_17287;
assign n_17933 = n_17798 ^ n_17926;
assign n_17934 = n_17927 ^ n_17240;
assign n_17935 = n_17928 ^ n_15988;
assign n_17936 = n_17929 ^ n_17928;
assign n_17937 = n_17929 ^ n_15988;
assign n_17938 = n_17931 & ~n_17930;
assign n_17939 = n_17931 ^ x81;
assign n_17940 = n_17932 ^ n_16030;
assign n_17941 = n_17934 ^ n_17315;
assign n_17942 = n_17935 & ~n_17936;
assign n_17943 = n_17937 ^ n_17928;
assign n_17944 = n_17938 ^ x81;
assign n_17945 = n_17923 & n_17939;
assign n_17946 = n_17261 ^ n_17941;
assign n_17947 = n_17941 & ~n_17321;
assign n_17948 = n_17942 ^ n_15988;
assign n_17949 = n_17943 ^ x80;
assign n_17950 = n_17944 ^ n_17943;
assign n_17951 = n_17946 ^ n_17309;
assign n_17952 = n_17817 ^ n_17946;
assign n_17953 = n_17947 ^ n_17261;
assign n_17954 = n_17932 ^ n_17948;
assign n_17955 = n_17950 & ~n_17949;
assign n_17956 = n_17950 ^ x80;
assign n_17957 = n_16836 & n_17951;
assign n_17958 = n_17953 ^ n_17335;
assign n_17959 = n_17954 ^ n_16030;
assign n_17960 = ~n_17954 & n_17940;
assign n_17961 = n_17955 ^ x80;
assign n_17962 = n_17956 & n_17945;
assign n_17963 = n_17945 ^ n_17956;
assign n_17964 = n_17957 ^ n_17309;
assign n_17965 = n_17283 ^ n_17958;
assign n_17966 = n_17958 & n_17343;
assign n_17967 = n_17959 ^ x95;
assign n_17968 = n_17960 ^ n_16030;
assign n_17969 = n_17961 ^ n_17959;
assign n_17970 = n_17961 ^ x95;
assign n_17971 = ~n_17417 & ~n_17963;
assign n_17972 = n_17963 ^ n_17417;
assign n_17973 = n_17964 ^ n_16068;
assign n_17974 = n_17965 ^ n_17335;
assign n_17975 = n_17839 ^ n_17965;
assign n_17976 = n_17966 ^ n_17283;
assign n_17977 = n_17968 ^ n_17964;
assign n_17978 = ~n_17967 & n_17969;
assign n_17979 = n_17970 ^ n_17959;
assign n_17980 = n_17443 ^ n_17971;
assign n_17981 = n_17972 ^ n_17410;
assign n_17982 = n_16878 & ~n_17974;
assign n_17983 = n_17976 ^ n_17356;
assign n_17984 = n_17977 ^ n_16068;
assign n_17985 = ~n_17977 & ~n_17973;
assign n_17986 = n_17978 ^ x95;
assign n_17987 = ~n_17962 & ~n_17979;
assign n_17988 = n_17979 ^ n_17962;
assign n_17989 = ~n_16454 & n_17981;
assign n_17990 = n_17982 ^ n_17335;
assign n_17991 = n_17304 ^ n_17983;
assign n_17992 = n_17983 & ~n_17364;
assign n_17993 = n_17984 ^ x94;
assign n_17994 = n_17985 ^ n_16068;
assign n_17995 = n_17986 ^ n_17984;
assign n_17996 = n_17971 ^ n_17988;
assign n_17997 = n_17980 ^ n_17988;
assign n_17998 = n_17989 ^ n_17410;
assign n_17999 = n_17990 ^ n_16108;
assign n_18000 = n_17991 ^ n_17356;
assign n_18001 = n_17860 ^ n_17991;
assign n_18002 = n_17992 ^ n_17304;
assign n_18003 = n_17994 ^ n_17990;
assign n_18004 = ~n_17995 & n_17993;
assign n_18005 = n_17995 ^ x94;
assign n_18006 = ~n_17996 & n_17980;
assign n_18007 = n_16476 & n_17996;
assign n_18008 = n_15935 & n_17998;
assign n_18009 = n_17998 ^ n_15935;
assign n_18010 = ~n_16922 & n_18000;
assign n_18011 = n_18002 ^ n_17385;
assign n_18012 = n_18002 ^ n_17377;
assign n_18013 = n_18003 ^ n_16108;
assign n_18014 = n_18003 & n_17999;
assign n_18015 = n_18004 ^ x94;
assign n_18016 = n_17987 & n_18005;
assign n_18017 = n_18005 ^ n_17987;
assign n_18018 = n_18006 ^ n_17443;
assign n_18019 = n_18007 ^ n_17443;
assign n_18020 = n_18008 ^ n_15962;
assign n_18021 = x231 & n_18009;
assign n_18022 = n_18009 ^ x231;
assign n_18023 = n_18010 ^ n_17356;
assign n_18024 = n_18011 ^ n_17377;
assign n_18025 = n_17881 ^ n_18011;
assign n_18026 = n_17385 & n_18012;
assign n_18027 = n_18013 ^ x93;
assign n_18028 = n_18014 ^ n_16108;
assign n_18029 = n_18015 ^ n_18013;
assign n_18030 = n_17483 ^ n_18017;
assign n_18031 = n_18017 ^ n_18018;
assign n_18032 = n_17483 ^ n_18018;
assign n_18033 = n_18019 ^ n_18008;
assign n_18034 = n_18019 ^ n_18020;
assign n_18035 = n_18021 ^ x230;
assign n_18036 = n_18023 ^ n_16150;
assign n_18037 = ~n_16965 & ~n_18024;
assign n_18038 = n_18026 ^ n_17324;
assign n_18039 = n_18028 ^ n_16150;
assign n_18040 = n_18028 ^ n_18023;
assign n_18041 = n_18029 ^ x93;
assign n_18042 = ~n_18029 & n_18027;
assign n_18043 = ~n_18031 & ~n_18030;
assign n_18044 = ~n_16518 & n_18031;
assign n_18045 = n_18032 ^ n_18017;
assign n_18046 = n_18020 & ~n_18033;
assign n_18047 = n_18034 ^ n_18021;
assign n_18048 = n_18034 ^ n_18035;
assign n_18049 = n_18037 ^ n_17377;
assign n_18050 = n_18038 ^ n_17400;
assign n_18051 = n_18039 ^ n_18023;
assign n_18052 = ~n_18036 & n_18040;
assign n_18053 = n_18041 ^ n_18016;
assign n_18054 = ~n_18016 & ~n_18041;
assign n_18055 = n_18042 ^ x93;
assign n_18056 = n_18043 ^ n_17483;
assign n_18057 = n_18044 ^ n_17483;
assign n_18058 = n_18046 ^ n_15962;
assign n_18059 = n_18035 & ~n_18047;
assign n_18060 = n_18022 & n_18048;
assign n_18061 = n_18048 ^ n_18022;
assign n_18062 = n_18049 ^ n_16192;
assign n_18063 = n_18050 ^ n_17346;
assign n_18064 = ~n_18050 & ~n_17408;
assign n_18065 = n_18051 ^ x92;
assign n_18066 = n_18052 ^ n_16150;
assign n_18067 = n_17507 ^ n_18053;
assign n_18068 = n_18055 ^ n_18051;
assign n_18069 = n_18053 ^ n_18056;
assign n_18070 = n_17507 ^ n_18056;
assign n_18071 = n_18057 ^ n_16011;
assign n_18072 = n_18058 ^ n_18057;
assign n_18073 = n_18058 ^ n_16011;
assign n_18074 = n_18059 ^ x230;
assign n_18075 = n_18063 ^ n_17393;
assign n_18076 = n_17902 ^ n_18063;
assign n_18077 = n_18064 ^ n_17346;
assign n_18078 = n_18066 ^ n_16192;
assign n_18079 = n_18066 ^ n_18049;
assign n_18080 = n_18068 ^ x92;
assign n_18081 = ~n_18068 & n_18065;
assign n_18082 = ~n_18069 & n_18067;
assign n_18083 = n_16553 & n_18069;
assign n_18084 = n_18070 ^ n_18053;
assign n_18085 = n_18071 & n_18072;
assign n_18086 = n_18073 ^ n_18057;
assign n_18087 = n_17008 & ~n_18075;
assign n_18088 = n_18077 ^ n_17422;
assign n_18089 = n_18078 ^ n_18049;
assign n_18090 = ~n_18062 & n_18079;
assign n_18091 = n_18054 ^ n_18080;
assign n_18092 = ~n_18080 & n_18054;
assign n_18093 = n_18081 ^ x92;
assign n_18094 = n_18082 ^ n_17507;
assign n_18095 = n_18083 ^ n_17507;
assign n_18096 = n_18085 ^ n_16011;
assign n_18097 = n_18074 ^ n_18086;
assign n_18098 = n_18086 ^ x229;
assign n_18099 = n_18087 ^ n_17393;
assign n_18100 = n_18088 ^ n_17367;
assign n_18101 = ~n_18088 & n_17431;
assign n_18102 = n_18089 ^ x91;
assign n_18103 = n_18090 ^ n_16192;
assign n_18104 = n_17529 ^ n_18091;
assign n_18105 = n_18093 ^ n_18089;
assign n_18106 = n_18094 ^ n_18091;
assign n_18107 = n_17529 ^ n_18094;
assign n_18108 = n_18095 ^ n_16053;
assign n_18109 = n_18096 ^ n_18095;
assign n_18110 = n_18096 ^ n_16053;
assign n_18111 = n_18097 ^ x229;
assign n_18112 = ~n_18097 & n_18098;
assign n_18113 = n_18099 ^ n_16234;
assign n_18114 = n_18100 ^ n_17422;
assign n_18115 = n_17924 ^ n_18100;
assign n_18116 = n_18101 ^ n_17367;
assign n_18117 = n_18103 ^ n_16234;
assign n_18118 = n_18103 ^ n_18099;
assign n_18119 = n_18105 ^ x91;
assign n_18120 = ~n_18105 & n_18102;
assign n_18121 = n_18106 & n_18104;
assign n_18122 = ~n_16603 & ~n_18106;
assign n_18123 = n_18107 ^ n_18091;
assign n_18124 = n_18108 & ~n_18109;
assign n_18125 = n_18110 ^ n_18095;
assign n_18126 = n_18060 & n_18111;
assign n_18127 = n_18111 ^ n_18060;
assign n_18128 = n_18112 ^ x229;
assign n_18129 = ~n_17051 & n_18114;
assign n_18130 = n_17449 ^ n_18116;
assign n_18131 = n_18117 ^ n_18099;
assign n_18132 = ~n_18113 & n_18118;
assign n_18133 = n_18092 ^ n_18119;
assign n_18134 = ~n_18119 & n_18092;
assign n_18135 = n_18120 ^ x91;
assign n_18136 = n_18121 ^ n_17529;
assign n_18137 = n_18122 ^ n_17529;
assign n_18138 = n_18124 ^ n_16053;
assign n_18139 = n_18125 ^ x228;
assign n_18140 = n_18128 ^ n_18125;
assign n_18141 = n_18129 ^ n_17422;
assign n_18142 = n_18130 ^ n_17388;
assign n_18143 = n_18131 ^ x90;
assign n_18144 = n_18132 ^ n_16234;
assign n_18145 = n_18133 ^ n_17540;
assign n_18146 = n_18135 ^ n_18131;
assign n_18147 = n_18136 ^ n_18133;
assign n_18148 = n_18136 ^ n_17540;
assign n_18149 = n_18137 ^ n_16092;
assign n_18150 = n_18138 ^ n_18137;
assign n_18151 = n_18138 ^ n_16092;
assign n_18152 = n_18140 & ~n_18139;
assign n_18153 = n_18140 ^ x228;
assign n_18154 = n_18141 ^ n_16276;
assign n_18155 = n_18142 ^ n_17449;
assign n_18156 = n_18142 ^ n_17939;
assign n_18157 = n_18144 ^ n_16276;
assign n_18158 = n_18141 ^ n_18144;
assign n_18159 = n_18146 ^ x90;
assign n_18160 = ~n_18146 & n_18143;
assign n_18161 = ~n_18147 & n_18145;
assign n_18162 = ~n_16640 & n_18147;
assign n_18163 = n_18148 ^ n_18133;
assign n_18164 = n_18149 & n_18150;
assign n_18165 = n_18151 ^ n_18137;
assign n_18166 = n_18152 ^ x228;
assign n_18167 = ~n_18126 & n_18153;
assign n_18168 = n_18153 ^ n_18126;
assign n_18169 = ~n_17079 & n_18155;
assign n_18170 = n_18156 ^ n_17923;
assign n_18171 = n_18141 ^ n_18157;
assign n_18172 = ~n_18154 & ~n_18158;
assign n_18173 = n_18159 ^ n_18134;
assign n_18174 = n_18134 & ~n_18159;
assign n_18175 = n_18160 ^ x90;
assign n_18176 = n_18161 ^ n_17540;
assign n_18177 = n_18162 ^ n_17540;
assign n_18178 = n_18164 ^ n_16092;
assign n_18179 = n_18165 ^ x227;
assign n_18180 = n_18166 ^ n_18165;
assign n_18181 = n_18169 ^ n_17449;
assign n_18182 = n_18171 ^ x89;
assign n_18183 = n_18172 ^ n_16276;
assign n_18184 = n_18173 ^ n_17563;
assign n_18185 = n_18175 ^ n_18171;
assign n_18186 = n_18176 ^ n_18173;
assign n_18187 = n_18176 ^ n_17563;
assign n_18188 = n_18177 ^ n_16131;
assign n_18189 = n_18178 ^ n_18177;
assign n_18190 = n_18178 ^ n_16131;
assign n_18191 = n_18180 & ~n_18179;
assign n_18192 = n_18180 ^ x227;
assign n_18193 = n_18181 ^ n_16318;
assign n_18194 = n_18183 ^ x88;
assign n_18195 = n_18185 ^ x89;
assign n_18196 = ~n_18185 & n_18182;
assign n_18197 = ~n_18186 & ~n_18184;
assign n_18198 = n_16692 & n_18186;
assign n_18199 = n_18187 ^ n_18173;
assign n_18200 = n_18188 & ~n_18189;
assign n_18201 = n_18190 ^ n_18177;
assign n_18202 = n_18191 ^ x227;
assign n_18203 = n_18167 & n_18192;
assign n_18204 = n_18192 ^ n_18167;
assign n_18205 = n_18194 ^ n_18193;
assign n_18206 = n_18195 ^ n_18174;
assign n_18207 = n_18174 & ~n_18195;
assign n_18208 = n_18196 ^ x89;
assign n_18209 = n_18197 ^ n_17563;
assign n_18210 = n_18198 ^ n_17563;
assign n_18211 = n_18200 ^ n_16131;
assign n_18212 = n_18201 ^ x226;
assign n_18213 = n_18202 ^ n_18201;
assign n_18214 = n_18206 ^ n_17581;
assign n_18215 = n_18208 ^ n_18205;
assign n_18216 = n_18209 ^ n_18206;
assign n_18217 = n_18209 ^ n_17581;
assign n_18218 = n_18210 ^ n_16173;
assign n_18219 = n_18211 ^ n_18210;
assign n_18220 = n_18211 ^ n_16173;
assign n_18221 = ~n_18213 & n_18212;
assign n_18222 = n_18213 ^ x226;
assign n_18223 = n_18215 ^ n_18207;
assign n_18224 = n_18216 & n_18214;
assign n_18225 = ~n_16732 & ~n_18216;
assign n_18226 = n_18217 ^ n_18206;
assign n_18227 = n_18218 & n_18219;
assign n_18228 = n_18220 ^ n_18210;
assign n_18229 = n_18221 ^ x226;
assign n_18230 = n_18222 & ~n_18203;
assign n_18231 = n_18203 ^ n_18222;
assign n_18232 = n_18223 ^ n_17596;
assign n_18233 = n_18224 ^ n_17581;
assign n_18234 = n_18225 ^ n_17581;
assign n_18235 = n_18227 ^ n_16173;
assign n_18236 = n_18228 ^ x225;
assign n_18237 = n_18229 ^ n_18228;
assign n_18238 = n_18233 ^ n_18223;
assign n_18239 = n_18233 ^ n_17596;
assign n_18240 = n_18235 ^ n_16215;
assign n_18241 = n_18234 ^ n_18235;
assign n_18242 = ~n_18237 & n_18236;
assign n_18243 = n_18237 ^ x225;
assign n_18244 = ~n_18238 & n_18232;
assign n_18245 = n_16772 & n_18238;
assign n_18246 = n_18239 ^ n_18223;
assign n_18247 = n_18234 ^ n_18240;
assign n_18248 = ~n_18240 & n_18241;
assign n_18249 = n_18242 ^ x225;
assign n_18250 = ~n_18230 & ~n_18243;
assign n_18251 = n_18243 ^ n_18230;
assign n_18252 = n_18244 ^ n_17596;
assign n_18253 = n_18245 ^ n_17596;
assign n_18254 = n_18247 ^ x224;
assign n_18255 = n_18248 ^ n_16215;
assign n_18256 = n_18249 ^ n_18247;
assign n_18257 = n_18252 ^ n_17613;
assign n_18258 = n_18253 ^ n_16257;
assign n_18259 = n_18255 ^ n_18253;
assign n_18260 = n_18255 ^ n_16257;
assign n_18261 = n_18256 & ~n_18254;
assign n_18262 = n_18256 ^ x224;
assign n_18263 = n_18257 & ~n_17620;
assign n_18264 = n_17461 ^ n_18257;
assign n_18265 = ~n_18258 & ~n_18259;
assign n_18266 = n_18260 ^ n_18253;
assign n_18267 = n_18261 ^ x224;
assign n_18268 = n_18250 & n_18262;
assign n_18269 = n_18262 ^ n_18250;
assign n_18270 = n_18263 ^ n_17461;
assign n_18271 = n_18264 ^ n_17613;
assign n_18272 = n_18265 ^ n_16257;
assign n_18273 = n_18266 ^ x239;
assign n_18274 = n_18267 ^ n_18266;
assign n_18275 = n_17633 ^ n_18270;
assign n_18276 = n_16815 & n_18271;
assign n_18277 = n_18272 ^ n_16299;
assign n_18278 = n_18274 & ~n_18273;
assign n_18279 = n_18274 ^ x239;
assign n_18280 = ~n_18275 & ~n_17640;
assign n_18281 = n_17481 ^ n_18275;
assign n_18282 = n_18276 ^ n_17613;
assign n_18283 = n_18278 ^ x239;
assign n_18284 = ~n_18268 & ~n_18279;
assign n_18285 = n_18279 ^ n_18268;
assign n_18286 = n_18280 ^ n_17481;
assign n_18287 = n_18281 ^ n_17628;
assign n_18288 = n_18282 ^ n_16299;
assign n_18289 = n_18272 ^ n_18282;
assign n_18290 = n_18277 ^ n_18282;
assign n_18291 = n_18286 ^ n_17655;
assign n_18292 = ~n_16858 & n_18287;
assign n_18293 = n_18288 & ~n_18289;
assign n_18294 = n_18283 ^ n_18290;
assign n_18295 = n_18290 ^ x238;
assign n_18296 = ~n_18291 & ~n_17661;
assign n_18297 = n_17517 ^ n_18291;
assign n_18298 = n_18292 ^ n_17628;
assign n_18299 = n_18293 ^ n_16299;
assign n_18300 = n_18294 ^ x238;
assign n_18301 = n_18294 & ~n_18295;
assign n_18302 = n_18296 ^ n_17517;
assign n_18303 = n_18297 ^ n_17655;
assign n_18304 = n_18298 ^ n_16338;
assign n_18305 = n_18299 ^ n_18298;
assign n_18306 = n_18300 & ~n_18284;
assign n_18307 = n_18284 ^ n_18300;
assign n_18308 = n_18301 ^ x238;
assign n_18309 = n_18302 ^ n_17674;
assign n_18310 = n_18302 ^ n_17681;
assign n_18311 = ~n_16902 & ~n_18303;
assign n_18312 = ~n_18305 & n_18304;
assign n_18313 = n_18305 ^ n_16338;
assign n_18314 = ~n_17681 & ~n_18309;
assign n_18315 = n_18310 ^ n_17666;
assign n_18316 = n_18311 ^ n_17655;
assign n_18317 = n_18312 ^ n_16338;
assign n_18318 = n_18308 ^ n_18313;
assign n_18319 = n_18313 ^ x237;
assign n_18320 = n_18314 ^ n_17535;
assign n_18321 = ~n_16945 & n_18315;
assign n_18322 = n_18316 ^ n_16374;
assign n_18323 = n_18317 ^ n_18316;
assign n_18324 = n_18317 ^ n_16374;
assign n_18325 = n_18318 ^ x237;
assign n_18326 = n_18318 & ~n_18319;
assign n_18327 = n_18320 ^ n_17697;
assign n_18328 = n_18321 ^ n_17666;
assign n_18329 = n_18322 & ~n_18323;
assign n_18330 = n_18324 ^ n_18316;
assign n_18331 = ~n_18306 & ~n_18325;
assign n_18332 = n_18325 ^ n_18306;
assign n_18333 = n_18326 ^ x237;
assign n_18334 = n_18327 & ~n_17703;
assign n_18335 = n_17558 ^ n_18327;
assign n_18336 = n_18329 ^ n_16374;
assign n_18337 = n_18330 ^ x236;
assign n_18338 = n_18333 ^ n_18330;
assign n_18339 = n_18334 ^ n_17558;
assign n_18340 = n_18335 ^ n_17697;
assign n_18341 = n_18336 ^ n_16401;
assign n_18342 = n_18328 ^ n_18336;
assign n_18343 = n_18338 & ~n_18337;
assign n_18344 = n_18338 ^ x236;
assign n_18345 = n_18339 ^ n_17716;
assign n_18346 = n_16988 & n_18340;
assign n_18347 = n_18328 ^ n_18341;
assign n_18348 = ~n_18341 & ~n_18342;
assign n_18349 = n_18343 ^ x236;
assign n_18350 = n_18331 & ~n_18344;
assign n_18351 = n_18344 ^ n_18331;
assign n_18352 = n_18345 & ~n_17723;
assign n_18353 = n_17576 ^ n_18345;
assign n_18354 = n_18346 ^ n_17697;
assign n_18355 = n_18347 ^ x235;
assign n_18356 = n_18348 ^ n_16401;
assign n_18357 = n_18349 ^ n_18347;
assign n_18358 = n_18352 ^ n_17576;
assign n_18359 = n_18353 ^ n_17716;
assign n_18360 = n_18022 ^ n_18353;
assign n_18361 = n_18354 ^ n_16422;
assign n_18362 = n_18356 ^ n_18354;
assign n_18363 = n_18356 ^ n_16422;
assign n_18364 = ~n_18357 & n_18355;
assign n_18365 = n_18357 ^ x235;
assign n_18366 = n_18358 ^ n_17737;
assign n_18367 = ~n_17030 & n_18359;
assign n_18368 = ~n_18361 & ~n_18362;
assign n_18369 = n_18363 ^ n_18354;
assign n_18370 = n_18364 ^ x235;
assign n_18371 = n_18350 & n_18365;
assign n_18372 = n_18365 ^ n_18350;
assign n_18373 = n_17598 ^ n_18366;
assign n_18374 = ~n_18366 & ~n_17744;
assign n_18375 = n_18367 ^ n_17716;
assign n_18376 = n_18368 ^ n_16422;
assign n_18377 = n_18370 ^ x234;
assign n_18378 = n_18369 ^ n_18370;
assign n_18379 = n_18373 ^ n_17737;
assign n_18380 = n_18061 ^ n_18373;
assign n_18381 = n_18374 ^ n_17598;
assign n_18382 = n_18375 ^ n_16435;
assign n_18383 = n_18376 ^ n_18375;
assign n_18384 = n_18376 ^ n_16435;
assign n_18385 = n_18369 ^ n_18377;
assign n_18386 = n_18377 & n_18378;
assign n_18387 = n_17070 & ~n_18379;
assign n_18388 = n_18381 ^ n_17751;
assign n_18389 = ~n_18382 & n_18383;
assign n_18390 = n_18384 ^ n_18375;
assign n_18391 = n_18371 & ~n_18385;
assign n_18392 = n_18385 ^ n_18371;
assign n_18393 = n_18386 ^ x234;
assign n_18394 = n_18387 ^ n_17737;
assign n_18395 = n_17625 ^ n_18388;
assign n_18396 = n_18388 & ~n_17760;
assign n_18397 = n_18389 ^ n_16435;
assign n_18398 = n_18390 ^ x233;
assign n_18399 = n_18393 ^ n_18390;
assign n_18400 = n_18394 ^ n_16463;
assign n_18401 = n_18395 ^ n_17751;
assign n_18402 = n_18127 ^ n_18395;
assign n_18403 = n_18396 ^ n_17625;
assign n_18404 = n_18397 ^ n_18394;
assign n_18405 = n_18397 ^ n_16463;
assign n_18406 = ~n_18399 & n_18398;
assign n_18407 = n_18399 ^ x233;
assign n_18408 = n_17107 & n_18401;
assign n_18409 = n_18403 ^ n_17652;
assign n_18410 = n_18403 ^ n_17781;
assign n_18411 = ~n_18400 & ~n_18404;
assign n_18412 = n_18405 ^ n_18394;
assign n_18413 = n_18406 ^ x233;
assign n_18414 = n_18391 & n_18407;
assign n_18415 = n_18407 ^ n_18391;
assign n_18416 = n_18408 ^ n_17751;
assign n_18417 = n_18409 ^ n_17781;
assign n_18418 = n_17788 & ~n_18410;
assign n_18419 = n_18411 ^ n_16463;
assign n_18420 = n_18412 ^ x232;
assign n_18421 = n_18413 ^ n_18412;
assign n_18422 = n_18416 ^ n_16489;
assign n_18423 = n_18417 ^ n_17773;
assign n_18424 = n_18168 ^ n_18417;
assign n_18425 = n_18418 ^ n_17652;
assign n_18426 = n_18419 ^ n_18416;
assign n_18427 = ~n_18421 & n_18420;
assign n_18428 = n_18421 ^ x232;
assign n_18429 = n_17142 & n_18423;
assign n_18430 = n_18425 ^ n_17800;
assign n_18431 = n_18426 ^ n_16489;
assign n_18432 = n_18426 & ~n_18422;
assign n_18433 = n_18427 ^ x232;
assign n_18434 = n_18428 & n_18414;
assign n_18435 = n_18414 ^ n_18428;
assign n_18436 = n_18429 ^ n_17773;
assign n_18437 = n_17673 ^ n_18430;
assign n_18438 = ~n_18430 & n_17807;
assign n_18439 = n_18431 ^ x247;
assign n_18440 = n_18432 ^ n_16489;
assign n_18441 = n_18433 ^ n_18431;
assign n_18442 = n_18433 ^ x247;
assign n_18443 = n_18436 ^ n_16523;
assign n_18444 = n_18437 ^ n_17800;
assign n_18445 = n_18204 ^ n_18437;
assign n_18446 = n_18438 ^ n_17673;
assign n_18447 = n_18440 ^ n_16523;
assign n_18448 = n_18440 ^ n_18436;
assign n_18449 = ~n_18439 & n_18441;
assign n_18450 = n_18442 ^ n_18431;
assign n_18451 = ~n_17171 & n_18444;
assign n_18452 = n_18446 ^ n_17820;
assign n_18453 = n_18447 ^ n_18436;
assign n_18454 = n_18443 & ~n_18448;
assign n_18455 = n_18449 ^ x247;
assign n_18456 = ~n_18434 & n_18450;
assign n_18457 = n_18450 ^ n_18434;
assign n_18458 = n_18451 ^ n_17800;
assign n_18459 = n_17695 ^ n_18452;
assign n_18460 = n_18452 & ~n_17827;
assign n_18461 = n_18453 ^ x246;
assign n_18462 = n_18454 ^ n_16523;
assign n_18463 = n_18455 ^ n_18453;
assign n_18464 = n_18458 ^ n_16558;
assign n_18465 = n_18459 ^ n_17820;
assign n_18466 = n_18231 ^ n_18459;
assign n_18467 = n_18460 ^ n_17695;
assign n_18468 = n_18462 ^ n_16558;
assign n_18469 = n_18462 ^ n_18458;
assign n_18470 = ~n_18463 & n_18461;
assign n_18471 = n_18463 ^ x246;
assign n_18472 = n_17189 & n_18465;
assign n_18473 = n_18467 ^ n_17841;
assign n_18474 = n_18468 ^ n_18458;
assign n_18475 = n_18464 & ~n_18469;
assign n_18476 = n_18470 ^ x246;
assign n_18477 = n_18456 & ~n_18471;
assign n_18478 = n_18472 ^ n_17820;
assign n_18479 = n_17714 ^ n_18473;
assign n_18480 = n_18473 & ~n_17848;
assign n_18481 = n_18474 ^ x245;
assign n_18482 = n_18475 ^ n_16558;
assign n_18483 = n_18476 ^ n_18474;
assign n_18484 = n_18478 ^ n_16596;
assign n_18485 = n_18479 ^ n_17841;
assign n_18486 = n_18251 ^ n_18479;
assign n_18487 = n_18480 ^ n_17714;
assign n_18488 = n_18482 ^ n_16596;
assign n_18489 = n_18482 ^ n_18478;
assign n_18490 = n_18483 ^ x245;
assign n_18491 = ~n_18483 & n_18481;
assign n_18492 = n_17204 & n_18485;
assign n_18493 = n_18487 ^ n_17862;
assign n_18494 = n_18488 ^ n_18478;
assign n_18495 = ~n_18484 & n_18489;
assign n_18496 = n_18490 ^ n_18477;
assign n_18497 = n_18477 & ~n_18490;
assign n_18498 = n_18491 ^ x245;
assign n_18499 = n_18492 ^ n_17841;
assign n_18500 = n_17735 ^ n_18493;
assign n_18501 = n_18493 & n_17869;
assign n_18502 = n_18494 ^ x244;
assign n_18503 = n_18495 ^ n_16596;
assign n_18504 = n_18496 ^ n_17972;
assign n_18505 = n_17972 & n_18496;
assign n_18506 = n_18498 ^ n_18494;
assign n_18507 = n_18499 ^ n_16634;
assign n_18508 = n_18500 ^ n_17862;
assign n_18509 = n_18269 ^ n_18500;
assign n_18510 = n_18501 ^ n_17735;
assign n_18511 = n_18503 ^ n_16634;
assign n_18512 = n_18503 ^ n_18499;
assign n_18513 = n_18504 ^ n_17963;
assign n_18514 = n_17997 ^ n_18505;
assign n_18515 = n_18506 ^ x244;
assign n_18516 = n_18506 & ~n_18502;
assign n_18517 = n_17230 & ~n_18508;
assign n_18518 = n_18510 ^ n_17883;
assign n_18519 = n_18511 ^ n_18499;
assign n_18520 = ~n_18507 & n_18512;
assign n_18521 = ~n_17417 & ~n_18513;
assign n_18522 = n_18515 ^ n_18497;
assign n_18523 = n_18497 & n_18515;
assign n_18524 = n_18516 ^ x244;
assign n_18525 = n_18517 ^ n_17862;
assign n_18526 = n_18518 ^ n_17757;
assign n_18527 = ~n_18518 & n_17890;
assign n_18528 = n_18519 ^ x243;
assign n_18529 = n_18520 ^ n_16634;
assign n_18530 = n_18521 ^ n_17963;
assign n_18531 = n_18522 ^ n_18505;
assign n_18532 = n_18514 ^ n_18522;
assign n_18533 = n_18524 ^ n_18519;
assign n_18534 = n_18525 ^ n_16669;
assign n_18535 = n_18526 ^ n_17883;
assign n_18536 = n_18285 ^ n_18526;
assign n_18537 = n_18527 ^ n_17757;
assign n_18538 = n_18529 ^ n_16669;
assign n_18539 = n_18529 ^ n_18525;
assign n_18540 = n_18530 ^ n_16454;
assign n_18541 = ~n_16454 & ~n_18530;
assign n_18542 = n_17443 & ~n_18531;
assign n_18543 = n_18531 & n_18514;
assign n_18544 = n_18533 ^ x243;
assign n_18545 = n_18533 & ~n_18528;
assign n_18546 = n_17250 & n_18535;
assign n_18547 = n_18537 ^ n_17904;
assign n_18548 = n_18538 ^ n_18525;
assign n_18549 = n_18534 & n_18539;
assign n_18550 = x391 & n_18540;
assign n_18551 = n_18540 ^ x391;
assign n_18552 = n_18541 ^ n_16476;
assign n_18553 = n_18542 ^ n_17997;
assign n_18554 = n_18543 ^ n_17997;
assign n_18555 = n_18544 ^ n_18523;
assign n_18556 = ~n_18523 & ~n_18544;
assign n_18557 = n_18545 ^ x243;
assign n_18558 = n_18546 ^ n_17883;
assign n_18559 = n_17779 ^ n_18547;
assign n_18560 = ~n_18547 & n_17911;
assign n_18561 = n_18548 ^ x242;
assign n_18562 = n_18549 ^ n_16669;
assign n_18563 = n_18550 ^ x390;
assign n_18564 = n_18553 ^ n_18552;
assign n_18565 = n_18553 ^ n_18541;
assign n_18566 = n_18045 ^ n_18554;
assign n_18567 = n_18554 ^ n_18555;
assign n_18568 = n_18045 ^ n_18555;
assign n_18569 = n_18557 ^ n_18548;
assign n_18570 = n_18558 ^ n_16710;
assign n_18571 = n_18559 ^ n_17904;
assign n_18572 = n_18307 ^ n_18559;
assign n_18573 = n_18560 ^ n_17779;
assign n_18574 = n_18562 ^ n_16710;
assign n_18575 = n_18562 ^ n_18558;
assign n_18576 = n_18564 ^ n_18550;
assign n_18577 = n_18564 ^ n_18563;
assign n_18578 = n_18552 & ~n_18565;
assign n_18579 = n_18566 ^ n_18555;
assign n_18580 = ~n_17483 & n_18567;
assign n_18581 = ~n_18567 & ~n_18568;
assign n_18582 = n_18569 ^ x242;
assign n_18583 = ~n_18569 & n_18561;
assign n_18584 = ~n_17271 & n_18571;
assign n_18585 = n_17926 ^ n_18573;
assign n_18586 = n_18574 ^ n_18558;
assign n_18587 = ~n_18570 & ~n_18575;
assign n_18588 = n_18563 & ~n_18576;
assign n_18589 = n_18578 ^ n_16476;
assign n_18590 = n_18580 ^ n_18045;
assign n_18591 = n_18581 ^ n_18045;
assign n_18592 = n_18582 ^ n_18556;
assign n_18593 = ~n_18556 & ~n_18582;
assign n_18594 = n_18583 ^ x242;
assign n_18595 = n_18584 ^ n_17904;
assign n_18596 = n_17798 ^ n_18585;
assign n_18597 = n_18585 & ~n_17933;
assign n_18598 = n_18586 ^ x241;
assign n_18599 = n_18587 ^ n_16710;
assign n_18600 = n_18588 ^ x390;
assign n_18601 = n_18589 ^ n_16518;
assign n_18602 = n_18590 ^ n_16518;
assign n_18603 = n_18589 ^ n_18590;
assign n_18604 = n_18084 ^ n_18591;
assign n_18605 = n_18591 ^ n_18592;
assign n_18606 = n_18084 ^ n_18592;
assign n_18607 = n_18594 ^ n_18586;
assign n_18608 = n_18595 ^ n_16748;
assign n_18609 = n_18596 ^ n_17917;
assign n_18610 = n_18332 ^ n_18596;
assign n_18611 = n_18597 ^ n_17798;
assign n_18612 = n_18594 ^ n_18598;
assign n_18613 = n_18595 ^ n_18599;
assign n_18614 = n_18601 ^ n_18590;
assign n_18615 = n_18602 & n_18603;
assign n_18616 = n_18604 ^ n_18592;
assign n_18617 = ~n_17507 & n_18605;
assign n_18618 = ~n_18605 & n_18606;
assign n_18619 = n_18598 & ~n_18607;
assign n_18620 = n_18608 ^ n_18599;
assign n_18621 = ~n_17287 & ~n_18609;
assign n_18622 = n_18611 ^ n_17817;
assign n_18623 = n_18611 ^ n_17946;
assign n_18624 = n_18593 ^ n_18612;
assign n_18625 = ~n_18612 & n_18593;
assign n_18626 = ~n_18608 & n_18613;
assign n_18627 = n_18600 ^ n_18614;
assign n_18628 = n_18614 ^ x389;
assign n_18629 = n_18615 ^ n_16518;
assign n_18630 = n_18617 ^ n_18084;
assign n_18631 = n_18618 ^ n_18084;
assign n_18632 = n_18619 ^ x241;
assign n_18633 = n_18620 ^ x240;
assign n_18634 = n_18621 ^ n_17917;
assign n_18635 = ~n_17315 & n_18622;
assign n_18636 = n_18622 ^ n_17946;
assign n_18637 = n_17952 & ~n_18623;
assign n_18638 = n_18123 ^ n_18624;
assign n_18639 = n_18626 ^ n_16748;
assign n_18640 = n_18627 ^ x389;
assign n_18641 = ~n_18627 & n_18628;
assign n_18642 = n_18629 ^ n_16553;
assign n_18643 = n_18630 ^ n_16553;
assign n_18644 = n_18629 ^ n_18630;
assign n_18645 = n_18631 ^ n_18624;
assign n_18646 = n_18123 ^ n_18631;
assign n_18647 = n_18632 ^ n_18620;
assign n_18648 = n_18634 ^ n_16792;
assign n_18649 = n_18635 ^ n_17946;
assign n_18650 = n_18351 ^ n_18636;
assign n_18651 = n_18637 ^ n_17817;
assign n_18652 = n_18639 ^ n_18634;
assign n_18653 = n_18640 & n_18577;
assign n_18654 = n_18577 ^ n_18640;
assign n_18655 = n_18641 ^ x389;
assign n_18656 = n_18642 ^ n_18630;
assign n_18657 = ~n_18643 & ~n_18644;
assign n_18658 = n_17529 & ~n_18645;
assign n_18659 = n_18645 & ~n_18638;
assign n_18660 = n_18646 ^ n_18624;
assign n_18661 = n_18647 ^ x240;
assign n_18662 = n_18647 & ~n_18633;
assign n_18663 = n_18649 ^ n_16836;
assign n_18664 = n_18651 ^ n_17965;
assign n_18665 = n_18652 ^ n_16792;
assign n_18666 = n_18652 & ~n_18648;
assign n_18667 = n_18655 ^ n_18656;
assign n_18668 = n_18656 ^ x388;
assign n_18669 = n_18657 ^ n_16553;
assign n_18670 = n_18658 ^ n_18123;
assign n_18671 = n_18659 ^ n_18123;
assign n_18672 = n_18625 ^ n_18661;
assign n_18673 = ~n_18661 & ~n_18625;
assign n_18674 = n_18662 ^ x240;
assign n_18675 = n_17839 ^ n_18664;
assign n_18676 = n_18664 & ~n_17975;
assign n_18677 = n_18665 ^ x255;
assign n_18678 = n_18666 ^ n_16792;
assign n_18679 = n_18667 ^ x388;
assign n_18680 = ~n_18667 & n_18668;
assign n_18681 = n_18669 ^ n_16603;
assign n_18682 = n_18670 ^ n_16603;
assign n_18683 = n_18669 ^ n_18670;
assign n_18684 = n_18163 ^ n_18671;
assign n_18685 = n_18671 ^ n_18672;
assign n_18686 = n_18163 ^ n_18672;
assign n_18687 = n_18674 ^ x255;
assign n_18688 = n_18665 ^ n_18674;
assign n_18689 = n_18675 ^ n_17965;
assign n_18690 = n_18372 ^ n_18675;
assign n_18691 = n_18676 ^ n_17839;
assign n_18692 = n_18678 ^ n_16836;
assign n_18693 = n_18678 ^ n_18649;
assign n_18694 = ~n_18653 & ~n_18679;
assign n_18695 = n_18679 ^ n_18653;
assign n_18696 = n_18680 ^ x388;
assign n_18697 = n_18681 ^ n_18670;
assign n_18698 = n_18682 & n_18683;
assign n_18699 = n_18684 ^ n_18672;
assign n_18700 = n_17540 & ~n_18685;
assign n_18701 = n_18685 & n_18686;
assign n_18702 = n_18665 ^ n_18687;
assign n_18703 = ~n_18677 & n_18688;
assign n_18704 = ~n_17335 & n_18689;
assign n_18705 = n_18691 ^ n_17991;
assign n_18706 = n_18692 ^ n_18649;
assign n_18707 = ~n_18663 & n_18693;
assign n_18708 = n_18696 ^ n_18697;
assign n_18709 = n_18697 ^ x387;
assign n_18710 = n_18698 ^ n_16603;
assign n_18711 = n_18700 ^ n_18163;
assign n_18712 = n_18701 ^ n_18163;
assign n_18713 = n_18673 ^ n_18702;
assign n_18714 = n_18702 & ~n_18673;
assign n_18715 = n_18703 ^ x255;
assign n_18716 = n_18704 ^ n_17965;
assign n_18717 = n_17860 ^ n_18705;
assign n_18718 = n_18705 & n_18001;
assign n_18719 = n_18706 ^ x254;
assign n_18720 = n_18707 ^ n_16836;
assign n_18721 = n_18708 ^ x387;
assign n_18722 = ~n_18708 & n_18709;
assign n_18723 = n_18710 ^ n_16640;
assign n_18724 = n_18711 ^ n_16640;
assign n_18725 = n_18710 ^ n_18711;
assign n_18726 = n_18199 ^ n_18712;
assign n_18727 = n_18712 ^ n_18713;
assign n_18728 = n_18199 ^ n_18713;
assign n_18729 = n_18715 ^ n_18706;
assign n_18730 = n_18716 ^ n_16878;
assign n_18731 = n_18717 ^ n_17991;
assign n_18732 = n_18392 ^ n_18717;
assign n_18733 = n_18718 ^ n_17860;
assign n_18734 = n_18720 ^ n_16878;
assign n_18735 = n_18720 ^ n_18716;
assign n_18736 = ~n_18694 & n_18721;
assign n_18737 = n_18721 ^ n_18694;
assign n_18738 = n_18722 ^ x387;
assign n_18739 = n_18723 ^ n_18711;
assign n_18740 = ~n_18724 & n_18725;
assign n_18741 = n_18726 ^ n_18713;
assign n_18742 = ~n_17563 & n_18727;
assign n_18743 = ~n_18727 & ~n_18728;
assign n_18744 = n_18729 ^ x254;
assign n_18745 = n_18729 & ~n_18719;
assign n_18746 = n_17356 & ~n_18731;
assign n_18747 = n_18733 ^ n_18011;
assign n_18748 = n_18734 ^ n_18716;
assign n_18749 = n_18730 & ~n_18735;
assign n_18750 = n_18738 ^ n_18739;
assign n_18751 = n_18739 ^ x386;
assign n_18752 = n_18740 ^ n_16640;
assign n_18753 = n_18742 ^ n_18199;
assign n_18754 = n_18743 ^ n_18199;
assign n_18755 = n_18744 ^ n_18714;
assign n_18756 = n_18714 & n_18744;
assign n_18757 = n_18745 ^ x254;
assign n_18758 = n_18746 ^ n_17991;
assign n_18759 = n_17881 ^ n_18747;
assign n_18760 = n_18747 & ~n_18025;
assign n_18761 = n_18748 ^ x253;
assign n_18762 = n_18749 ^ n_16878;
assign n_18763 = n_18750 ^ x386;
assign n_18764 = ~n_18750 & n_18751;
assign n_18765 = n_18752 ^ n_16692;
assign n_18766 = n_18753 ^ n_16692;
assign n_18767 = n_18752 ^ n_18753;
assign n_18768 = n_18226 ^ n_18754;
assign n_18769 = n_18754 ^ n_18755;
assign n_18770 = n_18226 ^ n_18755;
assign n_18771 = n_18757 ^ n_18748;
assign n_18772 = n_18758 ^ n_16922;
assign n_18773 = n_18759 ^ n_18011;
assign n_18774 = n_18415 ^ n_18759;
assign n_18775 = n_18760 ^ n_17881;
assign n_18776 = n_18762 ^ n_16922;
assign n_18777 = n_18762 ^ n_18758;
assign n_18778 = n_18736 & n_18763;
assign n_18779 = n_18763 ^ n_18736;
assign n_18780 = n_18764 ^ x386;
assign n_18781 = n_18765 ^ n_18753;
assign n_18782 = ~n_18766 & ~n_18767;
assign n_18783 = n_18768 ^ n_18755;
assign n_18784 = n_17581 & n_18769;
assign n_18785 = ~n_18769 & n_18770;
assign n_18786 = n_18771 ^ x253;
assign n_18787 = ~n_18771 & n_18761;
assign n_18788 = n_17377 & n_18773;
assign n_18789 = n_18775 ^ n_18063;
assign n_18790 = n_18776 ^ n_18758;
assign n_18791 = ~n_18772 & ~n_18777;
assign n_18792 = n_18780 ^ n_18781;
assign n_18793 = n_18781 ^ x385;
assign n_18794 = n_18782 ^ n_16692;
assign n_18795 = n_18784 ^ n_18226;
assign n_18796 = n_18785 ^ n_18226;
assign n_18797 = n_18786 ^ n_18756;
assign n_18798 = n_18756 & ~n_18786;
assign n_18799 = n_18787 ^ x253;
assign n_18800 = n_18788 ^ n_18011;
assign n_18801 = n_18789 ^ n_17902;
assign n_18802 = n_18789 & ~n_18076;
assign n_18803 = n_18790 ^ x252;
assign n_18804 = n_18791 ^ n_16922;
assign n_18805 = n_18792 ^ x385;
assign n_18806 = ~n_18792 & n_18793;
assign n_18807 = n_18794 ^ n_16732;
assign n_18808 = n_18795 ^ n_16732;
assign n_18809 = n_18794 ^ n_18795;
assign n_18810 = n_18246 ^ n_18796;
assign n_18811 = n_18796 ^ n_18797;
assign n_18812 = n_18246 ^ n_18797;
assign n_18813 = n_18799 ^ n_18790;
assign n_18814 = n_18800 ^ n_16965;
assign n_18815 = n_18801 ^ n_18063;
assign n_18816 = n_18435 ^ n_18801;
assign n_18817 = n_18802 ^ n_17902;
assign n_18818 = n_18804 ^ n_16965;
assign n_18819 = n_18804 ^ n_18800;
assign n_18820 = n_18805 & n_18778;
assign n_18821 = n_18778 ^ n_18805;
assign n_18822 = n_18806 ^ x385;
assign n_18823 = n_18807 ^ n_18795;
assign n_18824 = n_18808 & n_18809;
assign n_18825 = n_18810 ^ n_18797;
assign n_18826 = n_17596 & ~n_18811;
assign n_18827 = n_18811 & n_18812;
assign n_18828 = n_18813 ^ x252;
assign n_18829 = n_18813 & ~n_18803;
assign n_18830 = n_17400 & n_18815;
assign n_18831 = n_18817 ^ n_18100;
assign n_18832 = n_18818 ^ n_18800;
assign n_18833 = n_18814 & ~n_18819;
assign n_18834 = n_18822 ^ n_18823;
assign n_18835 = n_18823 ^ x384;
assign n_18836 = n_18824 ^ n_16732;
assign n_18837 = n_18826 ^ n_18246;
assign n_18838 = n_18827 ^ n_18246;
assign n_18839 = n_18828 ^ n_18798;
assign n_18840 = ~n_18798 & ~n_18828;
assign n_18841 = n_18829 ^ x252;
assign n_18842 = n_18830 ^ n_18063;
assign n_18843 = n_18831 ^ n_17924;
assign n_18844 = n_18831 & n_18115;
assign n_18845 = n_18832 ^ x251;
assign n_18846 = n_18833 ^ n_16965;
assign n_18847 = n_18834 ^ x384;
assign n_18848 = ~n_18834 & n_18835;
assign n_18849 = n_18836 ^ n_16772;
assign n_18850 = n_18837 ^ n_16772;
assign n_18851 = n_18836 ^ n_18837;
assign n_18852 = n_18838 ^ n_18264;
assign n_18853 = n_18839 ^ n_18838;
assign n_18854 = n_18839 ^ n_18264;
assign n_18855 = n_18841 ^ n_18832;
assign n_18856 = n_18842 ^ n_17008;
assign n_18857 = n_18843 ^ n_18100;
assign n_18858 = n_18457 ^ n_18843;
assign n_18859 = n_18844 ^ n_17924;
assign n_18860 = n_18846 ^ n_17008;
assign n_18861 = n_18846 ^ n_18842;
assign n_18862 = ~n_18820 & ~n_18847;
assign n_18863 = n_18847 ^ n_18820;
assign n_18864 = n_18848 ^ x384;
assign n_18865 = n_18849 ^ n_18837;
assign n_18866 = n_18850 & n_18851;
assign n_18867 = n_18852 ^ n_18839;
assign n_18868 = ~n_17613 & n_18853;
assign n_18869 = ~n_18853 & ~n_18854;
assign n_18870 = n_18855 ^ x251;
assign n_18871 = n_18855 & ~n_18845;
assign n_18872 = ~n_17422 & ~n_18857;
assign n_18873 = n_18859 ^ n_18170;
assign n_18874 = n_18860 ^ n_18842;
assign n_18875 = ~n_18856 & ~n_18861;
assign n_18876 = n_18864 ^ n_18865;
assign n_18877 = n_18865 ^ x399;
assign n_18878 = n_18866 ^ n_16772;
assign n_18879 = n_18868 ^ n_18264;
assign n_18880 = n_18869 ^ n_18264;
assign n_18881 = n_18870 ^ n_18840;
assign n_18882 = n_18840 & ~n_18870;
assign n_18883 = n_18871 ^ x251;
assign n_18884 = n_18872 ^ n_18100;
assign n_18885 = n_18873 ^ n_18142;
assign n_18886 = n_18873 ^ n_18456;
assign n_18887 = n_18874 ^ x250;
assign n_18888 = n_18875 ^ n_17008;
assign n_18889 = n_18876 ^ x399;
assign n_18890 = n_18876 & ~n_18877;
assign n_18891 = n_18878 ^ n_16815;
assign n_18892 = n_18879 ^ n_16815;
assign n_18893 = n_18878 ^ n_18879;
assign n_18894 = n_18880 ^ n_18281;
assign n_18895 = n_18881 ^ n_18880;
assign n_18896 = n_18881 ^ n_18281;
assign n_18897 = n_18883 ^ n_18874;
assign n_18898 = n_18884 ^ n_17051;
assign n_18899 = n_17449 & n_18885;
assign n_18900 = n_18886 ^ n_18471;
assign n_18901 = n_18888 ^ n_17051;
assign n_18902 = n_18884 ^ n_18888;
assign n_18903 = ~n_18862 & ~n_18889;
assign n_18904 = n_18889 ^ n_18862;
assign n_18905 = n_18890 ^ x399;
assign n_18906 = n_18891 ^ n_18879;
assign n_18907 = ~n_18892 & n_18893;
assign n_18908 = n_18894 ^ n_18881;
assign n_18909 = n_17633 & n_18895;
assign n_18910 = ~n_18895 & n_18896;
assign n_18911 = n_18897 ^ x250;
assign n_18912 = ~n_18897 & n_18887;
assign n_18913 = n_18899 ^ n_18142;
assign n_18914 = n_18884 ^ n_18901;
assign n_18915 = n_18898 & n_18902;
assign n_18916 = n_18905 ^ n_18906;
assign n_18917 = n_18906 ^ x398;
assign n_18918 = n_18907 ^ n_16815;
assign n_18919 = n_18909 ^ n_18281;
assign n_18920 = n_18910 ^ n_18281;
assign n_18921 = n_18882 ^ n_18911;
assign n_18922 = ~n_18911 & ~n_18882;
assign n_18923 = n_18912 ^ x250;
assign n_18924 = n_18913 ^ n_17079;
assign n_18925 = n_18914 ^ x249;
assign n_18926 = n_18915 ^ n_17051;
assign n_18927 = n_18916 ^ x398;
assign n_18928 = n_18916 & ~n_18917;
assign n_18929 = n_18918 ^ n_16858;
assign n_18930 = n_18919 ^ n_16858;
assign n_18931 = n_18919 ^ n_18918;
assign n_18932 = n_18920 ^ n_18921;
assign n_18933 = n_18921 ^ n_18297;
assign n_18934 = n_18923 ^ n_18914;
assign n_18935 = n_18926 ^ x248;
assign n_18936 = n_18903 & ~n_18927;
assign n_18937 = n_18927 ^ n_18903;
assign n_18938 = n_18928 ^ x398;
assign n_18939 = n_18919 ^ n_18929;
assign n_18940 = n_18930 & n_18931;
assign n_18941 = ~n_17655 & n_18932;
assign n_18942 = ~n_18932 & ~n_18933;
assign n_18943 = n_18933 ^ n_18920;
assign n_18944 = n_18934 ^ x249;
assign n_18945 = ~n_18934 & n_18925;
assign n_18946 = n_18935 ^ n_18924;
assign n_18947 = n_18938 ^ n_18939;
assign n_18948 = n_18939 ^ x397;
assign n_18949 = n_18940 ^ n_16858;
assign n_18950 = n_18941 ^ n_18297;
assign n_18951 = n_18942 ^ n_18297;
assign n_18952 = n_18944 ^ n_18922;
assign n_18953 = n_18922 & ~n_18944;
assign n_18954 = n_18945 ^ x249;
assign n_18955 = n_18947 ^ x397;
assign n_18956 = ~n_18947 & n_18948;
assign n_18957 = n_18949 ^ n_16902;
assign n_18958 = n_18949 ^ n_18950;
assign n_18959 = n_18951 ^ n_18310;
assign n_18960 = n_18951 ^ n_18952;
assign n_18961 = n_18952 ^ n_18310;
assign n_18962 = n_18954 ^ n_18946;
assign n_18963 = ~n_18955 & ~n_18936;
assign n_18964 = n_18936 ^ n_18955;
assign n_18965 = n_18956 ^ x397;
assign n_18966 = n_18957 ^ n_18950;
assign n_18967 = n_18957 & n_18958;
assign n_18968 = n_18959 ^ n_18952;
assign n_18969 = n_17674 & n_18960;
assign n_18970 = ~n_18960 & ~n_18961;
assign n_18971 = n_18962 ^ n_18953;
assign n_18972 = n_18965 ^ n_18966;
assign n_18973 = n_18966 ^ x396;
assign n_18974 = n_18967 ^ n_16902;
assign n_18975 = n_18969 ^ n_18310;
assign n_18976 = n_18970 ^ n_18310;
assign n_18977 = n_18971 ^ n_18335;
assign n_18978 = n_18972 ^ x396;
assign n_18979 = ~n_18972 & n_18973;
assign n_18980 = n_18974 ^ n_16945;
assign n_18981 = n_18975 ^ n_16945;
assign n_18982 = n_18975 ^ n_18974;
assign n_18983 = n_18976 ^ n_18971;
assign n_18984 = n_18976 ^ n_18335;
assign n_18985 = n_18963 & ~n_18978;
assign n_18986 = n_18979 ^ x396;
assign n_18987 = n_18975 ^ n_18980;
assign n_18988 = n_18981 & ~n_18982;
assign n_18989 = n_17697 & n_18983;
assign n_18990 = ~n_18983 & ~n_18977;
assign n_18991 = n_18984 ^ n_18971;
assign n_18992 = n_18986 ^ n_18987;
assign n_18993 = n_18987 ^ x395;
assign n_18994 = n_18988 ^ n_16945;
assign n_18995 = n_18989 ^ n_18335;
assign n_18996 = n_18990 ^ n_18335;
assign n_18997 = n_18992 ^ x395;
assign n_18998 = n_18992 & ~n_18993;
assign n_18999 = n_18994 ^ n_16988;
assign n_19000 = n_18995 ^ n_16988;
assign n_19001 = n_18994 ^ n_18995;
assign n_19002 = n_18996 ^ n_18022;
assign n_19003 = n_18360 ^ n_18996;
assign n_19004 = n_18997 ^ n_18985;
assign n_19005 = ~n_18985 & ~n_18997;
assign n_19006 = n_18998 ^ x395;
assign n_19007 = n_18999 ^ n_18995;
assign n_19008 = n_19000 & n_19001;
assign n_19009 = n_17716 & ~n_19002;
assign n_19010 = n_19002 & ~n_18360;
assign n_19011 = n_19004 ^ n_17963;
assign n_19012 = n_18504 & n_19004;
assign n_19013 = n_19004 ^ n_17972;
assign n_19014 = n_19004 ^ n_18504;
assign n_19015 = n_19006 ^ n_19007;
assign n_19016 = n_19007 ^ x394;
assign n_19017 = n_19008 ^ n_16988;
assign n_19018 = n_19009 ^ n_18353;
assign n_19019 = n_19010 ^ n_18353;
assign n_19020 = x167 & ~n_19011;
assign n_19021 = n_19011 ^ x167;
assign n_19022 = n_18532 ^ n_19012;
assign n_19023 = ~n_17417 & n_19013;
assign n_19024 = n_19015 ^ x394;
assign n_19025 = n_19015 & ~n_19016;
assign n_19026 = n_19017 ^ n_17030;
assign n_19027 = n_19018 ^ n_19017;
assign n_19028 = n_19019 ^ n_18373;
assign n_19029 = n_19020 ^ x166;
assign n_19030 = n_19023 ^ n_17443;
assign n_19031 = n_19005 ^ n_19024;
assign n_19032 = ~n_19024 & n_19005;
assign n_19033 = n_19025 ^ x394;
assign n_19034 = n_19018 ^ n_19026;
assign n_19035 = ~n_19026 & ~n_19027;
assign n_19036 = n_18061 ^ n_19028;
assign n_19037 = ~n_19028 & n_18380;
assign n_19038 = n_19031 ^ n_19012;
assign n_19039 = n_19022 ^ n_19031;
assign n_19040 = n_19033 ^ n_19034;
assign n_19041 = n_19034 ^ x393;
assign n_19042 = n_19035 ^ n_17030;
assign n_19043 = n_19036 ^ n_18373;
assign n_19044 = n_19037 ^ n_18061;
assign n_19045 = n_19038 ^ n_17997;
assign n_19046 = n_19038 & ~n_19022;
assign n_19047 = n_19040 ^ x393;
assign n_19048 = n_19040 & ~n_19041;
assign n_19049 = n_19042 ^ n_17070;
assign n_19050 = ~n_17737 & n_19043;
assign n_19051 = n_19044 ^ n_18127;
assign n_19052 = n_19044 ^ n_18395;
assign n_19053 = n_19045 ^ n_19023;
assign n_19054 = n_19046 ^ n_18532;
assign n_19055 = n_19047 ^ n_19032;
assign n_19056 = ~n_19032 & n_19047;
assign n_19057 = n_19048 ^ x393;
assign n_19058 = n_19050 ^ n_18373;
assign n_19059 = ~n_17751 & n_19051;
assign n_19060 = n_19051 ^ n_18395;
assign n_19061 = ~n_18402 & n_19052;
assign n_19062 = n_19053 ^ n_17443;
assign n_19063 = n_19053 & n_19030;
assign n_19064 = n_18579 ^ n_19054;
assign n_19065 = n_19054 ^ n_19055;
assign n_19066 = n_18579 ^ n_19055;
assign n_19067 = n_19057 ^ x392;
assign n_19068 = n_19049 ^ n_19058;
assign n_19069 = n_19058 ^ n_17070;
assign n_19070 = n_19042 ^ n_19058;
assign n_19071 = n_19059 ^ n_18395;
assign n_19072 = n_19061 ^ n_18127;
assign n_19073 = n_19062 ^ n_19020;
assign n_19074 = n_19062 ^ n_19029;
assign n_19075 = n_19063 ^ n_17443;
assign n_19076 = n_19064 ^ n_19055;
assign n_19077 = n_19065 ^ n_18045;
assign n_19078 = n_19065 & ~n_19066;
assign n_19079 = n_19057 ^ n_19068;
assign n_19080 = n_19069 & n_19070;
assign n_19081 = n_19071 ^ n_17107;
assign n_19082 = n_19072 ^ n_18168;
assign n_19083 = n_19072 ^ n_18417;
assign n_19084 = n_19029 & n_19073;
assign n_19085 = n_19075 ^ n_17483;
assign n_19086 = n_19077 ^ n_19075;
assign n_19087 = n_19078 ^ n_18579;
assign n_19088 = n_19079 ^ x392;
assign n_19089 = n_19079 & n_19067;
assign n_19090 = n_19080 ^ n_17070;
assign n_19091 = n_19082 ^ n_18417;
assign n_19092 = n_18424 & ~n_19083;
assign n_19093 = n_19084 ^ x166;
assign n_19094 = n_19077 ^ n_19085;
assign n_19095 = ~n_19085 & ~n_19086;
assign n_19096 = n_19056 ^ n_19088;
assign n_19097 = ~n_19088 & ~n_19056;
assign n_19098 = n_19089 ^ x392;
assign n_19099 = n_19090 ^ n_19071;
assign n_19100 = n_19091 ^ n_18409;
assign n_19101 = n_19092 ^ n_18168;
assign n_19102 = n_19093 ^ n_19094;
assign n_19103 = n_19094 ^ x165;
assign n_19104 = n_19095 ^ n_17483;
assign n_19105 = n_19087 ^ n_19096;
assign n_19106 = n_18616 ^ n_19096;
assign n_19107 = n_19098 ^ x407;
assign n_19108 = n_19099 ^ n_17107;
assign n_19109 = n_19099 & ~n_19081;
assign n_19110 = n_17781 & n_19100;
assign n_19111 = n_19101 ^ n_18437;
assign n_19112 = n_19102 ^ x165;
assign n_19113 = n_19102 & ~n_19103;
assign n_19114 = n_19104 ^ n_17507;
assign n_19115 = n_19105 ^ n_18084;
assign n_19116 = n_18616 ^ n_19105;
assign n_19117 = n_19105 & ~n_19106;
assign n_19118 = n_19107 ^ n_19108;
assign n_19119 = n_19108 ^ x407;
assign n_19120 = n_19098 ^ n_19108;
assign n_19121 = n_19109 ^ n_17107;
assign n_19122 = n_19110 ^ n_18409;
assign n_19123 = n_18204 ^ n_19111;
assign n_19124 = ~n_19111 & ~n_18445;
assign n_19125 = ~n_19112 & ~n_19074;
assign n_19126 = n_19074 ^ n_19112;
assign n_19127 = n_19113 ^ x165;
assign n_19128 = n_19114 ^ n_19115;
assign n_19129 = n_19115 ^ n_17507;
assign n_19130 = n_19104 ^ n_19115;
assign n_19131 = n_19117 ^ n_18616;
assign n_19132 = n_19097 ^ n_19118;
assign n_19133 = ~n_19118 & n_19097;
assign n_19134 = ~n_19119 & n_19120;
assign n_19135 = n_19121 ^ n_17142;
assign n_19136 = n_19122 ^ n_17142;
assign n_19137 = n_19121 ^ n_19122;
assign n_19138 = n_19123 ^ n_18437;
assign n_19139 = n_19124 ^ n_18204;
assign n_19140 = n_19127 ^ n_19128;
assign n_19141 = n_19128 ^ x164;
assign n_19142 = ~n_19129 & n_19130;
assign n_19143 = n_18660 ^ n_19131;
assign n_19144 = n_19131 ^ n_19132;
assign n_19145 = n_18660 ^ n_19132;
assign n_19146 = n_19134 ^ x407;
assign n_19147 = n_19135 ^ n_19122;
assign n_19148 = n_19136 & ~n_19137;
assign n_19149 = n_17800 & ~n_19138;
assign n_19150 = n_19139 ^ n_18459;
assign n_19151 = n_19140 ^ x164;
assign n_19152 = ~n_19140 & n_19141;
assign n_19153 = n_19142 ^ n_17507;
assign n_19154 = n_19143 ^ n_19132;
assign n_19155 = n_19144 ^ n_18123;
assign n_19156 = ~n_19144 & ~n_19145;
assign n_19157 = n_19146 ^ n_19147;
assign n_19158 = n_19147 ^ x406;
assign n_19159 = n_19148 ^ n_17142;
assign n_19160 = n_19149 ^ n_18437;
assign n_19161 = n_18231 ^ n_19150;
assign n_19162 = ~n_19150 & n_18466;
assign n_19163 = n_19151 & n_19125;
assign n_19164 = n_19125 ^ n_19151;
assign n_19165 = n_19152 ^ x164;
assign n_19166 = n_19153 ^ n_17529;
assign n_19167 = n_19021 ^ n_19154;
assign n_19168 = n_19155 ^ n_17529;
assign n_19169 = n_19153 ^ n_19155;
assign n_19170 = n_19156 ^ n_18660;
assign n_19171 = n_19157 ^ x406;
assign n_19172 = ~n_19157 & n_19158;
assign n_19173 = n_19159 ^ n_17171;
assign n_19174 = n_19160 ^ n_17171;
assign n_19175 = n_19159 ^ n_19160;
assign n_19176 = n_19161 ^ n_18459;
assign n_19177 = n_19162 ^ n_18231;
assign n_19178 = n_19165 ^ x163;
assign n_19179 = n_19166 ^ n_19155;
assign n_19180 = ~n_19168 & ~n_19169;
assign n_19181 = n_18699 ^ n_19170;
assign n_19182 = n_19133 ^ n_19171;
assign n_19183 = ~n_19171 & ~n_19133;
assign n_19184 = n_19172 ^ x406;
assign n_19185 = n_19173 ^ n_19160;
assign n_19186 = ~n_19174 & ~n_19175;
assign n_19187 = ~n_17820 & n_19176;
assign n_19188 = n_19177 ^ n_18479;
assign n_19189 = n_19165 ^ n_19179;
assign n_19190 = n_19180 ^ n_17529;
assign n_19191 = n_19182 ^ n_19170;
assign n_19192 = n_18699 ^ n_19182;
assign n_19193 = n_19181 ^ n_19182;
assign n_19194 = n_19184 ^ n_19185;
assign n_19195 = n_19185 ^ x405;
assign n_19196 = n_19186 ^ n_17171;
assign n_19197 = n_19187 ^ n_18459;
assign n_19198 = n_18251 ^ n_19188;
assign n_19199 = ~n_19188 & n_18486;
assign n_19200 = ~n_19189 & n_19178;
assign n_19201 = n_19189 ^ x163;
assign n_19202 = n_19190 ^ n_17540;
assign n_19203 = n_19191 ^ n_18163;
assign n_19204 = n_19191 & n_19192;
assign n_19205 = n_19193 ^ n_19074;
assign n_19206 = n_19194 ^ x405;
assign n_19207 = n_19194 & ~n_19195;
assign n_19208 = n_19196 ^ n_17189;
assign n_19209 = n_19197 ^ n_17189;
assign n_19210 = n_19196 ^ n_19197;
assign n_19211 = n_19198 ^ n_18479;
assign n_19212 = n_18551 ^ n_19198;
assign n_19213 = n_19199 ^ n_18251;
assign n_19214 = n_19200 ^ x163;
assign n_19215 = n_19163 & n_19201;
assign n_19216 = n_19201 ^ n_19163;
assign n_19217 = n_19202 ^ n_19203;
assign n_19218 = n_19203 ^ n_17540;
assign n_19219 = n_19190 ^ n_19203;
assign n_19220 = n_19204 ^ n_18699;
assign n_19221 = n_19183 ^ n_19206;
assign n_19222 = ~n_19206 & ~n_19183;
assign n_19223 = n_19207 ^ x405;
assign n_19224 = n_19208 ^ n_19197;
assign n_19225 = ~n_19209 & ~n_19210;
assign n_19226 = ~n_17841 & n_19211;
assign n_19227 = n_19213 ^ n_18500;
assign n_19228 = n_19214 ^ n_19217;
assign n_19229 = n_19217 ^ x162;
assign n_19230 = ~n_19218 & n_19219;
assign n_19231 = n_18741 ^ n_19220;
assign n_19232 = n_19220 ^ n_19221;
assign n_19233 = n_18741 ^ n_19221;
assign n_19234 = n_19223 ^ n_19224;
assign n_19235 = n_19224 ^ x404;
assign n_19236 = n_19225 ^ n_17189;
assign n_19237 = n_19226 ^ n_18479;
assign n_19238 = n_18269 ^ n_19227;
assign n_19239 = n_19227 & ~n_18509;
assign n_19240 = n_19228 ^ x162;
assign n_19241 = n_19228 & ~n_19229;
assign n_19242 = n_19230 ^ n_17540;
assign n_19243 = n_19231 ^ n_19221;
assign n_19244 = n_19232 ^ n_18199;
assign n_19245 = n_19232 & ~n_19233;
assign n_19246 = n_19234 ^ x404;
assign n_19247 = ~n_19234 & n_19235;
assign n_19248 = n_19236 ^ n_17204;
assign n_19249 = n_19237 ^ n_17204;
assign n_19250 = n_19236 ^ n_19237;
assign n_19251 = n_19238 ^ n_18500;
assign n_19252 = n_19238 ^ n_18577;
assign n_19253 = n_19239 ^ n_18269;
assign n_19254 = n_19215 & ~n_19240;
assign n_19255 = n_19240 ^ n_19215;
assign n_19256 = n_19241 ^ x162;
assign n_19257 = n_19242 ^ n_17563;
assign n_19258 = n_19126 ^ n_19243;
assign n_19259 = n_19244 ^ n_17563;
assign n_19260 = n_19242 ^ n_19244;
assign n_19261 = n_19245 ^ n_18741;
assign n_19262 = n_19222 ^ n_19246;
assign n_19263 = ~n_19246 & ~n_19222;
assign n_19264 = n_19247 ^ x404;
assign n_19265 = n_19248 ^ n_19237;
assign n_19266 = ~n_19249 & n_19250;
assign n_19267 = ~n_17862 & n_19251;
assign n_19268 = n_19253 ^ n_18526;
assign n_19269 = n_19257 ^ n_19244;
assign n_19270 = ~n_19259 & ~n_19260;
assign n_19271 = n_18783 ^ n_19261;
assign n_19272 = n_19261 ^ n_19262;
assign n_19273 = n_18783 ^ n_19262;
assign n_19274 = n_19264 ^ n_19265;
assign n_19275 = n_19265 ^ x403;
assign n_19276 = n_19266 ^ n_17204;
assign n_19277 = n_19267 ^ n_18500;
assign n_19278 = n_18285 ^ n_19268;
assign n_19279 = ~n_19268 & ~n_18536;
assign n_19280 = n_19256 ^ n_19269;
assign n_19281 = n_19269 ^ x161;
assign n_19282 = n_19270 ^ n_17563;
assign n_19283 = n_19271 ^ n_19262;
assign n_19284 = n_19272 ^ n_18226;
assign n_19285 = ~n_19272 & n_19273;
assign n_19286 = n_19274 ^ x403;
assign n_19287 = n_19274 & ~n_19275;
assign n_19288 = n_19276 ^ n_17230;
assign n_19289 = n_19277 ^ n_17230;
assign n_19290 = n_19276 ^ n_19277;
assign n_19291 = n_19278 ^ n_18526;
assign n_19292 = n_18654 ^ n_19278;
assign n_19293 = n_19279 ^ n_18285;
assign n_19294 = n_19280 ^ x161;
assign n_19295 = n_19280 & ~n_19281;
assign n_19296 = n_19282 ^ n_17581;
assign n_19297 = n_19164 ^ n_19283;
assign n_19298 = n_19284 ^ n_17581;
assign n_19299 = n_19282 ^ n_19284;
assign n_19300 = n_19285 ^ n_18783;
assign n_19301 = n_19286 ^ n_19263;
assign n_19302 = ~n_19263 & ~n_19286;
assign n_19303 = n_19287 ^ x403;
assign n_19304 = n_19288 ^ n_19277;
assign n_19305 = n_19289 & ~n_19290;
assign n_19306 = ~n_17883 & ~n_19291;
assign n_19307 = n_19293 ^ n_18559;
assign n_19308 = n_19294 & ~n_19254;
assign n_19309 = n_19254 ^ n_19294;
assign n_19310 = n_19295 ^ x161;
assign n_19311 = n_19296 ^ n_19284;
assign n_19312 = ~n_19298 & ~n_19299;
assign n_19313 = n_18825 ^ n_19300;
assign n_19314 = n_19301 ^ n_19300;
assign n_19315 = n_18825 ^ n_19301;
assign n_19316 = n_19303 ^ n_19304;
assign n_19317 = n_19304 ^ x402;
assign n_19318 = n_19305 ^ n_17230;
assign n_19319 = n_19306 ^ n_18526;
assign n_19320 = n_18307 ^ n_19307;
assign n_19321 = n_19307 & ~n_18572;
assign n_19322 = n_19310 ^ n_19311;
assign n_19323 = n_19311 ^ x160;
assign n_19324 = n_19312 ^ n_17581;
assign n_19325 = n_19313 ^ n_19301;
assign n_19326 = n_19314 ^ n_18246;
assign n_19327 = n_19314 & ~n_19315;
assign n_19328 = n_19316 ^ x402;
assign n_19329 = ~n_19316 & n_19317;
assign n_19330 = n_19318 ^ n_17250;
assign n_19331 = n_19319 ^ n_17250;
assign n_19332 = n_19318 ^ n_19319;
assign n_19333 = n_19320 ^ n_18559;
assign n_19334 = n_18695 ^ n_19320;
assign n_19335 = n_19321 ^ n_18307;
assign n_19336 = n_19322 ^ x160;
assign n_19337 = ~n_19322 & n_19323;
assign n_19338 = n_19324 ^ n_17596;
assign n_19339 = n_19216 ^ n_19325;
assign n_19340 = n_19326 ^ n_17596;
assign n_19341 = n_19324 ^ n_19326;
assign n_19342 = n_19327 ^ n_18825;
assign n_19343 = n_19302 ^ n_19328;
assign n_19344 = ~n_19328 & ~n_19302;
assign n_19345 = n_19329 ^ x402;
assign n_19346 = n_19330 ^ n_19319;
assign n_19347 = ~n_19331 & n_19332;
assign n_19348 = ~n_17904 & n_19333;
assign n_19349 = n_19335 ^ n_18332;
assign n_19350 = n_19335 ^ n_18596;
assign n_19351 = n_19336 & ~n_19308;
assign n_19352 = n_19308 ^ n_19336;
assign n_19353 = n_19337 ^ x160;
assign n_19354 = n_19338 ^ n_19326;
assign n_19355 = ~n_19340 & n_19341;
assign n_19356 = n_18867 ^ n_19342;
assign n_19357 = n_19342 ^ n_19343;
assign n_19358 = n_18867 ^ n_19343;
assign n_19359 = n_19345 ^ n_19346;
assign n_19360 = n_19346 ^ x401;
assign n_19361 = n_19347 ^ n_17250;
assign n_19362 = n_19348 ^ n_18559;
assign n_19363 = n_17926 & n_19349;
assign n_19364 = n_19349 ^ n_18596;
assign n_19365 = n_18610 & ~n_19350;
assign n_19366 = n_19353 ^ n_19354;
assign n_19367 = n_19354 ^ x175;
assign n_19368 = n_19355 ^ n_17596;
assign n_19369 = n_19356 ^ n_19343;
assign n_19370 = n_19357 ^ n_18264;
assign n_19371 = ~n_19357 & n_19358;
assign n_19372 = n_19359 ^ x401;
assign n_19373 = n_19359 & ~n_19360;
assign n_19374 = n_19361 ^ n_17271;
assign n_19375 = n_19362 ^ n_17271;
assign n_19376 = n_19361 ^ n_19362;
assign n_19377 = n_19363 ^ n_18596;
assign n_19378 = n_19364 ^ n_18737;
assign n_19379 = n_19365 ^ n_18332;
assign n_19380 = n_19366 ^ x175;
assign n_19381 = n_19366 & ~n_19367;
assign n_19382 = n_19368 ^ n_17613;
assign n_19383 = n_19255 ^ n_19369;
assign n_19384 = n_19370 ^ n_17613;
assign n_19385 = n_19368 ^ n_19370;
assign n_19386 = n_19371 ^ n_18867;
assign n_19387 = n_19344 ^ n_19372;
assign n_19388 = ~n_19372 & ~n_19344;
assign n_19389 = n_19373 ^ x401;
assign n_19390 = n_19374 ^ n_19362;
assign n_19391 = n_19375 & n_19376;
assign n_19392 = n_19377 ^ n_17287;
assign n_19393 = n_19379 ^ n_18351;
assign n_19394 = n_19379 ^ n_18636;
assign n_19395 = ~n_19351 & n_19380;
assign n_19396 = n_19380 ^ n_19351;
assign n_19397 = n_19381 ^ x175;
assign n_19398 = n_19382 ^ n_19370;
assign n_19399 = n_19384 & n_19385;
assign n_19400 = n_18908 ^ n_19386;
assign n_19401 = n_19386 ^ n_19387;
assign n_19402 = n_18908 ^ n_19387;
assign n_19403 = n_19389 ^ n_19390;
assign n_19404 = n_19390 ^ x400;
assign n_19405 = n_19391 ^ n_17271;
assign n_19406 = n_19393 ^ n_18636;
assign n_19407 = n_18650 & n_19394;
assign n_19408 = n_19397 ^ n_19398;
assign n_19409 = n_19398 ^ x174;
assign n_19410 = n_19399 ^ n_17613;
assign n_19411 = n_19400 ^ n_19387;
assign n_19412 = n_19401 ^ n_18281;
assign n_19413 = n_19401 & ~n_19402;
assign n_19414 = n_19403 ^ x400;
assign n_19415 = ~n_19403 & n_19404;
assign n_19416 = n_19405 ^ n_19377;
assign n_19417 = n_19406 ^ n_18622;
assign n_19418 = n_18779 ^ n_19406;
assign n_19419 = n_19407 ^ n_18351;
assign n_19420 = n_19408 ^ x174;
assign n_19421 = ~n_19408 & n_19409;
assign n_19422 = n_19410 ^ n_17633;
assign n_19423 = n_19309 ^ n_19411;
assign n_19424 = n_19412 ^ n_17633;
assign n_19425 = n_19410 ^ n_19412;
assign n_19426 = n_19413 ^ n_18908;
assign n_19427 = n_19414 ^ n_19388;
assign n_19428 = n_19388 & n_19414;
assign n_19429 = n_19415 ^ x400;
assign n_19430 = n_19416 ^ n_17287;
assign n_19431 = n_19416 & ~n_19392;
assign n_19432 = ~n_17946 & n_19417;
assign n_19433 = n_19419 ^ n_18675;
assign n_19434 = n_19420 & ~n_19395;
assign n_19435 = n_19395 ^ n_19420;
assign n_19436 = n_19421 ^ x174;
assign n_19437 = n_19422 ^ n_19412;
assign n_19438 = n_19424 & n_19425;
assign n_19439 = n_18943 ^ n_19426;
assign n_19440 = n_19426 ^ n_19427;
assign n_19441 = n_18943 ^ n_19427;
assign n_19442 = n_19429 ^ x415;
assign n_19443 = n_19430 ^ x415;
assign n_19444 = n_19429 ^ n_19430;
assign n_19445 = n_19431 ^ n_17287;
assign n_19446 = n_19432 ^ n_18622;
assign n_19447 = n_18372 ^ n_19433;
assign n_19448 = n_19433 & n_18690;
assign n_19449 = n_19436 ^ n_19437;
assign n_19450 = n_19437 ^ x173;
assign n_19451 = n_19438 ^ n_17633;
assign n_19452 = n_19439 ^ n_19427;
assign n_19453 = n_19440 ^ n_18297;
assign n_19454 = n_19440 & n_19441;
assign n_19455 = n_19442 ^ n_19430;
assign n_19456 = n_19443 & ~n_19444;
assign n_19457 = n_19445 ^ n_17315;
assign n_19458 = n_19446 ^ n_17315;
assign n_19459 = n_19445 ^ n_19446;
assign n_19460 = n_19447 ^ n_18675;
assign n_19461 = n_18821 ^ n_19447;
assign n_19462 = n_19448 ^ n_18372;
assign n_19463 = n_19449 ^ x173;
assign n_19464 = n_19449 & ~n_19450;
assign n_19465 = n_19451 ^ n_17655;
assign n_19466 = n_19352 ^ n_19452;
assign n_19467 = n_19453 ^ n_17655;
assign n_19468 = n_19451 ^ n_19453;
assign n_19469 = n_19454 ^ n_18943;
assign n_19470 = ~n_19428 & ~n_19455;
assign n_19471 = n_19455 ^ n_19428;
assign n_19472 = n_19456 ^ x415;
assign n_19473 = n_19457 ^ n_19446;
assign n_19474 = ~n_19458 & n_19459;
assign n_19475 = n_17965 & ~n_19460;
assign n_19476 = n_19462 ^ n_18717;
assign n_19477 = ~n_19463 & n_19434;
assign n_19478 = n_19434 ^ n_19463;
assign n_19479 = n_19464 ^ x173;
assign n_19480 = n_19465 ^ n_19453;
assign n_19481 = n_19467 & n_19468;
assign n_19482 = n_19469 ^ n_18968;
assign n_19483 = n_18968 ^ n_19471;
assign n_19484 = n_19469 ^ n_19471;
assign n_19485 = n_19472 ^ n_19473;
assign n_19486 = n_19473 ^ x414;
assign n_19487 = n_19474 ^ n_17315;
assign n_19488 = n_19475 ^ n_18675;
assign n_19489 = n_18392 ^ n_19476;
assign n_19490 = n_19476 & n_18732;
assign n_19491 = n_19479 ^ n_19480;
assign n_19492 = n_19480 ^ x172;
assign n_19493 = n_19481 ^ n_17655;
assign n_19494 = n_19482 ^ n_19471;
assign n_19495 = n_19483 & n_19484;
assign n_19496 = n_19484 ^ n_18310;
assign n_19497 = n_19485 ^ x414;
assign n_19498 = ~n_19485 & n_19486;
assign n_19499 = n_19487 ^ n_17335;
assign n_19500 = n_19488 ^ n_17335;
assign n_19501 = n_19487 ^ n_19488;
assign n_19502 = n_19489 ^ n_18717;
assign n_19503 = n_18863 ^ n_19489;
assign n_19504 = n_19490 ^ n_18392;
assign n_19505 = n_19491 ^ x172;
assign n_19506 = ~n_19491 & n_19492;
assign n_19507 = n_19493 ^ n_17674;
assign n_19508 = n_19396 ^ n_19494;
assign n_19509 = n_19495 ^ n_18968;
assign n_19510 = n_19496 ^ n_17674;
assign n_19511 = n_19493 ^ n_19496;
assign n_19512 = n_19497 ^ n_19470;
assign n_19513 = ~n_19470 & n_19497;
assign n_19514 = n_19498 ^ x414;
assign n_19515 = n_19499 ^ n_19488;
assign n_19516 = ~n_19500 & n_19501;
assign n_19517 = n_17991 & ~n_19502;
assign n_19518 = n_19504 ^ n_18759;
assign n_19519 = n_19477 ^ n_19505;
assign n_19520 = ~n_19505 & ~n_19477;
assign n_19521 = n_19506 ^ x172;
assign n_19522 = n_19507 ^ n_19496;
assign n_19523 = n_19509 ^ n_18991;
assign n_19524 = n_19510 & n_19511;
assign n_19525 = n_18991 ^ n_19512;
assign n_19526 = n_19509 ^ n_19512;
assign n_19527 = n_19514 ^ n_19515;
assign n_19528 = n_19515 ^ x413;
assign n_19529 = n_19516 ^ n_17335;
assign n_19530 = n_19517 ^ n_18717;
assign n_19531 = n_18415 ^ n_19518;
assign n_19532 = ~n_19518 & ~n_18774;
assign n_19533 = n_19521 ^ n_19522;
assign n_19534 = n_19522 ^ x171;
assign n_19535 = n_19523 ^ n_19512;
assign n_19536 = n_19524 ^ n_17674;
assign n_19537 = ~n_19525 & ~n_19526;
assign n_19538 = n_19526 ^ n_18335;
assign n_19539 = n_19527 ^ x413;
assign n_19540 = ~n_19527 & n_19528;
assign n_19541 = n_19529 ^ n_17356;
assign n_19542 = n_19530 ^ n_17356;
assign n_19543 = n_19529 ^ n_19530;
assign n_19544 = n_19531 ^ n_18759;
assign n_19545 = n_18904 ^ n_19531;
assign n_19546 = n_19532 ^ n_18415;
assign n_19547 = n_19533 ^ x171;
assign n_19548 = n_19533 & ~n_19534;
assign n_19549 = n_19435 ^ n_19535;
assign n_19550 = n_19536 ^ n_17697;
assign n_19551 = n_19537 ^ n_18991;
assign n_19552 = n_19538 ^ n_17697;
assign n_19553 = n_19536 ^ n_19538;
assign n_19554 = n_19539 ^ n_19513;
assign n_19555 = ~n_19513 & ~n_19539;
assign n_19556 = n_19540 ^ x413;
assign n_19557 = n_19541 ^ n_19530;
assign n_19558 = ~n_19542 & ~n_19543;
assign n_19559 = ~n_18011 & ~n_19544;
assign n_19560 = n_19546 ^ n_18801;
assign n_19561 = n_19520 & n_19547;
assign n_19562 = n_19547 ^ n_19520;
assign n_19563 = n_19548 ^ x171;
assign n_19564 = n_19550 ^ n_19538;
assign n_19565 = n_19551 ^ n_19003;
assign n_19566 = n_19552 & ~n_19553;
assign n_19567 = n_19003 ^ n_19554;
assign n_19568 = n_19551 ^ n_19554;
assign n_19569 = n_19556 ^ n_19557;
assign n_19570 = n_19557 ^ x412;
assign n_19571 = n_19558 ^ n_17356;
assign n_19572 = n_19559 ^ n_18759;
assign n_19573 = n_19560 ^ n_18435;
assign n_19574 = n_19560 & ~n_18816;
assign n_19575 = n_19563 ^ x170;
assign n_19576 = n_19564 ^ x170;
assign n_19577 = n_19563 ^ n_19564;
assign n_19578 = n_19565 ^ n_19554;
assign n_19579 = n_19566 ^ n_17697;
assign n_19580 = n_19567 & n_19568;
assign n_19581 = n_19568 ^ n_18353;
assign n_19582 = n_19569 ^ x412;
assign n_19583 = ~n_19569 & n_19570;
assign n_19584 = n_19571 ^ n_17377;
assign n_19585 = n_19572 ^ n_17377;
assign n_19586 = n_19571 ^ n_19572;
assign n_19587 = n_19573 ^ n_18801;
assign n_19588 = n_18937 ^ n_19573;
assign n_19589 = n_19574 ^ n_18435;
assign n_19590 = n_19575 ^ n_19564;
assign n_19591 = n_19576 & ~n_19577;
assign n_19592 = n_19478 ^ n_19578;
assign n_19593 = n_19579 ^ n_17716;
assign n_19594 = n_19580 ^ n_19003;
assign n_19595 = n_19581 ^ n_17716;
assign n_19596 = n_19579 ^ n_19581;
assign n_19597 = n_19555 ^ n_19582;
assign n_19598 = ~n_19582 & n_19555;
assign n_19599 = n_19583 ^ x412;
assign n_19600 = n_19584 ^ n_19572;
assign n_19601 = ~n_19585 & n_19586;
assign n_19602 = ~n_18063 & n_19587;
assign n_19603 = n_19589 ^ n_18843;
assign n_19604 = n_19561 & ~n_19590;
assign n_19605 = n_19590 ^ n_19561;
assign n_19606 = n_19591 ^ x170;
assign n_19607 = n_19593 ^ n_19581;
assign n_19608 = ~n_19595 & n_19596;
assign n_19609 = n_19594 ^ n_19597;
assign n_19610 = n_19597 ^ n_19036;
assign n_19611 = n_19599 ^ n_19600;
assign n_19612 = n_19600 ^ x411;
assign n_19613 = n_19601 ^ n_17377;
assign n_19614 = n_19602 ^ n_18801;
assign n_19615 = n_19603 ^ n_18457;
assign n_19616 = ~n_19603 & n_18858;
assign n_19617 = n_19606 ^ n_19607;
assign n_19618 = n_19607 ^ x169;
assign n_19619 = n_19608 ^ n_17716;
assign n_19620 = n_19609 ^ n_18373;
assign n_19621 = n_19609 ^ n_19036;
assign n_19622 = n_19609 & n_19610;
assign n_19623 = n_19611 ^ x411;
assign n_19624 = n_19611 & ~n_19612;
assign n_19625 = n_19613 ^ n_17400;
assign n_19626 = n_19614 ^ n_17400;
assign n_19627 = n_19613 ^ n_19614;
assign n_19628 = n_19615 ^ n_18843;
assign n_19629 = n_18964 ^ n_19615;
assign n_19630 = n_19616 ^ n_18457;
assign n_19631 = n_19617 ^ x169;
assign n_19632 = n_19617 & ~n_19618;
assign n_19633 = n_19619 ^ n_17737;
assign n_19634 = n_19620 ^ n_17737;
assign n_19635 = n_19619 ^ n_19620;
assign n_19636 = n_19519 ^ n_19621;
assign n_19637 = n_19622 ^ n_19036;
assign n_19638 = n_19598 ^ n_19623;
assign n_19639 = ~n_19623 & ~n_19598;
assign n_19640 = n_19624 ^ x411;
assign n_19641 = n_19625 ^ n_19614;
assign n_19642 = ~n_19626 & n_19627;
assign n_19643 = ~n_18100 & n_19628;
assign n_19644 = n_19630 ^ n_18900;
assign n_19645 = ~n_19604 & ~n_19631;
assign n_19646 = n_19631 ^ n_19604;
assign n_19647 = n_19632 ^ x169;
assign n_19648 = n_19633 ^ n_19620;
assign n_19649 = n_19634 & n_19635;
assign n_19650 = n_19060 ^ n_19637;
assign n_19651 = n_19637 ^ n_19638;
assign n_19652 = n_19060 ^ n_19638;
assign n_19653 = n_19640 ^ n_19641;
assign n_19654 = n_19641 ^ x410;
assign n_19655 = n_19642 ^ n_17400;
assign n_19656 = n_19643 ^ n_18843;
assign n_19657 = n_19644 ^ n_18873;
assign n_19658 = n_19644 ^ n_18963;
assign n_19659 = n_19647 ^ n_19648;
assign n_19660 = n_19648 ^ x168;
assign n_19661 = n_19649 ^ n_17737;
assign n_19662 = n_19650 ^ n_19638;
assign n_19663 = n_19651 ^ n_18395;
assign n_19664 = ~n_19651 & ~n_19652;
assign n_19665 = n_19653 ^ x410;
assign n_19666 = n_19653 & ~n_19654;
assign n_19667 = n_19655 ^ n_17422;
assign n_19668 = n_19656 ^ n_17422;
assign n_19669 = n_19656 ^ n_19655;
assign n_19670 = n_18142 & n_19657;
assign n_19671 = n_19658 ^ n_18978;
assign n_19672 = n_19659 ^ x168;
assign n_19673 = ~n_19659 & n_19660;
assign n_19674 = n_19562 ^ n_19662;
assign n_19675 = n_19661 ^ n_19663;
assign n_19676 = n_19663 ^ n_17751;
assign n_19677 = n_19664 ^ n_19060;
assign n_19678 = n_19639 ^ n_19665;
assign n_19679 = ~n_19665 & n_19639;
assign n_19680 = n_19666 ^ x410;
assign n_19681 = n_19656 ^ n_19667;
assign n_19682 = ~n_19668 & ~n_19669;
assign n_19683 = n_19670 ^ n_18873;
assign n_19684 = n_19645 & n_19672;
assign n_19685 = n_19672 ^ n_19645;
assign n_19686 = n_19673 ^ x168;
assign n_19687 = n_19675 ^ n_17751;
assign n_19688 = ~n_19675 & n_19676;
assign n_19689 = n_19677 ^ n_19678;
assign n_19690 = n_19678 ^ n_19091;
assign n_19691 = n_19680 ^ n_19681;
assign n_19692 = n_19681 ^ x409;
assign n_19693 = n_19682 ^ n_17422;
assign n_19694 = n_19683 ^ n_17449;
assign n_19695 = n_19686 ^ x183;
assign n_19696 = n_19687 ^ x183;
assign n_19697 = n_19686 ^ n_19687;
assign n_19698 = n_19688 ^ n_17751;
assign n_19699 = n_19689 ^ n_18417;
assign n_19700 = n_19689 ^ n_19091;
assign n_19701 = ~n_19689 & ~n_19690;
assign n_19702 = n_19691 ^ x409;
assign n_19703 = n_19691 & ~n_19692;
assign n_19704 = n_19693 ^ x408;
assign n_19705 = n_19695 ^ n_19687;
assign n_19706 = ~n_19696 & n_19697;
assign n_19707 = n_19698 ^ n_19699;
assign n_19708 = n_19699 ^ n_17781;
assign n_19709 = n_19605 ^ n_19700;
assign n_19710 = n_19701 ^ n_19091;
assign n_19711 = n_19679 ^ n_19702;
assign n_19712 = ~n_19702 & n_19679;
assign n_19713 = n_19703 ^ x409;
assign n_19714 = n_19704 ^ n_19694;
assign n_19715 = n_19684 & ~n_19705;
assign n_19716 = n_19705 ^ n_19684;
assign n_19717 = n_19706 ^ x183;
assign n_19718 = n_19707 ^ n_17781;
assign n_19719 = n_19707 & n_19708;
assign n_19720 = n_19710 ^ n_19711;
assign n_19721 = n_19711 ^ n_19123;
assign n_19722 = n_19713 ^ n_19714;
assign n_19723 = n_19717 ^ n_19718;
assign n_19724 = n_19718 ^ x182;
assign n_19725 = n_19719 ^ n_17781;
assign n_19726 = n_19720 ^ n_18437;
assign n_19727 = n_19720 ^ n_19123;
assign n_19728 = n_19720 & n_19721;
assign n_19729 = n_19722 ^ n_19712;
assign n_19730 = n_19723 ^ x182;
assign n_19731 = n_19723 & ~n_19724;
assign n_19732 = n_19725 ^ n_19726;
assign n_19733 = n_19726 ^ n_17800;
assign n_19734 = n_19646 ^ n_19727;
assign n_19735 = n_19728 ^ n_19123;
assign n_19736 = n_19729 ^ n_19161;
assign n_19737 = ~n_19715 & n_19730;
assign n_19738 = n_19730 ^ n_19715;
assign n_19739 = n_19731 ^ x182;
assign n_19740 = n_19732 ^ n_17800;
assign n_19741 = n_19732 & ~n_19733;
assign n_19742 = n_19735 ^ n_19729;
assign n_19743 = n_19735 ^ n_19161;
assign n_19744 = n_19739 ^ n_19740;
assign n_19745 = n_19740 ^ x181;
assign n_19746 = n_19741 ^ n_17800;
assign n_19747 = n_19742 & ~n_19736;
assign n_19748 = n_19742 ^ n_18459;
assign n_19749 = n_19743 ^ n_19729;
assign n_19750 = n_19744 ^ x181;
assign n_19751 = n_19744 & ~n_19745;
assign n_19752 = n_19746 ^ n_17820;
assign n_19753 = n_19747 ^ n_19161;
assign n_19754 = n_19748 ^ n_17820;
assign n_19755 = n_19748 ^ n_19746;
assign n_19756 = n_19685 ^ n_19749;
assign n_19757 = ~n_19750 & ~n_19737;
assign n_19758 = n_19737 ^ n_19750;
assign n_19759 = n_19751 ^ x181;
assign n_19760 = n_19748 ^ n_19752;
assign n_19761 = n_19753 ^ n_19198;
assign n_19762 = n_18551 ^ n_19753;
assign n_19763 = ~n_19754 & ~n_19755;
assign n_19764 = n_19759 ^ n_19760;
assign n_19765 = n_19760 ^ x180;
assign n_19766 = ~n_19212 & ~n_19761;
assign n_19767 = n_19762 ^ n_18479;
assign n_19768 = n_19762 ^ n_19198;
assign n_19769 = n_19763 ^ n_17820;
assign n_19770 = n_19764 ^ x180;
assign n_19771 = n_19764 & ~n_19765;
assign n_19772 = n_19766 ^ n_18551;
assign n_19773 = n_19767 ^ n_17841;
assign n_19774 = n_19716 ^ n_19768;
assign n_19775 = n_19767 ^ n_19769;
assign n_19776 = n_19769 ^ n_17841;
assign n_19777 = ~n_19757 & n_19770;
assign n_19778 = n_19770 ^ n_19757;
assign n_19779 = n_19771 ^ x180;
assign n_19780 = n_19772 ^ n_18577;
assign n_19781 = n_19252 ^ n_19772;
assign n_19782 = ~n_19773 & n_19775;
assign n_19783 = n_19767 ^ n_19776;
assign n_19784 = n_19780 & ~n_19252;
assign n_19785 = n_19780 ^ n_18500;
assign n_19786 = n_19738 ^ n_19781;
assign n_19787 = n_19782 ^ n_17841;
assign n_19788 = n_19779 ^ n_19783;
assign n_19789 = n_19783 ^ x179;
assign n_19790 = n_19784 ^ n_19238;
assign n_19791 = n_19787 ^ n_17862;
assign n_19792 = n_19787 ^ n_19785;
assign n_19793 = n_19788 ^ x179;
assign n_19794 = ~n_19788 & n_19789;
assign n_19795 = n_19790 ^ n_19278;
assign n_19796 = n_19791 ^ n_19785;
assign n_19797 = n_19791 & ~n_19792;
assign n_19798 = n_19777 & ~n_19793;
assign n_19799 = n_19793 ^ n_19777;
assign n_19800 = n_19794 ^ x179;
assign n_19801 = ~n_19795 & n_19292;
assign n_19802 = n_19795 ^ n_18654;
assign n_19803 = n_19796 ^ x178;
assign n_19804 = n_19797 ^ n_17862;
assign n_19805 = n_19800 ^ n_19796;
assign n_19806 = n_19801 ^ n_18654;
assign n_19807 = n_19802 ^ n_19278;
assign n_19808 = n_19758 ^ n_19802;
assign n_19809 = n_19804 ^ n_17883;
assign n_19810 = n_19805 & ~n_19803;
assign n_19811 = n_19805 ^ x178;
assign n_19812 = n_19806 ^ n_19320;
assign n_19813 = n_19807 ^ n_18526;
assign n_19814 = n_19810 ^ x178;
assign n_19815 = n_19798 & n_19811;
assign n_19816 = n_19811 ^ n_19798;
assign n_19817 = n_18695 ^ n_19812;
assign n_19818 = n_19812 & n_19334;
assign n_19819 = n_19813 ^ n_17883;
assign n_19820 = n_19813 ^ n_19804;
assign n_19821 = n_19813 ^ n_19809;
assign n_19822 = n_19814 ^ x177;
assign n_19823 = n_19817 ^ n_19320;
assign n_19824 = n_19778 ^ n_19817;
assign n_19825 = n_19818 ^ n_18695;
assign n_19826 = n_19819 & ~n_19820;
assign n_19827 = n_19814 ^ n_19821;
assign n_19828 = n_19823 ^ n_18559;
assign n_19829 = n_19825 ^ n_19378;
assign n_19830 = n_19825 ^ n_19364;
assign n_19831 = n_19826 ^ n_17883;
assign n_19832 = n_19827 & n_19822;
assign n_19833 = n_19827 ^ x177;
assign n_19834 = n_19828 ^ n_17904;
assign n_19835 = n_19829 ^ n_19364;
assign n_19836 = n_19799 ^ n_19829;
assign n_19837 = ~n_19378 & n_19830;
assign n_19838 = n_19828 ^ n_19831;
assign n_19839 = n_19831 ^ n_17904;
assign n_19840 = n_19832 ^ x177;
assign n_19841 = n_19815 & n_19833;
assign n_19842 = n_19833 ^ n_19815;
assign n_19843 = n_19835 ^ n_18596;
assign n_19844 = n_19837 ^ n_18737;
assign n_19845 = ~n_19834 & n_19838;
assign n_19846 = n_19828 ^ n_19839;
assign n_19847 = n_19843 ^ n_17926;
assign n_19848 = n_19844 ^ n_18779;
assign n_19849 = n_19844 ^ n_19406;
assign n_19850 = n_19845 ^ n_17904;
assign n_19851 = n_19840 ^ n_19846;
assign n_19852 = n_19846 ^ x176;
assign n_19853 = n_19848 ^ n_18636;
assign n_19854 = n_19848 ^ n_19406;
assign n_19855 = n_19418 & n_19849;
assign n_19856 = n_19850 ^ n_19843;
assign n_19857 = n_19851 ^ x176;
assign n_19858 = ~n_19851 & n_19852;
assign n_19859 = n_19853 ^ n_17946;
assign n_19860 = n_19816 ^ n_19854;
assign n_19861 = n_19855 ^ n_18779;
assign n_19862 = n_19856 ^ n_17926;
assign n_19863 = n_19856 & n_19847;
assign n_19864 = n_19841 & ~n_19857;
assign n_19865 = n_19857 ^ n_19841;
assign n_19866 = n_19858 ^ x176;
assign n_19867 = n_19861 ^ n_18821;
assign n_19868 = n_19861 ^ n_19447;
assign n_19869 = n_19862 ^ x191;
assign n_19870 = n_19863 ^ n_17926;
assign n_19871 = n_19862 ^ n_19866;
assign n_19872 = n_19866 ^ x191;
assign n_19873 = n_19867 ^ n_18675;
assign n_19874 = n_19867 ^ n_19447;
assign n_19875 = ~n_19461 & n_19868;
assign n_19876 = n_19870 ^ n_19853;
assign n_19877 = ~n_19869 & n_19871;
assign n_19878 = n_19862 ^ n_19872;
assign n_19879 = n_19873 ^ n_17965;
assign n_19880 = n_19842 ^ n_19874;
assign n_19881 = n_19875 ^ n_18821;
assign n_19882 = n_19876 ^ n_17946;
assign n_19883 = ~n_19876 & ~n_19859;
assign n_19884 = n_19877 ^ x191;
assign n_19885 = n_19864 & n_19878;
assign n_19886 = n_19878 ^ n_19864;
assign n_19887 = n_19881 ^ n_19489;
assign n_19888 = n_19882 ^ x190;
assign n_19889 = n_19883 ^ n_17946;
assign n_19890 = n_19884 ^ n_19882;
assign n_19891 = n_18863 ^ n_19887;
assign n_19892 = ~n_19887 & ~n_19503;
assign n_19893 = n_19889 ^ n_19873;
assign n_19894 = n_19890 & ~n_19888;
assign n_19895 = n_19890 ^ x190;
assign n_19896 = n_19891 ^ n_19489;
assign n_19897 = n_19865 ^ n_19891;
assign n_19898 = n_19892 ^ n_18863;
assign n_19899 = n_19893 ^ n_17965;
assign n_19900 = n_19893 & n_19879;
assign n_19901 = n_19894 ^ x190;
assign n_19902 = n_19885 & n_19895;
assign n_19903 = n_19895 ^ n_19885;
assign n_19904 = n_19896 ^ n_18717;
assign n_19905 = n_19898 ^ n_19531;
assign n_19906 = n_19899 ^ x189;
assign n_19907 = n_19900 ^ n_17965;
assign n_19908 = n_19901 ^ n_19899;
assign n_19909 = n_19904 ^ n_17991;
assign n_19910 = n_18904 ^ n_19905;
assign n_19911 = n_19905 & n_19545;
assign n_19912 = n_19907 ^ n_17991;
assign n_19913 = n_19907 ^ n_19904;
assign n_19914 = n_19908 & ~n_19906;
assign n_19915 = n_19908 ^ x189;
assign n_19916 = n_19910 ^ n_19531;
assign n_19917 = n_19886 ^ n_19910;
assign n_19918 = n_19911 ^ n_18904;
assign n_19919 = n_19912 ^ n_19904;
assign n_19920 = n_19909 & ~n_19913;
assign n_19921 = n_19914 ^ x189;
assign n_19922 = n_19902 & n_19915;
assign n_19923 = n_19915 ^ n_19902;
assign n_19924 = n_19916 ^ n_18759;
assign n_19925 = n_19918 ^ n_19573;
assign n_19926 = n_19919 ^ x188;
assign n_19927 = n_19920 ^ n_17991;
assign n_19928 = n_19921 ^ n_19919;
assign n_19929 = n_19924 ^ n_18011;
assign n_19930 = n_18937 ^ n_19925;
assign n_19931 = n_19925 & n_19588;
assign n_19932 = n_19927 ^ n_18011;
assign n_19933 = n_19927 ^ n_19924;
assign n_19934 = ~n_19928 & n_19926;
assign n_19935 = n_19928 ^ x188;
assign n_19936 = n_19930 ^ n_19573;
assign n_19937 = n_19903 ^ n_19930;
assign n_19938 = n_19931 ^ n_18937;
assign n_19939 = n_19932 ^ n_19924;
assign n_19940 = ~n_19929 & ~n_19933;
assign n_19941 = n_19934 ^ x188;
assign n_19942 = n_19922 & ~n_19935;
assign n_19943 = n_19935 ^ n_19922;
assign n_19944 = n_19936 ^ n_18801;
assign n_19945 = n_19938 ^ n_19615;
assign n_19946 = n_19939 ^ x187;
assign n_19947 = n_19940 ^ n_18011;
assign n_19948 = n_19941 ^ n_19939;
assign n_19949 = n_19944 ^ n_18063;
assign n_19950 = n_19945 ^ n_18964;
assign n_19951 = n_19945 & ~n_19629;
assign n_19952 = n_19947 ^ n_18063;
assign n_19953 = n_19947 ^ n_19944;
assign n_19954 = n_19948 & ~n_19946;
assign n_19955 = n_19948 ^ x187;
assign n_19956 = n_19950 ^ n_19615;
assign n_19957 = n_19923 ^ n_19950;
assign n_19958 = n_19951 ^ n_18964;
assign n_19959 = n_19952 ^ n_19944;
assign n_19960 = ~n_19949 & n_19953;
assign n_19961 = n_19954 ^ x187;
assign n_19962 = n_19942 & n_19955;
assign n_19963 = n_19955 ^ n_19942;
assign n_19964 = n_19956 ^ n_18843;
assign n_19965 = n_19958 ^ n_19671;
assign n_19966 = n_19959 ^ x186;
assign n_19967 = n_19960 ^ n_18063;
assign n_19968 = n_19961 ^ n_19959;
assign n_19969 = n_19014 & ~n_19963;
assign n_19970 = n_19963 ^ n_18496;
assign n_19971 = n_19963 ^ n_19014;
assign n_19972 = n_19964 ^ n_18100;
assign n_19973 = n_19965 ^ n_19644;
assign n_19974 = n_19943 ^ n_19965;
assign n_19975 = n_19967 ^ n_18100;
assign n_19976 = n_19967 ^ n_19964;
assign n_19977 = ~n_19968 & n_19966;
assign n_19978 = n_19968 ^ x186;
assign n_19979 = n_19039 ^ n_19969;
assign n_19980 = n_17972 & n_19970;
assign n_19981 = x263 & ~n_19970;
assign n_19982 = n_19970 ^ x263;
assign n_19983 = n_19973 ^ n_18873;
assign n_19984 = n_19975 ^ n_19964;
assign n_19985 = ~n_19972 & n_19976;
assign n_19986 = n_19977 ^ x186;
assign n_19987 = n_19962 & ~n_19978;
assign n_19988 = n_19978 ^ n_19962;
assign n_19989 = n_19980 ^ n_17997;
assign n_19990 = n_19981 ^ x262;
assign n_19991 = n_19983 ^ n_18142;
assign n_19992 = n_19984 ^ x185;
assign n_19993 = n_19985 ^ n_18100;
assign n_19994 = n_19986 ^ n_19984;
assign n_19995 = n_19988 ^ n_19969;
assign n_19996 = n_19988 ^ n_19979;
assign n_19997 = n_19993 ^ x184;
assign n_19998 = ~n_19994 & n_19992;
assign n_19999 = n_19994 ^ x185;
assign n_20000 = n_19979 & ~n_19995;
assign n_20001 = n_19996 ^ n_19038;
assign n_20002 = n_19997 ^ n_19991;
assign n_20003 = n_19998 ^ x185;
assign n_20004 = ~n_19999 & n_19987;
assign n_20005 = n_19987 ^ n_19999;
assign n_20006 = n_20000 ^ n_19039;
assign n_20007 = n_20001 ^ n_19980;
assign n_20008 = n_20001 ^ n_19989;
assign n_20009 = n_20003 ^ n_20002;
assign n_20010 = n_19076 ^ n_20005;
assign n_20011 = n_20006 ^ n_20005;
assign n_20012 = n_20006 ^ n_19076;
assign n_20013 = n_19989 & n_20007;
assign n_20014 = n_20008 ^ n_19981;
assign n_20015 = n_20008 ^ n_19990;
assign n_20016 = n_20009 ^ n_20004;
assign n_20017 = n_20010 & ~n_20011;
assign n_20018 = n_20012 ^ n_20005;
assign n_20019 = n_20013 ^ n_17997;
assign n_20020 = n_19990 & n_20014;
assign n_20021 = ~n_19982 & ~n_20015;
assign n_20022 = n_20015 ^ n_19982;
assign n_20023 = n_19116 ^ n_20016;
assign n_20024 = n_20017 ^ n_19076;
assign n_20025 = n_20018 ^ n_19065;
assign n_20026 = n_20019 ^ n_18045;
assign n_20027 = n_20020 ^ x262;
assign n_20028 = n_20024 ^ n_20016;
assign n_20029 = n_20024 ^ n_19116;
assign n_20030 = n_20025 ^ n_18045;
assign n_20031 = n_20019 ^ n_20025;
assign n_20032 = n_20026 ^ n_20025;
assign n_20033 = n_20023 & ~n_20028;
assign n_20034 = n_20029 ^ n_20016;
assign n_20035 = n_20030 & n_20031;
assign n_20036 = n_20027 ^ n_20032;
assign n_20037 = n_20032 ^ x261;
assign n_20038 = n_20033 ^ n_19116;
assign n_20039 = n_20034 ^ n_19105;
assign n_20040 = n_20035 ^ n_18045;
assign n_20041 = n_20036 ^ x261;
assign n_20042 = ~n_20036 & n_20037;
assign n_20043 = n_19154 ^ n_20038;
assign n_20044 = n_20039 ^ n_18084;
assign n_20045 = n_20040 ^ n_20039;
assign n_20046 = n_20040 ^ n_18084;
assign n_20047 = n_20021 & n_20041;
assign n_20048 = n_20041 ^ n_20021;
assign n_20049 = n_20042 ^ x261;
assign n_20050 = ~n_20043 & ~n_19167;
assign n_20051 = n_19021 ^ n_20043;
assign n_20052 = n_20044 & ~n_20045;
assign n_20053 = n_20046 ^ n_20039;
assign n_20054 = n_20050 ^ n_19021;
assign n_20055 = n_20051 ^ n_19144;
assign n_20056 = n_20052 ^ n_18084;
assign n_20057 = n_20049 ^ n_20053;
assign n_20058 = n_20053 ^ x260;
assign n_20059 = n_20054 ^ n_19074;
assign n_20060 = n_20054 ^ n_19193;
assign n_20061 = n_20055 ^ n_18123;
assign n_20062 = n_20056 ^ n_20055;
assign n_20063 = n_20056 ^ n_18123;
assign n_20064 = n_20057 ^ x260;
assign n_20065 = n_20057 & ~n_20058;
assign n_20066 = n_19205 & n_20059;
assign n_20067 = n_20060 ^ n_19074;
assign n_20068 = n_20061 & ~n_20062;
assign n_20069 = n_20063 ^ n_20055;
assign n_20070 = n_20047 & ~n_20064;
assign n_20071 = n_20064 ^ n_20047;
assign n_20072 = n_20065 ^ x260;
assign n_20073 = n_20066 ^ n_19193;
assign n_20074 = n_20067 ^ n_19191;
assign n_20075 = n_20068 ^ n_18123;
assign n_20076 = n_20069 ^ x259;
assign n_20077 = n_20072 ^ n_20069;
assign n_20078 = n_19243 ^ n_20073;
assign n_20079 = n_20075 ^ n_18163;
assign n_20080 = n_20074 ^ n_20075;
assign n_20081 = n_20077 & ~n_20076;
assign n_20082 = n_20077 ^ x259;
assign n_20083 = ~n_20078 & n_19258;
assign n_20084 = n_19126 ^ n_20078;
assign n_20085 = n_20074 ^ n_20079;
assign n_20086 = ~n_20079 & n_20080;
assign n_20087 = n_20081 ^ x259;
assign n_20088 = ~n_20082 & n_20070;
assign n_20089 = n_20070 ^ n_20082;
assign n_20090 = n_20083 ^ n_19126;
assign n_20091 = n_20084 ^ n_19232;
assign n_20092 = n_20085 ^ x258;
assign n_20093 = n_20086 ^ n_18163;
assign n_20094 = n_20087 ^ n_20085;
assign n_20095 = n_19283 ^ n_20090;
assign n_20096 = n_20091 ^ n_18199;
assign n_20097 = n_20093 ^ n_20091;
assign n_20098 = n_20093 ^ n_18199;
assign n_20099 = n_20094 & ~n_20092;
assign n_20100 = n_20094 ^ x258;
assign n_20101 = n_20095 & ~n_19297;
assign n_20102 = n_19164 ^ n_20095;
assign n_20103 = n_20096 & n_20097;
assign n_20104 = n_20098 ^ n_20091;
assign n_20105 = n_20099 ^ x258;
assign n_20106 = n_20088 & ~n_20100;
assign n_20107 = n_20100 ^ n_20088;
assign n_20108 = n_20101 ^ n_19164;
assign n_20109 = n_20102 ^ n_19272;
assign n_20110 = n_20103 ^ n_18199;
assign n_20111 = n_20105 ^ n_20104;
assign n_20112 = n_20105 ^ x257;
assign n_20113 = n_20108 ^ n_19325;
assign n_20114 = n_20108 ^ n_19216;
assign n_20115 = n_20109 ^ n_18226;
assign n_20116 = n_20110 ^ n_20109;
assign n_20117 = n_20110 ^ n_18226;
assign n_20118 = n_20111 ^ x257;
assign n_20119 = ~n_20111 & n_20112;
assign n_20120 = n_19339 & ~n_20113;
assign n_20121 = n_20114 ^ n_19325;
assign n_20122 = n_20115 & ~n_20116;
assign n_20123 = n_20117 ^ n_20109;
assign n_20124 = n_20118 & n_20106;
assign n_20125 = n_20106 ^ n_20118;
assign n_20126 = n_20119 ^ x257;
assign n_20127 = n_20120 ^ n_19216;
assign n_20128 = n_20121 ^ n_19314;
assign n_20129 = n_20122 ^ n_18226;
assign n_20130 = n_20123 ^ x256;
assign n_20131 = n_20126 ^ n_20123;
assign n_20132 = n_19369 ^ n_20127;
assign n_20133 = n_20128 ^ n_18246;
assign n_20134 = n_20129 ^ n_20128;
assign n_20135 = n_20129 ^ n_18246;
assign n_20136 = n_20131 & ~n_20130;
assign n_20137 = n_20131 ^ x256;
assign n_20138 = n_20132 & n_19383;
assign n_20139 = n_19255 ^ n_20132;
assign n_20140 = ~n_20133 & ~n_20134;
assign n_20141 = n_20135 ^ n_20128;
assign n_20142 = n_20136 ^ x256;
assign n_20143 = ~n_20124 & n_20137;
assign n_20144 = n_20137 ^ n_20124;
assign n_20145 = n_20138 ^ n_19255;
assign n_20146 = n_20139 ^ n_19357;
assign n_20147 = n_20140 ^ n_18246;
assign n_20148 = n_20141 ^ x271;
assign n_20149 = n_20142 ^ n_20141;
assign n_20150 = n_19411 ^ n_20145;
assign n_20151 = n_20146 ^ n_18264;
assign n_20152 = n_20147 ^ n_20146;
assign n_20153 = n_20147 ^ n_18264;
assign n_20154 = ~n_20149 & n_20148;
assign n_20155 = n_20149 ^ x271;
assign n_20156 = n_20150 & n_19423;
assign n_20157 = n_19309 ^ n_20150;
assign n_20158 = ~n_20151 & ~n_20152;
assign n_20159 = n_20153 ^ n_20146;
assign n_20160 = n_20154 ^ x271;
assign n_20161 = n_20155 & ~n_20143;
assign n_20162 = n_20143 ^ n_20155;
assign n_20163 = n_20156 ^ n_19309;
assign n_20164 = n_20157 ^ n_19401;
assign n_20165 = n_20158 ^ n_18264;
assign n_20166 = n_20159 ^ x270;
assign n_20167 = n_20160 ^ n_20159;
assign n_20168 = n_19452 ^ n_20163;
assign n_20169 = n_20164 ^ n_18281;
assign n_20170 = n_20165 ^ n_20164;
assign n_20171 = n_20165 ^ n_18281;
assign n_20172 = n_20167 & ~n_20166;
assign n_20173 = n_20167 ^ x270;
assign n_20174 = n_20168 & n_19466;
assign n_20175 = n_19352 ^ n_20168;
assign n_20176 = ~n_20169 & n_20170;
assign n_20177 = n_20171 ^ n_20164;
assign n_20178 = n_20172 ^ x270;
assign n_20179 = ~n_20161 & n_20173;
assign n_20180 = n_20173 ^ n_20161;
assign n_20181 = n_20174 ^ n_19352;
assign n_20182 = n_20175 ^ n_19440;
assign n_20183 = n_19982 ^ n_20175;
assign n_20184 = n_20176 ^ n_18281;
assign n_20185 = n_20177 ^ x269;
assign n_20186 = n_20178 ^ n_20177;
assign n_20187 = n_19494 ^ n_20181;
assign n_20188 = n_20182 ^ n_18297;
assign n_20189 = n_20184 ^ n_20182;
assign n_20190 = n_20184 ^ n_18297;
assign n_20191 = ~n_20186 & n_20185;
assign n_20192 = n_20186 ^ x269;
assign n_20193 = n_20187 & n_19508;
assign n_20194 = n_19396 ^ n_20187;
assign n_20195 = ~n_20188 & ~n_20189;
assign n_20196 = n_20190 ^ n_20182;
assign n_20197 = n_20191 ^ x269;
assign n_20198 = n_20179 & ~n_20192;
assign n_20199 = n_20192 ^ n_20179;
assign n_20200 = n_20193 ^ n_19396;
assign n_20201 = n_20194 ^ n_19484;
assign n_20202 = n_20022 ^ n_20194;
assign n_20203 = n_20195 ^ n_18297;
assign n_20204 = n_20196 ^ x268;
assign n_20205 = n_20197 ^ n_20196;
assign n_20206 = n_19535 ^ n_20200;
assign n_20207 = n_20201 ^ n_18310;
assign n_20208 = n_20203 ^ n_20201;
assign n_20209 = n_20203 ^ n_18310;
assign n_20210 = ~n_20205 & n_20204;
assign n_20211 = n_20205 ^ x268;
assign n_20212 = ~n_20206 & ~n_19549;
assign n_20213 = n_19435 ^ n_20206;
assign n_20214 = ~n_20207 & ~n_20208;
assign n_20215 = n_20209 ^ n_20201;
assign n_20216 = n_20210 ^ x268;
assign n_20217 = n_20211 & ~n_20198;
assign n_20218 = n_20198 ^ n_20211;
assign n_20219 = n_20212 ^ n_19435;
assign n_20220 = n_20213 ^ n_19526;
assign n_20221 = n_20048 ^ n_20213;
assign n_20222 = n_20214 ^ n_18310;
assign n_20223 = n_20215 ^ x267;
assign n_20224 = n_20216 ^ n_20215;
assign n_20225 = n_19578 ^ n_20219;
assign n_20226 = n_20220 ^ n_18335;
assign n_20227 = n_20222 ^ n_20220;
assign n_20228 = n_20222 ^ n_18335;
assign n_20229 = n_20224 & ~n_20223;
assign n_20230 = n_20224 ^ x267;
assign n_20231 = n_20225 & ~n_19592;
assign n_20232 = n_19478 ^ n_20225;
assign n_20233 = ~n_20226 & ~n_20227;
assign n_20234 = n_20228 ^ n_20220;
assign n_20235 = n_20229 ^ x267;
assign n_20236 = n_20230 & ~n_20217;
assign n_20237 = n_20217 ^ n_20230;
assign n_20238 = n_20231 ^ n_19478;
assign n_20239 = n_20232 ^ n_19568;
assign n_20240 = n_20232 ^ n_20071;
assign n_20241 = n_20233 ^ n_18335;
assign n_20242 = n_20234 ^ x266;
assign n_20243 = n_20235 ^ n_20234;
assign n_20244 = n_20238 ^ n_19621;
assign n_20245 = n_20239 ^ n_18353;
assign n_20246 = n_20241 ^ n_20239;
assign n_20247 = n_20241 ^ n_18353;
assign n_20248 = ~n_20243 & n_20242;
assign n_20249 = n_20243 ^ x266;
assign n_20250 = n_19519 ^ n_20244;
assign n_20251 = ~n_20244 & n_19636;
assign n_20252 = ~n_20245 & n_20246;
assign n_20253 = n_20247 ^ n_20239;
assign n_20254 = n_20248 ^ x266;
assign n_20255 = ~n_20249 & n_20236;
assign n_20256 = n_20236 ^ n_20249;
assign n_20257 = n_20250 ^ n_19609;
assign n_20258 = n_20089 ^ n_20250;
assign n_20259 = n_20251 ^ n_19519;
assign n_20260 = n_20252 ^ n_18353;
assign n_20261 = n_20253 ^ x265;
assign n_20262 = n_20254 ^ n_20253;
assign n_20263 = n_20257 ^ n_18373;
assign n_20264 = n_19662 ^ n_20259;
assign n_20265 = n_20260 ^ n_20257;
assign n_20266 = n_20260 ^ n_18373;
assign n_20267 = n_20262 & ~n_20261;
assign n_20268 = n_20262 ^ x265;
assign n_20269 = n_19562 ^ n_20264;
assign n_20270 = ~n_20264 & n_19674;
assign n_20271 = n_20263 & ~n_20265;
assign n_20272 = n_20266 ^ n_20257;
assign n_20273 = n_20267 ^ x265;
assign n_20274 = n_20268 & n_20255;
assign n_20275 = n_20255 ^ n_20268;
assign n_20276 = n_20269 ^ n_19651;
assign n_20277 = n_20269 ^ n_20107;
assign n_20278 = n_20270 ^ n_19562;
assign n_20279 = n_20271 ^ n_18373;
assign n_20280 = n_20272 ^ x264;
assign n_20281 = n_20273 ^ n_20272;
assign n_20282 = n_20273 ^ x264;
assign n_20283 = n_20276 ^ n_18395;
assign n_20284 = n_20278 ^ n_19700;
assign n_20285 = n_20279 ^ n_18395;
assign n_20286 = n_20279 ^ n_20276;
assign n_20287 = n_20280 & ~n_20281;
assign n_20288 = n_20282 ^ n_20272;
assign n_20289 = n_19605 ^ n_20284;
assign n_20290 = n_20284 & n_19709;
assign n_20291 = n_20285 ^ n_20276;
assign n_20292 = n_20283 & n_20286;
assign n_20293 = n_20287 ^ x264;
assign n_20294 = n_20274 & ~n_20288;
assign n_20295 = n_20288 ^ n_20274;
assign n_20296 = n_20289 ^ n_19689;
assign n_20297 = n_20289 ^ n_20125;
assign n_20298 = n_20290 ^ n_19605;
assign n_20299 = n_20291 ^ x279;
assign n_20300 = n_20292 ^ n_18395;
assign n_20301 = n_20293 ^ n_20291;
assign n_20302 = n_20293 ^ x279;
assign n_20303 = n_20296 ^ n_18417;
assign n_20304 = n_20298 ^ n_19727;
assign n_20305 = n_20300 ^ n_20296;
assign n_20306 = n_20299 & ~n_20301;
assign n_20307 = n_20302 ^ n_20291;
assign n_20308 = n_19646 ^ n_20304;
assign n_20309 = ~n_20304 & n_19734;
assign n_20310 = n_20305 ^ n_18417;
assign n_20311 = ~n_20305 & ~n_20303;
assign n_20312 = n_20306 ^ x279;
assign n_20313 = n_20294 & ~n_20307;
assign n_20314 = n_20307 ^ n_20294;
assign n_20315 = n_20308 ^ n_19720;
assign n_20316 = n_20144 ^ n_20308;
assign n_20317 = n_20309 ^ n_19646;
assign n_20318 = n_20310 ^ x278;
assign n_20319 = n_20311 ^ n_18417;
assign n_20320 = n_20312 ^ n_20310;
assign n_20321 = n_20315 ^ n_18437;
assign n_20322 = n_19749 ^ n_20317;
assign n_20323 = n_20319 ^ n_20315;
assign n_20324 = ~n_20320 & n_20318;
assign n_20325 = n_20320 ^ x278;
assign n_20326 = n_19685 ^ n_20322;
assign n_20327 = ~n_20322 & n_19756;
assign n_20328 = n_20323 ^ n_18437;
assign n_20329 = n_20323 & ~n_20321;
assign n_20330 = n_20324 ^ x278;
assign n_20331 = ~n_20313 & n_20325;
assign n_20332 = n_20325 ^ n_20313;
assign n_20333 = n_20326 ^ n_19742;
assign n_20334 = n_20326 ^ n_20162;
assign n_20335 = n_20327 ^ n_19685;
assign n_20336 = n_20328 ^ x277;
assign n_20337 = n_20329 ^ n_18437;
assign n_20338 = n_20330 ^ n_20328;
assign n_20339 = n_20333 ^ n_18459;
assign n_20340 = n_20335 ^ n_19768;
assign n_20341 = n_20337 ^ n_18459;
assign n_20342 = n_20337 ^ n_20333;
assign n_20343 = n_20338 & ~n_20336;
assign n_20344 = n_20338 ^ x277;
assign n_20345 = n_19716 ^ n_20340;
assign n_20346 = ~n_20340 & ~n_19774;
assign n_20347 = n_20341 ^ n_20333;
assign n_20348 = n_20339 & n_20342;
assign n_20349 = n_20343 ^ x277;
assign n_20350 = n_20331 & ~n_20344;
assign n_20351 = n_20344 ^ n_20331;
assign n_20352 = n_20345 ^ n_19762;
assign n_20353 = n_20180 ^ n_20345;
assign n_20354 = n_20346 ^ n_19716;
assign n_20355 = n_20347 ^ x276;
assign n_20356 = n_20348 ^ n_18459;
assign n_20357 = n_20349 ^ n_20347;
assign n_20358 = n_20352 ^ n_18479;
assign n_20359 = n_19781 ^ n_20354;
assign n_20360 = n_20356 ^ n_18479;
assign n_20361 = n_20356 ^ n_20352;
assign n_20362 = ~n_20357 & n_20355;
assign n_20363 = n_20357 ^ x276;
assign n_20364 = n_19738 ^ n_20359;
assign n_20365 = ~n_20359 & ~n_19786;
assign n_20366 = n_20360 ^ n_20352;
assign n_20367 = ~n_20358 & n_20361;
assign n_20368 = n_20362 ^ x276;
assign n_20369 = n_20350 & n_20363;
assign n_20370 = n_20363 ^ n_20350;
assign n_20371 = n_20364 ^ n_19780;
assign n_20372 = n_20199 ^ n_20364;
assign n_20373 = n_20365 ^ n_19738;
assign n_20374 = n_20366 ^ x275;
assign n_20375 = n_20367 ^ n_18479;
assign n_20376 = n_20368 ^ n_20366;
assign n_20377 = n_20371 ^ n_18500;
assign n_20378 = n_20373 ^ n_19758;
assign n_20379 = n_20373 ^ n_19802;
assign n_20380 = n_20375 ^ n_18500;
assign n_20381 = n_20375 ^ n_20371;
assign n_20382 = ~n_20376 & n_20374;
assign n_20383 = n_20376 ^ x275;
assign n_20384 = n_20378 ^ n_19802;
assign n_20385 = n_19808 & ~n_20379;
assign n_20386 = n_20380 ^ n_20371;
assign n_20387 = ~n_20377 & ~n_20381;
assign n_20388 = n_20382 ^ x275;
assign n_20389 = ~n_20369 & ~n_20383;
assign n_20390 = n_20383 ^ n_20369;
assign n_20391 = n_20384 ^ n_19807;
assign n_20392 = n_20218 ^ n_20384;
assign n_20393 = n_20385 ^ n_19758;
assign n_20394 = n_20386 ^ x274;
assign n_20395 = n_20387 ^ n_18500;
assign n_20396 = n_20388 ^ n_20386;
assign n_20397 = n_20391 ^ n_18526;
assign n_20398 = n_20393 ^ n_19817;
assign n_20399 = n_20395 ^ n_18526;
assign n_20400 = n_20395 ^ n_20391;
assign n_20401 = ~n_20396 & n_20394;
assign n_20402 = n_20396 ^ x274;
assign n_20403 = n_19778 ^ n_20398;
assign n_20404 = ~n_20398 & n_19824;
assign n_20405 = n_20399 ^ n_20391;
assign n_20406 = ~n_20397 & ~n_20400;
assign n_20407 = n_20401 ^ x274;
assign n_20408 = n_20389 & ~n_20402;
assign n_20409 = n_20402 ^ n_20389;
assign n_20410 = n_20403 ^ n_19823;
assign n_20411 = n_20237 ^ n_20403;
assign n_20412 = n_20404 ^ n_19778;
assign n_20413 = n_20405 ^ x273;
assign n_20414 = n_20406 ^ n_18526;
assign n_20415 = n_20407 ^ n_20405;
assign n_20416 = ~n_19971 & n_20409;
assign n_20417 = n_20409 ^ n_19014;
assign n_20418 = n_20409 ^ n_19004;
assign n_20419 = n_20409 ^ n_19971;
assign n_20420 = n_20410 ^ n_18559;
assign n_20421 = n_20412 ^ n_19829;
assign n_20422 = n_20414 ^ n_18559;
assign n_20423 = n_20414 ^ n_20410;
assign n_20424 = n_20415 ^ x273;
assign n_20425 = n_20415 & ~n_20413;
assign n_20426 = n_20416 ^ n_19996;
assign n_20427 = n_18504 & n_20417;
assign n_20428 = x359 & n_20418;
assign n_20429 = n_20418 ^ x359;
assign n_20430 = n_19799 ^ n_20421;
assign n_20431 = ~n_20421 & n_19836;
assign n_20432 = n_20422 ^ n_20410;
assign n_20433 = n_20420 & ~n_20423;
assign n_20434 = n_20424 ^ n_20408;
assign n_20435 = n_20408 & n_20424;
assign n_20436 = n_20425 ^ x273;
assign n_20437 = n_20427 ^ n_18532;
assign n_20438 = n_20428 ^ x358;
assign n_20439 = n_20430 ^ n_19835;
assign n_20440 = n_20430 ^ n_20256;
assign n_20441 = n_20431 ^ n_19799;
assign n_20442 = n_20432 ^ x272;
assign n_20443 = n_20433 ^ n_18559;
assign n_20444 = n_20434 ^ n_20416;
assign n_20445 = n_20426 ^ n_20434;
assign n_20446 = n_20436 ^ x272;
assign n_20447 = n_20436 ^ n_20432;
assign n_20448 = n_20439 ^ n_18596;
assign n_20449 = n_20441 ^ n_19854;
assign n_20450 = n_20443 ^ n_18596;
assign n_20451 = n_20443 ^ n_20439;
assign n_20452 = n_20444 & n_20426;
assign n_20453 = n_20444 ^ n_19039;
assign n_20454 = n_20446 ^ n_20432;
assign n_20455 = ~n_20442 & n_20447;
assign n_20456 = n_19816 ^ n_20449;
assign n_20457 = n_20449 & n_19860;
assign n_20458 = n_20450 ^ n_20439;
assign n_20459 = n_20448 & n_20451;
assign n_20460 = n_20452 ^ n_19996;
assign n_20461 = n_20453 ^ n_20427;
assign n_20462 = n_20435 ^ n_20454;
assign n_20463 = ~n_20454 & ~n_20435;
assign n_20464 = n_20455 ^ x272;
assign n_20465 = n_20456 ^ n_19848;
assign n_20466 = n_20275 ^ n_20456;
assign n_20467 = n_20457 ^ n_19816;
assign n_20468 = n_20458 ^ x287;
assign n_20469 = n_20459 ^ n_18596;
assign n_20470 = n_20460 ^ n_20018;
assign n_20471 = n_20461 & ~n_20437;
assign n_20472 = n_20461 ^ n_18532;
assign n_20473 = n_20460 ^ n_20462;
assign n_20474 = n_20462 ^ n_20018;
assign n_20475 = n_20464 ^ x287;
assign n_20476 = n_20464 ^ n_20458;
assign n_20477 = n_20465 ^ n_18636;
assign n_20478 = n_20467 ^ n_19874;
assign n_20479 = n_20469 ^ n_20465;
assign n_20480 = n_20470 ^ n_20462;
assign n_20481 = n_20471 ^ n_18532;
assign n_20482 = n_20472 ^ n_20428;
assign n_20483 = n_20473 ^ n_19076;
assign n_20484 = ~n_20473 & n_20474;
assign n_20485 = n_20475 ^ n_20458;
assign n_20486 = ~n_20468 & n_20476;
assign n_20487 = n_19842 ^ n_20478;
assign n_20488 = ~n_20478 & n_19880;
assign n_20489 = n_20479 ^ n_18636;
assign n_20490 = n_20479 & n_20477;
assign n_20491 = n_20481 ^ n_18579;
assign n_20492 = ~n_20482 & n_20438;
assign n_20493 = n_20482 ^ x358;
assign n_20494 = n_20483 ^ n_18579;
assign n_20495 = n_20481 ^ n_20483;
assign n_20496 = n_20484 ^ n_20018;
assign n_20497 = n_20485 ^ n_20463;
assign n_20498 = ~n_20463 & n_20485;
assign n_20499 = n_20486 ^ x287;
assign n_20500 = n_20487 ^ n_19867;
assign n_20501 = n_20295 ^ n_20487;
assign n_20502 = n_20488 ^ n_19842;
assign n_20503 = n_20489 ^ x286;
assign n_20504 = n_20490 ^ n_18636;
assign n_20505 = n_20491 ^ n_20483;
assign n_20506 = n_20492 ^ x358;
assign n_20507 = ~n_20494 & n_20495;
assign n_20508 = n_20496 ^ n_20034;
assign n_20509 = n_20496 ^ n_20497;
assign n_20510 = n_20497 ^ n_20034;
assign n_20511 = n_20499 ^ n_20489;
assign n_20512 = n_20500 ^ n_18675;
assign n_20513 = n_20502 ^ n_19891;
assign n_20514 = n_20504 ^ n_20500;
assign n_20515 = n_20506 ^ n_20505;
assign n_20516 = n_20506 ^ x357;
assign n_20517 = n_20507 ^ n_18579;
assign n_20518 = n_20508 ^ n_20497;
assign n_20519 = n_20509 ^ n_19116;
assign n_20520 = ~n_20509 & n_20510;
assign n_20521 = n_20511 ^ x286;
assign n_20522 = ~n_20511 & n_20503;
assign n_20523 = n_19865 ^ n_20513;
assign n_20524 = ~n_20513 & ~n_19897;
assign n_20525 = n_20514 ^ n_18675;
assign n_20526 = ~n_20514 & ~n_20512;
assign n_20527 = n_20515 ^ x357;
assign n_20528 = ~n_20515 & n_20516;
assign n_20529 = n_20517 ^ n_18616;
assign n_20530 = n_20519 ^ n_18616;
assign n_20531 = n_20517 ^ n_20519;
assign n_20532 = n_20520 ^ n_20034;
assign n_20533 = n_20521 ^ n_20498;
assign n_20534 = n_20498 & ~n_20521;
assign n_20535 = n_20522 ^ x286;
assign n_20536 = n_20523 ^ n_19896;
assign n_20537 = n_20314 ^ n_20523;
assign n_20538 = n_20524 ^ n_19865;
assign n_20539 = n_20525 ^ x285;
assign n_20540 = n_20526 ^ n_18675;
assign n_20541 = n_20527 & n_20493;
assign n_20542 = n_20493 ^ n_20527;
assign n_20543 = n_20528 ^ x357;
assign n_20544 = n_20529 ^ n_20519;
assign n_20545 = ~n_20530 & n_20531;
assign n_20546 = n_20532 ^ n_20051;
assign n_20547 = n_20532 ^ n_20533;
assign n_20548 = n_20533 ^ n_20051;
assign n_20549 = n_20535 ^ n_20525;
assign n_20550 = n_20536 ^ n_18717;
assign n_20551 = n_20538 ^ n_19910;
assign n_20552 = n_20540 ^ n_18717;
assign n_20553 = n_20540 ^ n_20536;
assign n_20554 = n_20543 ^ n_20544;
assign n_20555 = n_20544 ^ x356;
assign n_20556 = n_20545 ^ n_18616;
assign n_20557 = n_20546 ^ n_20533;
assign n_20558 = n_20547 ^ n_19154;
assign n_20559 = ~n_20547 & ~n_20548;
assign n_20560 = n_20549 ^ x285;
assign n_20561 = ~n_20549 & n_20539;
assign n_20562 = n_19886 ^ n_20551;
assign n_20563 = n_20551 & n_19917;
assign n_20564 = n_20552 ^ n_20536;
assign n_20565 = n_20550 & n_20553;
assign n_20566 = n_20554 ^ x356;
assign n_20567 = ~n_20554 & n_20555;
assign n_20568 = n_20556 ^ n_18660;
assign n_20569 = n_20558 ^ n_20556;
assign n_20570 = n_20559 ^ n_20051;
assign n_20571 = n_20560 ^ n_20534;
assign n_20572 = n_20534 & ~n_20560;
assign n_20573 = n_20561 ^ x285;
assign n_20574 = n_20562 ^ n_19916;
assign n_20575 = n_20332 ^ n_20562;
assign n_20576 = n_20563 ^ n_19886;
assign n_20577 = n_20564 ^ x284;
assign n_20578 = n_20565 ^ n_18717;
assign n_20579 = n_20541 & n_20566;
assign n_20580 = n_20566 ^ n_20541;
assign n_20581 = n_20567 ^ x356;
assign n_20582 = n_20558 ^ n_20568;
assign n_20583 = ~n_20568 & n_20569;
assign n_20584 = n_20570 ^ n_20067;
assign n_20585 = n_20570 ^ n_20571;
assign n_20586 = n_20571 ^ n_20067;
assign n_20587 = n_20573 ^ n_20564;
assign n_20588 = n_20574 ^ n_18759;
assign n_20589 = n_20576 ^ n_19930;
assign n_20590 = n_20578 ^ n_18759;
assign n_20591 = n_20578 ^ n_20574;
assign n_20592 = n_20581 ^ x355;
assign n_20593 = n_20581 ^ n_20582;
assign n_20594 = n_20583 ^ n_18660;
assign n_20595 = n_20584 ^ n_20571;
assign n_20596 = n_20585 ^ n_19193;
assign n_20597 = n_20585 & ~n_20586;
assign n_20598 = n_20587 ^ x284;
assign n_20599 = ~n_20587 & n_20577;
assign n_20600 = n_19903 ^ n_20589;
assign n_20601 = n_20589 & ~n_19937;
assign n_20602 = n_20590 ^ n_20574;
assign n_20603 = n_20588 & ~n_20591;
assign n_20604 = n_20593 & n_20592;
assign n_20605 = n_20593 ^ x355;
assign n_20606 = n_20594 ^ n_18699;
assign n_20607 = n_20596 ^ n_18699;
assign n_20608 = n_20594 ^ n_20596;
assign n_20609 = n_20597 ^ n_20067;
assign n_20610 = n_20598 ^ n_20572;
assign n_20611 = ~n_20572 & n_20598;
assign n_20612 = n_20599 ^ x284;
assign n_20613 = n_20600 ^ n_19936;
assign n_20614 = n_20351 ^ n_20600;
assign n_20615 = n_20601 ^ n_19903;
assign n_20616 = n_20602 ^ x283;
assign n_20617 = n_20603 ^ n_18759;
assign n_20618 = n_20604 ^ x355;
assign n_20619 = n_20579 & ~n_20605;
assign n_20620 = n_20605 ^ n_20579;
assign n_20621 = n_20606 ^ n_20596;
assign n_20622 = n_20607 & n_20608;
assign n_20623 = n_20609 ^ n_20084;
assign n_20624 = n_20609 ^ n_20610;
assign n_20625 = n_20610 ^ n_20084;
assign n_20626 = n_20612 ^ n_20602;
assign n_20627 = n_20613 ^ n_18801;
assign n_20628 = n_20615 ^ n_19950;
assign n_20629 = n_20617 ^ n_18801;
assign n_20630 = n_20617 ^ n_20613;
assign n_20631 = n_20618 ^ n_20621;
assign n_20632 = n_20621 ^ x354;
assign n_20633 = n_20622 ^ n_18699;
assign n_20634 = n_20623 ^ n_20610;
assign n_20635 = n_20624 ^ n_19243;
assign n_20636 = ~n_20624 & ~n_20625;
assign n_20637 = n_20626 ^ x283;
assign n_20638 = n_20626 & ~n_20616;
assign n_20639 = n_20628 ^ n_19923;
assign n_20640 = n_20628 & ~n_19957;
assign n_20641 = n_20629 ^ n_20613;
assign n_20642 = n_20627 & ~n_20630;
assign n_20643 = n_20631 ^ x354;
assign n_20644 = ~n_20631 & n_20632;
assign n_20645 = n_20633 ^ n_18741;
assign n_20646 = n_20635 ^ n_18741;
assign n_20647 = n_20633 ^ n_20635;
assign n_20648 = n_20636 ^ n_20084;
assign n_20649 = n_20637 ^ n_20611;
assign n_20650 = n_20611 & ~n_20637;
assign n_20651 = n_20638 ^ x283;
assign n_20652 = n_20639 ^ n_19956;
assign n_20653 = n_20370 ^ n_20639;
assign n_20654 = n_20640 ^ n_19923;
assign n_20655 = n_20641 ^ x282;
assign n_20656 = n_20642 ^ n_18801;
assign n_20657 = ~n_20619 & ~n_20643;
assign n_20658 = n_20643 ^ n_20619;
assign n_20659 = n_20644 ^ x354;
assign n_20660 = n_20645 ^ n_20635;
assign n_20661 = ~n_20646 & n_20647;
assign n_20662 = n_20648 ^ n_20102;
assign n_20663 = n_20648 ^ n_20649;
assign n_20664 = n_20649 ^ n_20102;
assign n_20665 = n_20651 ^ n_20641;
assign n_20666 = n_20652 ^ n_18843;
assign n_20667 = n_20654 ^ n_19974;
assign n_20668 = n_20656 ^ n_18843;
assign n_20669 = n_20656 ^ n_20652;
assign n_20670 = n_20659 ^ n_20660;
assign n_20671 = n_20660 ^ x353;
assign n_20672 = n_20661 ^ n_18741;
assign n_20673 = n_20662 ^ n_20649;
assign n_20674 = n_20663 ^ n_19283;
assign n_20675 = n_20663 & n_20664;
assign n_20676 = n_20665 ^ x282;
assign n_20677 = n_20665 & ~n_20655;
assign n_20678 = n_20667 ^ n_19983;
assign n_20679 = n_20390 ^ n_20667;
assign n_20680 = n_20668 ^ n_20652;
assign n_20681 = n_20666 & n_20669;
assign n_20682 = n_20670 ^ x353;
assign n_20683 = ~n_20670 & n_20671;
assign n_20684 = n_20672 ^ n_18783;
assign n_20685 = n_20674 ^ n_18783;
assign n_20686 = n_20672 ^ n_20674;
assign n_20687 = n_20675 ^ n_20102;
assign n_20688 = n_20676 ^ n_20650;
assign n_20689 = n_20650 & ~n_20676;
assign n_20690 = n_20677 ^ x282;
assign n_20691 = n_20680 ^ x281;
assign n_20692 = n_20681 ^ n_18843;
assign n_20693 = ~n_20657 & n_20682;
assign n_20694 = n_20682 ^ n_20657;
assign n_20695 = n_20683 ^ x353;
assign n_20696 = n_20684 ^ n_20674;
assign n_20697 = ~n_20685 & n_20686;
assign n_20698 = n_20687 ^ n_20121;
assign n_20699 = n_20687 ^ n_20688;
assign n_20700 = n_20688 ^ n_20121;
assign n_20701 = n_20690 ^ n_20680;
assign n_20702 = n_20692 ^ x280;
assign n_20703 = n_20695 ^ n_20696;
assign n_20704 = n_20696 ^ x352;
assign n_20705 = n_20697 ^ n_18783;
assign n_20706 = n_20698 ^ n_20688;
assign n_20707 = n_20699 ^ n_19325;
assign n_20708 = ~n_20699 & ~n_20700;
assign n_20709 = n_20701 ^ x281;
assign n_20710 = n_20701 & ~n_20691;
assign n_20711 = n_20702 ^ n_20678;
assign n_20712 = n_20703 ^ x352;
assign n_20713 = ~n_20703 & n_20704;
assign n_20714 = n_20705 ^ n_18825;
assign n_20715 = n_20707 ^ n_18825;
assign n_20716 = n_20705 ^ n_20707;
assign n_20717 = n_20708 ^ n_20121;
assign n_20718 = n_20709 ^ n_20689;
assign n_20719 = n_20689 & ~n_20709;
assign n_20720 = n_20710 ^ x281;
assign n_20721 = n_20693 & n_20712;
assign n_20722 = n_20712 ^ n_20693;
assign n_20723 = n_20713 ^ x352;
assign n_20724 = n_20714 ^ n_20707;
assign n_20725 = ~n_20715 & n_20716;
assign n_20726 = n_20717 ^ n_20139;
assign n_20727 = n_20717 ^ n_20718;
assign n_20728 = n_20718 ^ n_20139;
assign n_20729 = n_20720 ^ n_20711;
assign n_20730 = n_20723 ^ n_20724;
assign n_20731 = n_20724 ^ x367;
assign n_20732 = n_20725 ^ n_18825;
assign n_20733 = n_20726 ^ n_20718;
assign n_20734 = n_20727 ^ n_19369;
assign n_20735 = n_20727 & ~n_20728;
assign n_20736 = n_20729 ^ n_20719;
assign n_20737 = n_20730 ^ x367;
assign n_20738 = ~n_20730 & n_20731;
assign n_20739 = n_20732 ^ n_18867;
assign n_20740 = n_20734 ^ n_18867;
assign n_20741 = n_20732 ^ n_20734;
assign n_20742 = n_20735 ^ n_20139;
assign n_20743 = n_20736 ^ n_20157;
assign n_20744 = ~n_20721 & ~n_20737;
assign n_20745 = n_20737 ^ n_20721;
assign n_20746 = n_20738 ^ x367;
assign n_20747 = n_20739 ^ n_20734;
assign n_20748 = ~n_20740 & n_20741;
assign n_20749 = n_20742 ^ n_20736;
assign n_20750 = n_20742 ^ n_20157;
assign n_20751 = n_20746 ^ n_20747;
assign n_20752 = n_20747 ^ x366;
assign n_20753 = n_20748 ^ n_18867;
assign n_20754 = ~n_20749 & ~n_20743;
assign n_20755 = n_20749 ^ n_19411;
assign n_20756 = n_20750 ^ n_20736;
assign n_20757 = n_20751 ^ x366;
assign n_20758 = ~n_20751 & n_20752;
assign n_20759 = n_20753 ^ n_18908;
assign n_20760 = n_20754 ^ n_20157;
assign n_20761 = n_20755 ^ n_18908;
assign n_20762 = n_20753 ^ n_20755;
assign n_20763 = n_20757 & ~n_20744;
assign n_20764 = n_20744 ^ n_20757;
assign n_20765 = n_20758 ^ x366;
assign n_20766 = n_20759 ^ n_20755;
assign n_20767 = n_20760 ^ n_19982;
assign n_20768 = n_20183 ^ n_20760;
assign n_20769 = ~n_20761 & n_20762;
assign n_20770 = n_20765 ^ n_20766;
assign n_20771 = n_20766 ^ x365;
assign n_20772 = n_20767 & n_20183;
assign n_20773 = n_20767 ^ n_19452;
assign n_20774 = n_20769 ^ n_18908;
assign n_20775 = n_20770 ^ x365;
assign n_20776 = ~n_20770 & n_20771;
assign n_20777 = n_20772 ^ n_20175;
assign n_20778 = n_20774 ^ n_18943;
assign n_20779 = n_20773 ^ n_20774;
assign n_20780 = n_20763 & n_20775;
assign n_20781 = n_20775 ^ n_20763;
assign n_20782 = n_20776 ^ x365;
assign n_20783 = n_20777 ^ n_20194;
assign n_20784 = n_20773 ^ n_20778;
assign n_20785 = ~n_20778 & n_20779;
assign n_20786 = n_20783 & ~n_20202;
assign n_20787 = n_20022 ^ n_20783;
assign n_20788 = n_20782 ^ n_20784;
assign n_20789 = n_20784 ^ x364;
assign n_20790 = n_20785 ^ n_18943;
assign n_20791 = n_20786 ^ n_20022;
assign n_20792 = n_20787 ^ n_20194;
assign n_20793 = n_20788 ^ x364;
assign n_20794 = n_20788 & ~n_20789;
assign n_20795 = n_20790 ^ n_18968;
assign n_20796 = n_20791 ^ n_20213;
assign n_20797 = n_20792 ^ n_19494;
assign n_20798 = n_20780 & ~n_20793;
assign n_20799 = n_20793 ^ n_20780;
assign n_20800 = n_20794 ^ x364;
assign n_20801 = n_20796 & ~n_20221;
assign n_20802 = n_20048 ^ n_20796;
assign n_20803 = n_20797 ^ n_18968;
assign n_20804 = n_20790 ^ n_20797;
assign n_20805 = n_20795 ^ n_20797;
assign n_20806 = n_20800 ^ x363;
assign n_20807 = n_20801 ^ n_20048;
assign n_20808 = n_20802 ^ n_20213;
assign n_20809 = ~n_20803 & ~n_20804;
assign n_20810 = n_20800 ^ n_20805;
assign n_20811 = n_20807 ^ n_20071;
assign n_20812 = n_20807 ^ n_20232;
assign n_20813 = n_20808 ^ n_19535;
assign n_20814 = n_20809 ^ n_18968;
assign n_20815 = n_20810 & n_20806;
assign n_20816 = n_20810 ^ x363;
assign n_20817 = n_20811 ^ n_20232;
assign n_20818 = n_20811 ^ n_19578;
assign n_20819 = ~n_20240 & ~n_20812;
assign n_20820 = n_20813 ^ n_18991;
assign n_20821 = n_20814 ^ n_20813;
assign n_20822 = n_20814 ^ n_18991;
assign n_20823 = n_20815 ^ x363;
assign n_20824 = n_20798 & ~n_20816;
assign n_20825 = n_20816 ^ n_20798;
assign n_20826 = n_20818 ^ n_19003;
assign n_20827 = n_20819 ^ n_20071;
assign n_20828 = n_20820 & n_20821;
assign n_20829 = n_20822 ^ n_20813;
assign n_20830 = n_20827 ^ n_20250;
assign n_20831 = n_20828 ^ n_18991;
assign n_20832 = n_20823 ^ n_20829;
assign n_20833 = n_20829 ^ x362;
assign n_20834 = ~n_20830 & n_20258;
assign n_20835 = n_20089 ^ n_20830;
assign n_20836 = n_20831 ^ n_20818;
assign n_20837 = n_20831 ^ n_19003;
assign n_20838 = n_20832 ^ x362;
assign n_20839 = n_20832 & ~n_20833;
assign n_20840 = n_20834 ^ n_20089;
assign n_20841 = n_20835 ^ n_20250;
assign n_20842 = n_20826 & n_20836;
assign n_20843 = n_20837 ^ n_20818;
assign n_20844 = ~n_20824 & n_20838;
assign n_20845 = n_20838 ^ n_20824;
assign n_20846 = n_20839 ^ x362;
assign n_20847 = n_20840 ^ n_20269;
assign n_20848 = n_20840 ^ n_20277;
assign n_20849 = n_20841 ^ n_19621;
assign n_20850 = n_20842 ^ n_19003;
assign n_20851 = n_20843 ^ x361;
assign n_20852 = n_20846 ^ n_20843;
assign n_20853 = n_20277 & ~n_20847;
assign n_20854 = n_20848 ^ n_20269;
assign n_20855 = n_20429 ^ n_20848;
assign n_20856 = n_20849 ^ n_19036;
assign n_20857 = n_20850 ^ n_20849;
assign n_20858 = n_20850 ^ n_19036;
assign n_20859 = ~n_20852 & n_20851;
assign n_20860 = n_20852 ^ x361;
assign n_20861 = n_20853 ^ n_20107;
assign n_20862 = n_20854 ^ n_19662;
assign n_20863 = ~n_20856 & ~n_20857;
assign n_20864 = n_20858 ^ n_20849;
assign n_20865 = n_20859 ^ x361;
assign n_20866 = n_20844 & ~n_20860;
assign n_20867 = n_20860 ^ n_20844;
assign n_20868 = n_20861 ^ n_20289;
assign n_20869 = n_20861 ^ n_20125;
assign n_20870 = n_20862 ^ n_19060;
assign n_20871 = n_20863 ^ n_19036;
assign n_20872 = n_20864 ^ x360;
assign n_20873 = n_20865 ^ n_20864;
assign n_20874 = ~n_20297 & ~n_20868;
assign n_20875 = n_20869 ^ n_19700;
assign n_20876 = n_20869 ^ n_20289;
assign n_20877 = n_20871 ^ n_20862;
assign n_20878 = ~n_20873 & n_20872;
assign n_20879 = n_20873 ^ x360;
assign n_20880 = n_20874 ^ n_20125;
assign n_20881 = n_20875 ^ n_19091;
assign n_20882 = n_20876 ^ n_20493;
assign n_20883 = n_20877 & n_20870;
assign n_20884 = n_20877 ^ n_19060;
assign n_20885 = n_20878 ^ x360;
assign n_20886 = ~n_20866 & n_20879;
assign n_20887 = n_20879 ^ n_20866;
assign n_20888 = n_20880 ^ n_20308;
assign n_20889 = n_20883 ^ n_19060;
assign n_20890 = n_20884 ^ x375;
assign n_20891 = n_20885 ^ n_20884;
assign n_20892 = n_20885 ^ x375;
assign n_20893 = ~n_20888 & n_20316;
assign n_20894 = n_20144 ^ n_20888;
assign n_20895 = n_20889 ^ n_20875;
assign n_20896 = n_20890 & ~n_20891;
assign n_20897 = n_20892 ^ n_20884;
assign n_20898 = n_20893 ^ n_20144;
assign n_20899 = n_20894 ^ n_20308;
assign n_20900 = n_20542 ^ n_20894;
assign n_20901 = ~n_20895 & ~n_20881;
assign n_20902 = n_20895 ^ n_19091;
assign n_20903 = n_20896 ^ x375;
assign n_20904 = ~n_20897 & ~n_20886;
assign n_20905 = n_20886 ^ n_20897;
assign n_20906 = n_20898 ^ n_20326;
assign n_20907 = n_20898 ^ n_20162;
assign n_20908 = n_20899 ^ n_19727;
assign n_20909 = n_20901 ^ n_19091;
assign n_20910 = n_20902 ^ x374;
assign n_20911 = n_20903 ^ n_20902;
assign n_20912 = ~n_20905 & ~n_20419;
assign n_20913 = n_20905 ^ n_19971;
assign n_20914 = n_20905 ^ n_19963;
assign n_20915 = n_20419 ^ n_20905;
assign n_20916 = ~n_20334 & ~n_20906;
assign n_20917 = n_20907 ^ n_19749;
assign n_20918 = n_20907 ^ n_20326;
assign n_20919 = n_20908 ^ n_19123;
assign n_20920 = n_20909 ^ n_20908;
assign n_20921 = ~n_20911 & n_20910;
assign n_20922 = n_20911 ^ x374;
assign n_20923 = n_20445 ^ n_20912;
assign n_20924 = n_19014 & n_20913;
assign n_20925 = x455 & n_20914;
assign n_20926 = n_20914 ^ x455;
assign n_20927 = n_20916 ^ n_20162;
assign n_20928 = n_20917 ^ n_19161;
assign n_20929 = n_20580 ^ n_20918;
assign n_20930 = ~n_20920 & ~n_20919;
assign n_20931 = n_20920 ^ n_19123;
assign n_20932 = n_20921 ^ x374;
assign n_20933 = ~n_20904 & n_20922;
assign n_20934 = n_20922 ^ n_20904;
assign n_20935 = n_20924 ^ n_19039;
assign n_20936 = n_20925 ^ x454;
assign n_20937 = n_20927 ^ n_20345;
assign n_20938 = n_20930 ^ n_19123;
assign n_20939 = n_20931 ^ x373;
assign n_20940 = n_20932 ^ n_20931;
assign n_20941 = n_20934 ^ n_20912;
assign n_20942 = n_20934 ^ n_20923;
assign n_20943 = ~n_20937 & ~n_20353;
assign n_20944 = n_20180 ^ n_20937;
assign n_20945 = n_20938 ^ n_20917;
assign n_20946 = n_20938 ^ n_19161;
assign n_20947 = n_20940 & ~n_20939;
assign n_20948 = n_20940 ^ x373;
assign n_20949 = ~n_20923 & n_20941;
assign n_20950 = n_20942 ^ n_20444;
assign n_20951 = n_20943 ^ n_20180;
assign n_20952 = n_20944 ^ n_20345;
assign n_20953 = n_20620 ^ n_20944;
assign n_20954 = n_20928 & ~n_20945;
assign n_20955 = n_20946 ^ n_20917;
assign n_20956 = n_20947 ^ x373;
assign n_20957 = ~n_20933 & n_20948;
assign n_20958 = n_20948 ^ n_20933;
assign n_20959 = n_20949 ^ n_20445;
assign n_20960 = n_20950 ^ n_20924;
assign n_20961 = n_20951 ^ n_20364;
assign n_20962 = n_20952 ^ n_19768;
assign n_20963 = n_20954 ^ n_19161;
assign n_20964 = n_20955 ^ x372;
assign n_20965 = n_20956 ^ n_20955;
assign n_20966 = n_20480 ^ n_20958;
assign n_20967 = n_20959 ^ n_20958;
assign n_20968 = n_20959 ^ n_20480;
assign n_20969 = n_20960 & n_20935;
assign n_20970 = n_20960 ^ n_19039;
assign n_20971 = ~n_20961 & n_20372;
assign n_20972 = n_20199 ^ n_20961;
assign n_20973 = n_20962 ^ n_19198;
assign n_20974 = n_20963 ^ n_20962;
assign n_20975 = n_20963 ^ n_19198;
assign n_20976 = n_20965 & ~n_20964;
assign n_20977 = n_20965 ^ x372;
assign n_20978 = n_20966 & n_20967;
assign n_20979 = n_20968 ^ n_20958;
assign n_20980 = n_20969 ^ n_19039;
assign n_20981 = n_20970 ^ n_20925;
assign n_20982 = n_20970 ^ n_20936;
assign n_20983 = n_20971 ^ n_20199;
assign n_20984 = n_20972 ^ n_20364;
assign n_20985 = n_20658 ^ n_20972;
assign n_20986 = n_20973 & ~n_20974;
assign n_20987 = n_20975 ^ n_20962;
assign n_20988 = n_20976 ^ x372;
assign n_20989 = n_20977 & n_20957;
assign n_20990 = n_20957 ^ n_20977;
assign n_20991 = n_20978 ^ n_20480;
assign n_20992 = n_20979 ^ n_20473;
assign n_20993 = n_20980 ^ n_19076;
assign n_20994 = n_20936 & n_20981;
assign n_20995 = n_20983 ^ n_20384;
assign n_20996 = n_20984 ^ n_19781;
assign n_20997 = n_20986 ^ n_19198;
assign n_20998 = n_20987 ^ x371;
assign n_20999 = n_20988 ^ n_20987;
assign n_21000 = n_20518 ^ n_20990;
assign n_21001 = n_20991 ^ n_20990;
assign n_21002 = n_20991 ^ n_20518;
assign n_21003 = n_20992 ^ n_19076;
assign n_21004 = n_20980 ^ n_20992;
assign n_21005 = n_20993 ^ n_20992;
assign n_21006 = n_20994 ^ x454;
assign n_21007 = ~n_20995 & ~n_20392;
assign n_21008 = n_20218 ^ n_20995;
assign n_21009 = n_20996 ^ n_19238;
assign n_21010 = n_20997 ^ n_20996;
assign n_21011 = n_20997 ^ n_19238;
assign n_21012 = n_20999 & ~n_20998;
assign n_21013 = n_20999 ^ x371;
assign n_21014 = ~n_21000 & n_21001;
assign n_21015 = n_21002 ^ n_20990;
assign n_21016 = ~n_21003 & n_21004;
assign n_21017 = n_21005 ^ x453;
assign n_21018 = n_21006 ^ n_21005;
assign n_21019 = n_21007 ^ n_20218;
assign n_21020 = n_21008 ^ n_20384;
assign n_21021 = n_20694 ^ n_21008;
assign n_21022 = ~n_21009 & ~n_21010;
assign n_21023 = n_21011 ^ n_20996;
assign n_21024 = n_21012 ^ x371;
assign n_21025 = n_21013 & n_20989;
assign n_21026 = n_20989 ^ n_21013;
assign n_21027 = n_21014 ^ n_20518;
assign n_21028 = n_21015 ^ n_20509;
assign n_21029 = n_21016 ^ n_19076;
assign n_21030 = n_21018 & ~n_21017;
assign n_21031 = n_21018 ^ x453;
assign n_21032 = n_21019 ^ n_20403;
assign n_21033 = n_21020 ^ n_19802;
assign n_21034 = n_21022 ^ n_19238;
assign n_21035 = n_21023 ^ x370;
assign n_21036 = n_21024 ^ n_21023;
assign n_21037 = n_20557 ^ n_21026;
assign n_21038 = n_21027 ^ n_21026;
assign n_21039 = n_21027 ^ n_20557;
assign n_21040 = n_21028 ^ n_19116;
assign n_21041 = n_21029 ^ n_21028;
assign n_21042 = n_21029 ^ n_19116;
assign n_21043 = n_21030 ^ x453;
assign n_21044 = n_20237 ^ n_21032;
assign n_21045 = n_21032 & n_20411;
assign n_21046 = n_21033 ^ n_19278;
assign n_21047 = n_21034 ^ n_21033;
assign n_21048 = n_21034 ^ n_19278;
assign n_21049 = ~n_21036 & n_21035;
assign n_21050 = n_21036 ^ x370;
assign n_21051 = n_21037 & n_21038;
assign n_21052 = n_21039 ^ n_21026;
assign n_21053 = ~n_21040 & n_21041;
assign n_21054 = n_21042 ^ n_21028;
assign n_21055 = n_21044 ^ n_20403;
assign n_21056 = n_20722 ^ n_21044;
assign n_21057 = n_21045 ^ n_20237;
assign n_21058 = ~n_21046 & n_21047;
assign n_21059 = n_21048 ^ n_21033;
assign n_21060 = n_21049 ^ x370;
assign n_21061 = n_21050 & ~n_21025;
assign n_21062 = n_21025 ^ n_21050;
assign n_21063 = n_21051 ^ n_20557;
assign n_21064 = n_21052 ^ n_20547;
assign n_21065 = n_21053 ^ n_19116;
assign n_21066 = n_21043 ^ n_21054;
assign n_21067 = n_21054 ^ x452;
assign n_21068 = n_21055 ^ n_19817;
assign n_21069 = n_21057 ^ n_20440;
assign n_21070 = n_21057 ^ n_20430;
assign n_21071 = n_21058 ^ n_19278;
assign n_21072 = n_21059 ^ x369;
assign n_21073 = n_21060 ^ n_21059;
assign n_21074 = n_20595 ^ n_21062;
assign n_21075 = n_21063 ^ n_21062;
assign n_21076 = n_21063 ^ n_20595;
assign n_21077 = n_21064 ^ n_19154;
assign n_21078 = n_21065 ^ n_21064;
assign n_21079 = n_21065 ^ n_19154;
assign n_21080 = n_21066 ^ x452;
assign n_21081 = n_21066 & ~n_21067;
assign n_21082 = n_21068 ^ n_19320;
assign n_21083 = n_21069 ^ n_20430;
assign n_21084 = n_20745 ^ n_21069;
assign n_21085 = n_20440 & ~n_21070;
assign n_21086 = n_21071 ^ n_21068;
assign n_21087 = n_21071 ^ n_19320;
assign n_21088 = n_21073 & ~n_21072;
assign n_21089 = n_21073 ^ x369;
assign n_21090 = ~n_21074 & ~n_21075;
assign n_21091 = n_21076 ^ n_21062;
assign n_21092 = n_21077 & ~n_21078;
assign n_21093 = n_21079 ^ n_21064;
assign n_21094 = n_21031 & n_21080;
assign n_21095 = n_21080 ^ n_21031;
assign n_21096 = n_21081 ^ x452;
assign n_21097 = n_21083 ^ n_19829;
assign n_21098 = n_21085 ^ n_20256;
assign n_21099 = n_21082 & n_21086;
assign n_21100 = n_21087 ^ n_21068;
assign n_21101 = n_21088 ^ x369;
assign n_21102 = n_21061 & ~n_21089;
assign n_21103 = n_21089 ^ n_21061;
assign n_21104 = n_21090 ^ n_20595;
assign n_21105 = n_21091 ^ n_20585;
assign n_21106 = n_21092 ^ n_19154;
assign n_21107 = n_21093 ^ x451;
assign n_21108 = n_21096 ^ n_21093;
assign n_21109 = n_21097 ^ n_19364;
assign n_21110 = n_21098 ^ n_20275;
assign n_21111 = n_21098 ^ n_20456;
assign n_21112 = n_21099 ^ n_19320;
assign n_21113 = n_21100 ^ x368;
assign n_21114 = n_21101 ^ n_21100;
assign n_21115 = n_20634 ^ n_21103;
assign n_21116 = n_21104 ^ n_21103;
assign n_21117 = n_21104 ^ n_20634;
assign n_21118 = n_21105 ^ n_19193;
assign n_21119 = n_21106 ^ n_21105;
assign n_21120 = n_21106 ^ n_19193;
assign n_21121 = ~n_21108 & n_21107;
assign n_21122 = n_21108 ^ x451;
assign n_21123 = n_21110 ^ n_19854;
assign n_21124 = n_21110 ^ n_20456;
assign n_21125 = ~n_20466 & ~n_21111;
assign n_21126 = n_21112 ^ n_21097;
assign n_21127 = ~n_21114 & n_21113;
assign n_21128 = n_21114 ^ x368;
assign n_21129 = ~n_21115 & n_21116;
assign n_21130 = n_21117 ^ n_21103;
assign n_21131 = ~n_21118 & n_21119;
assign n_21132 = n_21120 ^ n_21105;
assign n_21133 = n_21121 ^ x451;
assign n_21134 = ~n_21094 & n_21122;
assign n_21135 = n_21122 ^ n_21094;
assign n_21136 = n_21123 ^ n_19406;
assign n_21137 = n_20764 ^ n_21124;
assign n_21138 = n_21125 ^ n_20275;
assign n_21139 = n_21126 ^ n_19364;
assign n_21140 = n_21126 & n_21109;
assign n_21141 = n_21127 ^ x368;
assign n_21142 = ~n_21128 & ~n_21102;
assign n_21143 = n_21102 ^ n_21128;
assign n_21144 = n_21129 ^ n_20634;
assign n_21145 = n_21130 ^ n_20624;
assign n_21146 = n_21131 ^ n_19193;
assign n_21147 = n_21132 ^ x450;
assign n_21148 = n_21133 ^ n_21132;
assign n_21149 = n_21138 ^ n_20487;
assign n_21150 = n_21139 ^ x383;
assign n_21151 = n_21140 ^ n_19364;
assign n_21152 = n_21141 ^ n_21139;
assign n_21153 = n_21141 ^ x383;
assign n_21154 = n_20673 ^ n_21143;
assign n_21155 = n_21144 ^ n_21143;
assign n_21156 = n_21144 ^ n_20673;
assign n_21157 = n_21145 ^ n_19243;
assign n_21158 = n_21146 ^ n_21145;
assign n_21159 = n_21146 ^ n_19243;
assign n_21160 = n_21148 & ~n_21147;
assign n_21161 = n_21148 ^ x450;
assign n_21162 = n_20295 ^ n_21149;
assign n_21163 = ~n_21149 & ~n_20501;
assign n_21164 = n_21151 ^ n_21123;
assign n_21165 = ~n_21150 & n_21152;
assign n_21166 = n_21153 ^ n_21139;
assign n_21167 = ~n_21154 & n_21155;
assign n_21168 = n_21156 ^ n_21143;
assign n_21169 = ~n_21157 & n_21158;
assign n_21170 = n_21159 ^ n_21145;
assign n_21171 = n_21160 ^ x450;
assign n_21172 = ~n_21161 & n_21134;
assign n_21173 = n_21134 ^ n_21161;
assign n_21174 = n_21162 ^ n_20487;
assign n_21175 = n_20781 ^ n_21162;
assign n_21176 = n_21163 ^ n_20295;
assign n_21177 = n_21164 ^ n_19406;
assign n_21178 = ~n_21164 & n_21136;
assign n_21179 = n_21165 ^ x383;
assign n_21180 = n_21166 & n_21142;
assign n_21181 = n_21142 ^ n_21166;
assign n_21182 = n_21167 ^ n_20673;
assign n_21183 = n_21168 ^ n_20663;
assign n_21184 = n_21169 ^ n_19243;
assign n_21185 = n_21170 ^ x449;
assign n_21186 = n_21171 ^ n_21170;
assign n_21187 = n_21174 ^ n_19874;
assign n_21188 = n_21176 ^ n_20523;
assign n_21189 = n_21177 ^ x382;
assign n_21190 = n_21178 ^ n_19406;
assign n_21191 = n_21179 ^ n_21177;
assign n_21192 = n_20706 ^ n_21181;
assign n_21193 = n_21182 ^ n_21181;
assign n_21194 = n_21182 ^ n_20706;
assign n_21195 = n_21183 ^ n_19283;
assign n_21196 = n_21184 ^ n_21183;
assign n_21197 = n_21184 ^ n_19283;
assign n_21198 = n_21186 & ~n_21185;
assign n_21199 = n_21186 ^ x449;
assign n_21200 = n_21187 ^ n_19447;
assign n_21201 = n_20314 ^ n_21188;
assign n_21202 = ~n_21188 & n_20537;
assign n_21203 = n_21190 ^ n_21187;
assign n_21204 = ~n_21191 & n_21189;
assign n_21205 = n_21191 ^ x382;
assign n_21206 = ~n_21192 & n_21193;
assign n_21207 = n_21194 ^ n_21181;
assign n_21208 = ~n_21195 & ~n_21196;
assign n_21209 = n_21197 ^ n_21183;
assign n_21210 = n_21198 ^ x449;
assign n_21211 = n_21172 & ~n_21199;
assign n_21212 = n_21199 ^ n_21172;
assign n_21213 = n_21201 ^ n_20523;
assign n_21214 = n_20799 ^ n_21201;
assign n_21215 = n_21202 ^ n_20314;
assign n_21216 = n_21203 ^ n_19447;
assign n_21217 = ~n_21203 & ~n_21200;
assign n_21218 = n_21204 ^ x382;
assign n_21219 = ~n_21180 & n_21205;
assign n_21220 = n_21205 ^ n_21180;
assign n_21221 = n_21206 ^ n_20706;
assign n_21222 = n_21207 ^ n_20699;
assign n_21223 = n_21208 ^ n_19283;
assign n_21224 = n_21209 ^ x448;
assign n_21225 = n_21210 ^ n_21209;
assign n_21226 = n_21213 ^ n_19891;
assign n_21227 = n_21215 ^ n_20562;
assign n_21228 = n_21216 ^ x381;
assign n_21229 = n_21217 ^ n_19447;
assign n_21230 = n_21218 ^ n_21216;
assign n_21231 = n_20733 ^ n_21220;
assign n_21232 = n_21221 ^ n_21220;
assign n_21233 = n_21221 ^ n_20733;
assign n_21234 = n_21222 ^ n_19325;
assign n_21235 = n_21223 ^ n_21222;
assign n_21236 = n_21223 ^ n_19325;
assign n_21237 = n_21225 & ~n_21224;
assign n_21238 = n_21225 ^ x448;
assign n_21239 = n_21226 ^ n_19489;
assign n_21240 = n_20332 ^ n_21227;
assign n_21241 = ~n_21227 & ~n_20575;
assign n_21242 = n_21229 ^ n_19489;
assign n_21243 = n_21229 ^ n_21226;
assign n_21244 = n_21230 & ~n_21228;
assign n_21245 = n_21230 ^ x381;
assign n_21246 = n_21231 & n_21232;
assign n_21247 = n_21233 ^ n_21220;
assign n_21248 = ~n_21234 & ~n_21235;
assign n_21249 = n_21236 ^ n_21222;
assign n_21250 = n_21237 ^ x448;
assign n_21251 = n_21211 & ~n_21238;
assign n_21252 = n_21238 ^ n_21211;
assign n_21253 = n_21240 ^ n_20562;
assign n_21254 = n_20825 ^ n_21240;
assign n_21255 = n_21241 ^ n_20332;
assign n_21256 = n_21242 ^ n_21226;
assign n_21257 = ~n_21239 & ~n_21243;
assign n_21258 = n_21244 ^ x381;
assign n_21259 = ~n_21219 & n_21245;
assign n_21260 = n_21245 ^ n_21219;
assign n_21261 = n_21246 ^ n_20733;
assign n_21262 = n_21247 ^ n_20727;
assign n_21263 = n_21248 ^ n_19325;
assign n_21264 = n_21249 ^ x463;
assign n_21265 = n_21250 ^ n_21249;
assign n_21266 = n_21253 ^ n_19910;
assign n_21267 = n_21255 ^ n_20600;
assign n_21268 = n_21256 ^ x380;
assign n_21269 = n_21257 ^ n_19489;
assign n_21270 = n_21258 ^ n_21256;
assign n_21271 = n_20756 ^ n_21260;
assign n_21272 = n_21261 ^ n_21260;
assign n_21273 = n_21261 ^ n_20756;
assign n_21274 = n_21262 ^ n_19369;
assign n_21275 = n_21263 ^ n_21262;
assign n_21276 = n_21263 ^ n_19369;
assign n_21277 = ~n_21265 & n_21264;
assign n_21278 = n_21265 ^ x463;
assign n_21279 = n_21266 ^ n_19531;
assign n_21280 = n_20351 ^ n_21267;
assign n_21281 = n_21267 & ~n_20614;
assign n_21282 = n_21269 ^ n_19531;
assign n_21283 = n_21269 ^ n_21266;
assign n_21284 = ~n_21270 & n_21268;
assign n_21285 = n_21270 ^ x380;
assign n_21286 = ~n_21271 & n_21272;
assign n_21287 = n_21273 ^ n_21260;
assign n_21288 = n_21274 & n_21275;
assign n_21289 = n_21276 ^ n_21262;
assign n_21290 = n_21277 ^ x463;
assign n_21291 = n_21251 & n_21278;
assign n_21292 = n_21280 ^ n_20600;
assign n_21293 = n_20845 ^ n_21280;
assign n_21294 = n_21281 ^ n_20351;
assign n_21295 = n_21282 ^ n_21266;
assign n_21296 = n_21279 & ~n_21283;
assign n_21297 = n_21284 ^ x380;
assign n_21298 = ~n_21285 & n_21259;
assign n_21299 = n_21259 ^ n_21285;
assign n_21300 = n_21286 ^ n_20756;
assign n_21301 = n_21287 ^ n_20749;
assign n_21302 = n_21288 ^ n_19369;
assign n_21303 = n_21289 ^ x462;
assign n_21304 = n_21290 ^ n_21289;
assign n_21305 = n_21292 ^ n_19930;
assign n_21306 = n_21294 ^ n_20639;
assign n_21307 = n_21295 ^ x379;
assign n_21308 = n_21296 ^ n_19531;
assign n_21309 = n_21297 ^ n_21295;
assign n_21310 = n_20768 ^ n_21299;
assign n_21311 = n_21300 ^ n_21299;
assign n_21312 = n_21300 ^ n_20768;
assign n_21313 = n_21301 ^ n_19411;
assign n_21314 = n_21302 ^ n_21301;
assign n_21315 = n_21302 ^ n_19411;
assign n_21316 = ~n_21304 & n_21303;
assign n_21317 = n_21304 ^ x462;
assign n_21318 = n_21305 ^ n_19573;
assign n_21319 = n_21306 ^ n_20370;
assign n_21320 = n_21306 & n_20653;
assign n_21321 = n_21308 ^ n_19573;
assign n_21322 = n_21308 ^ n_21305;
assign n_21323 = ~n_21309 & n_21307;
assign n_21324 = n_21309 ^ x379;
assign n_21325 = ~n_21310 & n_21311;
assign n_21326 = n_21312 ^ n_21299;
assign n_21327 = n_21313 & n_21314;
assign n_21328 = n_21315 ^ n_21301;
assign n_21329 = n_21316 ^ x462;
assign n_21330 = n_21317 & n_21291;
assign n_21331 = n_21291 ^ n_21317;
assign n_21332 = n_21319 ^ n_20639;
assign n_21333 = n_20867 ^ n_21319;
assign n_21334 = n_21320 ^ n_20370;
assign n_21335 = n_21321 ^ n_21305;
assign n_21336 = ~n_21318 & ~n_21322;
assign n_21337 = n_21323 ^ x379;
assign n_21338 = ~n_21298 & n_21324;
assign n_21339 = n_21324 ^ n_21298;
assign n_21340 = n_21325 ^ n_20768;
assign n_21341 = n_21326 ^ n_20767;
assign n_21342 = n_21327 ^ n_19411;
assign n_21343 = n_21328 ^ x461;
assign n_21344 = n_21329 ^ n_21328;
assign n_21345 = n_21331 & n_20915;
assign n_21346 = n_21331 ^ n_20419;
assign n_21347 = n_21331 ^ n_20409;
assign n_21348 = n_20915 ^ n_21331;
assign n_21349 = n_21332 ^ n_19950;
assign n_21350 = n_21334 ^ n_20679;
assign n_21351 = n_21335 ^ x378;
assign n_21352 = n_21336 ^ n_19573;
assign n_21353 = n_21337 ^ n_21335;
assign n_21354 = n_21339 ^ n_20787;
assign n_21355 = n_21340 ^ n_21339;
assign n_21356 = n_21340 ^ n_20787;
assign n_21357 = n_21341 ^ n_19452;
assign n_21358 = n_21342 ^ n_21341;
assign n_21359 = n_21342 ^ n_19452;
assign n_21360 = n_21344 & ~n_21343;
assign n_21361 = n_21344 ^ x461;
assign n_21362 = n_21345 ^ n_20942;
assign n_21363 = ~n_19971 & ~n_21346;
assign n_21364 = x39 & n_21347;
assign n_21365 = n_21347 ^ x39;
assign n_21366 = n_21349 ^ n_19615;
assign n_21367 = n_21350 ^ n_20667;
assign n_21368 = n_21352 ^ n_19615;
assign n_21369 = n_21352 ^ n_21349;
assign n_21370 = n_21353 & ~n_21351;
assign n_21371 = n_21353 ^ x378;
assign n_21372 = n_21354 & ~n_21355;
assign n_21373 = n_21356 ^ n_21339;
assign n_21374 = n_21357 & n_21358;
assign n_21375 = n_21359 ^ n_21341;
assign n_21376 = n_21360 ^ x461;
assign n_21377 = n_21330 & ~n_21361;
assign n_21378 = n_21361 ^ n_21330;
assign n_21379 = n_21363 ^ n_19996;
assign n_21380 = n_21364 ^ x38;
assign n_21381 = n_21367 ^ n_19965;
assign n_21382 = n_21368 ^ n_21349;
assign n_21383 = ~n_21366 & ~n_21369;
assign n_21384 = n_21370 ^ x378;
assign n_21385 = ~n_21338 & n_21371;
assign n_21386 = n_21371 ^ n_21338;
assign n_21387 = n_21372 ^ n_20787;
assign n_21388 = n_21373 ^ n_20792;
assign n_21389 = n_21374 ^ n_19452;
assign n_21390 = n_21375 ^ x460;
assign n_21391 = n_21376 ^ n_21375;
assign n_21392 = n_21378 ^ n_21345;
assign n_21393 = n_21362 ^ n_21378;
assign n_21394 = n_21381 ^ n_19644;
assign n_21395 = n_21382 ^ x377;
assign n_21396 = n_21383 ^ n_19615;
assign n_21397 = n_21384 ^ n_21382;
assign n_21398 = n_21386 ^ n_20802;
assign n_21399 = n_21387 ^ n_21386;
assign n_21400 = n_21387 ^ n_20802;
assign n_21401 = n_21388 ^ n_19494;
assign n_21402 = n_21389 ^ n_21388;
assign n_21403 = n_21389 ^ n_19494;
assign n_21404 = ~n_21391 & n_21390;
assign n_21405 = n_21391 ^ x460;
assign n_21406 = n_21392 & n_21362;
assign n_21407 = n_21392 ^ n_20445;
assign n_21408 = n_21396 ^ x376;
assign n_21409 = n_21397 ^ x377;
assign n_21410 = ~n_21397 & n_21395;
assign n_21411 = ~n_21398 & n_21399;
assign n_21412 = n_21400 ^ n_21386;
assign n_21413 = ~n_21401 & ~n_21402;
assign n_21414 = n_21403 ^ n_21388;
assign n_21415 = n_21404 ^ x460;
assign n_21416 = ~n_21377 & ~n_21405;
assign n_21417 = n_21405 ^ n_21377;
assign n_21418 = n_21406 ^ n_20942;
assign n_21419 = n_21407 ^ n_21363;
assign n_21420 = n_21408 ^ n_21394;
assign n_21421 = n_21409 ^ n_21385;
assign n_21422 = n_21385 & ~n_21409;
assign n_21423 = n_21410 ^ x377;
assign n_21424 = n_21411 ^ n_20802;
assign n_21425 = n_21412 ^ n_20808;
assign n_21426 = n_21413 ^ n_19494;
assign n_21427 = n_21414 ^ x459;
assign n_21428 = n_21415 ^ n_21414;
assign n_21429 = n_21417 ^ n_20979;
assign n_21430 = n_21418 ^ n_21417;
assign n_21431 = n_21418 ^ n_20979;
assign n_21432 = ~n_21419 & n_21379;
assign n_21433 = n_21419 ^ n_19996;
assign n_21434 = n_20817 ^ n_21421;
assign n_21435 = n_21423 ^ n_21420;
assign n_21436 = n_21424 ^ n_21421;
assign n_21437 = n_21424 ^ n_20817;
assign n_21438 = n_21425 ^ n_19535;
assign n_21439 = n_21426 ^ n_21425;
assign n_21440 = n_21426 ^ n_19535;
assign n_21441 = ~n_21428 & n_21427;
assign n_21442 = n_21428 ^ x459;
assign n_21443 = n_21430 & n_21429;
assign n_21444 = n_21430 ^ n_20480;
assign n_21445 = n_21431 ^ n_21417;
assign n_21446 = n_21432 ^ n_19996;
assign n_21447 = n_21364 ^ n_21433;
assign n_21448 = n_21380 ^ n_21433;
assign n_21449 = n_21435 ^ n_21422;
assign n_21450 = ~n_21434 & n_21436;
assign n_21451 = n_21437 ^ n_21421;
assign n_21452 = n_21438 & ~n_21439;
assign n_21453 = n_21440 ^ n_21425;
assign n_21454 = n_21441 ^ x459;
assign n_21455 = ~n_21442 & n_21416;
assign n_21456 = n_21416 ^ n_21442;
assign n_21457 = n_21443 ^ n_20979;
assign n_21458 = n_21444 ^ n_20018;
assign n_21459 = n_21446 ^ n_21444;
assign n_21460 = n_21446 ^ n_20018;
assign n_21461 = n_21380 & ~n_21447;
assign n_21462 = n_21449 ^ n_20835;
assign n_21463 = n_21450 ^ n_20817;
assign n_21464 = n_21451 ^ n_20811;
assign n_21465 = n_21452 ^ n_19535;
assign n_21466 = n_21453 ^ x458;
assign n_21467 = n_21454 ^ n_21453;
assign n_21468 = n_21456 ^ n_21015;
assign n_21469 = n_21456 ^ n_21457;
assign n_21470 = n_21457 ^ n_21015;
assign n_21471 = ~n_21458 & n_21459;
assign n_21472 = n_21460 ^ n_21444;
assign n_21473 = n_21461 ^ x38;
assign n_21474 = n_21463 ^ n_20835;
assign n_21475 = n_21463 ^ n_21449;
assign n_21476 = n_21464 ^ n_19578;
assign n_21477 = n_21465 ^ n_21464;
assign n_21478 = n_21465 ^ n_19578;
assign n_21479 = ~n_21467 & n_21466;
assign n_21480 = n_21467 ^ x458;
assign n_21481 = n_21469 & ~n_21468;
assign n_21482 = n_21469 ^ n_20518;
assign n_21483 = n_21470 ^ n_21456;
assign n_21484 = n_21471 ^ n_20018;
assign n_21485 = n_21472 ^ x37;
assign n_21486 = n_21473 ^ n_21472;
assign n_21487 = n_21474 ^ n_21449;
assign n_21488 = n_21462 & ~n_21475;
assign n_21489 = ~n_21476 & n_21477;
assign n_21490 = n_21478 ^ n_21464;
assign n_21491 = n_21479 ^ x458;
assign n_21492 = n_21455 & ~n_21480;
assign n_21493 = n_21480 ^ n_21455;
assign n_21494 = n_21481 ^ n_21015;
assign n_21495 = n_21482 ^ n_20034;
assign n_21496 = n_21484 ^ n_21482;
assign n_21497 = n_21484 ^ n_20034;
assign n_21498 = n_21486 & ~n_21485;
assign n_21499 = n_21486 ^ x37;
assign n_21500 = n_21487 ^ n_20841;
assign n_21501 = n_21488 ^ n_20835;
assign n_21502 = n_21489 ^ n_19578;
assign n_21503 = n_21490 ^ x457;
assign n_21504 = n_21491 ^ n_21490;
assign n_21505 = n_21493 ^ n_21052;
assign n_21506 = n_21494 ^ n_21493;
assign n_21507 = n_21494 ^ n_21052;
assign n_21508 = ~n_21495 & n_21496;
assign n_21509 = n_21497 ^ n_21482;
assign n_21510 = n_21498 ^ x37;
assign n_21511 = n_21500 ^ n_19621;
assign n_21512 = n_21501 ^ n_20855;
assign n_21513 = n_21501 ^ n_20848;
assign n_21514 = n_21502 ^ n_21500;
assign n_21515 = n_21502 ^ n_19621;
assign n_21516 = n_21504 & ~n_21503;
assign n_21517 = n_21504 ^ x457;
assign n_21518 = n_21506 & n_21505;
assign n_21519 = n_21506 ^ n_20557;
assign n_21520 = n_21507 ^ n_21493;
assign n_21521 = n_21508 ^ n_20034;
assign n_21522 = n_21509 ^ x36;
assign n_21523 = n_21510 ^ n_21509;
assign n_21524 = n_21512 ^ n_20854;
assign n_21525 = ~n_20855 & ~n_21513;
assign n_21526 = n_21511 & n_21514;
assign n_21527 = n_21515 ^ n_21500;
assign n_21528 = n_21516 ^ x457;
assign n_21529 = ~n_21492 & ~n_21517;
assign n_21530 = n_21517 ^ n_21492;
assign n_21531 = n_21518 ^ n_21052;
assign n_21532 = n_21519 ^ n_20051;
assign n_21533 = n_21365 ^ n_21520;
assign n_21534 = n_21521 ^ n_21519;
assign n_21535 = n_21521 ^ n_20051;
assign n_21536 = n_21523 & ~n_21522;
assign n_21537 = n_21523 ^ x36;
assign n_21538 = n_21524 ^ n_19662;
assign n_21539 = n_21525 ^ n_20429;
assign n_21540 = n_21526 ^ n_19621;
assign n_21541 = n_21527 ^ x456;
assign n_21542 = n_21528 ^ n_21527;
assign n_21543 = n_21530 ^ n_21091;
assign n_21544 = n_21531 ^ n_21530;
assign n_21545 = n_21531 ^ n_21091;
assign n_21546 = ~n_21532 & ~n_21534;
assign n_21547 = n_21535 ^ n_21519;
assign n_21548 = n_21536 ^ x36;
assign n_21549 = ~n_21499 & ~n_21537;
assign n_21550 = n_21537 ^ n_21499;
assign n_21551 = n_21539 ^ n_20493;
assign n_21552 = n_21539 ^ n_20876;
assign n_21553 = n_21540 ^ n_21524;
assign n_21554 = ~n_21542 & n_21541;
assign n_21555 = n_21542 ^ x456;
assign n_21556 = ~n_21544 & n_21543;
assign n_21557 = n_21544 ^ n_20595;
assign n_21558 = n_21545 ^ n_21530;
assign n_21559 = n_21546 ^ n_20051;
assign n_21560 = n_21547 ^ x35;
assign n_21561 = n_21548 ^ n_21547;
assign n_21562 = n_21551 ^ n_20876;
assign n_21563 = ~n_20882 & ~n_21552;
assign n_21564 = n_21553 ^ n_19662;
assign n_21565 = n_21553 & ~n_21538;
assign n_21566 = n_21554 ^ x456;
assign n_21567 = n_21529 & n_21555;
assign n_21568 = n_21555 ^ n_21529;
assign n_21569 = n_21556 ^ n_21091;
assign n_21570 = n_21557 ^ n_20067;
assign n_21571 = n_21558 ^ n_21448;
assign n_21572 = n_21559 ^ n_21557;
assign n_21573 = n_21559 ^ n_20067;
assign n_21574 = n_21561 & ~n_21560;
assign n_21575 = n_21561 ^ x35;
assign n_21576 = n_21562 ^ n_20869;
assign n_21577 = n_21563 ^ n_20493;
assign n_21578 = n_21564 ^ x471;
assign n_21579 = n_21565 ^ n_19662;
assign n_21580 = n_21566 ^ n_21564;
assign n_21581 = n_21566 ^ x471;
assign n_21582 = n_21568 ^ n_21130;
assign n_21583 = n_21568 ^ n_21569;
assign n_21584 = n_21569 ^ n_21130;
assign n_21585 = ~n_21570 & n_21572;
assign n_21586 = n_21573 ^ n_21557;
assign n_21587 = n_21574 ^ x35;
assign n_21588 = n_21549 & ~n_21575;
assign n_21589 = n_21575 ^ n_21549;
assign n_21590 = n_21576 ^ n_19700;
assign n_21591 = n_21577 ^ n_20542;
assign n_21592 = n_21577 ^ n_20894;
assign n_21593 = n_21579 ^ n_21576;
assign n_21594 = n_21578 & ~n_21580;
assign n_21595 = n_21581 ^ n_21564;
assign n_21596 = ~n_21583 & ~n_21582;
assign n_21597 = n_21583 ^ n_20634;
assign n_21598 = n_21584 ^ n_21568;
assign n_21599 = n_21585 ^ n_20067;
assign n_21600 = n_21586 ^ x34;
assign n_21601 = n_21587 ^ n_21586;
assign n_21602 = n_21591 ^ n_20894;
assign n_21603 = n_20900 & n_21592;
assign n_21604 = n_21593 ^ n_19700;
assign n_21605 = n_21593 & n_21590;
assign n_21606 = n_21594 ^ x471;
assign n_21607 = ~n_21567 & ~n_21595;
assign n_21608 = n_21595 ^ n_21567;
assign n_21609 = n_21596 ^ n_21130;
assign n_21610 = n_21597 ^ n_20084;
assign n_21611 = n_21598 ^ n_21499;
assign n_21612 = n_21599 ^ n_21597;
assign n_21613 = n_21599 ^ n_20084;
assign n_21614 = ~n_21601 & n_21600;
assign n_21615 = n_21601 ^ x34;
assign n_21616 = n_21602 ^ n_20899;
assign n_21617 = n_21603 ^ n_20542;
assign n_21618 = n_21604 ^ x470;
assign n_21619 = n_21605 ^ n_19700;
assign n_21620 = n_21606 ^ n_21604;
assign n_21621 = n_21608 ^ n_21168;
assign n_21622 = n_21609 ^ n_21608;
assign n_21623 = n_21609 ^ n_21168;
assign n_21624 = n_21610 & n_21612;
assign n_21625 = n_21613 ^ n_21597;
assign n_21626 = n_21614 ^ x34;
assign n_21627 = n_21588 & n_21615;
assign n_21628 = n_21615 ^ n_21588;
assign n_21629 = n_21616 ^ n_19727;
assign n_21630 = n_21617 ^ n_20918;
assign n_21631 = n_21619 ^ n_21616;
assign n_21632 = n_21620 & ~n_21618;
assign n_21633 = n_21620 ^ x470;
assign n_21634 = ~n_21622 & n_21621;
assign n_21635 = n_21622 ^ n_20673;
assign n_21636 = n_21623 ^ n_21608;
assign n_21637 = n_21624 ^ n_20084;
assign n_21638 = n_21625 ^ x33;
assign n_21639 = n_21626 ^ n_21625;
assign n_21640 = n_20580 ^ n_21630;
assign n_21641 = n_21630 & ~n_20929;
assign n_21642 = n_21631 ^ n_19727;
assign n_21643 = n_21631 & ~n_21629;
assign n_21644 = n_21632 ^ x470;
assign n_21645 = ~n_21607 & ~n_21633;
assign n_21646 = n_21633 ^ n_21607;
assign n_21647 = n_21634 ^ n_21168;
assign n_21648 = n_21635 ^ n_20102;
assign n_21649 = n_21550 ^ n_21636;
assign n_21650 = n_21637 ^ n_21635;
assign n_21651 = n_21637 ^ n_20102;
assign n_21652 = n_21639 & ~n_21638;
assign n_21653 = n_21639 ^ x33;
assign n_21654 = n_21640 ^ n_20907;
assign n_21655 = n_21641 ^ n_20580;
assign n_21656 = n_21642 ^ x469;
assign n_21657 = n_21643 ^ n_19727;
assign n_21658 = n_21644 ^ n_21642;
assign n_21659 = n_21646 ^ n_21207;
assign n_21660 = n_21647 ^ n_21646;
assign n_21661 = n_21647 ^ n_21207;
assign n_21662 = ~n_21648 & ~n_21650;
assign n_21663 = n_21651 ^ n_21635;
assign n_21664 = n_21652 ^ x33;
assign n_21665 = ~n_21627 & n_21653;
assign n_21666 = n_21653 ^ n_21627;
assign n_21667 = n_21654 ^ n_19749;
assign n_21668 = n_21655 ^ n_20620;
assign n_21669 = n_21655 ^ n_20944;
assign n_21670 = n_21657 ^ n_19749;
assign n_21671 = n_21657 ^ n_21654;
assign n_21672 = n_21658 & ~n_21656;
assign n_21673 = n_21658 ^ x469;
assign n_21674 = n_21660 & ~n_21659;
assign n_21675 = n_21660 ^ n_20706;
assign n_21676 = n_21661 ^ n_21646;
assign n_21677 = n_21662 ^ n_20102;
assign n_21678 = n_21663 ^ x32;
assign n_21679 = n_21664 ^ n_21663;
assign n_21680 = n_21668 ^ n_20944;
assign n_21681 = ~n_20953 & ~n_21669;
assign n_21682 = n_21670 ^ n_21654;
assign n_21683 = n_21667 & ~n_21671;
assign n_21684 = n_21672 ^ x469;
assign n_21685 = ~n_21645 & n_21673;
assign n_21686 = n_21673 ^ n_21645;
assign n_21687 = n_21674 ^ n_21207;
assign n_21688 = n_21675 ^ n_20121;
assign n_21689 = n_21589 ^ n_21676;
assign n_21690 = n_21677 ^ n_21675;
assign n_21691 = n_21677 ^ n_20121;
assign n_21692 = n_21679 & ~n_21678;
assign n_21693 = n_21679 ^ x32;
assign n_21694 = n_21680 ^ n_20952;
assign n_21695 = n_21681 ^ n_20620;
assign n_21696 = n_21682 ^ x468;
assign n_21697 = n_21683 ^ n_19749;
assign n_21698 = n_21684 ^ n_21682;
assign n_21699 = n_21686 ^ n_21247;
assign n_21700 = n_21686 ^ n_21687;
assign n_21701 = n_21687 ^ n_21247;
assign n_21702 = ~n_21688 & ~n_21690;
assign n_21703 = n_21691 ^ n_21675;
assign n_21704 = n_21692 ^ x32;
assign n_21705 = ~n_21665 & ~n_21693;
assign n_21706 = n_21693 ^ n_21665;
assign n_21707 = n_21694 ^ n_19768;
assign n_21708 = n_21695 ^ n_20972;
assign n_21709 = n_21697 ^ n_19768;
assign n_21710 = n_21697 ^ n_21694;
assign n_21711 = ~n_21698 & n_21696;
assign n_21712 = n_21698 ^ x468;
assign n_21713 = n_21700 & n_21699;
assign n_21714 = n_21700 ^ n_20733;
assign n_21715 = n_21701 ^ n_21686;
assign n_21716 = n_21702 ^ n_20121;
assign n_21717 = n_21703 ^ x47;
assign n_21718 = n_21704 ^ n_21703;
assign n_21719 = n_20658 ^ n_21708;
assign n_21720 = n_21708 & ~n_20985;
assign n_21721 = n_21709 ^ n_21694;
assign n_21722 = n_21707 & ~n_21710;
assign n_21723 = n_21711 ^ x468;
assign n_21724 = ~n_21685 & n_21712;
assign n_21725 = n_21712 ^ n_21685;
assign n_21726 = n_21713 ^ n_21247;
assign n_21727 = n_21714 ^ n_20139;
assign n_21728 = n_21628 ^ n_21715;
assign n_21729 = n_21716 ^ n_21714;
assign n_21730 = n_21716 ^ n_20139;
assign n_21731 = ~n_21718 & n_21717;
assign n_21732 = n_21718 ^ x47;
assign n_21733 = n_21719 ^ n_20984;
assign n_21734 = n_21720 ^ n_20658;
assign n_21735 = n_21721 ^ x467;
assign n_21736 = n_21722 ^ n_19768;
assign n_21737 = n_21723 ^ n_21721;
assign n_21738 = n_21725 ^ n_21287;
assign n_21739 = n_21726 ^ n_21725;
assign n_21740 = n_21726 ^ n_21287;
assign n_21741 = n_21727 & ~n_21729;
assign n_21742 = n_21730 ^ n_21714;
assign n_21743 = n_21731 ^ x47;
assign n_21744 = n_21705 & n_21732;
assign n_21745 = n_21732 ^ n_21705;
assign n_21746 = n_21733 ^ n_19781;
assign n_21747 = n_21734 ^ n_21008;
assign n_21748 = n_21736 ^ n_19781;
assign n_21749 = n_21736 ^ n_21733;
assign n_21750 = ~n_21737 & n_21735;
assign n_21751 = n_21737 ^ x467;
assign n_21752 = n_21739 & ~n_21738;
assign n_21753 = n_21739 ^ n_20756;
assign n_21754 = n_21740 ^ n_21725;
assign n_21755 = n_21741 ^ n_20139;
assign n_21756 = n_21742 ^ x46;
assign n_21757 = n_21743 ^ n_21742;
assign n_21758 = n_20694 ^ n_21747;
assign n_21759 = ~n_21747 & n_21021;
assign n_21760 = n_21748 ^ n_21733;
assign n_21761 = ~n_21746 & ~n_21749;
assign n_21762 = n_21750 ^ x467;
assign n_21763 = n_21724 & n_21751;
assign n_21764 = n_21751 ^ n_21724;
assign n_21765 = n_21752 ^ n_21287;
assign n_21766 = n_21753 ^ n_20157;
assign n_21767 = n_21666 ^ n_21754;
assign n_21768 = n_21755 ^ n_21753;
assign n_21769 = n_21755 ^ n_20157;
assign n_21770 = ~n_21757 & n_21756;
assign n_21771 = n_21757 ^ x46;
assign n_21772 = n_21758 ^ n_21020;
assign n_21773 = n_21759 ^ n_20694;
assign n_21774 = n_21760 ^ x466;
assign n_21775 = n_21761 ^ n_19781;
assign n_21776 = n_21762 ^ n_21760;
assign n_21777 = n_21764 ^ n_21326;
assign n_21778 = n_21765 ^ n_21764;
assign n_21779 = n_21765 ^ n_21326;
assign n_21780 = ~n_21766 & ~n_21768;
assign n_21781 = n_21769 ^ n_21753;
assign n_21782 = n_21770 ^ x46;
assign n_21783 = ~n_21744 & ~n_21771;
assign n_21784 = n_21771 ^ n_21744;
assign n_21785 = n_21772 ^ n_19802;
assign n_21786 = n_21773 ^ n_21044;
assign n_21787 = n_21775 ^ n_19802;
assign n_21788 = n_21775 ^ n_21772;
assign n_21789 = n_21776 & ~n_21774;
assign n_21790 = n_21776 ^ x466;
assign n_21791 = ~n_21778 & n_21777;
assign n_21792 = n_21778 ^ n_20768;
assign n_21793 = n_21779 ^ n_21764;
assign n_21794 = n_21780 ^ n_20157;
assign n_21795 = n_21781 ^ x45;
assign n_21796 = n_21782 ^ n_21781;
assign n_21797 = n_20722 ^ n_21786;
assign n_21798 = ~n_21786 & ~n_21056;
assign n_21799 = n_21787 ^ n_21772;
assign n_21800 = n_21785 & n_21788;
assign n_21801 = n_21789 ^ x466;
assign n_21802 = ~n_21763 & n_21790;
assign n_21803 = n_21790 ^ n_21763;
assign n_21804 = n_21791 ^ n_21326;
assign n_21805 = n_21792 ^ n_20175;
assign n_21806 = n_21706 ^ n_21793;
assign n_21807 = n_21794 ^ n_21792;
assign n_21808 = n_21794 ^ n_20175;
assign n_21809 = n_21796 & ~n_21795;
assign n_21810 = n_21796 ^ x45;
assign n_21811 = n_21797 ^ n_21055;
assign n_21812 = n_20926 ^ n_21797;
assign n_21813 = n_21798 ^ n_20722;
assign n_21814 = n_21799 ^ x465;
assign n_21815 = n_21800 ^ n_19802;
assign n_21816 = n_21801 ^ n_21799;
assign n_21817 = n_21803 ^ n_21373;
assign n_21818 = n_21804 ^ n_21803;
assign n_21819 = n_21804 ^ n_21373;
assign n_21820 = ~n_21805 & ~n_21807;
assign n_21821 = n_21808 ^ n_21792;
assign n_21822 = n_21809 ^ x45;
assign n_21823 = ~n_21783 & ~n_21810;
assign n_21824 = n_21810 ^ n_21783;
assign n_21825 = n_21811 ^ n_19817;
assign n_21826 = n_21813 ^ n_21069;
assign n_21827 = n_21815 ^ n_19817;
assign n_21828 = n_21815 ^ n_21811;
assign n_21829 = n_21816 & ~n_21814;
assign n_21830 = n_21816 ^ x465;
assign n_21831 = ~n_21817 & ~n_21818;
assign n_21832 = n_21818 ^ n_20787;
assign n_21833 = n_21819 ^ n_21803;
assign n_21834 = n_21820 ^ n_20175;
assign n_21835 = n_21821 ^ x44;
assign n_21836 = n_21822 ^ n_21821;
assign n_21837 = n_20745 ^ n_21826;
assign n_21838 = ~n_21826 & ~n_21084;
assign n_21839 = n_21827 ^ n_21811;
assign n_21840 = ~n_21825 & n_21828;
assign n_21841 = n_21829 ^ x465;
assign n_21842 = n_21802 & n_21830;
assign n_21843 = n_21830 ^ n_21802;
assign n_21844 = n_21831 ^ n_21373;
assign n_21845 = n_21832 ^ n_20194;
assign n_21846 = n_21745 ^ n_21833;
assign n_21847 = n_21834 ^ n_21832;
assign n_21848 = n_21834 ^ n_20194;
assign n_21849 = ~n_21836 & n_21835;
assign n_21850 = n_21836 ^ x44;
assign n_21851 = n_21837 ^ n_21083;
assign n_21852 = n_20982 ^ n_21837;
assign n_21853 = n_21838 ^ n_20745;
assign n_21854 = n_21839 ^ x464;
assign n_21855 = n_21840 ^ n_19817;
assign n_21856 = n_21841 ^ n_21839;
assign n_21857 = n_21843 ^ n_21412;
assign n_21858 = n_21844 ^ n_21843;
assign n_21859 = n_21844 ^ n_21412;
assign n_21860 = n_21845 & n_21847;
assign n_21861 = n_21848 ^ n_21832;
assign n_21862 = n_21849 ^ x44;
assign n_21863 = ~n_21823 & ~n_21850;
assign n_21864 = n_21850 ^ n_21823;
assign n_21865 = n_21851 ^ n_19829;
assign n_21866 = n_21853 ^ n_20764;
assign n_21867 = n_21853 ^ n_21124;
assign n_21868 = n_21855 ^ n_21851;
assign n_21869 = n_21856 ^ x464;
assign n_21870 = n_21856 & ~n_21854;
assign n_21871 = ~n_21857 & ~n_21858;
assign n_21872 = n_21858 ^ n_20802;
assign n_21873 = n_21859 ^ n_21843;
assign n_21874 = n_21860 ^ n_20194;
assign n_21875 = n_21861 ^ x43;
assign n_21876 = n_21862 ^ n_21861;
assign n_21877 = n_21866 ^ n_21124;
assign n_21878 = n_21137 & ~n_21867;
assign n_21879 = n_21868 ^ n_19829;
assign n_21880 = n_21868 & ~n_21865;
assign n_21881 = n_21869 ^ n_21842;
assign n_21882 = n_21842 & n_21869;
assign n_21883 = n_21870 ^ x464;
assign n_21884 = n_21871 ^ n_21412;
assign n_21885 = n_21872 ^ n_20213;
assign n_21886 = n_21784 ^ n_21873;
assign n_21887 = n_21874 ^ n_21872;
assign n_21888 = n_21874 ^ n_20213;
assign n_21889 = ~n_21876 & n_21875;
assign n_21890 = n_21876 ^ x43;
assign n_21891 = n_21877 ^ n_21110;
assign n_21892 = n_21877 ^ n_21031;
assign n_21893 = n_21878 ^ n_20764;
assign n_21894 = n_21879 ^ x479;
assign n_21895 = n_21880 ^ n_19829;
assign n_21896 = n_21881 ^ n_21451;
assign n_21897 = n_21883 ^ x479;
assign n_21898 = n_21883 ^ n_21879;
assign n_21899 = n_21884 ^ n_21881;
assign n_21900 = n_21884 ^ n_21451;
assign n_21901 = n_21885 & ~n_21887;
assign n_21902 = n_21888 ^ n_21872;
assign n_21903 = n_21889 ^ x43;
assign n_21904 = ~n_21863 & n_21890;
assign n_21905 = n_21890 ^ n_21863;
assign n_21906 = n_21891 ^ n_19854;
assign n_21907 = n_21893 ^ n_21162;
assign n_21908 = n_21895 ^ n_21891;
assign n_21909 = n_21897 ^ n_21879;
assign n_21910 = ~n_21894 & n_21898;
assign n_21911 = ~n_21896 & n_21899;
assign n_21912 = n_21899 ^ n_20817;
assign n_21913 = n_21900 ^ n_21881;
assign n_21914 = n_21901 ^ n_20213;
assign n_21915 = n_21902 ^ x42;
assign n_21916 = n_21903 ^ n_21902;
assign n_21917 = n_20781 ^ n_21907;
assign n_21918 = n_21907 & n_21175;
assign n_21919 = n_21908 ^ n_19854;
assign n_21920 = ~n_21908 & ~n_21906;
assign n_21921 = n_21909 ^ n_21882;
assign n_21922 = n_21882 & n_21909;
assign n_21923 = n_21910 ^ x479;
assign n_21924 = n_21911 ^ n_21451;
assign n_21925 = n_21912 ^ n_20232;
assign n_21926 = n_21824 ^ n_21913;
assign n_21927 = n_21914 ^ n_21912;
assign n_21928 = n_21914 ^ n_20232;
assign n_21929 = n_21916 & ~n_21915;
assign n_21930 = n_21916 ^ x42;
assign n_21931 = n_21917 ^ n_21174;
assign n_21932 = n_21095 ^ n_21917;
assign n_21933 = n_21918 ^ n_20781;
assign n_21934 = n_21919 ^ x478;
assign n_21935 = n_21920 ^ n_19854;
assign n_21936 = n_21921 ^ n_21487;
assign n_21937 = n_21923 ^ n_21919;
assign n_21938 = n_21924 ^ n_21921;
assign n_21939 = n_21924 ^ n_21487;
assign n_21940 = n_21925 & n_21927;
assign n_21941 = n_21928 ^ n_21912;
assign n_21942 = n_21929 ^ x42;
assign n_21943 = n_21930 & ~n_21904;
assign n_21944 = n_21904 ^ n_21930;
assign n_21945 = n_21931 ^ n_19874;
assign n_21946 = n_21933 ^ n_21201;
assign n_21947 = n_21935 ^ n_21931;
assign n_21948 = n_21937 ^ x478;
assign n_21949 = n_21937 & ~n_21934;
assign n_21950 = n_21938 ^ n_20835;
assign n_21951 = n_21938 & n_21936;
assign n_21952 = n_21939 ^ n_21921;
assign n_21953 = n_21940 ^ n_20232;
assign n_21954 = n_21941 ^ x41;
assign n_21955 = n_21942 ^ n_21941;
assign n_21956 = n_20799 ^ n_21946;
assign n_21957 = ~n_21946 & ~n_21214;
assign n_21958 = n_21947 ^ n_19874;
assign n_21959 = n_21947 & ~n_21945;
assign n_21960 = n_21948 ^ n_21922;
assign n_21961 = ~n_21922 & ~n_21948;
assign n_21962 = n_21949 ^ x478;
assign n_21963 = n_21950 ^ n_20250;
assign n_21964 = n_21951 ^ n_21487;
assign n_21965 = n_21864 ^ n_21952;
assign n_21966 = n_21953 ^ n_21950;
assign n_21967 = n_21953 ^ n_20250;
assign n_21968 = n_21955 & ~n_21954;
assign n_21969 = n_21955 ^ x41;
assign n_21970 = n_21956 ^ n_21213;
assign n_21971 = n_21135 ^ n_21956;
assign n_21972 = n_21957 ^ n_20799;
assign n_21973 = n_21958 ^ x477;
assign n_21974 = n_21959 ^ n_19874;
assign n_21975 = n_21960 ^ n_21512;
assign n_21976 = n_21962 ^ n_21958;
assign n_21977 = n_21964 ^ n_21960;
assign n_21978 = ~n_21963 & ~n_21966;
assign n_21979 = n_21967 ^ n_21950;
assign n_21980 = n_21968 ^ x41;
assign n_21981 = n_21943 & n_21969;
assign n_21982 = n_21969 ^ n_21943;
assign n_21983 = n_21970 ^ n_19891;
assign n_21984 = n_21972 ^ n_21240;
assign n_21985 = n_21974 ^ n_19891;
assign n_21986 = n_21974 ^ n_21970;
assign n_21987 = n_21975 ^ n_21964;
assign n_21988 = n_21976 ^ x477;
assign n_21989 = ~n_21976 & n_21973;
assign n_21990 = n_21977 ^ n_20848;
assign n_21991 = n_21977 & n_21975;
assign n_21992 = n_21978 ^ n_20250;
assign n_21993 = n_21979 ^ x40;
assign n_21994 = n_21980 ^ n_21979;
assign n_21995 = n_20825 ^ n_21984;
assign n_21996 = ~n_21984 & n_21254;
assign n_21997 = n_21985 ^ n_21970;
assign n_21998 = n_21983 & ~n_21986;
assign n_21999 = n_21987 ^ n_21905;
assign n_22000 = n_21961 ^ n_21988;
assign n_22001 = ~n_21988 & ~n_21961;
assign n_22002 = n_21989 ^ x477;
assign n_22003 = n_21990 ^ n_20269;
assign n_22004 = n_21991 ^ n_21512;
assign n_22005 = n_21992 ^ n_20269;
assign n_22006 = n_21992 ^ n_21990;
assign n_22007 = n_21994 & ~n_21993;
assign n_22008 = n_21994 ^ x40;
assign n_22009 = n_21995 ^ n_21253;
assign n_22010 = n_21995 ^ n_21173;
assign n_22011 = n_21996 ^ n_20825;
assign n_22012 = n_21997 ^ x476;
assign n_22013 = n_21998 ^ n_19891;
assign n_22014 = n_22000 ^ n_21562;
assign n_22015 = n_22002 ^ n_21997;
assign n_22016 = n_22004 ^ n_22000;
assign n_22017 = n_22005 ^ n_21990;
assign n_22018 = ~n_22003 & n_22006;
assign n_22019 = n_22007 ^ x40;
assign n_22020 = n_21981 & n_22008;
assign n_22021 = n_22008 ^ n_21981;
assign n_22022 = n_22009 ^ n_19910;
assign n_22023 = n_22011 ^ n_21280;
assign n_22024 = n_22013 ^ n_19910;
assign n_22025 = n_22013 ^ n_22009;
assign n_22026 = n_22015 ^ x476;
assign n_22027 = n_22015 & ~n_22012;
assign n_22028 = n_22016 ^ n_20876;
assign n_22029 = n_22016 & n_22014;
assign n_22030 = n_22016 ^ n_21562;
assign n_22031 = n_22017 ^ x55;
assign n_22032 = n_22018 ^ n_20269;
assign n_22033 = n_22019 ^ n_22017;
assign n_22034 = n_22019 ^ x55;
assign n_22035 = n_20845 ^ n_22023;
assign n_22036 = n_22023 & n_21293;
assign n_22037 = n_22024 ^ n_22009;
assign n_22038 = ~n_22022 & n_22025;
assign n_22039 = n_22026 ^ n_22001;
assign n_22040 = n_22001 & n_22026;
assign n_22041 = n_22027 ^ x476;
assign n_22042 = n_22028 ^ n_20289;
assign n_22043 = n_22029 ^ n_21562;
assign n_22044 = n_21944 ^ n_22030;
assign n_22045 = n_22032 ^ n_22028;
assign n_22046 = n_22031 & ~n_22033;
assign n_22047 = n_22034 ^ n_22017;
assign n_22048 = n_22035 ^ n_21292;
assign n_22049 = n_21212 ^ n_22035;
assign n_22050 = n_22036 ^ n_20845;
assign n_22051 = n_22037 ^ x475;
assign n_22052 = n_22038 ^ n_19910;
assign n_22053 = n_22039 ^ n_21602;
assign n_22054 = n_22041 ^ n_22037;
assign n_22055 = n_22043 ^ n_22039;
assign n_22056 = n_22043 ^ n_21602;
assign n_22057 = n_22045 ^ n_20289;
assign n_22058 = ~n_22045 & n_22042;
assign n_22059 = n_22046 ^ x55;
assign n_22060 = ~n_22020 & n_22047;
assign n_22061 = n_22047 ^ n_22020;
assign n_22062 = n_22048 ^ n_19930;
assign n_22063 = n_22050 ^ n_21319;
assign n_22064 = n_22052 ^ n_19930;
assign n_22065 = n_22052 ^ n_22048;
assign n_22066 = n_22054 ^ x475;
assign n_22067 = ~n_22054 & n_22051;
assign n_22068 = n_22055 ^ n_20894;
assign n_22069 = ~n_22055 & n_22053;
assign n_22070 = n_22056 ^ n_22039;
assign n_22071 = n_22057 ^ x54;
assign n_22072 = n_22058 ^ n_20289;
assign n_22073 = n_22059 ^ n_22057;
assign n_22074 = n_22063 ^ n_20867;
assign n_22075 = n_22063 & ~n_21333;
assign n_22076 = n_22064 ^ n_22048;
assign n_22077 = ~n_22062 & ~n_22065;
assign n_22078 = n_22066 ^ n_22040;
assign n_22079 = n_22040 & ~n_22066;
assign n_22080 = n_22067 ^ x475;
assign n_22081 = n_22068 ^ n_20308;
assign n_22082 = n_22069 ^ n_21602;
assign n_22083 = n_21982 ^ n_22070;
assign n_22084 = n_22072 ^ n_22068;
assign n_22085 = n_22073 & ~n_22071;
assign n_22086 = n_22073 ^ x54;
assign n_22087 = n_22074 ^ n_21332;
assign n_22088 = n_21252 ^ n_22074;
assign n_22089 = n_22075 ^ n_20867;
assign n_22090 = n_22076 ^ x474;
assign n_22091 = n_22077 ^ n_19930;
assign n_22092 = n_22078 ^ n_21640;
assign n_22093 = n_22080 ^ n_22076;
assign n_22094 = n_22082 ^ n_22078;
assign n_22095 = n_22082 ^ n_21640;
assign n_22096 = n_22084 ^ n_20308;
assign n_22097 = n_22084 & n_22081;
assign n_22098 = n_22085 ^ x54;
assign n_22099 = ~n_22060 & n_22086;
assign n_22100 = n_22086 ^ n_22060;
assign n_22101 = n_22087 ^ n_19950;
assign n_22102 = n_22089 ^ n_21350;
assign n_22103 = n_22091 ^ n_19950;
assign n_22104 = n_22091 ^ n_22087;
assign n_22105 = n_22093 ^ x474;
assign n_22106 = ~n_22093 & n_22090;
assign n_22107 = n_22094 ^ n_20918;
assign n_22108 = n_22094 & ~n_22092;
assign n_22109 = n_22095 ^ n_22078;
assign n_22110 = n_22096 ^ x53;
assign n_22111 = n_22097 ^ n_20308;
assign n_22112 = n_22098 ^ n_22096;
assign n_22113 = n_22102 ^ n_20887;
assign n_22114 = n_22103 ^ n_22087;
assign n_22115 = n_22101 & ~n_22104;
assign n_22116 = n_22105 ^ n_22079;
assign n_22117 = n_22079 & ~n_22105;
assign n_22118 = n_22106 ^ x474;
assign n_22119 = n_22107 ^ n_20326;
assign n_22120 = n_22108 ^ n_21640;
assign n_22121 = n_22021 ^ n_22109;
assign n_22122 = n_22111 ^ n_20326;
assign n_22123 = n_22111 ^ n_22107;
assign n_22124 = n_22112 & ~n_22110;
assign n_22125 = n_22112 ^ x53;
assign n_22126 = n_22113 ^ n_21381;
assign n_22127 = n_22113 ^ n_21251;
assign n_22128 = n_22114 ^ x473;
assign n_22129 = n_22115 ^ n_19950;
assign n_22130 = n_22116 ^ n_21680;
assign n_22131 = n_22118 ^ n_22114;
assign n_22132 = n_22120 ^ n_22116;
assign n_22133 = n_22120 ^ n_21680;
assign n_22134 = n_22122 ^ n_22107;
assign n_22135 = n_22119 & ~n_22123;
assign n_22136 = n_22124 ^ x53;
assign n_22137 = n_22099 & n_22125;
assign n_22138 = n_22125 ^ n_22099;
assign n_22139 = n_22127 ^ n_21278;
assign n_22140 = n_22129 ^ x472;
assign n_22141 = n_22131 ^ x473;
assign n_22142 = ~n_22131 & n_22128;
assign n_22143 = n_22132 ^ n_20944;
assign n_22144 = n_22132 & ~n_22130;
assign n_22145 = n_22133 ^ n_22116;
assign n_22146 = n_22134 ^ x52;
assign n_22147 = n_22135 ^ n_20326;
assign n_22148 = n_22136 ^ n_22134;
assign n_22149 = n_22140 ^ n_22126;
assign n_22150 = n_22141 ^ n_22117;
assign n_22151 = n_22117 & ~n_22141;
assign n_22152 = n_22142 ^ x473;
assign n_22153 = n_22143 ^ n_20345;
assign n_22154 = n_22144 ^ n_21680;
assign n_22155 = n_22061 ^ n_22145;
assign n_22156 = n_22147 ^ n_20345;
assign n_22157 = n_22147 ^ n_22143;
assign n_22158 = ~n_22148 & n_22146;
assign n_22159 = n_22148 ^ x52;
assign n_22160 = n_22150 ^ n_21719;
assign n_22161 = n_22152 ^ n_22149;
assign n_22162 = n_22154 ^ n_22150;
assign n_22163 = n_22154 ^ n_21719;
assign n_22164 = n_22156 ^ n_22143;
assign n_22165 = n_22153 & n_22157;
assign n_22166 = n_22158 ^ x52;
assign n_22167 = n_22137 & ~n_22159;
assign n_22168 = n_22159 ^ n_22137;
assign n_22169 = n_22161 ^ n_22151;
assign n_22170 = n_22162 ^ n_20972;
assign n_22171 = n_22162 & n_22160;
assign n_22172 = n_22163 ^ n_22150;
assign n_22173 = n_22164 ^ x51;
assign n_22174 = n_22165 ^ n_20345;
assign n_22175 = n_22166 ^ n_22164;
assign n_22176 = n_22169 ^ n_21758;
assign n_22177 = n_22170 ^ n_20364;
assign n_22178 = n_22171 ^ n_21719;
assign n_22179 = n_22100 ^ n_22172;
assign n_22180 = n_22174 ^ n_20364;
assign n_22181 = n_22174 ^ n_22170;
assign n_22182 = n_22175 ^ x51;
assign n_22183 = ~n_22175 & n_22173;
assign n_22184 = n_22178 ^ n_22169;
assign n_22185 = n_22178 ^ n_21758;
assign n_22186 = n_22180 ^ n_22170;
assign n_22187 = ~n_22177 & ~n_22181;
assign n_22188 = ~n_22182 & n_22167;
assign n_22189 = n_22167 ^ n_22182;
assign n_22190 = n_22183 ^ x51;
assign n_22191 = n_22184 ^ n_21008;
assign n_22192 = ~n_22184 & ~n_22176;
assign n_22193 = n_22185 ^ n_22169;
assign n_22194 = n_22186 ^ x50;
assign n_22195 = n_22187 ^ n_20364;
assign n_22196 = n_22190 ^ n_22186;
assign n_22197 = n_22191 ^ n_20384;
assign n_22198 = n_22192 ^ n_21758;
assign n_22199 = n_22138 ^ n_22193;
assign n_22200 = n_22195 ^ n_20384;
assign n_22201 = n_22195 ^ n_22191;
assign n_22202 = n_22196 ^ x50;
assign n_22203 = ~n_22196 & n_22194;
assign n_22204 = n_22198 ^ n_21797;
assign n_22205 = n_22200 ^ n_22191;
assign n_22206 = ~n_22197 & n_22201;
assign n_22207 = n_22188 & ~n_22202;
assign n_22208 = n_22202 ^ n_22188;
assign n_22209 = n_22203 ^ x50;
assign n_22210 = n_20926 ^ n_22204;
assign n_22211 = n_22204 & n_21812;
assign n_22212 = n_22205 ^ x49;
assign n_22213 = n_22206 ^ n_20384;
assign n_22214 = n_22209 ^ n_22205;
assign n_22215 = n_22210 ^ n_21797;
assign n_22216 = n_22168 ^ n_22210;
assign n_22217 = n_22211 ^ n_20926;
assign n_22218 = n_22213 ^ n_20403;
assign n_22219 = n_22214 ^ x49;
assign n_22220 = n_22214 & ~n_22212;
assign n_22221 = n_22215 ^ n_21044;
assign n_22222 = n_22217 ^ n_21837;
assign n_22223 = ~n_22207 & ~n_22219;
assign n_22224 = n_22219 ^ n_22207;
assign n_22225 = n_22220 ^ x49;
assign n_22226 = n_22218 ^ n_22221;
assign n_22227 = n_22221 ^ n_20403;
assign n_22228 = n_22213 ^ n_22221;
assign n_22229 = n_20982 ^ n_22222;
assign n_22230 = n_22222 & n_21852;
assign n_22231 = n_22225 ^ n_22226;
assign n_22232 = n_22226 ^ x48;
assign n_22233 = n_22227 & ~n_22228;
assign n_22234 = n_22229 ^ n_21837;
assign n_22235 = n_22189 ^ n_22229;
assign n_22236 = n_22230 ^ n_20982;
assign n_22237 = n_22231 ^ x48;
assign n_22238 = ~n_22231 & n_22232;
assign n_22239 = n_22233 ^ n_20403;
assign n_22240 = n_22234 ^ n_21069;
assign n_22241 = n_22236 ^ n_21031;
assign n_22242 = n_22236 ^ n_21877;
assign n_22243 = ~n_22223 & ~n_22237;
assign n_22244 = n_22237 ^ n_22223;
assign n_22245 = n_22238 ^ x48;
assign n_22246 = n_22239 ^ n_22240;
assign n_22247 = n_22240 ^ n_20430;
assign n_22248 = n_22241 ^ n_21124;
assign n_22249 = n_22241 ^ n_21877;
assign n_22250 = ~n_21892 & ~n_22242;
assign n_22251 = n_22245 ^ x63;
assign n_22252 = n_22246 ^ n_20430;
assign n_22253 = n_22246 & ~n_22247;
assign n_22254 = n_22248 ^ n_20456;
assign n_22255 = n_22208 ^ n_22249;
assign n_22256 = n_22250 ^ n_21031;
assign n_22257 = n_22251 ^ n_22252;
assign n_22258 = n_22252 ^ x63;
assign n_22259 = n_22245 ^ n_22252;
assign n_22260 = n_22253 ^ n_20430;
assign n_22261 = n_22256 ^ n_21917;
assign n_22262 = ~n_22243 & ~n_22257;
assign n_22263 = n_22257 ^ n_22243;
assign n_22264 = ~n_22258 & n_22259;
assign n_22265 = n_22260 ^ n_22248;
assign n_22266 = n_21095 ^ n_22261;
assign n_22267 = n_22261 & n_21932;
assign n_22268 = n_22264 ^ x63;
assign n_22269 = n_22265 ^ n_20456;
assign n_22270 = ~n_22265 & n_22254;
assign n_22271 = n_22266 ^ n_21917;
assign n_22272 = n_22224 ^ n_22266;
assign n_22273 = n_22267 ^ n_21095;
assign n_22274 = n_22268 ^ n_22269;
assign n_22275 = n_22269 ^ x62;
assign n_22276 = n_22270 ^ n_20456;
assign n_22277 = n_22271 ^ n_21162;
assign n_22278 = n_22273 ^ n_21956;
assign n_22279 = n_22274 ^ x62;
assign n_22280 = ~n_22274 & n_22275;
assign n_22281 = n_22276 ^ n_22277;
assign n_22282 = n_22277 ^ n_20487;
assign n_22283 = n_21135 ^ n_22278;
assign n_22284 = ~n_22278 & n_21971;
assign n_22285 = n_22262 & n_22279;
assign n_22286 = n_22279 ^ n_22262;
assign n_22287 = n_22280 ^ x62;
assign n_22288 = n_22281 ^ n_20487;
assign n_22289 = n_22281 & n_22282;
assign n_22290 = n_22283 ^ n_21956;
assign n_22291 = n_22244 ^ n_22283;
assign n_22292 = n_22284 ^ n_21135;
assign n_22293 = n_22287 ^ n_22288;
assign n_22294 = n_22288 ^ x61;
assign n_22295 = n_22289 ^ n_20487;
assign n_22296 = n_22290 ^ n_21201;
assign n_22297 = n_22292 ^ n_21173;
assign n_22298 = n_22292 ^ n_21995;
assign n_22299 = n_22293 ^ x61;
assign n_22300 = ~n_22293 & n_22294;
assign n_22301 = n_22295 ^ n_20523;
assign n_22302 = n_22296 ^ n_20523;
assign n_22303 = n_22295 ^ n_22296;
assign n_22304 = n_22297 ^ n_21240;
assign n_22305 = n_22297 ^ n_21995;
assign n_22306 = n_22010 & ~n_22298;
assign n_22307 = ~n_22285 & ~n_22299;
assign n_22308 = n_22299 ^ n_22285;
assign n_22309 = n_22300 ^ x61;
assign n_22310 = n_22301 ^ n_22296;
assign n_22311 = n_22302 & n_22303;
assign n_22312 = n_22304 ^ n_20562;
assign n_22313 = n_22263 ^ n_22305;
assign n_22314 = n_22306 ^ n_21173;
assign n_22315 = n_22309 ^ n_22310;
assign n_22316 = n_22310 ^ x60;
assign n_22317 = n_22311 ^ n_20523;
assign n_22318 = n_22314 ^ n_22035;
assign n_22319 = n_22315 ^ x60;
assign n_22320 = n_22315 & ~n_22316;
assign n_22321 = n_22317 ^ n_20562;
assign n_22322 = n_22317 ^ n_22304;
assign n_22323 = n_21212 ^ n_22318;
assign n_22324 = ~n_22318 & n_22049;
assign n_22325 = ~n_22307 & ~n_22319;
assign n_22326 = n_22320 ^ x60;
assign n_22327 = n_22321 ^ n_22304;
assign n_22328 = ~n_22312 & n_22322;
assign n_22329 = n_22323 ^ n_22035;
assign n_22330 = n_22286 ^ n_22323;
assign n_22331 = n_22324 ^ n_21212;
assign n_22332 = n_22326 ^ n_22327;
assign n_22333 = n_22327 ^ x59;
assign n_22334 = n_22328 ^ n_20562;
assign n_22335 = n_22329 ^ n_21280;
assign n_22336 = n_22331 ^ n_21252;
assign n_22337 = n_22331 ^ n_22074;
assign n_22338 = n_22332 ^ x59;
assign n_22339 = n_22332 & ~n_22333;
assign n_22340 = n_22334 ^ n_20600;
assign n_22341 = n_22335 ^ n_20600;
assign n_22342 = n_22334 ^ n_22335;
assign n_22343 = n_22336 ^ n_21319;
assign n_22344 = n_22336 ^ n_22074;
assign n_22345 = n_22088 & ~n_22337;
assign n_22346 = n_22325 ^ n_22338;
assign n_22347 = ~n_22338 & n_22325;
assign n_22348 = n_22339 ^ x59;
assign n_22349 = n_22340 ^ n_22335;
assign n_22350 = n_22341 & ~n_22342;
assign n_22351 = n_22343 ^ n_20639;
assign n_22352 = n_22308 ^ n_22344;
assign n_22353 = n_22345 ^ n_21252;
assign n_22354 = n_22346 ^ n_20905;
assign n_22355 = ~n_22346 & n_21348;
assign n_22356 = n_22346 ^ n_20915;
assign n_22357 = n_22348 ^ n_22349;
assign n_22358 = n_22349 ^ x58;
assign n_22359 = n_22350 ^ n_20600;
assign n_22360 = n_22353 ^ n_22139;
assign n_22361 = x135 & n_22354;
assign n_22362 = n_22354 ^ x135;
assign n_22363 = n_21393 ^ n_22355;
assign n_22364 = ~n_20419 & ~n_22356;
assign n_22365 = n_22356 ^ n_21331;
assign n_22366 = n_22357 ^ x58;
assign n_22367 = ~n_22357 & n_22358;
assign n_22368 = n_22359 ^ n_20639;
assign n_22369 = n_22359 ^ n_22343;
assign n_22370 = n_22360 ^ n_22113;
assign n_22371 = n_22360 ^ n_22307;
assign n_22372 = n_22361 ^ x134;
assign n_22373 = n_22364 ^ n_20445;
assign n_22374 = n_22366 ^ n_22347;
assign n_22375 = ~n_22347 & ~n_22366;
assign n_22376 = n_22367 ^ x58;
assign n_22377 = n_22368 ^ n_22343;
assign n_22378 = ~n_22351 & n_22369;
assign n_22379 = n_22370 ^ n_21350;
assign n_22380 = n_22371 ^ n_22319;
assign n_22381 = n_22374 ^ n_22363;
assign n_22382 = n_22374 ^ n_22355;
assign n_22383 = n_22376 ^ n_22377;
assign n_22384 = n_22377 ^ x57;
assign n_22385 = n_22378 ^ n_20639;
assign n_22386 = n_22379 ^ n_20667;
assign n_22387 = n_22381 ^ n_21392;
assign n_22388 = ~n_22363 & n_22382;
assign n_22389 = n_22383 ^ x57;
assign n_22390 = n_22383 & ~n_22384;
assign n_22391 = n_22385 ^ x56;
assign n_22392 = n_22387 ^ n_22373;
assign n_22393 = n_22387 ^ n_22364;
assign n_22394 = n_22388 ^ n_21393;
assign n_22395 = n_22389 ^ n_22375;
assign n_22396 = ~n_22375 & ~n_22389;
assign n_22397 = n_22390 ^ x57;
assign n_22398 = n_22391 ^ n_22386;
assign n_22399 = n_22392 ^ n_22361;
assign n_22400 = n_22392 ^ n_22372;
assign n_22401 = ~n_22373 & n_22393;
assign n_22402 = n_22394 ^ n_21445;
assign n_22403 = n_21445 ^ n_22395;
assign n_22404 = n_22394 ^ n_22395;
assign n_22405 = n_22397 ^ n_22398;
assign n_22406 = n_22372 & ~n_22399;
assign n_22407 = n_22362 & n_22400;
assign n_22408 = n_22400 ^ n_22362;
assign n_22409 = n_22401 ^ n_20445;
assign n_22410 = n_22402 ^ n_22395;
assign n_22411 = n_22403 & n_22404;
assign n_22412 = n_22405 ^ n_22396;
assign n_22413 = n_22406 ^ x134;
assign n_22414 = n_22410 ^ n_21430;
assign n_22415 = n_22411 ^ n_21445;
assign n_22416 = n_21483 ^ n_22412;
assign n_22417 = n_22409 ^ n_22414;
assign n_22418 = n_22414 ^ n_20480;
assign n_22419 = n_22415 ^ n_21483;
assign n_22420 = n_22415 ^ n_22412;
assign n_22421 = n_22417 ^ n_20480;
assign n_22422 = n_22417 & n_22418;
assign n_22423 = n_22419 ^ n_22412;
assign n_22424 = ~n_22416 & n_22420;
assign n_22425 = n_22413 ^ n_22421;
assign n_22426 = n_22421 ^ x133;
assign n_22427 = n_22422 ^ n_20480;
assign n_22428 = n_22423 ^ n_21469;
assign n_22429 = n_22424 ^ n_21483;
assign n_22430 = n_22425 ^ x133;
assign n_22431 = n_22425 & ~n_22426;
assign n_22432 = n_22427 ^ n_20518;
assign n_22433 = n_22428 ^ n_20518;
assign n_22434 = n_22427 ^ n_22428;
assign n_22435 = n_21520 ^ n_22429;
assign n_22436 = n_22407 & ~n_22430;
assign n_22437 = n_22430 ^ n_22407;
assign n_22438 = n_22431 ^ x133;
assign n_22439 = n_22432 ^ n_22428;
assign n_22440 = n_22433 & ~n_22434;
assign n_22441 = n_21365 ^ n_22435;
assign n_22442 = n_22435 & ~n_21533;
assign n_22443 = n_22438 ^ n_22439;
assign n_22444 = n_22439 ^ x132;
assign n_22445 = n_22440 ^ n_20518;
assign n_22446 = n_22441 ^ n_21506;
assign n_22447 = n_22442 ^ n_21365;
assign n_22448 = n_22443 ^ x132;
assign n_22449 = ~n_22443 & n_22444;
assign n_22450 = n_22445 ^ n_20557;
assign n_22451 = n_22446 ^ n_20557;
assign n_22452 = n_22445 ^ n_22446;
assign n_22453 = n_21558 ^ n_22447;
assign n_22454 = ~n_22436 & ~n_22448;
assign n_22455 = n_22448 ^ n_22436;
assign n_22456 = n_22449 ^ x132;
assign n_22457 = n_22450 ^ n_22446;
assign n_22458 = ~n_22451 & ~n_22452;
assign n_22459 = n_22453 ^ n_21448;
assign n_22460 = ~n_22453 & n_21571;
assign n_22461 = n_22456 ^ n_22457;
assign n_22462 = n_22457 ^ x131;
assign n_22463 = n_22458 ^ n_20557;
assign n_22464 = n_22459 ^ n_21544;
assign n_22465 = n_22460 ^ n_21448;
assign n_22466 = n_22461 ^ x131;
assign n_22467 = n_22461 & ~n_22462;
assign n_22468 = n_22463 ^ n_20595;
assign n_22469 = n_22464 ^ n_20595;
assign n_22470 = n_22463 ^ n_22464;
assign n_22471 = n_22465 ^ n_21611;
assign n_22472 = n_22465 ^ n_21499;
assign n_22473 = ~n_22454 & ~n_22466;
assign n_22474 = n_22466 ^ n_22454;
assign n_22475 = n_22467 ^ x131;
assign n_22476 = n_22468 ^ n_22464;
assign n_22477 = n_22469 & n_22470;
assign n_22478 = n_22471 ^ n_21583;
assign n_22479 = ~n_21611 & ~n_22472;
assign n_22480 = n_22475 ^ n_22476;
assign n_22481 = n_22476 ^ x130;
assign n_22482 = n_22477 ^ n_20595;
assign n_22483 = n_22479 ^ n_21598;
assign n_22484 = n_22480 ^ x130;
assign n_22485 = n_22480 & ~n_22481;
assign n_22486 = n_22482 ^ n_20634;
assign n_22487 = n_22478 ^ n_22482;
assign n_22488 = n_21636 ^ n_22483;
assign n_22489 = n_22484 & ~n_22473;
assign n_22490 = n_22473 ^ n_22484;
assign n_22491 = n_22485 ^ x130;
assign n_22492 = n_22478 ^ n_22486;
assign n_22493 = n_22486 & n_22487;
assign n_22494 = n_21550 ^ n_22488;
assign n_22495 = ~n_22488 & ~n_21649;
assign n_22496 = n_22491 ^ n_22492;
assign n_22497 = n_22492 ^ x129;
assign n_22498 = n_22493 ^ n_20634;
assign n_22499 = n_22494 ^ n_21622;
assign n_22500 = n_22495 ^ n_21550;
assign n_22501 = n_22496 ^ x129;
assign n_22502 = n_22496 & ~n_22497;
assign n_22503 = n_22498 ^ n_20673;
assign n_22504 = n_22499 ^ n_20673;
assign n_22505 = n_22498 ^ n_22499;
assign n_22506 = n_21676 ^ n_22500;
assign n_22507 = ~n_22501 & ~n_22489;
assign n_22508 = n_22489 ^ n_22501;
assign n_22509 = n_22502 ^ x129;
assign n_22510 = n_22503 ^ n_22499;
assign n_22511 = n_22504 & ~n_22505;
assign n_22512 = n_21589 ^ n_22506;
assign n_22513 = ~n_22506 & ~n_21689;
assign n_22514 = n_22509 ^ x128;
assign n_22515 = n_22509 ^ n_22510;
assign n_22516 = n_22511 ^ n_20673;
assign n_22517 = n_22512 ^ n_21660;
assign n_22518 = n_22513 ^ n_21589;
assign n_22519 = ~n_22515 & n_22514;
assign n_22520 = n_22515 ^ x128;
assign n_22521 = n_22516 ^ n_20706;
assign n_22522 = n_22517 ^ n_20706;
assign n_22523 = n_22516 ^ n_22517;
assign n_22524 = n_22518 ^ n_21628;
assign n_22525 = n_22518 ^ n_21715;
assign n_22526 = n_22519 ^ x128;
assign n_22527 = ~n_22520 & ~n_22507;
assign n_22528 = n_22507 ^ n_22520;
assign n_22529 = n_22521 ^ n_22517;
assign n_22530 = n_22522 & ~n_22523;
assign n_22531 = n_22524 ^ n_21715;
assign n_22532 = ~n_21728 & ~n_22525;
assign n_22533 = n_22526 ^ n_22529;
assign n_22534 = n_22529 ^ x143;
assign n_22535 = n_22530 ^ n_20706;
assign n_22536 = n_22531 ^ n_21700;
assign n_22537 = n_22532 ^ n_21628;
assign n_22538 = n_22533 ^ x143;
assign n_22539 = ~n_22533 & n_22534;
assign n_22540 = n_22535 ^ n_20733;
assign n_22541 = n_22536 ^ n_20733;
assign n_22542 = n_22535 ^ n_22536;
assign n_22543 = n_21754 ^ n_22537;
assign n_22544 = ~n_22538 & n_22527;
assign n_22545 = n_22527 ^ n_22538;
assign n_22546 = n_22539 ^ x143;
assign n_22547 = n_22540 ^ n_22536;
assign n_22548 = n_22541 & n_22542;
assign n_22549 = n_21666 ^ n_22543;
assign n_22550 = n_22543 & ~n_21767;
assign n_22551 = n_22546 ^ n_22547;
assign n_22552 = n_22547 ^ x142;
assign n_22553 = n_22548 ^ n_20733;
assign n_22554 = n_22549 ^ n_21739;
assign n_22555 = n_22550 ^ n_21666;
assign n_22556 = n_22551 ^ x142;
assign n_22557 = ~n_22551 & n_22552;
assign n_22558 = n_22553 ^ n_20756;
assign n_22559 = n_22554 ^ n_20756;
assign n_22560 = n_22553 ^ n_22554;
assign n_22561 = n_21793 ^ n_22555;
assign n_22562 = ~n_22556 & n_22544;
assign n_22563 = n_22544 ^ n_22556;
assign n_22564 = n_22557 ^ x142;
assign n_22565 = n_22558 ^ n_22554;
assign n_22566 = ~n_22559 & n_22560;
assign n_22567 = n_21706 ^ n_22561;
assign n_22568 = ~n_22561 & n_21806;
assign n_22569 = n_22564 ^ n_22565;
assign n_22570 = n_22565 ^ x141;
assign n_22571 = n_22566 ^ n_20756;
assign n_22572 = n_22567 ^ n_21778;
assign n_22573 = n_22567 ^ n_22362;
assign n_22574 = n_22568 ^ n_21706;
assign n_22575 = n_22569 ^ x141;
assign n_22576 = ~n_22569 & n_22570;
assign n_22577 = n_22571 ^ n_20768;
assign n_22578 = n_22572 ^ n_20768;
assign n_22579 = n_22571 ^ n_22572;
assign n_22580 = n_21833 ^ n_22574;
assign n_22581 = n_22562 & ~n_22575;
assign n_22582 = n_22575 ^ n_22562;
assign n_22583 = n_22576 ^ x141;
assign n_22584 = n_22577 ^ n_22572;
assign n_22585 = ~n_22578 & n_22579;
assign n_22586 = n_21745 ^ n_22580;
assign n_22587 = n_22580 & ~n_21846;
assign n_22588 = n_22583 ^ n_22584;
assign n_22589 = n_22584 ^ x140;
assign n_22590 = n_22585 ^ n_20768;
assign n_22591 = n_22586 ^ n_21818;
assign n_22592 = n_22408 ^ n_22586;
assign n_22593 = n_22587 ^ n_21745;
assign n_22594 = n_22588 ^ x140;
assign n_22595 = ~n_22588 & n_22589;
assign n_22596 = n_22590 ^ n_20787;
assign n_22597 = n_22591 ^ n_20787;
assign n_22598 = n_22590 ^ n_22591;
assign n_22599 = n_21873 ^ n_22593;
assign n_22600 = n_22581 & ~n_22594;
assign n_22601 = n_22594 ^ n_22581;
assign n_22602 = n_22595 ^ x140;
assign n_22603 = n_22596 ^ n_22591;
assign n_22604 = n_22597 & ~n_22598;
assign n_22605 = ~n_22599 & ~n_21886;
assign n_22606 = n_21784 ^ n_22599;
assign n_22607 = n_22602 ^ n_22603;
assign n_22608 = n_22603 ^ x139;
assign n_22609 = n_22604 ^ n_20787;
assign n_22610 = n_22605 ^ n_21784;
assign n_22611 = n_22606 ^ n_21858;
assign n_22612 = n_22437 ^ n_22606;
assign n_22613 = n_22607 ^ x139;
assign n_22614 = n_22607 & ~n_22608;
assign n_22615 = n_22609 ^ n_20802;
assign n_22616 = n_21913 ^ n_22610;
assign n_22617 = n_22611 ^ n_20802;
assign n_22618 = n_22609 ^ n_22611;
assign n_22619 = n_22600 ^ n_22613;
assign n_22620 = ~n_22613 & ~n_22600;
assign n_22621 = n_22614 ^ x139;
assign n_22622 = n_22615 ^ n_22611;
assign n_22623 = ~n_22616 & ~n_21926;
assign n_22624 = n_21824 ^ n_22616;
assign n_22625 = n_22617 & ~n_22618;
assign n_22626 = n_22621 ^ n_22622;
assign n_22627 = n_22622 ^ x138;
assign n_22628 = n_22623 ^ n_21824;
assign n_22629 = n_22624 ^ n_21899;
assign n_22630 = n_22455 ^ n_22624;
assign n_22631 = n_22625 ^ n_20802;
assign n_22632 = n_22626 ^ x138;
assign n_22633 = n_22626 & ~n_22627;
assign n_22634 = n_21952 ^ n_22628;
assign n_22635 = n_22629 ^ n_20817;
assign n_22636 = n_22631 ^ n_22629;
assign n_22637 = n_22631 ^ n_20817;
assign n_22638 = n_22620 & ~n_22632;
assign n_22639 = n_22632 ^ n_22620;
assign n_22640 = n_22633 ^ x138;
assign n_22641 = ~n_22634 & ~n_21965;
assign n_22642 = n_21864 ^ n_22634;
assign n_22643 = n_22635 & ~n_22636;
assign n_22644 = n_22637 ^ n_22629;
assign n_22645 = n_22641 ^ n_21864;
assign n_22646 = n_22642 ^ n_21938;
assign n_22647 = n_22474 ^ n_22642;
assign n_22648 = n_22643 ^ n_20817;
assign n_22649 = n_22640 ^ n_22644;
assign n_22650 = n_22644 ^ x137;
assign n_22651 = n_22645 ^ n_21987;
assign n_22652 = n_22645 ^ n_21999;
assign n_22653 = n_22646 ^ n_20835;
assign n_22654 = n_22648 ^ n_22646;
assign n_22655 = n_22648 ^ n_20835;
assign n_22656 = n_22649 ^ x137;
assign n_22657 = n_22649 & ~n_22650;
assign n_22658 = n_21999 & ~n_22651;
assign n_22659 = n_22652 ^ n_22490;
assign n_22660 = n_22652 ^ n_21977;
assign n_22661 = ~n_22653 & n_22654;
assign n_22662 = n_22655 ^ n_22646;
assign n_22663 = n_22656 & ~n_22638;
assign n_22664 = n_22638 ^ n_22656;
assign n_22665 = n_22657 ^ x137;
assign n_22666 = n_22658 ^ n_21905;
assign n_22667 = n_22660 ^ n_20848;
assign n_22668 = n_22661 ^ n_20835;
assign n_22669 = n_22662 ^ x136;
assign n_22670 = n_22665 ^ n_22662;
assign n_22671 = n_22666 ^ n_21944;
assign n_22672 = n_22666 ^ n_22030;
assign n_22673 = n_22668 ^ n_22660;
assign n_22674 = ~n_22670 & n_22669;
assign n_22675 = n_22670 ^ x136;
assign n_22676 = n_22671 ^ n_22030;
assign n_22677 = n_22044 & n_22672;
assign n_22678 = n_22673 ^ n_20848;
assign n_22679 = n_22673 & ~n_22667;
assign n_22680 = n_22674 ^ x136;
assign n_22681 = n_22663 & ~n_22675;
assign n_22682 = n_22675 ^ n_22663;
assign n_22683 = n_22676 ^ n_22508;
assign n_22684 = n_22676 ^ n_22016;
assign n_22685 = n_22677 ^ n_21944;
assign n_22686 = n_22678 ^ x151;
assign n_22687 = n_22679 ^ n_20848;
assign n_22688 = n_22680 ^ n_22678;
assign n_22689 = n_22680 ^ x151;
assign n_22690 = n_22684 ^ n_20876;
assign n_22691 = n_22070 ^ n_22685;
assign n_22692 = n_22687 ^ n_22684;
assign n_22693 = n_22686 & ~n_22688;
assign n_22694 = n_22689 ^ n_22678;
assign n_22695 = n_21982 ^ n_22691;
assign n_22696 = n_22691 & n_22083;
assign n_22697 = n_22692 ^ n_20876;
assign n_22698 = n_22692 & n_22690;
assign n_22699 = n_22693 ^ x151;
assign n_22700 = ~n_22681 & n_22694;
assign n_22701 = n_22694 ^ n_22681;
assign n_22702 = n_22695 ^ n_22055;
assign n_22703 = n_22528 ^ n_22695;
assign n_22704 = n_22696 ^ n_21982;
assign n_22705 = n_22697 ^ x150;
assign n_22706 = n_22698 ^ n_20876;
assign n_22707 = n_22699 ^ n_22697;
assign n_22708 = n_22702 ^ n_20894;
assign n_22709 = n_22109 ^ n_22704;
assign n_22710 = n_22706 ^ n_22702;
assign n_22711 = n_22707 & ~n_22705;
assign n_22712 = n_22707 ^ x150;
assign n_22713 = n_22021 ^ n_22709;
assign n_22714 = n_22709 & ~n_22121;
assign n_22715 = n_22710 ^ n_20894;
assign n_22716 = ~n_22710 & n_22708;
assign n_22717 = n_22711 ^ x150;
assign n_22718 = ~n_22700 & n_22712;
assign n_22719 = n_22712 ^ n_22700;
assign n_22720 = n_22713 ^ n_22094;
assign n_22721 = n_22545 ^ n_22713;
assign n_22722 = n_22714 ^ n_22021;
assign n_22723 = n_22715 ^ x149;
assign n_22724 = n_22716 ^ n_20894;
assign n_22725 = n_22717 ^ n_22715;
assign n_22726 = n_22720 ^ n_20918;
assign n_22727 = n_22145 ^ n_22722;
assign n_22728 = n_22724 ^ n_20918;
assign n_22729 = n_22724 ^ n_22720;
assign n_22730 = ~n_22725 & n_22723;
assign n_22731 = n_22725 ^ x149;
assign n_22732 = n_22061 ^ n_22727;
assign n_22733 = n_22727 & ~n_22155;
assign n_22734 = n_22728 ^ n_22720;
assign n_22735 = n_22726 & n_22729;
assign n_22736 = n_22730 ^ x149;
assign n_22737 = n_22718 & ~n_22731;
assign n_22738 = n_22731 ^ n_22718;
assign n_22739 = n_22732 ^ n_22132;
assign n_22740 = n_22563 ^ n_22732;
assign n_22741 = n_22733 ^ n_22061;
assign n_22742 = n_22734 ^ x148;
assign n_22743 = n_22735 ^ n_20918;
assign n_22744 = n_22736 ^ n_22734;
assign n_22745 = n_22739 ^ n_20944;
assign n_22746 = n_22172 ^ n_22741;
assign n_22747 = n_22743 ^ n_20944;
assign n_22748 = n_22743 ^ n_22739;
assign n_22749 = ~n_22744 & n_22742;
assign n_22750 = n_22744 ^ x148;
assign n_22751 = n_22100 ^ n_22746;
assign n_22752 = ~n_22746 & ~n_22179;
assign n_22753 = n_22747 ^ n_22739;
assign n_22754 = ~n_22745 & ~n_22748;
assign n_22755 = n_22749 ^ x148;
assign n_22756 = n_22737 & ~n_22750;
assign n_22757 = n_22750 ^ n_22737;
assign n_22758 = n_22751 ^ n_22162;
assign n_22759 = n_22582 ^ n_22751;
assign n_22760 = n_22752 ^ n_22100;
assign n_22761 = n_22753 ^ x147;
assign n_22762 = n_22754 ^ n_20944;
assign n_22763 = n_22755 ^ n_22753;
assign n_22764 = n_22758 ^ n_20972;
assign n_22765 = n_22193 ^ n_22760;
assign n_22766 = n_22762 ^ n_20972;
assign n_22767 = n_22762 ^ n_22758;
assign n_22768 = ~n_22763 & n_22761;
assign n_22769 = n_22763 ^ x147;
assign n_22770 = n_22138 ^ n_22765;
assign n_22771 = n_22765 & n_22199;
assign n_22772 = n_22766 ^ n_22758;
assign n_22773 = ~n_22764 & n_22767;
assign n_22774 = n_22768 ^ x147;
assign n_22775 = n_22756 & ~n_22769;
assign n_22776 = n_22770 ^ n_22184;
assign n_22777 = n_22601 ^ n_22770;
assign n_22778 = n_22771 ^ n_22138;
assign n_22779 = n_22772 ^ x146;
assign n_22780 = n_22773 ^ n_20972;
assign n_22781 = n_22774 ^ n_22772;
assign n_22782 = n_22776 ^ n_21008;
assign n_22783 = n_22778 ^ n_22210;
assign n_22784 = n_22780 ^ n_21008;
assign n_22785 = n_22780 ^ n_22776;
assign n_22786 = n_22781 & ~n_22779;
assign n_22787 = n_22781 ^ x146;
assign n_22788 = n_22168 ^ n_22783;
assign n_22789 = ~n_22783 & ~n_22216;
assign n_22790 = n_22784 ^ n_22776;
assign n_22791 = ~n_22782 & ~n_22785;
assign n_22792 = n_22786 ^ x146;
assign n_22793 = ~n_22775 & ~n_22787;
assign n_22794 = n_22787 ^ n_22775;
assign n_22795 = n_22788 ^ n_22215;
assign n_22796 = n_22619 ^ n_22788;
assign n_22797 = n_22789 ^ n_22168;
assign n_22798 = n_22790 ^ x145;
assign n_22799 = n_22791 ^ n_21008;
assign n_22800 = n_22792 ^ n_22790;
assign n_22801 = ~n_22365 & n_22794;
assign n_22802 = n_22794 ^ n_21331;
assign n_22803 = n_22795 ^ n_21044;
assign n_22804 = n_22797 ^ n_22235;
assign n_22805 = n_22797 ^ n_22229;
assign n_22806 = n_22799 ^ n_21044;
assign n_22807 = n_22799 ^ n_22795;
assign n_22808 = n_22800 ^ x145;
assign n_22809 = n_22800 & ~n_22798;
assign n_22810 = n_22801 ^ n_22381;
assign n_22811 = n_20915 & ~n_22802;
assign n_22812 = x231 & n_22802;
assign n_22813 = n_22802 ^ n_22356;
assign n_22814 = n_22802 ^ x231;
assign n_22815 = n_22804 ^ n_22234;
assign n_22816 = n_22639 ^ n_22804;
assign n_22817 = n_22235 & ~n_22805;
assign n_22818 = n_22806 ^ n_22795;
assign n_22819 = n_22803 & ~n_22807;
assign n_22820 = n_22808 ^ n_22793;
assign n_22821 = ~n_22793 & n_22808;
assign n_22822 = n_22809 ^ x145;
assign n_22823 = n_22811 ^ n_20942;
assign n_22824 = n_22812 ^ x230;
assign n_22825 = n_22815 ^ n_21069;
assign n_22826 = n_22817 ^ n_22189;
assign n_22827 = n_22818 ^ x144;
assign n_22828 = n_22819 ^ n_21044;
assign n_22829 = n_22820 ^ n_22801;
assign n_22830 = n_22810 ^ n_22820;
assign n_22831 = n_22822 ^ n_22818;
assign n_22832 = n_22826 ^ n_22249;
assign n_22833 = n_22828 ^ n_22815;
assign n_22834 = ~n_22829 & n_22810;
assign n_22835 = n_22829 ^ n_21393;
assign n_22836 = n_22831 ^ x144;
assign n_22837 = n_22831 & ~n_22827;
assign n_22838 = n_22208 ^ n_22832;
assign n_22839 = ~n_22832 & n_22255;
assign n_22840 = n_22833 ^ n_21069;
assign n_22841 = ~n_22833 & ~n_22825;
assign n_22842 = n_22834 ^ n_22381;
assign n_22843 = n_22835 ^ n_22811;
assign n_22844 = n_22835 ^ n_22823;
assign n_22845 = n_22821 ^ n_22836;
assign n_22846 = n_22836 & n_22821;
assign n_22847 = n_22837 ^ x144;
assign n_22848 = n_22838 ^ n_22241;
assign n_22849 = n_22664 ^ n_22838;
assign n_22850 = n_22839 ^ n_22208;
assign n_22851 = n_22840 ^ x159;
assign n_22852 = n_22841 ^ n_21069;
assign n_22853 = n_22842 ^ n_22410;
assign n_22854 = n_22823 & n_22843;
assign n_22855 = n_22844 ^ n_22812;
assign n_22856 = n_22842 ^ n_22845;
assign n_22857 = n_22845 ^ n_22410;
assign n_22858 = n_22847 ^ x159;
assign n_22859 = n_22847 ^ n_22840;
assign n_22860 = n_22848 ^ n_21124;
assign n_22861 = n_22850 ^ n_22224;
assign n_22862 = n_22850 ^ n_22266;
assign n_22863 = n_22852 ^ n_22848;
assign n_22864 = n_22853 ^ n_22845;
assign n_22865 = n_22854 ^ n_20942;
assign n_22866 = n_22855 & n_22824;
assign n_22867 = n_22855 ^ x230;
assign n_22868 = n_22856 ^ n_21445;
assign n_22869 = n_22856 & n_22857;
assign n_22870 = n_22858 ^ n_22840;
assign n_22871 = n_22851 & ~n_22859;
assign n_22872 = n_22861 ^ n_22266;
assign n_22873 = n_22272 & ~n_22862;
assign n_22874 = n_22863 ^ n_21124;
assign n_22875 = n_22863 & n_22860;
assign n_22876 = n_22865 ^ n_20979;
assign n_22877 = n_22866 ^ x230;
assign n_22878 = n_22868 ^ n_20979;
assign n_22879 = n_22865 ^ n_22868;
assign n_22880 = n_22869 ^ n_22410;
assign n_22881 = n_22870 ^ n_22846;
assign n_22882 = n_22846 & ~n_22870;
assign n_22883 = n_22871 ^ x159;
assign n_22884 = n_22872 ^ n_22271;
assign n_22885 = n_22682 ^ n_22872;
assign n_22886 = n_22873 ^ n_22224;
assign n_22887 = n_22874 ^ x158;
assign n_22888 = n_22875 ^ n_21124;
assign n_22889 = n_22876 ^ n_22868;
assign n_22890 = n_22878 & n_22879;
assign n_22891 = n_22880 ^ n_22423;
assign n_22892 = n_22880 ^ n_22881;
assign n_22893 = n_22881 ^ n_22423;
assign n_22894 = n_22883 ^ n_22874;
assign n_22895 = n_22884 ^ n_21162;
assign n_22896 = n_22886 ^ n_22283;
assign n_22897 = n_22888 ^ n_22884;
assign n_22898 = n_22877 ^ n_22889;
assign n_22899 = n_22889 ^ x229;
assign n_22900 = n_22890 ^ n_20979;
assign n_22901 = n_22891 ^ n_22881;
assign n_22902 = n_22892 ^ n_21483;
assign n_22903 = n_22892 & ~n_22893;
assign n_22904 = n_22894 ^ x158;
assign n_22905 = ~n_22894 & n_22887;
assign n_22906 = n_22244 ^ n_22896;
assign n_22907 = n_22896 & n_22291;
assign n_22908 = n_22897 ^ n_21162;
assign n_22909 = ~n_22897 & ~n_22895;
assign n_22910 = n_22898 ^ x229;
assign n_22911 = ~n_22898 & n_22899;
assign n_22912 = n_22900 ^ n_21015;
assign n_22913 = n_22902 ^ n_21015;
assign n_22914 = n_22900 ^ n_22902;
assign n_22915 = n_22903 ^ n_22423;
assign n_22916 = n_22882 ^ n_22904;
assign n_22917 = ~n_22904 & n_22882;
assign n_22918 = n_22905 ^ x158;
assign n_22919 = n_22906 ^ n_22290;
assign n_22920 = n_22701 ^ n_22906;
assign n_22921 = n_22907 ^ n_22244;
assign n_22922 = n_22908 ^ x157;
assign n_22923 = n_22909 ^ n_21162;
assign n_22924 = n_22911 ^ x229;
assign n_22925 = n_22912 ^ n_22902;
assign n_22926 = n_22913 & ~n_22914;
assign n_22927 = n_22915 ^ n_22441;
assign n_22928 = n_22915 ^ n_22916;
assign n_22929 = n_22916 ^ n_22441;
assign n_22930 = n_22918 ^ n_22908;
assign n_22931 = n_22919 ^ n_21201;
assign n_22932 = n_22921 ^ n_22305;
assign n_22933 = n_22923 ^ n_21201;
assign n_22934 = n_22923 ^ n_22919;
assign n_22935 = n_22924 ^ n_22925;
assign n_22936 = n_22925 ^ x228;
assign n_22937 = n_22926 ^ n_21015;
assign n_22938 = n_22927 ^ n_22916;
assign n_22939 = n_22928 ^ n_21520;
assign n_22940 = n_22928 & ~n_22929;
assign n_22941 = n_22930 ^ x157;
assign n_22942 = ~n_22930 & n_22922;
assign n_22943 = n_22263 ^ n_22932;
assign n_22944 = ~n_22932 & ~n_22313;
assign n_22945 = n_22933 ^ n_22919;
assign n_22946 = n_22931 & ~n_22934;
assign n_22947 = n_22935 ^ x228;
assign n_22948 = n_22935 & ~n_22936;
assign n_22949 = n_22937 ^ n_21052;
assign n_22950 = n_22939 ^ n_21052;
assign n_22951 = n_22937 ^ n_22939;
assign n_22952 = n_22940 ^ n_22441;
assign n_22953 = n_22941 ^ n_22917;
assign n_22954 = ~n_22917 & n_22941;
assign n_22955 = n_22942 ^ x157;
assign n_22956 = n_22943 ^ n_22297;
assign n_22957 = n_22719 ^ n_22943;
assign n_22958 = n_22944 ^ n_22263;
assign n_22959 = n_22945 ^ x156;
assign n_22960 = n_22946 ^ n_21201;
assign n_22961 = n_22948 ^ x228;
assign n_22962 = n_22949 ^ n_22939;
assign n_22963 = n_22950 & n_22951;
assign n_22964 = n_22952 ^ n_22459;
assign n_22965 = n_22952 ^ n_22953;
assign n_22966 = n_22953 ^ n_22459;
assign n_22967 = n_22955 ^ n_22945;
assign n_22968 = n_22956 ^ n_21240;
assign n_22969 = n_22958 ^ n_22323;
assign n_22970 = n_22960 ^ n_21240;
assign n_22971 = n_22960 ^ n_22956;
assign n_22972 = n_22961 ^ n_22962;
assign n_22973 = n_22962 ^ x227;
assign n_22974 = n_22963 ^ n_21052;
assign n_22975 = n_22964 ^ n_22953;
assign n_22976 = n_22965 ^ n_21558;
assign n_22977 = ~n_22965 & ~n_22966;
assign n_22978 = n_22967 ^ x156;
assign n_22979 = ~n_22967 & n_22959;
assign n_22980 = n_22286 ^ n_22969;
assign n_22981 = n_22969 & ~n_22330;
assign n_22982 = n_22970 ^ n_22956;
assign n_22983 = ~n_22968 & ~n_22971;
assign n_22984 = n_22972 ^ x227;
assign n_22985 = n_22972 & ~n_22973;
assign n_22986 = n_22974 ^ n_21091;
assign n_22987 = n_22976 ^ n_21091;
assign n_22988 = n_22974 ^ n_22976;
assign n_22989 = n_22977 ^ n_22459;
assign n_22990 = n_22954 ^ n_22978;
assign n_22991 = ~n_22978 & ~n_22954;
assign n_22992 = n_22979 ^ x156;
assign n_22993 = n_22980 ^ n_22329;
assign n_22994 = n_22738 ^ n_22980;
assign n_22995 = n_22981 ^ n_22286;
assign n_22996 = n_22982 ^ x155;
assign n_22997 = n_22983 ^ n_21240;
assign n_22998 = n_22985 ^ x227;
assign n_22999 = n_22986 ^ n_22976;
assign n_23000 = n_22987 & ~n_22988;
assign n_23001 = n_22989 ^ n_22471;
assign n_23002 = n_22989 ^ n_22990;
assign n_23003 = n_22990 ^ n_22471;
assign n_23004 = n_22992 ^ n_22982;
assign n_23005 = n_22993 ^ n_21280;
assign n_23006 = n_22995 ^ n_22344;
assign n_23007 = n_22997 ^ n_21280;
assign n_23008 = n_22997 ^ n_22993;
assign n_23009 = n_22998 ^ n_22999;
assign n_23010 = n_22999 ^ x226;
assign n_23011 = n_23000 ^ n_21091;
assign n_23012 = n_23001 ^ n_22990;
assign n_23013 = n_23002 ^ n_21598;
assign n_23014 = n_23002 & n_23003;
assign n_23015 = n_23004 ^ x155;
assign n_23016 = n_23004 & ~n_22996;
assign n_23017 = n_22308 ^ n_23006;
assign n_23018 = n_23006 & n_22352;
assign n_23019 = n_23007 ^ n_22993;
assign n_23020 = ~n_23005 & ~n_23008;
assign n_23021 = n_23009 ^ x226;
assign n_23022 = ~n_23009 & n_23010;
assign n_23023 = n_23011 ^ n_21130;
assign n_23024 = n_23013 ^ n_21130;
assign n_23025 = n_23011 ^ n_23013;
assign n_23026 = n_23014 ^ n_22471;
assign n_23027 = n_22991 ^ n_23015;
assign n_23028 = ~n_23015 & ~n_22991;
assign n_23029 = n_23016 ^ x155;
assign n_23030 = n_23017 ^ n_22336;
assign n_23031 = n_22757 ^ n_23017;
assign n_23032 = n_23018 ^ n_22308;
assign n_23033 = n_23019 ^ x154;
assign n_23034 = n_23020 ^ n_21280;
assign n_23035 = n_23022 ^ x226;
assign n_23036 = n_23023 ^ n_23013;
assign n_23037 = ~n_23024 & ~n_23025;
assign n_23038 = n_23026 ^ n_22494;
assign n_23039 = n_23026 ^ n_23027;
assign n_23040 = n_23027 ^ n_22494;
assign n_23041 = n_23029 ^ n_23019;
assign n_23042 = n_23030 ^ n_21319;
assign n_23043 = n_23032 ^ n_22380;
assign n_23044 = n_23034 ^ n_21319;
assign n_23045 = n_23034 ^ n_23030;
assign n_23046 = n_23035 ^ n_23036;
assign n_23047 = n_23036 ^ x225;
assign n_23048 = n_23037 ^ n_21130;
assign n_23049 = n_23038 ^ n_23027;
assign n_23050 = n_23039 ^ n_21636;
assign n_23051 = n_23039 & n_23040;
assign n_23052 = n_23041 ^ x154;
assign n_23053 = ~n_23041 & n_23033;
assign n_23054 = n_23043 ^ n_22379;
assign n_23055 = n_22769 ^ n_23043;
assign n_23056 = n_23044 ^ n_23030;
assign n_23057 = ~n_23042 & ~n_23045;
assign n_23058 = n_23046 ^ x225;
assign n_23059 = n_23046 & ~n_23047;
assign n_23060 = n_23048 ^ n_21168;
assign n_23061 = n_23050 ^ n_21168;
assign n_23062 = n_23048 ^ n_23050;
assign n_23063 = n_23051 ^ n_22494;
assign n_23064 = n_23028 ^ n_23052;
assign n_23065 = n_23052 & n_23028;
assign n_23066 = n_23053 ^ x154;
assign n_23067 = n_23055 ^ n_22756;
assign n_23068 = n_23056 ^ x153;
assign n_23069 = n_23057 ^ n_21319;
assign n_23070 = ~n_23021 & n_23058;
assign n_23071 = n_23058 ^ n_23021;
assign n_23072 = n_23059 ^ x225;
assign n_23073 = n_23060 ^ n_23050;
assign n_23074 = ~n_23061 & n_23062;
assign n_23075 = n_23063 ^ n_22512;
assign n_23076 = n_23063 ^ n_23064;
assign n_23077 = n_23064 ^ n_22512;
assign n_23078 = n_23066 ^ n_23056;
assign n_23079 = n_23069 ^ x152;
assign n_23080 = n_23072 ^ n_23073;
assign n_23081 = n_23073 ^ x224;
assign n_23082 = n_23074 ^ n_21168;
assign n_23083 = n_23075 ^ n_23064;
assign n_23084 = n_23076 ^ n_21676;
assign n_23085 = ~n_23076 & ~n_23077;
assign n_23086 = n_23078 ^ x153;
assign n_23087 = n_23078 & ~n_23068;
assign n_23088 = n_23079 ^ n_23054;
assign n_23089 = n_23080 ^ x224;
assign n_23090 = ~n_23080 & n_23081;
assign n_23091 = n_23082 ^ n_21207;
assign n_23092 = n_23084 ^ n_21207;
assign n_23093 = n_23082 ^ n_23084;
assign n_23094 = n_23085 ^ n_22512;
assign n_23095 = n_23065 ^ n_23086;
assign n_23096 = n_23086 & ~n_23065;
assign n_23097 = n_23087 ^ x153;
assign n_23098 = ~n_23070 & n_23089;
assign n_23099 = n_23089 ^ n_23070;
assign n_23100 = n_23090 ^ x224;
assign n_23101 = n_23091 ^ n_23084;
assign n_23102 = ~n_23092 & n_23093;
assign n_23103 = n_23094 ^ n_22531;
assign n_23104 = n_23094 ^ n_23095;
assign n_23105 = n_23095 ^ n_22531;
assign n_23106 = n_23097 ^ n_23096;
assign n_23107 = n_23100 ^ n_23101;
assign n_23108 = n_23101 ^ x239;
assign n_23109 = n_23102 ^ n_21207;
assign n_23110 = n_23103 ^ n_23095;
assign n_23111 = n_23104 ^ n_21715;
assign n_23112 = n_23104 & n_23105;
assign n_23113 = n_23106 ^ n_23088;
assign n_23114 = n_23107 ^ x239;
assign n_23115 = ~n_23107 & n_23108;
assign n_23116 = n_23109 ^ n_21247;
assign n_23117 = n_23111 ^ n_21247;
assign n_23118 = n_23109 ^ n_23111;
assign n_23119 = n_23112 ^ n_22531;
assign n_23120 = n_23113 ^ n_22549;
assign n_23121 = ~n_23098 & ~n_23114;
assign n_23122 = n_23114 ^ n_23098;
assign n_23123 = n_23115 ^ x239;
assign n_23124 = n_23116 ^ n_23111;
assign n_23125 = n_23117 & n_23118;
assign n_23126 = n_23119 ^ n_23113;
assign n_23127 = n_23119 ^ n_22549;
assign n_23128 = n_23123 ^ n_23124;
assign n_23129 = n_23124 ^ x238;
assign n_23130 = n_23125 ^ n_21247;
assign n_23131 = ~n_23126 & ~n_23120;
assign n_23132 = n_23126 ^ n_21754;
assign n_23133 = n_23127 ^ n_23113;
assign n_23134 = n_23128 ^ x238;
assign n_23135 = n_23128 & ~n_23129;
assign n_23136 = n_23130 ^ n_21287;
assign n_23137 = n_23131 ^ n_22549;
assign n_23138 = n_23132 ^ n_21287;
assign n_23139 = n_23130 ^ n_23132;
assign n_23140 = n_23121 & n_23134;
assign n_23141 = n_23134 ^ n_23121;
assign n_23142 = n_23135 ^ x238;
assign n_23143 = n_23136 ^ n_23132;
assign n_23144 = n_23137 ^ n_22362;
assign n_23145 = n_22573 ^ n_23137;
assign n_23146 = ~n_23138 & n_23139;
assign n_23147 = n_23142 ^ n_23143;
assign n_23148 = n_23143 ^ x237;
assign n_23149 = ~n_23144 & ~n_22573;
assign n_23150 = n_23144 ^ n_21793;
assign n_23151 = n_23146 ^ n_21287;
assign n_23152 = n_23147 ^ x237;
assign n_23153 = n_23147 & ~n_23148;
assign n_23154 = n_23149 ^ n_22567;
assign n_23155 = n_23151 ^ n_21326;
assign n_23156 = n_23150 ^ n_23151;
assign n_23157 = ~n_23140 & ~n_23152;
assign n_23158 = n_23152 ^ n_23140;
assign n_23159 = n_23153 ^ x237;
assign n_23160 = n_23154 ^ n_22586;
assign n_23161 = n_23150 ^ n_23155;
assign n_23162 = n_23155 & ~n_23156;
assign n_23163 = n_23160 & ~n_22592;
assign n_23164 = n_22408 ^ n_23160;
assign n_23165 = n_23159 ^ n_23161;
assign n_23166 = n_23161 ^ x236;
assign n_23167 = n_23162 ^ n_21326;
assign n_23168 = n_23163 ^ n_22408;
assign n_23169 = n_23164 ^ n_22586;
assign n_23170 = n_23165 ^ x236;
assign n_23171 = ~n_23165 & n_23166;
assign n_23172 = n_23167 ^ n_21373;
assign n_23173 = n_23168 ^ n_22606;
assign n_23174 = n_23169 ^ n_21833;
assign n_23175 = ~n_23157 & ~n_23170;
assign n_23176 = n_23170 ^ n_23157;
assign n_23177 = n_23171 ^ x236;
assign n_23178 = n_23173 & n_22612;
assign n_23179 = n_22437 ^ n_23173;
assign n_23180 = n_23174 ^ n_21373;
assign n_23181 = n_23167 ^ n_23174;
assign n_23182 = n_23172 ^ n_23174;
assign n_23183 = n_23177 ^ x235;
assign n_23184 = n_23178 ^ n_22437;
assign n_23185 = n_23179 ^ n_22606;
assign n_23186 = n_23180 & n_23181;
assign n_23187 = n_23177 ^ n_23182;
assign n_23188 = n_23184 ^ n_22624;
assign n_23189 = n_23185 ^ n_21873;
assign n_23190 = n_23186 ^ n_21373;
assign n_23191 = ~n_23187 & n_23183;
assign n_23192 = n_23187 ^ x235;
assign n_23193 = n_23188 & ~n_22630;
assign n_23194 = n_22455 ^ n_23188;
assign n_23195 = n_23189 ^ n_21412;
assign n_23196 = n_23190 ^ n_23189;
assign n_23197 = n_23190 ^ n_21412;
assign n_23198 = n_23191 ^ x235;
assign n_23199 = ~n_23175 & n_23192;
assign n_23200 = n_23192 ^ n_23175;
assign n_23201 = n_23193 ^ n_22455;
assign n_23202 = n_23194 ^ n_22624;
assign n_23203 = ~n_23195 & ~n_23196;
assign n_23204 = n_23197 ^ n_23189;
assign n_23205 = n_23201 ^ n_22642;
assign n_23206 = n_23202 ^ n_21913;
assign n_23207 = n_23203 ^ n_21412;
assign n_23208 = n_23198 ^ n_23204;
assign n_23209 = n_23204 ^ x234;
assign n_23210 = ~n_23205 & ~n_22647;
assign n_23211 = n_22474 ^ n_23205;
assign n_23212 = n_23206 ^ n_21451;
assign n_23213 = n_23207 ^ n_23206;
assign n_23214 = n_23207 ^ n_21451;
assign n_23215 = n_23208 ^ x234;
assign n_23216 = ~n_23208 & n_23209;
assign n_23217 = n_23210 ^ n_22474;
assign n_23218 = n_23211 ^ n_22642;
assign n_23219 = ~n_23212 & n_23213;
assign n_23220 = n_23214 ^ n_23206;
assign n_23221 = n_23199 & n_23215;
assign n_23222 = n_23215 ^ n_23199;
assign n_23223 = n_23216 ^ x234;
assign n_23224 = n_23217 ^ n_22652;
assign n_23225 = n_23217 ^ n_22659;
assign n_23226 = n_23218 ^ n_21952;
assign n_23227 = n_23219 ^ n_21451;
assign n_23228 = n_23220 ^ x233;
assign n_23229 = n_23223 ^ n_23220;
assign n_23230 = ~n_22659 & n_23224;
assign n_23231 = n_23225 ^ n_22652;
assign n_23232 = n_22814 ^ n_23225;
assign n_23233 = n_23226 ^ n_21487;
assign n_23234 = n_23227 ^ n_23226;
assign n_23235 = n_23227 ^ n_21487;
assign n_23236 = n_23229 & ~n_23228;
assign n_23237 = n_23229 ^ x233;
assign n_23238 = n_23230 ^ n_22490;
assign n_23239 = n_23231 ^ n_21987;
assign n_23240 = n_23233 & n_23234;
assign n_23241 = n_23235 ^ n_23226;
assign n_23242 = n_23236 ^ x233;
assign n_23243 = ~n_23221 & n_23237;
assign n_23244 = n_23237 ^ n_23221;
assign n_23245 = n_23238 ^ n_22676;
assign n_23246 = n_23238 ^ n_22508;
assign n_23247 = n_23239 ^ n_21512;
assign n_23248 = n_23240 ^ n_21487;
assign n_23249 = n_23241 ^ x232;
assign n_23250 = n_23242 ^ n_23241;
assign n_23251 = ~n_22683 & n_23245;
assign n_23252 = n_23246 ^ n_22030;
assign n_23253 = n_23246 ^ n_22676;
assign n_23254 = n_23248 ^ n_23239;
assign n_23255 = ~n_23250 & n_23249;
assign n_23256 = n_23250 ^ x232;
assign n_23257 = n_23251 ^ n_22508;
assign n_23258 = n_23252 ^ n_21562;
assign n_23259 = n_22867 ^ n_23253;
assign n_23260 = ~n_23254 & ~n_23247;
assign n_23261 = n_23254 ^ n_21512;
assign n_23262 = n_23255 ^ x232;
assign n_23263 = ~n_23243 & n_23256;
assign n_23264 = n_23257 ^ n_22695;
assign n_23265 = n_23260 ^ n_21512;
assign n_23266 = n_23261 ^ x247;
assign n_23267 = n_23262 ^ n_23261;
assign n_23268 = n_23262 ^ x247;
assign n_23269 = ~n_23264 & ~n_22703;
assign n_23270 = n_22528 ^ n_23264;
assign n_23271 = n_23265 ^ n_23252;
assign n_23272 = n_23266 & ~n_23267;
assign n_23273 = n_23268 ^ n_23261;
assign n_23274 = n_23269 ^ n_22528;
assign n_23275 = n_23270 ^ n_22695;
assign n_23276 = n_22910 ^ n_23270;
assign n_23277 = ~n_23271 & ~n_23258;
assign n_23278 = n_23271 ^ n_21562;
assign n_23279 = n_23272 ^ x247;
assign n_23280 = ~n_23263 & ~n_23273;
assign n_23281 = n_23273 ^ n_23263;
assign n_23282 = n_23274 ^ n_22713;
assign n_23283 = n_23275 ^ n_22070;
assign n_23284 = n_23277 ^ n_21562;
assign n_23285 = n_23278 ^ x246;
assign n_23286 = n_23279 ^ n_23278;
assign n_23287 = n_23279 ^ x246;
assign n_23288 = ~n_23281 & ~n_22813;
assign n_23289 = n_23281 ^ n_22365;
assign n_23290 = n_23281 ^ n_22346;
assign n_23291 = n_22813 ^ n_23281;
assign n_23292 = n_23282 & n_22721;
assign n_23293 = n_22545 ^ n_23282;
assign n_23294 = n_23283 ^ n_21602;
assign n_23295 = n_23284 ^ n_23283;
assign n_23296 = ~n_23285 & n_23286;
assign n_23297 = n_23287 ^ n_23278;
assign n_23298 = n_22830 ^ n_23288;
assign n_23299 = n_21348 & n_23289;
assign n_23300 = x327 & n_23290;
assign n_23301 = n_23290 ^ x327;
assign n_23302 = n_23292 ^ n_22545;
assign n_23303 = n_23293 ^ n_22713;
assign n_23304 = n_22947 ^ n_23293;
assign n_23305 = n_23295 & ~n_23294;
assign n_23306 = n_23295 ^ n_21602;
assign n_23307 = n_23296 ^ x246;
assign n_23308 = n_23280 & n_23297;
assign n_23309 = n_23297 ^ n_23280;
assign n_23310 = n_23299 ^ n_21393;
assign n_23311 = n_23300 ^ x326;
assign n_23312 = n_23302 ^ n_22732;
assign n_23313 = n_23303 ^ n_22109;
assign n_23314 = n_23305 ^ n_21602;
assign n_23315 = n_23306 ^ x245;
assign n_23316 = n_23307 ^ n_23306;
assign n_23317 = n_23309 ^ n_23288;
assign n_23318 = n_23309 ^ n_23298;
assign n_23319 = ~n_23312 & n_22740;
assign n_23320 = n_22563 ^ n_23312;
assign n_23321 = n_23313 ^ n_21640;
assign n_23322 = n_23314 ^ n_23313;
assign n_23323 = n_23314 ^ n_21640;
assign n_23324 = ~n_23316 & n_23315;
assign n_23325 = n_23316 ^ x245;
assign n_23326 = n_23298 & n_23317;
assign n_23327 = n_23318 ^ n_22829;
assign n_23328 = n_23319 ^ n_22563;
assign n_23329 = n_23320 ^ n_22732;
assign n_23330 = n_22984 ^ n_23320;
assign n_23331 = n_23321 & ~n_23322;
assign n_23332 = n_23323 ^ n_23313;
assign n_23333 = n_23324 ^ x245;
assign n_23334 = n_23325 & ~n_23308;
assign n_23335 = n_23308 ^ n_23325;
assign n_23336 = n_23326 ^ n_22830;
assign n_23337 = n_23327 ^ n_23299;
assign n_23338 = n_23328 ^ n_22751;
assign n_23339 = n_23329 ^ n_22145;
assign n_23340 = n_23331 ^ n_21640;
assign n_23341 = n_23332 ^ x244;
assign n_23342 = n_23333 ^ n_23332;
assign n_23343 = n_22864 ^ n_23335;
assign n_23344 = n_23336 ^ n_23335;
assign n_23345 = n_23336 ^ n_22864;
assign n_23346 = n_23337 & ~n_23310;
assign n_23347 = n_23337 ^ n_21393;
assign n_23348 = ~n_23338 & n_22759;
assign n_23349 = n_22582 ^ n_23338;
assign n_23350 = n_23339 ^ n_21680;
assign n_23351 = n_23340 ^ n_23339;
assign n_23352 = n_23340 ^ n_21680;
assign n_23353 = n_23342 & ~n_23341;
assign n_23354 = n_23342 ^ x244;
assign n_23355 = ~n_23343 & n_23344;
assign n_23356 = n_23345 ^ n_23335;
assign n_23357 = n_23346 ^ n_21393;
assign n_23358 = n_23347 ^ n_23300;
assign n_23359 = n_23347 ^ n_23311;
assign n_23360 = n_23348 ^ n_22582;
assign n_23361 = n_23349 ^ n_22751;
assign n_23362 = n_23349 ^ n_23021;
assign n_23363 = ~n_23350 & n_23351;
assign n_23364 = n_23352 ^ n_23339;
assign n_23365 = n_23353 ^ x244;
assign n_23366 = n_23354 & ~n_23334;
assign n_23367 = n_23334 ^ n_23354;
assign n_23368 = n_23355 ^ n_22864;
assign n_23369 = n_23356 ^ n_22856;
assign n_23370 = n_23357 ^ n_21445;
assign n_23371 = n_23311 & ~n_23358;
assign n_23372 = n_23360 ^ n_22770;
assign n_23373 = n_23361 ^ n_22172;
assign n_23374 = n_23363 ^ n_21680;
assign n_23375 = n_23364 ^ x243;
assign n_23376 = n_23365 ^ n_23364;
assign n_23377 = n_22901 ^ n_23367;
assign n_23378 = n_23368 ^ n_23367;
assign n_23379 = n_23368 ^ n_22901;
assign n_23380 = n_23369 ^ n_21445;
assign n_23381 = n_23357 ^ n_23369;
assign n_23382 = n_23370 ^ n_23369;
assign n_23383 = n_23371 ^ x326;
assign n_23384 = ~n_23372 & n_22777;
assign n_23385 = n_22601 ^ n_23372;
assign n_23386 = n_23373 ^ n_21719;
assign n_23387 = n_23374 ^ n_23373;
assign n_23388 = n_23374 ^ n_21719;
assign n_23389 = ~n_23376 & n_23375;
assign n_23390 = n_23376 ^ x243;
assign n_23391 = n_23377 & ~n_23378;
assign n_23392 = n_23379 ^ n_23367;
assign n_23393 = n_23380 & n_23381;
assign n_23394 = n_23382 ^ x325;
assign n_23395 = n_23383 ^ n_23382;
assign n_23396 = n_23384 ^ n_22601;
assign n_23397 = n_23385 ^ n_22770;
assign n_23398 = n_23071 ^ n_23385;
assign n_23399 = ~n_23386 & ~n_23387;
assign n_23400 = n_23388 ^ n_23373;
assign n_23401 = n_23389 ^ x243;
assign n_23402 = ~n_23390 & n_23366;
assign n_23403 = n_23366 ^ n_23390;
assign n_23404 = n_23391 ^ n_22901;
assign n_23405 = n_23392 ^ n_22892;
assign n_23406 = n_23393 ^ n_21445;
assign n_23407 = n_23395 & ~n_23394;
assign n_23408 = n_23395 ^ x325;
assign n_23409 = n_23396 ^ n_22788;
assign n_23410 = n_23397 ^ n_22193;
assign n_23411 = n_23399 ^ n_21719;
assign n_23412 = n_23400 ^ x242;
assign n_23413 = n_23401 ^ n_23400;
assign n_23414 = n_22938 ^ n_23403;
assign n_23415 = n_23404 ^ n_23403;
assign n_23416 = n_23404 ^ n_22938;
assign n_23417 = n_23405 ^ n_21483;
assign n_23418 = n_23406 ^ n_23405;
assign n_23419 = n_23406 ^ n_21483;
assign n_23420 = n_23407 ^ x325;
assign n_23421 = n_22619 ^ n_23409;
assign n_23422 = ~n_23409 & n_22796;
assign n_23423 = n_23410 ^ n_21758;
assign n_23424 = n_23411 ^ n_23410;
assign n_23425 = n_23411 ^ n_21758;
assign n_23426 = ~n_23413 & n_23412;
assign n_23427 = n_23413 ^ x242;
assign n_23428 = n_23414 & ~n_23415;
assign n_23429 = n_23416 ^ n_23403;
assign n_23430 = ~n_23417 & n_23418;
assign n_23431 = n_23419 ^ n_23405;
assign n_23432 = n_23421 ^ n_22788;
assign n_23433 = n_23099 ^ n_23421;
assign n_23434 = n_23422 ^ n_22619;
assign n_23435 = n_23423 & n_23424;
assign n_23436 = n_23425 ^ n_23410;
assign n_23437 = n_23426 ^ x242;
assign n_23438 = n_23402 & ~n_23427;
assign n_23439 = n_23427 ^ n_23402;
assign n_23440 = n_23428 ^ n_22938;
assign n_23441 = n_23429 ^ n_22928;
assign n_23442 = n_23430 ^ n_21483;
assign n_23443 = n_23420 ^ n_23431;
assign n_23444 = n_23431 ^ x324;
assign n_23445 = n_23432 ^ n_22210;
assign n_23446 = n_23434 ^ n_22816;
assign n_23447 = n_23434 ^ n_22804;
assign n_23448 = n_23435 ^ n_21758;
assign n_23449 = n_23436 ^ x241;
assign n_23450 = n_23437 ^ n_23436;
assign n_23451 = n_22975 ^ n_23439;
assign n_23452 = n_23440 ^ n_23439;
assign n_23453 = n_23440 ^ n_22975;
assign n_23454 = n_23441 ^ n_21520;
assign n_23455 = n_23442 ^ n_23441;
assign n_23456 = n_23442 ^ n_21520;
assign n_23457 = n_23443 ^ x324;
assign n_23458 = n_23443 & ~n_23444;
assign n_23459 = n_23445 ^ n_21797;
assign n_23460 = n_23446 ^ n_22804;
assign n_23461 = n_23122 ^ n_23446;
assign n_23462 = ~n_22816 & ~n_23447;
assign n_23463 = n_23448 ^ n_23445;
assign n_23464 = n_23448 ^ n_21797;
assign n_23465 = ~n_23450 & n_23449;
assign n_23466 = n_23450 ^ x241;
assign n_23467 = n_23451 & ~n_23452;
assign n_23468 = n_23453 ^ n_23439;
assign n_23469 = n_23454 & n_23455;
assign n_23470 = n_23456 ^ n_23441;
assign n_23471 = n_23458 ^ x324;
assign n_23472 = n_23460 ^ n_22229;
assign n_23473 = n_23462 ^ n_22639;
assign n_23474 = ~n_23459 & ~n_23463;
assign n_23475 = n_23464 ^ n_23445;
assign n_23476 = n_23465 ^ x241;
assign n_23477 = n_23466 & ~n_23438;
assign n_23478 = n_23438 ^ n_23466;
assign n_23479 = n_23467 ^ n_22975;
assign n_23480 = n_23468 ^ n_22965;
assign n_23481 = n_23469 ^ n_21520;
assign n_23482 = n_23470 ^ x323;
assign n_23483 = n_23471 ^ n_23470;
assign n_23484 = n_23472 ^ n_21837;
assign n_23485 = n_23473 ^ n_22664;
assign n_23486 = n_23473 ^ n_22838;
assign n_23487 = n_23474 ^ n_21797;
assign n_23488 = n_23475 ^ x240;
assign n_23489 = n_23476 ^ n_23475;
assign n_23490 = n_23012 ^ n_23478;
assign n_23491 = n_23479 ^ n_23478;
assign n_23492 = n_23479 ^ n_23012;
assign n_23493 = n_23480 ^ n_21558;
assign n_23494 = n_23481 ^ n_23480;
assign n_23495 = n_23481 ^ n_21558;
assign n_23496 = ~n_23483 & n_23482;
assign n_23497 = n_23483 ^ x323;
assign n_23498 = n_23485 ^ n_22249;
assign n_23499 = n_23485 ^ n_22838;
assign n_23500 = n_22849 & n_23486;
assign n_23501 = n_23487 ^ n_23472;
assign n_23502 = ~n_23489 & n_23488;
assign n_23503 = n_23489 ^ x240;
assign n_23504 = ~n_23490 & n_23491;
assign n_23505 = n_23492 ^ n_23478;
assign n_23506 = n_23493 & n_23494;
assign n_23507 = n_23495 ^ n_23480;
assign n_23508 = n_23496 ^ x323;
assign n_23509 = n_23498 ^ n_21877;
assign n_23510 = n_23141 ^ n_23499;
assign n_23511 = n_23500 ^ n_22664;
assign n_23512 = n_23501 ^ n_21837;
assign n_23513 = n_23501 & n_23484;
assign n_23514 = n_23502 ^ x240;
assign n_23515 = ~n_23477 & ~n_23503;
assign n_23516 = n_23503 ^ n_23477;
assign n_23517 = n_23504 ^ n_23012;
assign n_23518 = n_23505 ^ n_23002;
assign n_23519 = n_23506 ^ n_21558;
assign n_23520 = n_23507 ^ x322;
assign n_23521 = n_23508 ^ n_23507;
assign n_23522 = n_23511 ^ n_22872;
assign n_23523 = n_23512 ^ x255;
assign n_23524 = n_23513 ^ n_21837;
assign n_23525 = n_23514 ^ n_23512;
assign n_23526 = n_23514 ^ x255;
assign n_23527 = n_23049 ^ n_23516;
assign n_23528 = n_23517 ^ n_23516;
assign n_23529 = n_23517 ^ n_23049;
assign n_23530 = n_23518 ^ n_21598;
assign n_23531 = n_23519 ^ n_23518;
assign n_23532 = n_23519 ^ n_21598;
assign n_23533 = n_23521 & ~n_23520;
assign n_23534 = n_23521 ^ x322;
assign n_23535 = n_22682 ^ n_23522;
assign n_23536 = ~n_23522 & n_22885;
assign n_23537 = n_23524 ^ n_23498;
assign n_23538 = n_23523 & ~n_23525;
assign n_23539 = n_23526 ^ n_23512;
assign n_23540 = n_23527 & n_23528;
assign n_23541 = n_23529 ^ n_23516;
assign n_23542 = ~n_23530 & ~n_23531;
assign n_23543 = n_23532 ^ n_23518;
assign n_23544 = n_23533 ^ x322;
assign n_23545 = ~n_23497 & n_23534;
assign n_23546 = n_23534 ^ n_23497;
assign n_23547 = n_23535 ^ n_22872;
assign n_23548 = n_23158 ^ n_23535;
assign n_23549 = n_23536 ^ n_22682;
assign n_23550 = n_23537 ^ n_21877;
assign n_23551 = ~n_23537 & n_23509;
assign n_23552 = n_23538 ^ x255;
assign n_23553 = ~n_23515 & n_23539;
assign n_23554 = n_23539 ^ n_23515;
assign n_23555 = n_23540 ^ n_23049;
assign n_23556 = n_23541 ^ n_23039;
assign n_23557 = n_23542 ^ n_21598;
assign n_23558 = n_23543 ^ x321;
assign n_23559 = n_23544 ^ n_23543;
assign n_23560 = n_23547 ^ n_22266;
assign n_23561 = n_23549 ^ n_22906;
assign n_23562 = n_23550 ^ x254;
assign n_23563 = n_23551 ^ n_21877;
assign n_23564 = n_23552 ^ n_23550;
assign n_23565 = n_23083 ^ n_23554;
assign n_23566 = n_23555 ^ n_23554;
assign n_23567 = n_23555 ^ n_23083;
assign n_23568 = n_23556 ^ n_21636;
assign n_23569 = n_23557 ^ n_23556;
assign n_23570 = n_23557 ^ n_21636;
assign n_23571 = n_23559 & ~n_23558;
assign n_23572 = n_23559 ^ x321;
assign n_23573 = n_23560 ^ n_21917;
assign n_23574 = n_22701 ^ n_23561;
assign n_23575 = ~n_23561 & ~n_22920;
assign n_23576 = n_23563 ^ n_23560;
assign n_23577 = n_23564 & ~n_23562;
assign n_23578 = n_23564 ^ x254;
assign n_23579 = n_23565 & ~n_23566;
assign n_23580 = n_23567 ^ n_23554;
assign n_23581 = n_23568 & ~n_23569;
assign n_23582 = n_23570 ^ n_23556;
assign n_23583 = n_23571 ^ x321;
assign n_23584 = n_23572 & n_23545;
assign n_23585 = n_23545 ^ n_23572;
assign n_23586 = n_23574 ^ n_22906;
assign n_23587 = n_23176 ^ n_23574;
assign n_23588 = n_23575 ^ n_22701;
assign n_23589 = n_23576 ^ n_21917;
assign n_23590 = n_23576 & ~n_23573;
assign n_23591 = n_23577 ^ x254;
assign n_23592 = n_23578 & ~n_23553;
assign n_23593 = n_23553 ^ n_23578;
assign n_23594 = n_23579 ^ n_23083;
assign n_23595 = n_23580 ^ n_23076;
assign n_23596 = n_23581 ^ n_21636;
assign n_23597 = n_23582 ^ x320;
assign n_23598 = n_23583 ^ n_23582;
assign n_23599 = n_23586 ^ n_22283;
assign n_23600 = n_23588 ^ n_22943;
assign n_23601 = n_23589 ^ x253;
assign n_23602 = n_23590 ^ n_21917;
assign n_23603 = n_23591 ^ n_23589;
assign n_23604 = n_23110 ^ n_23593;
assign n_23605 = n_23594 ^ n_23593;
assign n_23606 = n_23594 ^ n_23110;
assign n_23607 = n_23595 ^ n_21676;
assign n_23608 = n_23596 ^ n_23595;
assign n_23609 = n_23596 ^ n_21676;
assign n_23610 = n_23598 & ~n_23597;
assign n_23611 = n_23598 ^ x320;
assign n_23612 = n_23599 ^ n_21956;
assign n_23613 = n_22719 ^ n_23600;
assign n_23614 = n_23600 & n_22957;
assign n_23615 = n_23602 ^ n_21956;
assign n_23616 = n_23602 ^ n_23599;
assign n_23617 = ~n_23603 & n_23601;
assign n_23618 = n_23603 ^ x253;
assign n_23619 = ~n_23604 & n_23605;
assign n_23620 = n_23606 ^ n_23593;
assign n_23621 = ~n_23607 & ~n_23608;
assign n_23622 = n_23609 ^ n_23595;
assign n_23623 = n_23610 ^ x320;
assign n_23624 = ~n_23584 & ~n_23611;
assign n_23625 = n_23611 ^ n_23584;
assign n_23626 = n_23613 ^ n_22943;
assign n_23627 = n_23200 ^ n_23613;
assign n_23628 = n_23614 ^ n_22719;
assign n_23629 = n_23615 ^ n_23599;
assign n_23630 = ~n_23612 & n_23616;
assign n_23631 = n_23617 ^ x253;
assign n_23632 = ~n_23618 & n_23592;
assign n_23633 = n_23592 ^ n_23618;
assign n_23634 = n_23619 ^ n_23110;
assign n_23635 = n_23620 ^ n_23104;
assign n_23636 = n_23621 ^ n_21676;
assign n_23637 = n_23622 ^ x335;
assign n_23638 = n_23623 ^ n_23622;
assign n_23639 = n_23626 ^ n_22305;
assign n_23640 = n_23628 ^ n_22980;
assign n_23641 = n_23629 ^ x252;
assign n_23642 = n_23630 ^ n_21956;
assign n_23643 = n_23631 ^ n_23629;
assign n_23644 = n_23133 ^ n_23633;
assign n_23645 = n_23634 ^ n_23633;
assign n_23646 = n_23634 ^ n_23133;
assign n_23647 = n_23635 ^ n_21715;
assign n_23648 = n_23636 ^ n_23635;
assign n_23649 = n_23636 ^ n_21715;
assign n_23650 = ~n_23638 & n_23637;
assign n_23651 = n_23638 ^ x335;
assign n_23652 = n_23639 ^ n_21995;
assign n_23653 = n_22738 ^ n_23640;
assign n_23654 = n_23640 & ~n_22994;
assign n_23655 = n_23642 ^ n_21995;
assign n_23656 = n_23642 ^ n_23639;
assign n_23657 = ~n_23643 & n_23641;
assign n_23658 = n_23643 ^ x252;
assign n_23659 = ~n_23644 & n_23645;
assign n_23660 = n_23646 ^ n_23633;
assign n_23661 = n_23647 & n_23648;
assign n_23662 = n_23649 ^ n_23635;
assign n_23663 = n_23650 ^ x335;
assign n_23664 = n_23624 & n_23651;
assign n_23665 = n_23653 ^ n_22980;
assign n_23666 = n_23222 ^ n_23653;
assign n_23667 = n_23654 ^ n_22738;
assign n_23668 = n_23655 ^ n_23639;
assign n_23669 = ~n_23652 & n_23656;
assign n_23670 = n_23657 ^ x252;
assign n_23671 = ~n_23632 & n_23658;
assign n_23672 = n_23658 ^ n_23632;
assign n_23673 = n_23659 ^ n_23133;
assign n_23674 = n_23660 ^ n_23126;
assign n_23675 = n_23661 ^ n_21715;
assign n_23676 = n_23662 ^ x334;
assign n_23677 = n_23663 ^ n_23662;
assign n_23678 = n_23665 ^ n_22323;
assign n_23679 = n_23667 ^ n_23017;
assign n_23680 = n_23668 ^ x251;
assign n_23681 = n_23669 ^ n_21995;
assign n_23682 = n_23670 ^ n_23668;
assign n_23683 = n_23145 ^ n_23672;
assign n_23684 = n_23673 ^ n_23672;
assign n_23685 = n_23673 ^ n_23145;
assign n_23686 = n_23674 ^ n_21754;
assign n_23687 = n_23675 ^ n_23674;
assign n_23688 = n_23675 ^ n_21754;
assign n_23689 = ~n_23677 & n_23676;
assign n_23690 = n_23677 ^ x334;
assign n_23691 = n_23678 ^ n_22035;
assign n_23692 = n_22757 ^ n_23679;
assign n_23693 = ~n_23679 & n_23031;
assign n_23694 = n_23681 ^ n_22035;
assign n_23695 = n_23681 ^ n_23678;
assign n_23696 = ~n_23682 & n_23680;
assign n_23697 = n_23682 ^ x251;
assign n_23698 = ~n_23683 & ~n_23684;
assign n_23699 = n_23685 ^ n_23672;
assign n_23700 = ~n_23686 & n_23687;
assign n_23701 = n_23688 ^ n_23674;
assign n_23702 = n_23689 ^ x334;
assign n_23703 = n_23664 & n_23690;
assign n_23704 = n_23690 ^ n_23664;
assign n_23705 = n_23692 ^ n_23017;
assign n_23706 = n_23244 ^ n_23692;
assign n_23707 = n_23693 ^ n_22757;
assign n_23708 = n_23694 ^ n_23678;
assign n_23709 = n_23691 & ~n_23695;
assign n_23710 = n_23696 ^ x251;
assign n_23711 = ~n_23697 & ~n_23671;
assign n_23712 = n_23671 ^ n_23697;
assign n_23713 = n_23698 ^ n_23145;
assign n_23714 = n_23699 ^ n_23144;
assign n_23715 = n_23700 ^ n_21754;
assign n_23716 = n_23701 ^ x333;
assign n_23717 = n_23702 ^ n_23701;
assign n_23718 = n_23704 & n_23291;
assign n_23719 = n_23704 ^ n_22813;
assign n_23720 = n_23704 ^ n_22794;
assign n_23721 = n_23291 ^ n_23704;
assign n_23722 = n_23705 ^ n_22344;
assign n_23723 = n_23707 ^ n_23067;
assign n_23724 = n_23708 ^ x250;
assign n_23725 = n_23709 ^ n_22035;
assign n_23726 = n_23710 ^ n_23708;
assign n_23727 = n_23712 ^ n_23164;
assign n_23728 = n_23713 ^ n_23712;
assign n_23729 = n_23713 ^ n_23164;
assign n_23730 = n_23714 ^ n_21793;
assign n_23731 = n_23715 ^ n_23714;
assign n_23732 = n_23715 ^ n_21793;
assign n_23733 = ~n_23717 & n_23716;
assign n_23734 = n_23717 ^ x333;
assign n_23735 = n_23718 ^ n_23318;
assign n_23736 = ~n_22365 & ~n_23719;
assign n_23737 = x423 & n_23720;
assign n_23738 = n_23720 ^ x423;
assign n_23739 = n_23722 ^ n_22074;
assign n_23740 = n_23723 ^ n_23043;
assign n_23741 = n_23723 ^ n_23243;
assign n_23742 = n_23725 ^ n_22074;
assign n_23743 = n_23725 ^ n_23722;
assign n_23744 = n_23726 ^ x250;
assign n_23745 = n_23726 & ~n_23724;
assign n_23746 = n_23727 & n_23728;
assign n_23747 = n_23729 ^ n_23712;
assign n_23748 = n_23730 & n_23731;
assign n_23749 = n_23732 ^ n_23714;
assign n_23750 = n_23733 ^ x333;
assign n_23751 = ~n_23703 & ~n_23734;
assign n_23752 = n_23734 ^ n_23703;
assign n_23753 = n_23736 ^ n_22381;
assign n_23754 = n_23737 ^ x422;
assign n_23755 = n_23740 ^ n_22360;
assign n_23756 = n_23741 ^ n_23256;
assign n_23757 = n_23742 ^ n_23722;
assign n_23758 = n_23739 & ~n_23743;
assign n_23759 = n_23744 & n_23711;
assign n_23760 = n_23711 ^ n_23744;
assign n_23761 = n_23745 ^ x250;
assign n_23762 = n_23746 ^ n_23164;
assign n_23763 = n_23747 ^ n_23169;
assign n_23764 = n_23748 ^ n_21793;
assign n_23765 = n_23749 ^ x332;
assign n_23766 = n_23750 ^ n_23749;
assign n_23767 = n_23752 ^ n_23718;
assign n_23768 = n_23735 ^ n_23752;
assign n_23769 = n_23755 ^ n_22113;
assign n_23770 = n_23757 ^ x249;
assign n_23771 = n_23758 ^ n_22074;
assign n_23772 = n_23760 ^ n_23179;
assign n_23773 = n_23761 ^ n_23757;
assign n_23774 = n_23762 ^ n_23760;
assign n_23775 = n_23762 ^ n_23179;
assign n_23776 = n_23763 ^ n_21833;
assign n_23777 = n_23764 ^ n_23763;
assign n_23778 = n_23764 ^ n_21833;
assign n_23779 = n_23766 & ~n_23765;
assign n_23780 = n_23766 ^ x332;
assign n_23781 = n_23767 & ~n_23735;
assign n_23782 = n_23767 ^ n_22830;
assign n_23783 = n_23771 ^ x248;
assign n_23784 = n_23773 ^ x249;
assign n_23785 = n_23773 & ~n_23770;
assign n_23786 = ~n_23772 & ~n_23774;
assign n_23787 = n_23775 ^ n_23760;
assign n_23788 = ~n_23776 & ~n_23777;
assign n_23789 = n_23778 ^ n_23763;
assign n_23790 = n_23779 ^ x332;
assign n_23791 = n_23751 & n_23780;
assign n_23792 = n_23780 ^ n_23751;
assign n_23793 = n_23781 ^ n_23318;
assign n_23794 = n_23782 ^ n_23736;
assign n_23795 = n_23783 ^ n_23769;
assign n_23796 = n_23759 ^ n_23784;
assign n_23797 = n_23784 & n_23759;
assign n_23798 = n_23785 ^ x249;
assign n_23799 = n_23786 ^ n_23179;
assign n_23800 = n_23787 ^ n_23185;
assign n_23801 = n_23788 ^ n_21833;
assign n_23802 = n_23789 ^ x331;
assign n_23803 = n_23790 ^ n_23789;
assign n_23804 = n_23792 ^ n_23356;
assign n_23805 = n_23793 ^ n_23792;
assign n_23806 = n_23793 ^ n_23356;
assign n_23807 = n_23794 & n_23753;
assign n_23808 = n_23794 ^ n_22381;
assign n_23809 = n_23796 ^ n_23194;
assign n_23810 = n_23798 ^ n_23797;
assign n_23811 = n_23799 ^ n_23796;
assign n_23812 = n_23799 ^ n_23194;
assign n_23813 = n_23800 ^ n_21873;
assign n_23814 = n_23801 ^ n_23800;
assign n_23815 = n_23801 ^ n_21873;
assign n_23816 = n_23803 & ~n_23802;
assign n_23817 = n_23803 ^ x331;
assign n_23818 = ~n_23805 & n_23804;
assign n_23819 = n_23805 ^ n_22864;
assign n_23820 = n_23806 ^ n_23792;
assign n_23821 = n_23807 ^ n_22381;
assign n_23822 = n_23808 ^ n_23737;
assign n_23823 = n_23808 ^ n_23754;
assign n_23824 = n_23810 ^ n_23795;
assign n_23825 = ~n_23809 & n_23811;
assign n_23826 = n_23812 ^ n_23796;
assign n_23827 = ~n_23813 & ~n_23814;
assign n_23828 = n_23815 ^ n_23800;
assign n_23829 = n_23816 ^ x331;
assign n_23830 = n_23817 & n_23791;
assign n_23831 = n_23791 ^ n_23817;
assign n_23832 = n_23818 ^ n_23356;
assign n_23833 = n_23819 ^ n_22410;
assign n_23834 = n_23821 ^ n_23819;
assign n_23835 = n_23821 ^ n_22410;
assign n_23836 = n_23754 & n_23822;
assign n_23837 = n_23824 ^ n_23211;
assign n_23838 = n_23825 ^ n_23194;
assign n_23839 = n_23826 ^ n_23202;
assign n_23840 = n_23827 ^ n_21873;
assign n_23841 = n_23828 ^ x330;
assign n_23842 = n_23829 ^ n_23828;
assign n_23843 = n_23831 ^ n_23392;
assign n_23844 = n_23832 ^ n_23831;
assign n_23845 = n_23832 ^ n_23392;
assign n_23846 = ~n_23833 & ~n_23834;
assign n_23847 = n_23835 ^ n_23819;
assign n_23848 = n_23836 ^ x422;
assign n_23849 = n_23838 ^ n_23211;
assign n_23850 = n_23838 ^ n_23824;
assign n_23851 = n_23839 ^ n_21913;
assign n_23852 = n_23840 ^ n_23839;
assign n_23853 = n_23840 ^ n_21913;
assign n_23854 = ~n_23842 & n_23841;
assign n_23855 = n_23842 ^ x330;
assign n_23856 = ~n_23844 & ~n_23843;
assign n_23857 = n_23844 ^ n_22901;
assign n_23858 = n_23845 ^ n_23831;
assign n_23859 = n_23846 ^ n_22410;
assign n_23860 = n_23847 ^ x421;
assign n_23861 = n_23848 ^ n_23847;
assign n_23862 = n_23849 ^ n_23824;
assign n_23863 = n_23837 & ~n_23850;
assign n_23864 = n_23851 & n_23852;
assign n_23865 = n_23853 ^ n_23839;
assign n_23866 = n_23854 ^ x330;
assign n_23867 = ~n_23855 & n_23830;
assign n_23868 = n_23830 ^ n_23855;
assign n_23869 = n_23856 ^ n_23392;
assign n_23870 = n_23857 ^ n_22423;
assign n_23871 = n_23859 ^ n_23857;
assign n_23872 = n_23859 ^ n_22423;
assign n_23873 = n_23861 & ~n_23860;
assign n_23874 = n_23861 ^ x421;
assign n_23875 = n_23862 ^ n_23218;
assign n_23876 = n_23863 ^ n_23211;
assign n_23877 = n_23864 ^ n_21913;
assign n_23878 = n_23865 ^ x329;
assign n_23879 = n_23866 ^ n_23865;
assign n_23880 = n_23868 ^ n_23429;
assign n_23881 = n_23869 ^ n_23868;
assign n_23882 = n_23869 ^ n_23429;
assign n_23883 = ~n_23870 & n_23871;
assign n_23884 = n_23872 ^ n_23857;
assign n_23885 = n_23873 ^ x421;
assign n_23886 = n_23874 & n_23823;
assign n_23887 = n_23823 ^ n_23874;
assign n_23888 = n_23875 ^ n_21952;
assign n_23889 = n_23876 ^ n_23232;
assign n_23890 = n_23876 ^ n_23225;
assign n_23891 = n_23877 ^ n_23875;
assign n_23892 = n_23877 ^ n_21952;
assign n_23893 = ~n_23879 & n_23878;
assign n_23894 = n_23879 ^ x329;
assign n_23895 = ~n_23881 & n_23880;
assign n_23896 = n_23881 ^ n_22938;
assign n_23897 = n_23882 ^ n_23868;
assign n_23898 = n_23883 ^ n_22423;
assign n_23899 = n_23884 ^ x420;
assign n_23900 = n_23885 ^ n_23884;
assign n_23901 = n_23889 ^ n_23231;
assign n_23902 = ~n_23232 & n_23890;
assign n_23903 = ~n_23888 & ~n_23891;
assign n_23904 = n_23892 ^ n_23875;
assign n_23905 = n_23893 ^ x329;
assign n_23906 = n_23894 & ~n_23867;
assign n_23907 = n_23867 ^ n_23894;
assign n_23908 = n_23895 ^ n_23429;
assign n_23909 = n_23738 ^ n_23897;
assign n_23910 = n_23898 ^ n_22441;
assign n_23911 = n_23896 ^ n_23898;
assign n_23912 = ~n_23900 & n_23899;
assign n_23913 = n_23900 ^ x420;
assign n_23914 = n_23901 ^ n_21987;
assign n_23915 = n_23902 ^ n_22814;
assign n_23916 = n_23903 ^ n_21952;
assign n_23917 = n_23904 ^ x328;
assign n_23918 = n_23905 ^ n_23904;
assign n_23919 = n_23907 ^ n_23468;
assign n_23920 = n_23908 ^ n_23907;
assign n_23921 = n_23908 ^ n_23468;
assign n_23922 = n_23896 ^ n_23910;
assign n_23923 = n_23910 & n_23911;
assign n_23924 = n_23912 ^ x420;
assign n_23925 = ~n_23886 & n_23913;
assign n_23926 = n_23913 ^ n_23886;
assign n_23927 = n_23915 ^ n_22867;
assign n_23928 = n_23915 ^ n_23253;
assign n_23929 = n_23916 ^ n_23901;
assign n_23930 = ~n_23918 & n_23917;
assign n_23931 = n_23918 ^ x328;
assign n_23932 = n_23920 & ~n_23919;
assign n_23933 = n_23920 ^ n_22975;
assign n_23934 = n_23921 ^ n_23907;
assign n_23935 = n_23922 ^ x419;
assign n_23936 = n_23923 ^ n_22441;
assign n_23937 = n_23924 ^ n_23922;
assign n_23938 = n_23927 ^ n_23253;
assign n_23939 = n_23259 & n_23928;
assign n_23940 = n_23929 ^ n_21987;
assign n_23941 = n_23929 & n_23914;
assign n_23942 = n_23930 ^ x328;
assign n_23943 = ~n_23931 & ~n_23906;
assign n_23944 = n_23906 ^ n_23931;
assign n_23945 = n_23932 ^ n_23468;
assign n_23946 = n_23933 ^ n_22459;
assign n_23947 = n_23934 ^ n_23823;
assign n_23948 = n_23936 ^ n_23933;
assign n_23949 = n_23936 ^ n_22459;
assign n_23950 = ~n_23937 & n_23935;
assign n_23951 = n_23937 ^ x419;
assign n_23952 = n_23938 ^ n_23246;
assign n_23953 = n_23939 ^ n_22867;
assign n_23954 = n_23940 ^ x343;
assign n_23955 = n_23941 ^ n_21987;
assign n_23956 = n_23942 ^ n_23940;
assign n_23957 = n_23942 ^ x343;
assign n_23958 = n_23944 ^ n_23505;
assign n_23959 = n_23945 ^ n_23944;
assign n_23960 = n_23945 ^ n_23505;
assign n_23961 = ~n_23946 & ~n_23948;
assign n_23962 = n_23949 ^ n_23933;
assign n_23963 = n_23950 ^ x419;
assign n_23964 = n_23925 & n_23951;
assign n_23965 = n_23951 ^ n_23925;
assign n_23966 = n_23952 ^ n_22030;
assign n_23967 = n_23953 ^ n_22910;
assign n_23968 = n_23953 ^ n_23270;
assign n_23969 = n_23955 ^ n_23952;
assign n_23970 = n_23954 & ~n_23956;
assign n_23971 = n_23957 ^ n_23940;
assign n_23972 = n_23959 & n_23958;
assign n_23973 = n_23959 ^ n_23012;
assign n_23974 = n_23960 ^ n_23944;
assign n_23975 = n_23961 ^ n_22459;
assign n_23976 = n_23963 ^ n_23962;
assign n_23977 = n_23963 ^ x418;
assign n_23978 = n_23967 ^ n_23270;
assign n_23979 = ~n_23276 & ~n_23968;
assign n_23980 = n_23969 ^ n_22030;
assign n_23981 = n_23969 & n_23966;
assign n_23982 = n_23970 ^ x343;
assign n_23983 = ~n_23971 & n_23943;
assign n_23984 = n_23943 ^ n_23971;
assign n_23985 = n_23972 ^ n_23505;
assign n_23986 = n_23973 ^ n_22471;
assign n_23987 = n_23887 ^ n_23974;
assign n_23988 = n_23975 ^ n_23973;
assign n_23989 = n_23975 ^ n_22471;
assign n_23990 = n_23976 ^ x418;
assign n_23991 = ~n_23976 & n_23977;
assign n_23992 = n_23978 ^ n_23275;
assign n_23993 = n_23979 ^ n_22910;
assign n_23994 = n_23980 ^ x342;
assign n_23995 = n_23981 ^ n_22030;
assign n_23996 = n_23982 ^ n_23980;
assign n_23997 = n_23984 ^ n_23541;
assign n_23998 = n_23985 ^ n_23984;
assign n_23999 = n_23985 ^ n_23541;
assign n_24000 = n_23986 & n_23988;
assign n_24001 = n_23989 ^ n_23973;
assign n_24002 = n_23964 & n_23990;
assign n_24003 = n_23990 ^ n_23964;
assign n_24004 = n_23991 ^ x418;
assign n_24005 = n_23992 ^ n_22070;
assign n_24006 = n_23993 ^ n_23293;
assign n_24007 = n_23995 ^ n_23992;
assign n_24008 = n_23996 & ~n_23994;
assign n_24009 = n_23996 ^ x342;
assign n_24010 = n_23998 & n_23997;
assign n_24011 = n_23998 ^ n_23049;
assign n_24012 = n_23999 ^ n_23984;
assign n_24013 = n_24000 ^ n_22471;
assign n_24014 = n_24001 ^ x417;
assign n_24015 = n_24004 ^ n_24001;
assign n_24016 = n_22947 ^ n_24006;
assign n_24017 = n_24006 & n_23304;
assign n_24018 = n_24007 ^ n_22070;
assign n_24019 = n_24007 & n_24005;
assign n_24020 = n_24008 ^ x342;
assign n_24021 = n_23983 & n_24009;
assign n_24022 = n_24009 ^ n_23983;
assign n_24023 = n_24010 ^ n_23541;
assign n_24024 = n_24011 ^ n_22494;
assign n_24025 = n_23926 ^ n_24012;
assign n_24026 = n_24013 ^ n_24011;
assign n_24027 = n_24013 ^ n_22494;
assign n_24028 = ~n_24015 & n_24014;
assign n_24029 = n_24015 ^ x417;
assign n_24030 = n_24016 ^ n_23303;
assign n_24031 = n_24017 ^ n_22947;
assign n_24032 = n_24018 ^ x341;
assign n_24033 = n_24019 ^ n_22070;
assign n_24034 = n_24020 ^ n_24018;
assign n_24035 = n_24022 ^ n_23580;
assign n_24036 = n_24023 ^ n_24022;
assign n_24037 = n_24023 ^ n_23580;
assign n_24038 = n_24024 & n_24026;
assign n_24039 = n_24027 ^ n_24011;
assign n_24040 = n_24028 ^ x417;
assign n_24041 = ~n_24002 & ~n_24029;
assign n_24042 = n_24029 ^ n_24002;
assign n_24043 = n_24030 ^ n_22109;
assign n_24044 = n_24031 ^ n_23320;
assign n_24045 = n_24033 ^ n_22109;
assign n_24046 = n_24033 ^ n_24030;
assign n_24047 = ~n_24034 & n_24032;
assign n_24048 = n_24034 ^ x341;
assign n_24049 = n_24036 & n_24035;
assign n_24050 = n_24036 ^ n_23083;
assign n_24051 = n_24037 ^ n_24022;
assign n_24052 = n_24038 ^ n_22494;
assign n_24053 = n_24039 ^ x416;
assign n_24054 = n_24040 ^ n_24039;
assign n_24055 = n_22984 ^ n_24044;
assign n_24056 = n_24044 & ~n_23330;
assign n_24057 = n_24045 ^ n_24030;
assign n_24058 = ~n_24043 & ~n_24046;
assign n_24059 = n_24047 ^ x341;
assign n_24060 = n_24021 & ~n_24048;
assign n_24061 = n_24048 ^ n_24021;
assign n_24062 = n_24049 ^ n_23580;
assign n_24063 = n_24050 ^ n_22512;
assign n_24064 = n_23965 ^ n_24051;
assign n_24065 = n_24052 ^ n_24050;
assign n_24066 = n_24052 ^ n_22512;
assign n_24067 = n_24054 & ~n_24053;
assign n_24068 = n_24054 ^ x416;
assign n_24069 = n_24055 ^ n_23329;
assign n_24070 = n_24056 ^ n_22984;
assign n_24071 = n_24057 ^ x340;
assign n_24072 = n_24058 ^ n_22109;
assign n_24073 = n_24059 ^ n_24057;
assign n_24074 = n_24061 ^ n_23620;
assign n_24075 = n_24062 ^ n_24061;
assign n_24076 = n_24062 ^ n_23620;
assign n_24077 = ~n_24063 & ~n_24065;
assign n_24078 = n_24066 ^ n_24050;
assign n_24079 = n_24067 ^ x416;
assign n_24080 = n_24041 & n_24068;
assign n_24081 = n_24068 ^ n_24041;
assign n_24082 = n_24069 ^ n_22145;
assign n_24083 = n_24070 ^ n_23362;
assign n_24084 = n_24070 ^ n_23021;
assign n_24085 = n_24072 ^ n_22145;
assign n_24086 = n_24072 ^ n_24069;
assign n_24087 = ~n_24073 & n_24071;
assign n_24088 = n_24073 ^ x340;
assign n_24089 = n_24075 & n_24074;
assign n_24090 = n_24075 ^ n_23110;
assign n_24091 = n_24076 ^ n_24061;
assign n_24092 = n_24077 ^ n_22512;
assign n_24093 = n_24078 ^ x431;
assign n_24094 = n_24079 ^ n_24078;
assign n_24095 = n_24083 ^ n_23361;
assign n_24096 = ~n_23362 & ~n_24084;
assign n_24097 = n_24085 ^ n_24069;
assign n_24098 = n_24082 & ~n_24086;
assign n_24099 = n_24087 ^ x340;
assign n_24100 = n_24060 & ~n_24088;
assign n_24101 = n_24088 ^ n_24060;
assign n_24102 = n_24089 ^ n_23620;
assign n_24103 = n_24090 ^ n_22531;
assign n_24104 = n_24003 ^ n_24091;
assign n_24105 = n_24092 ^ n_24090;
assign n_24106 = n_24092 ^ n_22531;
assign n_24107 = n_24094 & ~n_24093;
assign n_24108 = n_24094 ^ x431;
assign n_24109 = n_24096 ^ n_23349;
assign n_24110 = n_24097 ^ x339;
assign n_24111 = n_24098 ^ n_22145;
assign n_24112 = n_24099 ^ n_24097;
assign n_24113 = n_24101 ^ n_23660;
assign n_24114 = n_24102 ^ n_24101;
assign n_24115 = n_24102 ^ n_23660;
assign n_24116 = n_24103 & n_24105;
assign n_24117 = n_24106 ^ n_24090;
assign n_24118 = n_24107 ^ x431;
assign n_24119 = ~n_24080 & ~n_24108;
assign n_24120 = n_24108 ^ n_24080;
assign n_24121 = n_24109 ^ n_23385;
assign n_24122 = n_24111 ^ n_22172;
assign n_24123 = n_24095 ^ n_24111;
assign n_24124 = ~n_24112 & n_24110;
assign n_24125 = n_24112 ^ x339;
assign n_24126 = ~n_24114 & n_24113;
assign n_24127 = n_24114 ^ n_23133;
assign n_24128 = n_24115 ^ n_24101;
assign n_24129 = n_24116 ^ n_22531;
assign n_24130 = n_24117 ^ x430;
assign n_24131 = n_24118 ^ n_24117;
assign n_24132 = n_23071 ^ n_24121;
assign n_24133 = ~n_24121 & n_23398;
assign n_24134 = n_24095 ^ n_24122;
assign n_24135 = ~n_24122 & ~n_24123;
assign n_24136 = n_24124 ^ x339;
assign n_24137 = ~n_24125 & n_24100;
assign n_24138 = n_24100 ^ n_24125;
assign n_24139 = n_24126 ^ n_23660;
assign n_24140 = n_24127 ^ n_22549;
assign n_24141 = n_24042 ^ n_24128;
assign n_24142 = n_24129 ^ n_24127;
assign n_24143 = n_24129 ^ n_22549;
assign n_24144 = n_24131 & ~n_24130;
assign n_24145 = n_24131 ^ x430;
assign n_24146 = n_24132 ^ n_23397;
assign n_24147 = n_24133 ^ n_23071;
assign n_24148 = n_24134 ^ x338;
assign n_24149 = n_24135 ^ n_22172;
assign n_24150 = n_24136 ^ n_24134;
assign n_24151 = n_24138 ^ n_23699;
assign n_24152 = n_24139 ^ n_24138;
assign n_24153 = n_24139 ^ n_23699;
assign n_24154 = n_24140 & n_24142;
assign n_24155 = n_24143 ^ n_24127;
assign n_24156 = n_24144 ^ x430;
assign n_24157 = n_24145 & ~n_24119;
assign n_24158 = n_24119 ^ n_24145;
assign n_24159 = n_24146 ^ n_22193;
assign n_24160 = n_24147 ^ n_23421;
assign n_24161 = n_24149 ^ n_22193;
assign n_24162 = n_24149 ^ n_24146;
assign n_24163 = n_24150 & ~n_24148;
assign n_24164 = n_24150 ^ x338;
assign n_24165 = ~n_24152 & n_24151;
assign n_24166 = n_24152 ^ n_23145;
assign n_24167 = n_24153 ^ n_24138;
assign n_24168 = n_24154 ^ n_22549;
assign n_24169 = n_24155 ^ x429;
assign n_24170 = n_24156 ^ n_24155;
assign n_24171 = n_23099 ^ n_24160;
assign n_24172 = ~n_24160 & ~n_23433;
assign n_24173 = n_24161 ^ n_24146;
assign n_24174 = ~n_24159 & n_24162;
assign n_24175 = n_24163 ^ x338;
assign n_24176 = n_24164 & n_24137;
assign n_24177 = n_24137 ^ n_24164;
assign n_24178 = n_24165 ^ n_23699;
assign n_24179 = n_24166 ^ n_22567;
assign n_24180 = n_24081 ^ n_24167;
assign n_24181 = n_24168 ^ n_24166;
assign n_24182 = n_24168 ^ n_22567;
assign n_24183 = ~n_24170 & n_24169;
assign n_24184 = n_24170 ^ x429;
assign n_24185 = n_24171 ^ n_23432;
assign n_24186 = n_23301 ^ n_24171;
assign n_24187 = n_24172 ^ n_23099;
assign n_24188 = n_24174 ^ n_22193;
assign n_24189 = n_24175 ^ n_24173;
assign n_24190 = n_24175 ^ x337;
assign n_24191 = n_24177 ^ n_23747;
assign n_24192 = n_24178 ^ n_24177;
assign n_24193 = n_24178 ^ n_23747;
assign n_24194 = n_24179 & n_24181;
assign n_24195 = n_24182 ^ n_24166;
assign n_24196 = n_24183 ^ x429;
assign n_24197 = ~n_24184 & n_24157;
assign n_24198 = n_24157 ^ n_24184;
assign n_24199 = n_24185 ^ n_22210;
assign n_24200 = n_24187 ^ n_23446;
assign n_24201 = n_24188 ^ n_22210;
assign n_24202 = n_24188 ^ n_24185;
assign n_24203 = n_24189 ^ x337;
assign n_24204 = ~n_24189 & n_24190;
assign n_24205 = ~n_24191 & n_24192;
assign n_24206 = n_24192 ^ n_23164;
assign n_24207 = n_24193 ^ n_24177;
assign n_24208 = n_24194 ^ n_22567;
assign n_24209 = n_24195 ^ x428;
assign n_24210 = n_24196 ^ n_24195;
assign n_24211 = n_23122 ^ n_24200;
assign n_24212 = ~n_24200 & n_23461;
assign n_24213 = n_24201 ^ n_24185;
assign n_24214 = n_24199 & ~n_24202;
assign n_24215 = ~n_24176 & n_24203;
assign n_24216 = n_24203 ^ n_24176;
assign n_24217 = n_24204 ^ x337;
assign n_24218 = n_24205 ^ n_23747;
assign n_24219 = n_24206 ^ n_22586;
assign n_24220 = n_24120 ^ n_24207;
assign n_24221 = n_24208 ^ n_24206;
assign n_24222 = n_24208 ^ n_22586;
assign n_24223 = n_24210 & ~n_24209;
assign n_24224 = n_24210 ^ x428;
assign n_24225 = n_24211 ^ n_23460;
assign n_24226 = n_23359 ^ n_24211;
assign n_24227 = n_24212 ^ n_23122;
assign n_24228 = n_24213 ^ x336;
assign n_24229 = n_24214 ^ n_22210;
assign n_24230 = n_24216 ^ n_23787;
assign n_24231 = n_24217 ^ n_24213;
assign n_24232 = n_24218 ^ n_24216;
assign n_24233 = n_24218 ^ n_23787;
assign n_24234 = ~n_24219 & ~n_24221;
assign n_24235 = n_24222 ^ n_24206;
assign n_24236 = n_24223 ^ x428;
assign n_24237 = n_24197 & n_24224;
assign n_24238 = n_24224 ^ n_24197;
assign n_24239 = n_24225 ^ n_22229;
assign n_24240 = n_24227 ^ n_23141;
assign n_24241 = n_24227 ^ n_23499;
assign n_24242 = n_24229 ^ n_24225;
assign n_24243 = n_24231 ^ x336;
assign n_24244 = n_24231 & ~n_24228;
assign n_24245 = ~n_24230 & n_24232;
assign n_24246 = n_24232 ^ n_23179;
assign n_24247 = n_24233 ^ n_24216;
assign n_24248 = n_24234 ^ n_22586;
assign n_24249 = n_24235 ^ x427;
assign n_24250 = n_24236 ^ n_24235;
assign n_24251 = n_24240 ^ n_23499;
assign n_24252 = n_23510 & ~n_24241;
assign n_24253 = n_24242 ^ n_22229;
assign n_24254 = n_24242 & n_24239;
assign n_24255 = n_24243 ^ n_24215;
assign n_24256 = ~n_24215 & n_24243;
assign n_24257 = n_24244 ^ x336;
assign n_24258 = n_24245 ^ n_23787;
assign n_24259 = n_24246 ^ n_22606;
assign n_24260 = n_24158 ^ n_24247;
assign n_24261 = n_24248 ^ n_24246;
assign n_24262 = n_24248 ^ n_22606;
assign n_24263 = n_24250 & ~n_24249;
assign n_24264 = n_24250 ^ x427;
assign n_24265 = n_24251 ^ n_23485;
assign n_24266 = n_24251 ^ n_23408;
assign n_24267 = n_24252 ^ n_23141;
assign n_24268 = n_24253 ^ x351;
assign n_24269 = n_24254 ^ n_22229;
assign n_24270 = n_24255 ^ n_23826;
assign n_24271 = n_24257 ^ x351;
assign n_24272 = n_24257 ^ n_24253;
assign n_24273 = n_24258 ^ n_24255;
assign n_24274 = n_24258 ^ n_23826;
assign n_24275 = n_24259 & ~n_24261;
assign n_24276 = n_24262 ^ n_24246;
assign n_24277 = n_24263 ^ x427;
assign n_24278 = n_24264 & n_24237;
assign n_24279 = n_24237 ^ n_24264;
assign n_24280 = n_24265 ^ n_22249;
assign n_24281 = n_24267 ^ n_23158;
assign n_24282 = n_24267 ^ n_23535;
assign n_24283 = n_24269 ^ n_24265;
assign n_24284 = n_24271 ^ n_24253;
assign n_24285 = ~n_24268 & n_24272;
assign n_24286 = ~n_24270 & ~n_24273;
assign n_24287 = n_24273 ^ n_23194;
assign n_24288 = n_24274 ^ n_24255;
assign n_24289 = n_24275 ^ n_22606;
assign n_24290 = n_24276 ^ x426;
assign n_24291 = n_24277 ^ n_24276;
assign n_24292 = n_24281 ^ n_23535;
assign n_24293 = n_23548 & n_24282;
assign n_24294 = n_24283 ^ n_22249;
assign n_24295 = ~n_24283 & n_24280;
assign n_24296 = n_24284 ^ n_24256;
assign n_24297 = ~n_24256 & ~n_24284;
assign n_24298 = n_24285 ^ x351;
assign n_24299 = n_24286 ^ n_23826;
assign n_24300 = n_24287 ^ n_22624;
assign n_24301 = n_24198 ^ n_24288;
assign n_24302 = n_24289 ^ n_24287;
assign n_24303 = n_24289 ^ n_22624;
assign n_24304 = n_24291 & ~n_24290;
assign n_24305 = n_24291 ^ x426;
assign n_24306 = n_24292 ^ n_23547;
assign n_24307 = n_24292 ^ n_23457;
assign n_24308 = n_24293 ^ n_23158;
assign n_24309 = n_24294 ^ x350;
assign n_24310 = n_24295 ^ n_22249;
assign n_24311 = n_24296 ^ n_23862;
assign n_24312 = n_24298 ^ n_24294;
assign n_24313 = n_24299 ^ n_24296;
assign n_24314 = n_24299 ^ n_23862;
assign n_24315 = n_24300 & n_24302;
assign n_24316 = n_24303 ^ n_24287;
assign n_24317 = n_24304 ^ x426;
assign n_24318 = n_24278 & n_24305;
assign n_24319 = n_24305 ^ n_24278;
assign n_24320 = n_24306 ^ n_22266;
assign n_24321 = n_24308 ^ n_23574;
assign n_24322 = n_24310 ^ n_24306;
assign n_24323 = n_24312 ^ x350;
assign n_24324 = ~n_24312 & n_24309;
assign n_24325 = n_24313 ^ n_23211;
assign n_24326 = n_24313 & n_24311;
assign n_24327 = n_24314 ^ n_24296;
assign n_24328 = n_24315 ^ n_22624;
assign n_24329 = n_24316 ^ x425;
assign n_24330 = n_24317 ^ n_24316;
assign n_24331 = n_23176 ^ n_24321;
assign n_24332 = n_24321 & n_23587;
assign n_24333 = n_24322 ^ n_22266;
assign n_24334 = n_24322 & ~n_24320;
assign n_24335 = n_24297 ^ n_24323;
assign n_24336 = ~n_24323 & ~n_24297;
assign n_24337 = n_24324 ^ x350;
assign n_24338 = n_24325 ^ n_22642;
assign n_24339 = n_24326 ^ n_23862;
assign n_24340 = n_24238 ^ n_24327;
assign n_24341 = n_24325 ^ n_24328;
assign n_24342 = n_24328 ^ n_22642;
assign n_24343 = n_24330 & ~n_24329;
assign n_24344 = n_24330 ^ x425;
assign n_24345 = n_24331 ^ n_23586;
assign n_24346 = n_23497 ^ n_24331;
assign n_24347 = n_24332 ^ n_23176;
assign n_24348 = n_24333 ^ x349;
assign n_24349 = n_24334 ^ n_22266;
assign n_24350 = n_24335 ^ n_23889;
assign n_24351 = n_24337 ^ n_24333;
assign n_24352 = n_24339 ^ n_24335;
assign n_24353 = n_24339 ^ n_23889;
assign n_24354 = n_24338 & n_24341;
assign n_24355 = n_24325 ^ n_24342;
assign n_24356 = n_24343 ^ x425;
assign n_24357 = n_24318 & n_24344;
assign n_24358 = n_24344 ^ n_24318;
assign n_24359 = n_24345 ^ n_22283;
assign n_24360 = n_24347 ^ n_23613;
assign n_24361 = n_24349 ^ n_22283;
assign n_24362 = n_24349 ^ n_24345;
assign n_24363 = n_24351 ^ x349;
assign n_24364 = n_24351 & ~n_24348;
assign n_24365 = n_24352 ^ n_23225;
assign n_24366 = n_24352 & n_24350;
assign n_24367 = n_24353 ^ n_24335;
assign n_24368 = n_24354 ^ n_22642;
assign n_24369 = n_24355 ^ x424;
assign n_24370 = n_24356 ^ n_24355;
assign n_24371 = n_23200 ^ n_24360;
assign n_24372 = ~n_24360 & n_23627;
assign n_24373 = n_24361 ^ n_24345;
assign n_24374 = n_24359 & n_24362;
assign n_24375 = n_24336 ^ n_24363;
assign n_24376 = n_24363 & n_24336;
assign n_24377 = n_24364 ^ x349;
assign n_24378 = n_24365 ^ n_22652;
assign n_24379 = n_24366 ^ n_23889;
assign n_24380 = n_24367 ^ n_24279;
assign n_24381 = n_24368 ^ n_24365;
assign n_24382 = ~n_24370 & n_24369;
assign n_24383 = n_24370 ^ x424;
assign n_24384 = n_24371 ^ n_23626;
assign n_24385 = n_23546 ^ n_24371;
assign n_24386 = n_24372 ^ n_23200;
assign n_24387 = n_24373 ^ x348;
assign n_24388 = n_24374 ^ n_22283;
assign n_24389 = n_24375 ^ n_23938;
assign n_24390 = n_24377 ^ n_24373;
assign n_24391 = n_24379 ^ n_24375;
assign n_24392 = n_24379 ^ n_23938;
assign n_24393 = n_24381 ^ n_22652;
assign n_24394 = n_24381 & ~n_24378;
assign n_24395 = n_24382 ^ x424;
assign n_24396 = ~n_24357 & n_24383;
assign n_24397 = n_24383 ^ n_24357;
assign n_24398 = n_24384 ^ n_22305;
assign n_24399 = n_24386 ^ n_23653;
assign n_24400 = n_24388 ^ n_22305;
assign n_24401 = n_24388 ^ n_24384;
assign n_24402 = n_24390 ^ x348;
assign n_24403 = ~n_24390 & n_24387;
assign n_24404 = n_24391 ^ n_23253;
assign n_24405 = ~n_24391 & ~n_24389;
assign n_24406 = n_24392 ^ n_24375;
assign n_24407 = n_24393 ^ x439;
assign n_24408 = n_24394 ^ n_22652;
assign n_24409 = n_24395 ^ x439;
assign n_24410 = n_24393 ^ n_24395;
assign n_24411 = n_23222 ^ n_24399;
assign n_24412 = ~n_24399 & ~n_23666;
assign n_24413 = n_24400 ^ n_24384;
assign n_24414 = ~n_24398 & n_24401;
assign n_24415 = n_24376 ^ n_24402;
assign n_24416 = ~n_24402 & n_24376;
assign n_24417 = n_24403 ^ x348;
assign n_24418 = n_24404 ^ n_22676;
assign n_24419 = n_24405 ^ n_23938;
assign n_24420 = n_24319 ^ n_24406;
assign n_24421 = n_24408 ^ n_24404;
assign n_24422 = n_24393 ^ n_24409;
assign n_24423 = n_24407 & ~n_24410;
assign n_24424 = n_24411 ^ n_23665;
assign n_24425 = n_23585 ^ n_24411;
assign n_24426 = n_24412 ^ n_23222;
assign n_24427 = n_24413 ^ x347;
assign n_24428 = n_24414 ^ n_22305;
assign n_24429 = n_24415 ^ n_23978;
assign n_24430 = n_24417 ^ n_24413;
assign n_24431 = n_24419 ^ n_24415;
assign n_24432 = n_24419 ^ n_23978;
assign n_24433 = n_24421 ^ n_22676;
assign n_24434 = ~n_24421 & n_24418;
assign n_24435 = ~n_24422 & ~n_24396;
assign n_24436 = n_24396 ^ n_24422;
assign n_24437 = n_24423 ^ x439;
assign n_24438 = n_24424 ^ n_22323;
assign n_24439 = n_24426 ^ n_23692;
assign n_24440 = n_24428 ^ n_22323;
assign n_24441 = n_24428 ^ n_24424;
assign n_24442 = n_24430 ^ x347;
assign n_24443 = ~n_24430 & n_24427;
assign n_24444 = n_24431 ^ n_23270;
assign n_24445 = ~n_24431 & n_24429;
assign n_24446 = n_24432 ^ n_24415;
assign n_24447 = n_24433 ^ x438;
assign n_24448 = n_24434 ^ n_22676;
assign n_24449 = n_24437 ^ n_24433;
assign n_24450 = n_24439 ^ n_23244;
assign n_24451 = ~n_24439 & n_23706;
assign n_24452 = n_24440 ^ n_24424;
assign n_24453 = ~n_24438 & n_24441;
assign n_24454 = n_24416 ^ n_24442;
assign n_24455 = ~n_24442 & n_24416;
assign n_24456 = n_24443 ^ x347;
assign n_24457 = n_24444 ^ n_22695;
assign n_24458 = n_24445 ^ n_23978;
assign n_24459 = n_24358 ^ n_24446;
assign n_24460 = n_24448 ^ n_24444;
assign n_24461 = n_24449 ^ x438;
assign n_24462 = n_24449 & ~n_24447;
assign n_24463 = n_24450 ^ n_23705;
assign n_24464 = n_23625 ^ n_24450;
assign n_24465 = n_24451 ^ n_23244;
assign n_24466 = n_24452 ^ x346;
assign n_24467 = n_24453 ^ n_22323;
assign n_24468 = n_24454 ^ n_24016;
assign n_24469 = n_24456 ^ n_24452;
assign n_24470 = n_24458 ^ n_24454;
assign n_24471 = n_24458 ^ n_24016;
assign n_24472 = n_24460 ^ n_22695;
assign n_24473 = ~n_24460 & ~n_24457;
assign n_24474 = n_24435 & n_24461;
assign n_24475 = n_24461 ^ n_24435;
assign n_24476 = n_24462 ^ x438;
assign n_24477 = n_24463 ^ n_22344;
assign n_24478 = n_24465 ^ n_23756;
assign n_24479 = n_24467 ^ n_22344;
assign n_24480 = n_24467 ^ n_24463;
assign n_24481 = n_24469 ^ x346;
assign n_24482 = ~n_24469 & n_24466;
assign n_24483 = n_24470 ^ n_23293;
assign n_24484 = ~n_24470 & n_24468;
assign n_24485 = n_24471 ^ n_24454;
assign n_24486 = n_24472 ^ x437;
assign n_24487 = n_24473 ^ n_22695;
assign n_24488 = n_24476 ^ n_24472;
assign n_24489 = n_24478 ^ n_23755;
assign n_24490 = n_24478 ^ n_23624;
assign n_24491 = n_24479 ^ n_24463;
assign n_24492 = ~n_24477 & n_24480;
assign n_24493 = n_24455 ^ n_24481;
assign n_24494 = ~n_24481 & n_24455;
assign n_24495 = n_24482 ^ x346;
assign n_24496 = n_24483 ^ n_22713;
assign n_24497 = n_24484 ^ n_24016;
assign n_24498 = n_24397 ^ n_24485;
assign n_24499 = n_24487 ^ n_22713;
assign n_24500 = n_24483 ^ n_24487;
assign n_24501 = n_24488 ^ x437;
assign n_24502 = ~n_24488 & n_24486;
assign n_24503 = n_24490 ^ n_23651;
assign n_24504 = n_24491 ^ x345;
assign n_24505 = n_24492 ^ n_22344;
assign n_24506 = n_24493 ^ n_24055;
assign n_24507 = n_24495 ^ n_24491;
assign n_24508 = n_24497 ^ n_24493;
assign n_24509 = n_24497 ^ n_24055;
assign n_24510 = n_24483 ^ n_24499;
assign n_24511 = ~n_24496 & n_24500;
assign n_24512 = ~n_24474 & n_24501;
assign n_24513 = n_24501 ^ n_24474;
assign n_24514 = n_24502 ^ x437;
assign n_24515 = n_24505 ^ x344;
assign n_24516 = n_24507 ^ x345;
assign n_24517 = ~n_24507 & n_24504;
assign n_24518 = n_24508 ^ n_23320;
assign n_24519 = ~n_24508 & n_24506;
assign n_24520 = n_24509 ^ n_24493;
assign n_24521 = n_24510 ^ x436;
assign n_24522 = n_24511 ^ n_22713;
assign n_24523 = n_24514 ^ n_24510;
assign n_24524 = n_24515 ^ n_24489;
assign n_24525 = n_24494 ^ n_24516;
assign n_24526 = n_24516 & ~n_24494;
assign n_24527 = n_24517 ^ x345;
assign n_24528 = n_24518 ^ n_22732;
assign n_24529 = n_24519 ^ n_24055;
assign n_24530 = n_24436 ^ n_24520;
assign n_24531 = n_24522 ^ n_22732;
assign n_24532 = n_24518 ^ n_24522;
assign n_24533 = n_24523 ^ x436;
assign n_24534 = n_24523 & ~n_24521;
assign n_24535 = n_24525 ^ n_24083;
assign n_24536 = n_24527 ^ n_24524;
assign n_24537 = n_24529 ^ n_24525;
assign n_24538 = n_24529 ^ n_24083;
assign n_24539 = n_24518 ^ n_24531;
assign n_24540 = n_24528 & ~n_24532;
assign n_24541 = ~n_24512 & n_24533;
assign n_24542 = n_24533 ^ n_24512;
assign n_24543 = n_24534 ^ x436;
assign n_24544 = n_24536 ^ n_24526;
assign n_24545 = n_24537 ^ n_23349;
assign n_24546 = n_24537 & ~n_24535;
assign n_24547 = n_24538 ^ n_24525;
assign n_24548 = n_24539 ^ x435;
assign n_24549 = n_24540 ^ n_22732;
assign n_24550 = n_24543 ^ n_24539;
assign n_24551 = n_24544 ^ n_24132;
assign n_24552 = n_24545 ^ n_22751;
assign n_24553 = n_24546 ^ n_24083;
assign n_24554 = n_24475 ^ n_24547;
assign n_24555 = n_24549 ^ n_22751;
assign n_24556 = n_24545 ^ n_24549;
assign n_24557 = n_24550 ^ x435;
assign n_24558 = ~n_24550 & n_24548;
assign n_24559 = n_24553 ^ n_24544;
assign n_24560 = n_24553 ^ n_24132;
assign n_24561 = n_24545 ^ n_24555;
assign n_24562 = ~n_24552 & n_24556;
assign n_24563 = n_24541 & ~n_24557;
assign n_24564 = n_24557 ^ n_24541;
assign n_24565 = n_24558 ^ x435;
assign n_24566 = n_24559 ^ n_23385;
assign n_24567 = ~n_24559 & n_24551;
assign n_24568 = n_24560 ^ n_24544;
assign n_24569 = n_24561 ^ x434;
assign n_24570 = n_24562 ^ n_22751;
assign n_24571 = n_24565 ^ n_24561;
assign n_24572 = n_24566 ^ n_22770;
assign n_24573 = n_24567 ^ n_24132;
assign n_24574 = n_24513 ^ n_24568;
assign n_24575 = n_24570 ^ n_22770;
assign n_24576 = n_24570 ^ n_24566;
assign n_24577 = n_24571 ^ x434;
assign n_24578 = n_24571 & ~n_24569;
assign n_24579 = n_24573 ^ n_24171;
assign n_24580 = n_24575 ^ n_24566;
assign n_24581 = n_24572 & ~n_24576;
assign n_24582 = ~n_24563 & ~n_24577;
assign n_24583 = n_24577 ^ n_24563;
assign n_24584 = n_24578 ^ x434;
assign n_24585 = n_23301 ^ n_24579;
assign n_24586 = n_24579 & ~n_24186;
assign n_24587 = n_24580 ^ x433;
assign n_24588 = n_24581 ^ n_22770;
assign n_24589 = n_24584 ^ n_24580;
assign n_24590 = n_24585 ^ n_24171;
assign n_24591 = n_24542 ^ n_24585;
assign n_24592 = n_24586 ^ n_23301;
assign n_24593 = n_24588 ^ n_22788;
assign n_24594 = n_24589 ^ x433;
assign n_24595 = ~n_24589 & n_24587;
assign n_24596 = n_24590 ^ n_23421;
assign n_24597 = n_24592 ^ n_24211;
assign n_24598 = n_24582 & n_24594;
assign n_24599 = n_24594 ^ n_24582;
assign n_24600 = n_24595 ^ x433;
assign n_24601 = n_24593 ^ n_24596;
assign n_24602 = n_24596 ^ n_22788;
assign n_24603 = n_24588 ^ n_24596;
assign n_24604 = n_23359 ^ n_24597;
assign n_24605 = n_24597 & ~n_24226;
assign n_24606 = n_24600 ^ n_24601;
assign n_24607 = n_24601 ^ x432;
assign n_24608 = n_24602 & ~n_24603;
assign n_24609 = n_24604 ^ n_24211;
assign n_24610 = n_24604 ^ n_24564;
assign n_24611 = n_24605 ^ n_23359;
assign n_24612 = n_24606 ^ x432;
assign n_24613 = ~n_24606 & n_24607;
assign n_24614 = n_24608 ^ n_22788;
assign n_24615 = n_24609 ^ n_23446;
assign n_24616 = n_24611 ^ n_23408;
assign n_24617 = n_24611 ^ n_24251;
assign n_24618 = ~n_24598 & ~n_24612;
assign n_24619 = n_24612 ^ n_24598;
assign n_24620 = n_24613 ^ x432;
assign n_24621 = n_24614 ^ n_24615;
assign n_24622 = n_24615 ^ n_22804;
assign n_24623 = n_24616 ^ n_23499;
assign n_24624 = n_24616 ^ n_24251;
assign n_24625 = n_24266 & n_24617;
assign n_24626 = n_24620 ^ x447;
assign n_24627 = n_24621 ^ n_22804;
assign n_24628 = n_24621 & ~n_24622;
assign n_24629 = n_24623 ^ n_22838;
assign n_24630 = n_24583 ^ n_24624;
assign n_24631 = n_24625 ^ n_23408;
assign n_24632 = n_24626 ^ n_24627;
assign n_24633 = n_24627 ^ x447;
assign n_24634 = n_24620 ^ n_24627;
assign n_24635 = n_24628 ^ n_22804;
assign n_24636 = n_24631 ^ n_23457;
assign n_24637 = n_24631 ^ n_24292;
assign n_24638 = ~n_24618 & ~n_24632;
assign n_24639 = n_24632 ^ n_24618;
assign n_24640 = ~n_24633 & n_24634;
assign n_24641 = n_24635 ^ n_24623;
assign n_24642 = n_24636 ^ n_23535;
assign n_24643 = n_24636 ^ n_24292;
assign n_24644 = n_24307 & ~n_24637;
assign n_24645 = n_24640 ^ x447;
assign n_24646 = n_24641 ^ n_22838;
assign n_24647 = ~n_24641 & n_24629;
assign n_24648 = n_24642 ^ n_22872;
assign n_24649 = n_24599 ^ n_24643;
assign n_24650 = n_24644 ^ n_23457;
assign n_24651 = n_24645 ^ n_24646;
assign n_24652 = n_24646 ^ x446;
assign n_24653 = n_24647 ^ n_22838;
assign n_24654 = n_24650 ^ n_24346;
assign n_24655 = n_24650 ^ n_24331;
assign n_24656 = n_24651 ^ x446;
assign n_24657 = ~n_24651 & n_24652;
assign n_24658 = n_24653 ^ n_24642;
assign n_24659 = n_24654 ^ n_24331;
assign n_24660 = n_24619 ^ n_24654;
assign n_24661 = ~n_24346 & n_24655;
assign n_24662 = n_24638 & n_24656;
assign n_24663 = n_24656 ^ n_24638;
assign n_24664 = n_24657 ^ x446;
assign n_24665 = n_24658 ^ n_22872;
assign n_24666 = ~n_24658 & n_24648;
assign n_24667 = n_24659 ^ n_23574;
assign n_24668 = n_24661 ^ n_23497;
assign n_24669 = n_24664 ^ n_24665;
assign n_24670 = n_24665 ^ x445;
assign n_24671 = n_24666 ^ n_22872;
assign n_24672 = n_24668 ^ n_24371;
assign n_24673 = n_24669 ^ x445;
assign n_24674 = ~n_24669 & n_24670;
assign n_24675 = n_24671 ^ n_22906;
assign n_24676 = n_24667 ^ n_24671;
assign n_24677 = n_23546 ^ n_24672;
assign n_24678 = ~n_24672 & ~n_24385;
assign n_24679 = n_24662 & n_24673;
assign n_24680 = n_24673 ^ n_24662;
assign n_24681 = n_24674 ^ x445;
assign n_24682 = n_24667 ^ n_24675;
assign n_24683 = n_24675 & n_24676;
assign n_24684 = n_24677 ^ n_24371;
assign n_24685 = n_24639 ^ n_24677;
assign n_24686 = n_24678 ^ n_23546;
assign n_24687 = n_24681 ^ n_24682;
assign n_24688 = n_24682 ^ x444;
assign n_24689 = n_24683 ^ n_22906;
assign n_24690 = n_24684 ^ n_23613;
assign n_24691 = n_24686 ^ n_24411;
assign n_24692 = n_24687 ^ x444;
assign n_24693 = n_24687 & ~n_24688;
assign n_24694 = n_24689 ^ n_22943;
assign n_24695 = n_24690 ^ n_22943;
assign n_24696 = n_24689 ^ n_24690;
assign n_24697 = n_23585 ^ n_24691;
assign n_24698 = ~n_24691 & ~n_24425;
assign n_24699 = ~n_24679 & n_24692;
assign n_24700 = n_24692 ^ n_24679;
assign n_24701 = n_24693 ^ x444;
assign n_24702 = n_24694 ^ n_24690;
assign n_24703 = n_24695 & ~n_24696;
assign n_24704 = n_24697 ^ n_24411;
assign n_24705 = n_24663 ^ n_24697;
assign n_24706 = n_24698 ^ n_23585;
assign n_24707 = n_24701 ^ n_24702;
assign n_24708 = n_24702 ^ x443;
assign n_24709 = n_24703 ^ n_22943;
assign n_24710 = n_24704 ^ n_23653;
assign n_24711 = n_24706 ^ n_23625;
assign n_24712 = n_24706 ^ n_24450;
assign n_24713 = n_24707 ^ x443;
assign n_24714 = ~n_24707 & n_24708;
assign n_24715 = n_24709 ^ n_22980;
assign n_24716 = n_24710 ^ n_22980;
assign n_24717 = n_24709 ^ n_24710;
assign n_24718 = n_24711 ^ n_23692;
assign n_24719 = n_24711 ^ n_24450;
assign n_24720 = n_24464 & n_24712;
assign n_24721 = n_24699 ^ n_24713;
assign n_24722 = n_24713 & ~n_24699;
assign n_24723 = n_24714 ^ x443;
assign n_24724 = n_24715 ^ n_24710;
assign n_24725 = ~n_24716 & ~n_24717;
assign n_24726 = n_24718 ^ n_23017;
assign n_24727 = n_24719 ^ n_24680;
assign n_24728 = n_24720 ^ n_23625;
assign n_24729 = n_24721 ^ n_23281;
assign n_24730 = ~n_24721 & n_23721;
assign n_24731 = n_24721 ^ n_23291;
assign n_24732 = n_23721 ^ n_24721;
assign n_24733 = n_24723 ^ n_24724;
assign n_24734 = n_24724 ^ x442;
assign n_24735 = n_24725 ^ n_22980;
assign n_24736 = n_24728 ^ n_24503;
assign n_24737 = x7 & n_24729;
assign n_24738 = n_24729 ^ x7;
assign n_24739 = n_23768 ^ n_24730;
assign n_24740 = ~n_22813 & ~n_24731;
assign n_24741 = n_24733 ^ x442;
assign n_24742 = n_24733 & ~n_24734;
assign n_24743 = n_24735 ^ n_23017;
assign n_24744 = n_24735 ^ n_24718;
assign n_24745 = n_24736 ^ n_24478;
assign n_24746 = n_24737 ^ x6;
assign n_24747 = n_24740 ^ n_22830;
assign n_24748 = n_24722 ^ n_24741;
assign n_24749 = n_24741 & ~n_24722;
assign n_24750 = n_24742 ^ x442;
assign n_24751 = n_24743 ^ n_24718;
assign n_24752 = ~n_24726 & ~n_24744;
assign n_24753 = n_24745 ^ n_23723;
assign n_24754 = n_24748 ^ n_24739;
assign n_24755 = n_24748 ^ n_24730;
assign n_24756 = n_24750 ^ n_24751;
assign n_24757 = n_24751 ^ x441;
assign n_24758 = n_24752 ^ n_23017;
assign n_24759 = n_24753 ^ n_23043;
assign n_24760 = n_24754 ^ n_23767;
assign n_24761 = n_24739 & ~n_24755;
assign n_24762 = n_24756 ^ x441;
assign n_24763 = ~n_24756 & n_24757;
assign n_24764 = n_24758 ^ x440;
assign n_24765 = n_24760 ^ n_24740;
assign n_24766 = n_24761 ^ n_23768;
assign n_24767 = n_24762 ^ n_24749;
assign n_24768 = ~n_24749 & n_24762;
assign n_24769 = n_24763 ^ x441;
assign n_24770 = n_24764 ^ n_24759;
assign n_24771 = n_24765 ^ n_22830;
assign n_24772 = n_24765 & n_24747;
assign n_24773 = n_24766 ^ n_23820;
assign n_24774 = n_23820 ^ n_24767;
assign n_24775 = n_24766 ^ n_24767;
assign n_24776 = n_24769 ^ n_24770;
assign n_24777 = n_24771 ^ n_24737;
assign n_24778 = n_24771 ^ n_24746;
assign n_24779 = n_24772 ^ n_22830;
assign n_24780 = n_24773 ^ n_24767;
assign n_24781 = n_24774 & n_24775;
assign n_24782 = n_24776 ^ n_24768;
assign n_24783 = n_24746 & n_24777;
assign n_24784 = n_24779 ^ n_22864;
assign n_24785 = n_24780 ^ n_23805;
assign n_24786 = n_24781 ^ n_23820;
assign n_24787 = n_23858 ^ n_24782;
assign n_24788 = n_24783 ^ x6;
assign n_24789 = n_24784 ^ n_24785;
assign n_24790 = n_24785 ^ n_22864;
assign n_24791 = n_24779 ^ n_24785;
assign n_24792 = n_24786 ^ n_23858;
assign n_24793 = n_24786 ^ n_24782;
assign n_24794 = n_24788 ^ n_24789;
assign n_24795 = n_24789 ^ x5;
assign n_24796 = n_24790 & ~n_24791;
assign n_24797 = n_24792 ^ n_24782;
assign n_24798 = n_24787 & n_24793;
assign n_24799 = n_24794 ^ x5;
assign n_24800 = ~n_24794 & n_24795;
assign n_24801 = n_24796 ^ n_22864;
assign n_24802 = n_24797 ^ n_23844;
assign n_24803 = n_24798 ^ n_23858;
assign n_24804 = n_24799 & ~n_24778;
assign n_24805 = n_24778 ^ n_24799;
assign n_24806 = n_24800 ^ x5;
assign n_24807 = n_24801 ^ n_22901;
assign n_24808 = n_24802 ^ n_24801;
assign n_24809 = n_23897 ^ n_24803;
assign n_24810 = n_24802 ^ n_24807;
assign n_24811 = n_24807 & n_24808;
assign n_24812 = n_23738 ^ n_24809;
assign n_24813 = ~n_24809 & n_23909;
assign n_24814 = n_24806 ^ n_24810;
assign n_24815 = n_24810 ^ x4;
assign n_24816 = n_24811 ^ n_22901;
assign n_24817 = n_24812 ^ n_23881;
assign n_24818 = n_24813 ^ n_23738;
assign n_24819 = n_24814 ^ x4;
assign n_24820 = n_24814 & ~n_24815;
assign n_24821 = n_24816 ^ n_22938;
assign n_24822 = n_24817 ^ n_22938;
assign n_24823 = n_24816 ^ n_24817;
assign n_24824 = n_24818 ^ n_23947;
assign n_24825 = n_24818 ^ n_23823;
assign n_24826 = n_24819 & ~n_24804;
assign n_24827 = n_24804 ^ n_24819;
assign n_24828 = n_24820 ^ x4;
assign n_24829 = n_24821 ^ n_24817;
assign n_24830 = n_24822 & ~n_24823;
assign n_24831 = n_24824 ^ n_23920;
assign n_24832 = ~n_23947 & ~n_24825;
assign n_24833 = n_24828 ^ n_24829;
assign n_24834 = n_24829 ^ x3;
assign n_24835 = n_24830 ^ n_22938;
assign n_24836 = n_24832 ^ n_23934;
assign n_24837 = n_24833 ^ x3;
assign n_24838 = ~n_24833 & n_24834;
assign n_24839 = n_24835 ^ n_22975;
assign n_24840 = n_24831 ^ n_24835;
assign n_24841 = n_23974 ^ n_24836;
assign n_24842 = n_24826 & ~n_24837;
assign n_24843 = n_24837 ^ n_24826;
assign n_24844 = n_24838 ^ x3;
assign n_24845 = n_24831 ^ n_24839;
assign n_24846 = n_24839 & ~n_24840;
assign n_24847 = n_23887 ^ n_24841;
assign n_24848 = n_24841 & ~n_23987;
assign n_24849 = n_24844 ^ x2;
assign n_24850 = n_24844 ^ n_24845;
assign n_24851 = n_24846 ^ n_22975;
assign n_24852 = n_24847 ^ n_23959;
assign n_24853 = n_24848 ^ n_23887;
assign n_24854 = ~n_24850 & n_24849;
assign n_24855 = n_24850 ^ x2;
assign n_24856 = n_24851 ^ n_23012;
assign n_24857 = n_24852 ^ n_23012;
assign n_24858 = n_24851 ^ n_24852;
assign n_24859 = n_24012 ^ n_24853;
assign n_24860 = n_24854 ^ x2;
assign n_24861 = n_24842 & ~n_24855;
assign n_24862 = n_24855 ^ n_24842;
assign n_24863 = n_24856 ^ n_24852;
assign n_24864 = ~n_24857 & n_24858;
assign n_24865 = n_23926 ^ n_24859;
assign n_24866 = ~n_24859 & n_24025;
assign n_24867 = n_24860 ^ x1;
assign n_24868 = n_24860 ^ n_24863;
assign n_24869 = n_24864 ^ n_23012;
assign n_24870 = n_24865 ^ n_23998;
assign n_24871 = n_24866 ^ n_23926;
assign n_24872 = n_24868 & n_24867;
assign n_24873 = n_24868 ^ x1;
assign n_24874 = n_24869 ^ n_23049;
assign n_24875 = n_24870 ^ n_23049;
assign n_24876 = n_24869 ^ n_24870;
assign n_24877 = n_24051 ^ n_24871;
assign n_24878 = n_24872 ^ x1;
assign n_24879 = n_24873 & n_24861;
assign n_24880 = n_24861 ^ n_24873;
assign n_24881 = n_24874 ^ n_24870;
assign n_24882 = ~n_24875 & ~n_24876;
assign n_24883 = n_23965 ^ n_24877;
assign n_24884 = n_24877 & n_24064;
assign n_24885 = n_24878 ^ n_24881;
assign n_24886 = n_24881 ^ x0;
assign n_24887 = n_24882 ^ n_23049;
assign n_24888 = n_24883 ^ n_24036;
assign n_24889 = n_24884 ^ n_23965;
assign n_24890 = n_24885 ^ x0;
assign n_24891 = n_24885 & ~n_24886;
assign n_24892 = n_24887 ^ n_23083;
assign n_24893 = n_24888 ^ n_23083;
assign n_24894 = n_24887 ^ n_24888;
assign n_24895 = n_24091 ^ n_24889;
assign n_24896 = n_24890 & n_24879;
assign n_24897 = n_24879 ^ n_24890;
assign n_24898 = n_24891 ^ x0;
assign n_24899 = n_24892 ^ n_24888;
assign n_24900 = ~n_24893 & n_24894;
assign n_24901 = n_24003 ^ n_24895;
assign n_24902 = n_24895 & ~n_24104;
assign n_24903 = n_24898 ^ n_24899;
assign n_24904 = n_24899 ^ x15;
assign n_24905 = n_24900 ^ n_23083;
assign n_24906 = n_24901 ^ n_24075;
assign n_24907 = n_24902 ^ n_24003;
assign n_24908 = n_24903 ^ x15;
assign n_24909 = ~n_24903 & n_24904;
assign n_24910 = n_24905 ^ n_23110;
assign n_24911 = n_24906 ^ n_23110;
assign n_24912 = n_24905 ^ n_24906;
assign n_24913 = n_24128 ^ n_24907;
assign n_24914 = n_24896 & ~n_24908;
assign n_24915 = n_24908 ^ n_24896;
assign n_24916 = n_24909 ^ x15;
assign n_24917 = n_24910 ^ n_24906;
assign n_24918 = ~n_24911 & n_24912;
assign n_24919 = n_24042 ^ n_24913;
assign n_24920 = ~n_24913 & ~n_24141;
assign n_24921 = n_24916 ^ n_24917;
assign n_24922 = n_24917 ^ x14;
assign n_24923 = n_24918 ^ n_23110;
assign n_24924 = n_24919 ^ n_24114;
assign n_24925 = n_24920 ^ n_24042;
assign n_24926 = n_24921 ^ x14;
assign n_24927 = ~n_24921 & n_24922;
assign n_24928 = n_24923 ^ n_23133;
assign n_24929 = n_24924 ^ n_23133;
assign n_24930 = n_24923 ^ n_24924;
assign n_24931 = n_24167 ^ n_24925;
assign n_24932 = n_24914 & ~n_24926;
assign n_24933 = n_24926 ^ n_24914;
assign n_24934 = n_24927 ^ x14;
assign n_24935 = n_24928 ^ n_24924;
assign n_24936 = n_24929 & ~n_24930;
assign n_24937 = n_24081 ^ n_24931;
assign n_24938 = n_24931 & ~n_24180;
assign n_24939 = n_24934 ^ n_24935;
assign n_24940 = n_24935 ^ x13;
assign n_24941 = n_24936 ^ n_23133;
assign n_24942 = n_24937 ^ n_24152;
assign n_24943 = n_24738 ^ n_24937;
assign n_24944 = n_24938 ^ n_24081;
assign n_24945 = n_24939 ^ x13;
assign n_24946 = n_24939 & ~n_24940;
assign n_24947 = n_24941 ^ n_23145;
assign n_24948 = n_24942 ^ n_23145;
assign n_24949 = n_24941 ^ n_24942;
assign n_24950 = n_24207 ^ n_24944;
assign n_24951 = n_24932 & n_24945;
assign n_24952 = n_24945 ^ n_24932;
assign n_24953 = n_24946 ^ x13;
assign n_24954 = n_24947 ^ n_24942;
assign n_24955 = n_24948 & n_24949;
assign n_24956 = n_24120 ^ n_24950;
assign n_24957 = ~n_24950 & ~n_24220;
assign n_24958 = n_24953 ^ n_24954;
assign n_24959 = n_24954 ^ x12;
assign n_24960 = n_24955 ^ n_23145;
assign n_24961 = n_24956 ^ n_24192;
assign n_24962 = n_24778 ^ n_24956;
assign n_24963 = n_24957 ^ n_24120;
assign n_24964 = n_24958 ^ x12;
assign n_24965 = n_24958 & ~n_24959;
assign n_24966 = n_24960 ^ n_23164;
assign n_24967 = n_24961 ^ n_23164;
assign n_24968 = n_24960 ^ n_24961;
assign n_24969 = n_24247 ^ n_24963;
assign n_24970 = ~n_24951 & ~n_24964;
assign n_24971 = n_24964 ^ n_24951;
assign n_24972 = n_24965 ^ x12;
assign n_24973 = n_24966 ^ n_24961;
assign n_24974 = n_24967 & n_24968;
assign n_24975 = n_24158 ^ n_24969;
assign n_24976 = n_24969 & ~n_24260;
assign n_24977 = n_24972 ^ n_24973;
assign n_24978 = n_24973 ^ x11;
assign n_24979 = n_24974 ^ n_23164;
assign n_24980 = n_24975 ^ n_24232;
assign n_24981 = n_24805 ^ n_24975;
assign n_24982 = n_24976 ^ n_24158;
assign n_24983 = n_24977 ^ x11;
assign n_24984 = ~n_24977 & n_24978;
assign n_24985 = n_24979 ^ n_23179;
assign n_24986 = n_24980 ^ n_23179;
assign n_24987 = n_24979 ^ n_24980;
assign n_24988 = n_24288 ^ n_24982;
assign n_24989 = n_24983 & n_24970;
assign n_24990 = n_24970 ^ n_24983;
assign n_24991 = n_24984 ^ x11;
assign n_24992 = n_24985 ^ n_24980;
assign n_24993 = n_24986 & n_24987;
assign n_24994 = n_24198 ^ n_24988;
assign n_24995 = n_24988 & ~n_24301;
assign n_24996 = n_24991 ^ n_24992;
assign n_24997 = n_24992 ^ x10;
assign n_24998 = n_24993 ^ n_23179;
assign n_24999 = n_24994 ^ n_24273;
assign n_25000 = n_24827 ^ n_24994;
assign n_25001 = n_24995 ^ n_24198;
assign n_25002 = n_24996 ^ x10;
assign n_25003 = n_24996 & ~n_24997;
assign n_25004 = n_24998 ^ n_23194;
assign n_25005 = n_24999 ^ n_23194;
assign n_25006 = n_24998 ^ n_24999;
assign n_25007 = n_24327 ^ n_25001;
assign n_25008 = ~n_24989 & n_25002;
assign n_25009 = n_25002 ^ n_24989;
assign n_25010 = n_25003 ^ x10;
assign n_25011 = n_25004 ^ n_24999;
assign n_25012 = ~n_25005 & n_25006;
assign n_25013 = n_24238 ^ n_25007;
assign n_25014 = n_25007 & n_24340;
assign n_25015 = n_25010 ^ n_25011;
assign n_25016 = n_25011 ^ x9;
assign n_25017 = n_25012 ^ n_23194;
assign n_25018 = n_25013 ^ n_24313;
assign n_25019 = n_24843 ^ n_25013;
assign n_25020 = n_25014 ^ n_24238;
assign n_25021 = n_25015 ^ x9;
assign n_25022 = n_25015 & ~n_25016;
assign n_25023 = n_25017 ^ n_23211;
assign n_25024 = n_25018 ^ n_23211;
assign n_25025 = n_25017 ^ n_25018;
assign n_25026 = n_25020 ^ n_24380;
assign n_25027 = n_25020 ^ n_24367;
assign n_25028 = ~n_25021 & ~n_25008;
assign n_25029 = n_25008 ^ n_25021;
assign n_25030 = n_25022 ^ x9;
assign n_25031 = n_25023 ^ n_25018;
assign n_25032 = ~n_25024 & n_25025;
assign n_25033 = n_25026 ^ n_24352;
assign n_25034 = n_24862 ^ n_25026;
assign n_25035 = ~n_24380 & n_25027;
assign n_25036 = n_25030 ^ n_25031;
assign n_25037 = n_25031 ^ x8;
assign n_25038 = n_25032 ^ n_23211;
assign n_25039 = n_25033 ^ n_23225;
assign n_25040 = n_25035 ^ n_24279;
assign n_25041 = n_25036 ^ x8;
assign n_25042 = n_25036 & ~n_25037;
assign n_25043 = n_25038 ^ n_25033;
assign n_25044 = n_25040 ^ n_24319;
assign n_25045 = n_25040 ^ n_24406;
assign n_25046 = n_25028 & ~n_25041;
assign n_25047 = n_25041 ^ n_25028;
assign n_25048 = n_25042 ^ x8;
assign n_25049 = n_25043 ^ n_23225;
assign n_25050 = n_25043 & n_25039;
assign n_25051 = n_25044 ^ n_24406;
assign n_25052 = ~n_24420 & n_25045;
assign n_25053 = n_25048 ^ x23;
assign n_25054 = n_25049 ^ x23;
assign n_25055 = n_25048 ^ n_25049;
assign n_25056 = n_25050 ^ n_23225;
assign n_25057 = n_25051 ^ n_24391;
assign n_25058 = n_24880 ^ n_25051;
assign n_25059 = n_25052 ^ n_24319;
assign n_25060 = n_25053 ^ n_25049;
assign n_25061 = n_25054 & ~n_25055;
assign n_25062 = n_25056 ^ n_25057;
assign n_25063 = n_25057 ^ n_23253;
assign n_25064 = n_24446 ^ n_25059;
assign n_25065 = ~n_25046 & ~n_25060;
assign n_25066 = n_25060 ^ n_25046;
assign n_25067 = n_25061 ^ x23;
assign n_25068 = n_25062 ^ n_23253;
assign n_25069 = n_25062 & ~n_25063;
assign n_25070 = n_24358 ^ n_25064;
assign n_25071 = n_25064 & ~n_24459;
assign n_25072 = n_25067 ^ n_25068;
assign n_25073 = n_25068 ^ x22;
assign n_25074 = n_25069 ^ n_23253;
assign n_25075 = n_25070 ^ n_24431;
assign n_25076 = n_24897 ^ n_25070;
assign n_25077 = n_25071 ^ n_24358;
assign n_25078 = n_25072 ^ x22;
assign n_25079 = ~n_25072 & n_25073;
assign n_25080 = n_25074 ^ n_25075;
assign n_25081 = n_25075 ^ n_23270;
assign n_25082 = n_24485 ^ n_25077;
assign n_25083 = ~n_25065 & n_25078;
assign n_25084 = n_25078 ^ n_25065;
assign n_25085 = n_25079 ^ x22;
assign n_25086 = n_25080 ^ n_23270;
assign n_25087 = n_25080 & ~n_25081;
assign n_25088 = n_24397 ^ n_25082;
assign n_25089 = n_25082 & ~n_24498;
assign n_25090 = n_25085 ^ n_25086;
assign n_25091 = n_25086 ^ x21;
assign n_25092 = n_25087 ^ n_23270;
assign n_25093 = n_25088 ^ n_24470;
assign n_25094 = n_24915 ^ n_25088;
assign n_25095 = n_25089 ^ n_24397;
assign n_25096 = n_25090 ^ x21;
assign n_25097 = ~n_25090 & n_25091;
assign n_25098 = n_25092 ^ n_23293;
assign n_25099 = n_25093 ^ n_23293;
assign n_25100 = n_25092 ^ n_25093;
assign n_25101 = n_24520 ^ n_25095;
assign n_25102 = n_25083 & n_25096;
assign n_25103 = n_25096 ^ n_25083;
assign n_25104 = n_25097 ^ x21;
assign n_25105 = n_25098 ^ n_25093;
assign n_25106 = ~n_25099 & n_25100;
assign n_25107 = n_24436 ^ n_25101;
assign n_25108 = n_25101 & ~n_24530;
assign n_25109 = n_25104 ^ n_25105;
assign n_25110 = n_25105 ^ x20;
assign n_25111 = n_25106 ^ n_23293;
assign n_25112 = n_25107 ^ n_24508;
assign n_25113 = n_24933 ^ n_25107;
assign n_25114 = n_25108 ^ n_24436;
assign n_25115 = n_25109 ^ x20;
assign n_25116 = ~n_25109 & n_25110;
assign n_25117 = n_25111 ^ n_23320;
assign n_25118 = n_25112 ^ n_23320;
assign n_25119 = n_25111 ^ n_25112;
assign n_25120 = n_24547 ^ n_25114;
assign n_25121 = n_25102 & n_25115;
assign n_25122 = n_25115 ^ n_25102;
assign n_25123 = n_25116 ^ x20;
assign n_25124 = n_25117 ^ n_25112;
assign n_25125 = n_25118 & n_25119;
assign n_25126 = n_24475 ^ n_25120;
assign n_25127 = ~n_25120 & n_24554;
assign n_25128 = n_25123 ^ n_25124;
assign n_25129 = n_25124 ^ x19;
assign n_25130 = n_25125 ^ n_23320;
assign n_25131 = n_25126 ^ n_24537;
assign n_25132 = n_24952 ^ n_25126;
assign n_25133 = n_25127 ^ n_24475;
assign n_25134 = n_25128 ^ x19;
assign n_25135 = n_25128 & ~n_25129;
assign n_25136 = n_25130 ^ n_23349;
assign n_25137 = n_25131 ^ n_23349;
assign n_25138 = n_25130 ^ n_25131;
assign n_25139 = n_24568 ^ n_25133;
assign n_25140 = n_25121 & ~n_25134;
assign n_25141 = n_25134 ^ n_25121;
assign n_25142 = n_25135 ^ x19;
assign n_25143 = n_25136 ^ n_25131;
assign n_25144 = n_25137 & ~n_25138;
assign n_25145 = n_24513 ^ n_25139;
assign n_25146 = n_25139 & ~n_24574;
assign n_25147 = n_25142 ^ n_25143;
assign n_25148 = n_25143 ^ x18;
assign n_25149 = n_25144 ^ n_23349;
assign n_25150 = n_25145 ^ n_24559;
assign n_25151 = n_24971 ^ n_25145;
assign n_25152 = n_25146 ^ n_24513;
assign n_25153 = n_25147 ^ x18;
assign n_25154 = ~n_25147 & n_25148;
assign n_25155 = n_25149 ^ n_23385;
assign n_25156 = n_25150 ^ n_23385;
assign n_25157 = n_25149 ^ n_25150;
assign n_25158 = n_25152 ^ n_24585;
assign n_25159 = n_25140 ^ n_25153;
assign n_25160 = ~n_25153 & ~n_25140;
assign n_25161 = n_25154 ^ x18;
assign n_25162 = n_25155 ^ n_25150;
assign n_25163 = n_25156 & ~n_25157;
assign n_25164 = n_24542 ^ n_25158;
assign n_25165 = ~n_25158 & ~n_24591;
assign n_25166 = n_25159 ^ n_23704;
assign n_25167 = ~n_25159 & ~n_24732;
assign n_25168 = n_24732 ^ n_25159;
assign n_25169 = n_25161 ^ n_25162;
assign n_25170 = n_25162 ^ x17;
assign n_25171 = n_25163 ^ n_23385;
assign n_25172 = n_25164 ^ n_24590;
assign n_25173 = n_24990 ^ n_25164;
assign n_25174 = n_25165 ^ n_24542;
assign n_25175 = x103 & ~n_25166;
assign n_25176 = n_23291 & n_25166;
assign n_25177 = n_25166 ^ x103;
assign n_25178 = n_25167 ^ n_24754;
assign n_25179 = n_25169 ^ x17;
assign n_25180 = ~n_25169 & n_25170;
assign n_25181 = n_25171 ^ n_23421;
assign n_25182 = n_25172 ^ n_23421;
assign n_25183 = n_25171 ^ n_25172;
assign n_25184 = n_25174 ^ n_24610;
assign n_25185 = n_25174 ^ n_24604;
assign n_25186 = n_25175 ^ x102;
assign n_25187 = n_25176 ^ n_23318;
assign n_25188 = n_25179 ^ n_25160;
assign n_25189 = ~n_25160 & n_25179;
assign n_25190 = n_25180 ^ x17;
assign n_25191 = n_25181 ^ n_25172;
assign n_25192 = n_25182 & ~n_25183;
assign n_25193 = n_25184 ^ n_24609;
assign n_25194 = n_25009 ^ n_25184;
assign n_25195 = ~n_24610 & n_25185;
assign n_25196 = n_25188 ^ n_25167;
assign n_25197 = n_25178 ^ n_25188;
assign n_25198 = n_25190 ^ n_25191;
assign n_25199 = n_25191 ^ x16;
assign n_25200 = n_25192 ^ n_23421;
assign n_25201 = n_25193 ^ n_23446;
assign n_25202 = n_25195 ^ n_24564;
assign n_25203 = n_25196 ^ n_23768;
assign n_25204 = n_25196 & n_25178;
assign n_25205 = n_25198 ^ x16;
assign n_25206 = ~n_25198 & n_25199;
assign n_25207 = n_25200 ^ n_25193;
assign n_25208 = n_25202 ^ n_24583;
assign n_25209 = n_25202 ^ n_24624;
assign n_25210 = n_25203 ^ n_25187;
assign n_25211 = n_25203 ^ n_25176;
assign n_25212 = n_25204 ^ n_24754;
assign n_25213 = n_25205 ^ n_25189;
assign n_25214 = ~n_25189 & ~n_25205;
assign n_25215 = n_25206 ^ x16;
assign n_25216 = n_25207 ^ n_23446;
assign n_25217 = n_25207 & n_25201;
assign n_25218 = n_25208 ^ n_24624;
assign n_25219 = n_24630 & ~n_25209;
assign n_25220 = n_25210 ^ n_25175;
assign n_25221 = n_25210 ^ n_25186;
assign n_25222 = ~n_25187 & n_25211;
assign n_25223 = n_25212 ^ n_24780;
assign n_25224 = n_25212 ^ n_25213;
assign n_25225 = n_25213 ^ n_24780;
assign n_25226 = n_25215 ^ x31;
assign n_25227 = n_25216 ^ x31;
assign n_25228 = n_25215 ^ n_25216;
assign n_25229 = n_25217 ^ n_23446;
assign n_25230 = n_25218 ^ n_24616;
assign n_25231 = n_25029 ^ n_25218;
assign n_25232 = n_25219 ^ n_24583;
assign n_25233 = n_25186 & ~n_25220;
assign n_25234 = ~n_25177 & n_25221;
assign n_25235 = n_25221 ^ n_25177;
assign n_25236 = n_25222 ^ n_23318;
assign n_25237 = n_25223 ^ n_25213;
assign n_25238 = n_25224 ^ n_23820;
assign n_25239 = n_25224 & ~n_25225;
assign n_25240 = n_25226 ^ n_25216;
assign n_25241 = n_25227 & ~n_25228;
assign n_25242 = n_25229 ^ n_25230;
assign n_25243 = n_25230 ^ n_23499;
assign n_25244 = n_25232 ^ n_24643;
assign n_25245 = n_25233 ^ x102;
assign n_25246 = n_25236 ^ n_23356;
assign n_25247 = n_25238 ^ n_23356;
assign n_25248 = n_25236 ^ n_25238;
assign n_25249 = n_25239 ^ n_24780;
assign n_25250 = n_25240 ^ n_25214;
assign n_25251 = ~n_25214 & n_25240;
assign n_25252 = n_25241 ^ x31;
assign n_25253 = n_25242 ^ n_23499;
assign n_25254 = ~n_25242 & n_25243;
assign n_25255 = n_24599 ^ n_25244;
assign n_25256 = n_25244 & ~n_24649;
assign n_25257 = n_25246 ^ n_25238;
assign n_25258 = ~n_25247 & n_25248;
assign n_25259 = n_25249 ^ n_24797;
assign n_25260 = n_25249 ^ n_25250;
assign n_25261 = n_25250 ^ n_24797;
assign n_25262 = n_25252 ^ n_25253;
assign n_25263 = n_25253 ^ x30;
assign n_25264 = n_25254 ^ n_23499;
assign n_25265 = n_25255 ^ n_24636;
assign n_25266 = n_25047 ^ n_25255;
assign n_25267 = n_25256 ^ n_24599;
assign n_25268 = n_25245 ^ n_25257;
assign n_25269 = n_25257 ^ x101;
assign n_25270 = n_25258 ^ n_23356;
assign n_25271 = n_25259 ^ n_25250;
assign n_25272 = n_25260 ^ n_23858;
assign n_25273 = n_25260 & n_25261;
assign n_25274 = n_25262 ^ x30;
assign n_25275 = n_25262 & ~n_25263;
assign n_25276 = n_25264 ^ n_25265;
assign n_25277 = n_25265 ^ n_23535;
assign n_25278 = n_25267 ^ n_24654;
assign n_25279 = n_25268 ^ x101;
assign n_25280 = ~n_25268 & n_25269;
assign n_25281 = n_25270 ^ n_23392;
assign n_25282 = n_25272 ^ n_23392;
assign n_25283 = n_25270 ^ n_25272;
assign n_25284 = n_25273 ^ n_24797;
assign n_25285 = n_25274 ^ n_25251;
assign n_25286 = ~n_25251 & n_25274;
assign n_25287 = n_25275 ^ x30;
assign n_25288 = n_25276 ^ n_23535;
assign n_25289 = ~n_25276 & ~n_25277;
assign n_25290 = n_24619 ^ n_25278;
assign n_25291 = ~n_25278 & ~n_24660;
assign n_25292 = ~n_25234 & ~n_25279;
assign n_25293 = n_25279 ^ n_25234;
assign n_25294 = n_25280 ^ x101;
assign n_25295 = n_25281 ^ n_25272;
assign n_25296 = ~n_25282 & ~n_25283;
assign n_25297 = n_25284 ^ n_24812;
assign n_25298 = n_25284 ^ n_25285;
assign n_25299 = n_25285 ^ n_24812;
assign n_25300 = n_25287 ^ n_25288;
assign n_25301 = n_25288 ^ x29;
assign n_25302 = n_25289 ^ n_23535;
assign n_25303 = n_25290 ^ n_24659;
assign n_25304 = n_25066 ^ n_25290;
assign n_25305 = n_25291 ^ n_24619;
assign n_25306 = n_25294 ^ n_25295;
assign n_25307 = n_25295 ^ x100;
assign n_25308 = n_25296 ^ n_23392;
assign n_25309 = n_25297 ^ n_25285;
assign n_25310 = n_25298 ^ n_23897;
assign n_25311 = n_25298 & n_25299;
assign n_25312 = n_25300 ^ x29;
assign n_25313 = ~n_25300 & n_25301;
assign n_25314 = n_25302 ^ n_23574;
assign n_25315 = n_25303 ^ n_23574;
assign n_25316 = n_25302 ^ n_25303;
assign n_25317 = n_25305 ^ n_24677;
assign n_25318 = n_25306 ^ x100;
assign n_25319 = ~n_25306 & n_25307;
assign n_25320 = n_25308 ^ n_23429;
assign n_25321 = n_25310 ^ n_23429;
assign n_25322 = n_25308 ^ n_25310;
assign n_25323 = n_25311 ^ n_24812;
assign n_25324 = n_25286 ^ n_25312;
assign n_25325 = n_25312 & ~n_25286;
assign n_25326 = n_25313 ^ x29;
assign n_25327 = n_25314 ^ n_25303;
assign n_25328 = n_25315 & n_25316;
assign n_25329 = n_24639 ^ n_25317;
assign n_25330 = n_25317 & n_24685;
assign n_25331 = ~n_25292 & n_25318;
assign n_25332 = n_25318 ^ n_25292;
assign n_25333 = n_25319 ^ x100;
assign n_25334 = n_25320 ^ n_25310;
assign n_25335 = ~n_25321 & n_25322;
assign n_25336 = n_25323 ^ n_24824;
assign n_25337 = n_25323 ^ n_25324;
assign n_25338 = n_25324 ^ n_24824;
assign n_25339 = n_25326 ^ n_25327;
assign n_25340 = n_25327 ^ x28;
assign n_25341 = n_25328 ^ n_23574;
assign n_25342 = n_25329 ^ n_24684;
assign n_25343 = n_25084 ^ n_25329;
assign n_25344 = n_25330 ^ n_24639;
assign n_25345 = n_25333 ^ n_25334;
assign n_25346 = n_25334 ^ x99;
assign n_25347 = n_25335 ^ n_23429;
assign n_25348 = n_25336 ^ n_25324;
assign n_25349 = n_25337 ^ n_23934;
assign n_25350 = n_25337 & n_25338;
assign n_25351 = n_25339 ^ x28;
assign n_25352 = ~n_25339 & n_25340;
assign n_25353 = n_25341 ^ n_23613;
assign n_25354 = n_25342 ^ n_23613;
assign n_25355 = n_25341 ^ n_25342;
assign n_25356 = n_25344 ^ n_24697;
assign n_25357 = n_25345 ^ x99;
assign n_25358 = n_25345 & ~n_25346;
assign n_25359 = n_25347 ^ n_23468;
assign n_25360 = n_25349 ^ n_23468;
assign n_25361 = n_25347 ^ n_25349;
assign n_25362 = n_25350 ^ n_24824;
assign n_25363 = n_25325 ^ n_25351;
assign n_25364 = ~n_25351 & ~n_25325;
assign n_25365 = n_25352 ^ x28;
assign n_25366 = n_25353 ^ n_25342;
assign n_25367 = ~n_25354 & n_25355;
assign n_25368 = n_24663 ^ n_25356;
assign n_25369 = n_25356 & ~n_24705;
assign n_25370 = n_25331 & ~n_25357;
assign n_25371 = n_25357 ^ n_25331;
assign n_25372 = n_25358 ^ x99;
assign n_25373 = n_25359 ^ n_25349;
assign n_25374 = n_25360 & ~n_25361;
assign n_25375 = n_25362 ^ n_24847;
assign n_25376 = n_25362 ^ n_25363;
assign n_25377 = n_25363 ^ n_24847;
assign n_25378 = n_25365 ^ n_25366;
assign n_25379 = n_25366 ^ x27;
assign n_25380 = n_25367 ^ n_23613;
assign n_25381 = n_25368 ^ n_24704;
assign n_25382 = n_25103 ^ n_25368;
assign n_25383 = n_25369 ^ n_24663;
assign n_25384 = n_25372 ^ n_25373;
assign n_25385 = n_25373 ^ x98;
assign n_25386 = n_25374 ^ n_23468;
assign n_25387 = n_25375 ^ n_25363;
assign n_25388 = n_25376 ^ n_23974;
assign n_25389 = ~n_25376 & ~n_25377;
assign n_25390 = n_25378 ^ x27;
assign n_25391 = ~n_25378 & n_25379;
assign n_25392 = n_25380 ^ n_23653;
assign n_25393 = n_25381 ^ n_23653;
assign n_25394 = n_25380 ^ n_25381;
assign n_25395 = n_25383 ^ n_24719;
assign n_25396 = n_25384 ^ x98;
assign n_25397 = ~n_25384 & n_25385;
assign n_25398 = n_25386 ^ n_23505;
assign n_25399 = n_25388 ^ n_23505;
assign n_25400 = n_25386 ^ n_25388;
assign n_25401 = n_25389 ^ n_24847;
assign n_25402 = n_25364 ^ n_25390;
assign n_25403 = n_25390 & ~n_25364;
assign n_25404 = n_25391 ^ x27;
assign n_25405 = n_25392 ^ n_25381;
assign n_25406 = ~n_25393 & n_25394;
assign n_25407 = n_25395 ^ n_24680;
assign n_25408 = n_25395 & ~n_24727;
assign n_25409 = n_25396 & n_25370;
assign n_25410 = n_25370 ^ n_25396;
assign n_25411 = n_25397 ^ x98;
assign n_25412 = n_25398 ^ n_25388;
assign n_25413 = ~n_25399 & ~n_25400;
assign n_25414 = n_25401 ^ n_24865;
assign n_25415 = n_25401 ^ n_25402;
assign n_25416 = n_25402 ^ n_24865;
assign n_25417 = n_25404 ^ n_25405;
assign n_25418 = n_25405 ^ x26;
assign n_25419 = n_25406 ^ n_23653;
assign n_25420 = n_25407 ^ n_24711;
assign n_25421 = n_25122 ^ n_25407;
assign n_25422 = n_25408 ^ n_24680;
assign n_25423 = n_25411 ^ n_25412;
assign n_25424 = n_25412 ^ x97;
assign n_25425 = n_25413 ^ n_23505;
assign n_25426 = n_25414 ^ n_25402;
assign n_25427 = n_25415 ^ n_24012;
assign n_25428 = n_25415 & n_25416;
assign n_25429 = n_25417 ^ x26;
assign n_25430 = ~n_25417 & n_25418;
assign n_25431 = n_25419 ^ n_23692;
assign n_25432 = n_25420 ^ n_23692;
assign n_25433 = n_25419 ^ n_25420;
assign n_25434 = n_25422 ^ n_24736;
assign n_25435 = n_25423 ^ x97;
assign n_25436 = n_25423 & ~n_25424;
assign n_25437 = n_25425 ^ n_23541;
assign n_25438 = n_25427 ^ n_23541;
assign n_25439 = n_25425 ^ n_25427;
assign n_25440 = n_25428 ^ n_24865;
assign n_25441 = ~n_25429 & ~n_25403;
assign n_25442 = n_25403 ^ n_25429;
assign n_25443 = n_25430 ^ x26;
assign n_25444 = n_25431 ^ n_25420;
assign n_25445 = n_25432 & n_25433;
assign n_25446 = n_25434 ^ n_24700;
assign n_25447 = n_25409 & ~n_25435;
assign n_25448 = n_25435 ^ n_25409;
assign n_25449 = n_25436 ^ x97;
assign n_25450 = n_25437 ^ n_25427;
assign n_25451 = n_25438 & n_25439;
assign n_25452 = n_25440 ^ n_24883;
assign n_25453 = n_25440 ^ n_25442;
assign n_25454 = n_25442 ^ n_24883;
assign n_25455 = n_25443 ^ n_25444;
assign n_25456 = n_25444 ^ x25;
assign n_25457 = n_25445 ^ n_23692;
assign n_25458 = n_25446 ^ n_24753;
assign n_25459 = n_25449 ^ n_25450;
assign n_25460 = n_25450 ^ x96;
assign n_25461 = n_25451 ^ n_23541;
assign n_25462 = n_25452 ^ n_25442;
assign n_25463 = n_25453 ^ n_24051;
assign n_25464 = ~n_25453 & n_25454;
assign n_25465 = n_25455 ^ x25;
assign n_25466 = n_25455 & ~n_25456;
assign n_25467 = n_25457 ^ x24;
assign n_25468 = n_25459 ^ x96;
assign n_25469 = n_25459 & ~n_25460;
assign n_25470 = n_25461 ^ n_23580;
assign n_25471 = n_25463 ^ n_23580;
assign n_25472 = n_25461 ^ n_25463;
assign n_25473 = n_25464 ^ n_24883;
assign n_25474 = n_25465 & n_25441;
assign n_25475 = n_25441 ^ n_25465;
assign n_25476 = n_25466 ^ x25;
assign n_25477 = n_25467 ^ n_25458;
assign n_25478 = n_25447 ^ n_25468;
assign n_25479 = n_25468 & ~n_25447;
assign n_25480 = n_25469 ^ x96;
assign n_25481 = n_25470 ^ n_25463;
assign n_25482 = ~n_25471 & ~n_25472;
assign n_25483 = n_25473 ^ n_24901;
assign n_25484 = n_25475 ^ n_25473;
assign n_25485 = n_25475 ^ n_24901;
assign n_25486 = n_25476 ^ n_25477;
assign n_25487 = n_25480 ^ n_25481;
assign n_25488 = n_25481 ^ x111;
assign n_25489 = n_25482 ^ n_23580;
assign n_25490 = n_25483 ^ n_25475;
assign n_25491 = n_25484 ^ n_24091;
assign n_25492 = ~n_25484 & n_25485;
assign n_25493 = n_25486 ^ n_25474;
assign n_25494 = n_25487 ^ x111;
assign n_25495 = n_25487 & ~n_25488;
assign n_25496 = n_25489 ^ n_23620;
assign n_25497 = n_25491 ^ n_23620;
assign n_25498 = n_25489 ^ n_25491;
assign n_25499 = n_25492 ^ n_24901;
assign n_25500 = n_25493 ^ n_24919;
assign n_25501 = ~n_25479 & ~n_25494;
assign n_25502 = n_25494 ^ n_25479;
assign n_25503 = n_25495 ^ x111;
assign n_25504 = n_25496 ^ n_25491;
assign n_25505 = ~n_25497 & ~n_25498;
assign n_25506 = n_25493 ^ n_25499;
assign n_25507 = n_25499 ^ n_24919;
assign n_25508 = n_25503 ^ n_25504;
assign n_25509 = n_25504 ^ x110;
assign n_25510 = n_25505 ^ n_23620;
assign n_25511 = ~n_25506 & n_25500;
assign n_25512 = n_25506 ^ n_24128;
assign n_25513 = n_25507 ^ n_25493;
assign n_25514 = n_25508 ^ x110;
assign n_25515 = ~n_25508 & n_25509;
assign n_25516 = n_25510 ^ n_23660;
assign n_25517 = n_25511 ^ n_24919;
assign n_25518 = n_25512 ^ n_23660;
assign n_25519 = n_25510 ^ n_25512;
assign n_25520 = n_25501 & n_25514;
assign n_25521 = n_25514 ^ n_25501;
assign n_25522 = n_25515 ^ x110;
assign n_25523 = n_25516 ^ n_25512;
assign n_25524 = n_25517 ^ n_24937;
assign n_25525 = n_25518 & ~n_25519;
assign n_25526 = n_25522 ^ n_25523;
assign n_25527 = n_25523 ^ x109;
assign n_25528 = n_25524 & n_24943;
assign n_25529 = n_24738 ^ n_25524;
assign n_25530 = n_25525 ^ n_23660;
assign n_25531 = n_25526 ^ x109;
assign n_25532 = ~n_25526 & n_25527;
assign n_25533 = n_25528 ^ n_24738;
assign n_25534 = n_25529 ^ n_24937;
assign n_25535 = n_25530 ^ n_23699;
assign n_25536 = n_25520 & n_25531;
assign n_25537 = n_25531 ^ n_25520;
assign n_25538 = n_25532 ^ x109;
assign n_25539 = n_25533 ^ n_24956;
assign n_25540 = n_25534 ^ n_24167;
assign n_25541 = ~n_25539 & n_24962;
assign n_25542 = n_25539 ^ n_24778;
assign n_25543 = n_25540 ^ n_23699;
assign n_25544 = n_25530 ^ n_25540;
assign n_25545 = n_25535 ^ n_25540;
assign n_25546 = n_25541 ^ n_24778;
assign n_25547 = n_25542 ^ n_24956;
assign n_25548 = ~n_25543 & n_25544;
assign n_25549 = n_25538 ^ n_25545;
assign n_25550 = n_25545 ^ x108;
assign n_25551 = n_25546 ^ n_24975;
assign n_25552 = n_25547 ^ n_24207;
assign n_25553 = n_25548 ^ n_23699;
assign n_25554 = n_25549 ^ x108;
assign n_25555 = n_25549 & ~n_25550;
assign n_25556 = n_25551 & n_24981;
assign n_25557 = n_24805 ^ n_25551;
assign n_25558 = n_25553 ^ n_23747;
assign n_25559 = n_25552 ^ n_25553;
assign n_25560 = ~n_25554 & n_25536;
assign n_25561 = n_25536 ^ n_25554;
assign n_25562 = n_25555 ^ x108;
assign n_25563 = n_25556 ^ n_24805;
assign n_25564 = n_25557 ^ n_24975;
assign n_25565 = n_25552 ^ n_25558;
assign n_25566 = n_25558 & n_25559;
assign n_25567 = n_25563 ^ n_24994;
assign n_25568 = n_25564 ^ n_24247;
assign n_25569 = n_25562 ^ n_25565;
assign n_25570 = n_25565 ^ x107;
assign n_25571 = n_25566 ^ n_23747;
assign n_25572 = ~n_25567 & ~n_25000;
assign n_25573 = n_24827 ^ n_25567;
assign n_25574 = n_25568 ^ n_23787;
assign n_25575 = n_25569 ^ x107;
assign n_25576 = n_25569 & ~n_25570;
assign n_25577 = n_25571 ^ n_25568;
assign n_25578 = n_25571 ^ n_23787;
assign n_25579 = n_25572 ^ n_24827;
assign n_25580 = n_25573 ^ n_24994;
assign n_25581 = ~n_25560 & n_25575;
assign n_25582 = n_25575 ^ n_25560;
assign n_25583 = n_25576 ^ x107;
assign n_25584 = n_25574 & ~n_25577;
assign n_25585 = n_25578 ^ n_25568;
assign n_25586 = n_25579 ^ n_25013;
assign n_25587 = n_25580 ^ n_24288;
assign n_25588 = n_25583 ^ x106;
assign n_25589 = n_25584 ^ n_23787;
assign n_25590 = n_25583 ^ n_25585;
assign n_25591 = ~n_25586 & n_25019;
assign n_25592 = n_24843 ^ n_25586;
assign n_25593 = n_25587 ^ n_23826;
assign n_25594 = n_25589 ^ n_25587;
assign n_25595 = n_25589 ^ n_23826;
assign n_25596 = ~n_25590 & n_25588;
assign n_25597 = n_25590 ^ x106;
assign n_25598 = n_25591 ^ n_24843;
assign n_25599 = n_25592 ^ n_25013;
assign n_25600 = ~n_25593 & ~n_25594;
assign n_25601 = n_25595 ^ n_25587;
assign n_25602 = n_25596 ^ x106;
assign n_25603 = n_25581 & ~n_25597;
assign n_25604 = n_25597 ^ n_25581;
assign n_25605 = n_25598 ^ n_25026;
assign n_25606 = n_25598 ^ n_25034;
assign n_25607 = n_25599 ^ n_24327;
assign n_25608 = n_25600 ^ n_23826;
assign n_25609 = n_25601 ^ x105;
assign n_25610 = n_25602 ^ n_25601;
assign n_25611 = n_25034 & ~n_25605;
assign n_25612 = n_25606 ^ n_25177;
assign n_25613 = n_25606 ^ n_25026;
assign n_25614 = n_25607 ^ n_23862;
assign n_25615 = n_25608 ^ n_25607;
assign n_25616 = n_25608 ^ n_23862;
assign n_25617 = n_25610 & ~n_25609;
assign n_25618 = n_25610 ^ x105;
assign n_25619 = n_25611 ^ n_24862;
assign n_25620 = n_25613 ^ n_24367;
assign n_25621 = ~n_25614 & ~n_25615;
assign n_25622 = n_25616 ^ n_25607;
assign n_25623 = n_25617 ^ x105;
assign n_25624 = ~n_25603 & ~n_25618;
assign n_25625 = n_25618 ^ n_25603;
assign n_25626 = n_25619 ^ n_25051;
assign n_25627 = n_25619 ^ n_24880;
assign n_25628 = n_25620 ^ n_23889;
assign n_25629 = n_25621 ^ n_23862;
assign n_25630 = n_25622 ^ x104;
assign n_25631 = n_25623 ^ n_25622;
assign n_25632 = ~n_25058 & ~n_25626;
assign n_25633 = n_25627 ^ n_25051;
assign n_25634 = n_25627 ^ n_24406;
assign n_25635 = n_25629 ^ n_25620;
assign n_25636 = ~n_25631 & n_25630;
assign n_25637 = n_25631 ^ x104;
assign n_25638 = n_25632 ^ n_24880;
assign n_25639 = n_25235 ^ n_25633;
assign n_25640 = n_25634 ^ n_23938;
assign n_25641 = ~n_25635 & ~n_25628;
assign n_25642 = n_25635 ^ n_23889;
assign n_25643 = n_25636 ^ x104;
assign n_25644 = n_25624 & n_25637;
assign n_25645 = n_25637 ^ n_25624;
assign n_25646 = n_25638 ^ n_25070;
assign n_25647 = n_25641 ^ n_23889;
assign n_25648 = n_25642 ^ x119;
assign n_25649 = n_25643 ^ n_25642;
assign n_25650 = n_25643 ^ x119;
assign n_25651 = n_25646 & ~n_25076;
assign n_25652 = n_24897 ^ n_25646;
assign n_25653 = n_25647 ^ n_25634;
assign n_25654 = ~n_25648 & n_25649;
assign n_25655 = n_25650 ^ n_25642;
assign n_25656 = n_25651 ^ n_24897;
assign n_25657 = n_25652 ^ n_25070;
assign n_25658 = n_25293 ^ n_25652;
assign n_25659 = ~n_25653 & ~n_25640;
assign n_25660 = n_25653 ^ n_23938;
assign n_25661 = n_25654 ^ x119;
assign n_25662 = ~n_25644 & n_25655;
assign n_25663 = n_25655 ^ n_25644;
assign n_25664 = n_25656 ^ n_25088;
assign n_25665 = n_25657 ^ n_24446;
assign n_25666 = n_25659 ^ n_23938;
assign n_25667 = n_25660 ^ x118;
assign n_25668 = n_25661 ^ n_25660;
assign n_25669 = n_25663 & n_25168;
assign n_25670 = n_25663 ^ n_24732;
assign n_25671 = n_25663 ^ n_24721;
assign n_25672 = n_25664 & n_25094;
assign n_25673 = n_24915 ^ n_25664;
assign n_25674 = n_25665 ^ n_23978;
assign n_25675 = n_25666 ^ n_25665;
assign n_25676 = ~n_25668 & n_25667;
assign n_25677 = n_25668 ^ x118;
assign n_25678 = n_25197 ^ n_25669;
assign n_25679 = n_23721 & ~n_25670;
assign n_25680 = n_25670 ^ n_25159;
assign n_25681 = x199 & ~n_25671;
assign n_25682 = n_25671 ^ x199;
assign n_25683 = n_25672 ^ n_24915;
assign n_25684 = n_25673 ^ n_25088;
assign n_25685 = n_25332 ^ n_25673;
assign n_25686 = ~n_25675 & n_25674;
assign n_25687 = n_25675 ^ n_23978;
assign n_25688 = n_25676 ^ x118;
assign n_25689 = n_25662 & ~n_25677;
assign n_25690 = n_25677 ^ n_25662;
assign n_25691 = n_25679 ^ n_23768;
assign n_25692 = n_25681 ^ x198;
assign n_25693 = n_25683 ^ n_25107;
assign n_25694 = n_25684 ^ n_24485;
assign n_25695 = n_25686 ^ n_23978;
assign n_25696 = n_25687 ^ x117;
assign n_25697 = n_25688 ^ n_25687;
assign n_25698 = n_25690 ^ n_25669;
assign n_25699 = n_25690 ^ n_25678;
assign n_25700 = ~n_25693 & n_25113;
assign n_25701 = n_24933 ^ n_25693;
assign n_25702 = n_25694 ^ n_24016;
assign n_25703 = n_25695 ^ n_25694;
assign n_25704 = n_25695 ^ n_24016;
assign n_25705 = ~n_25697 & n_25696;
assign n_25706 = n_25697 ^ x117;
assign n_25707 = ~n_25678 & ~n_25698;
assign n_25708 = n_25699 ^ n_25196;
assign n_25709 = n_25700 ^ n_24933;
assign n_25710 = n_25701 ^ n_25107;
assign n_25711 = n_25371 ^ n_25701;
assign n_25712 = ~n_25702 & n_25703;
assign n_25713 = n_25704 ^ n_25694;
assign n_25714 = n_25705 ^ x117;
assign n_25715 = n_25689 & ~n_25706;
assign n_25716 = n_25706 ^ n_25689;
assign n_25717 = n_25707 ^ n_25197;
assign n_25718 = n_25708 ^ n_25679;
assign n_25719 = n_25708 ^ n_25691;
assign n_25720 = n_25709 ^ n_25126;
assign n_25721 = n_25710 ^ n_24520;
assign n_25722 = n_25712 ^ n_24016;
assign n_25723 = n_25713 ^ x116;
assign n_25724 = n_25714 ^ n_25713;
assign n_25725 = n_25237 ^ n_25717;
assign n_25726 = n_25716 ^ n_25717;
assign n_25727 = n_25691 & ~n_25718;
assign n_25728 = n_25719 ^ n_25681;
assign n_25729 = n_25719 ^ n_25692;
assign n_25730 = n_24952 ^ n_25720;
assign n_25731 = n_25720 & n_25132;
assign n_25732 = n_25721 ^ n_24055;
assign n_25733 = n_25722 ^ n_25721;
assign n_25734 = n_25722 ^ n_24055;
assign n_25735 = n_25724 & ~n_25723;
assign n_25736 = n_25724 ^ x116;
assign n_25737 = n_25716 ^ n_25725;
assign n_25738 = n_25725 & n_25726;
assign n_25739 = n_25727 ^ n_23768;
assign n_25740 = n_25692 & ~n_25728;
assign n_25741 = ~n_25682 & n_25729;
assign n_25742 = n_25729 ^ n_25682;
assign n_25743 = n_25730 ^ n_25410;
assign n_25744 = n_25730 ^ n_25126;
assign n_25745 = n_25731 ^ n_24952;
assign n_25746 = n_25732 & ~n_25733;
assign n_25747 = n_25734 ^ n_25721;
assign n_25748 = n_25735 ^ x116;
assign n_25749 = n_25736 & n_25715;
assign n_25750 = n_25715 ^ n_25736;
assign n_25751 = n_25737 ^ n_25224;
assign n_25752 = n_25738 ^ n_25237;
assign n_25753 = n_25739 ^ n_23820;
assign n_25754 = n_25740 ^ x198;
assign n_25755 = n_25744 ^ n_24547;
assign n_25756 = n_25745 ^ n_25145;
assign n_25757 = n_25746 ^ n_24055;
assign n_25758 = n_25747 ^ x115;
assign n_25759 = n_25748 ^ n_25747;
assign n_25760 = n_25271 ^ n_25750;
assign n_25761 = n_25751 ^ n_23820;
assign n_25762 = n_25739 ^ n_25751;
assign n_25763 = n_25752 ^ n_25750;
assign n_25764 = n_25752 ^ n_25271;
assign n_25765 = n_25753 ^ n_25751;
assign n_25766 = n_25755 ^ n_24083;
assign n_25767 = n_25756 & n_25151;
assign n_25768 = n_24971 ^ n_25756;
assign n_25769 = n_25757 ^ n_25755;
assign n_25770 = n_25757 ^ n_24083;
assign n_25771 = ~n_25759 & n_25758;
assign n_25772 = n_25759 ^ x115;
assign n_25773 = n_25761 & n_25762;
assign n_25774 = ~n_25760 & ~n_25763;
assign n_25775 = n_25764 ^ n_25750;
assign n_25776 = n_25754 ^ n_25765;
assign n_25777 = n_25765 ^ x197;
assign n_25778 = n_25767 ^ n_24971;
assign n_25779 = n_25768 ^ n_25145;
assign n_25780 = n_25448 ^ n_25768;
assign n_25781 = n_25766 & ~n_25769;
assign n_25782 = n_25770 ^ n_25755;
assign n_25783 = n_25771 ^ x115;
assign n_25784 = n_25772 & ~n_25749;
assign n_25785 = n_25749 ^ n_25772;
assign n_25786 = n_25773 ^ n_23820;
assign n_25787 = n_25774 ^ n_25271;
assign n_25788 = n_25775 ^ n_25260;
assign n_25789 = n_25776 ^ x197;
assign n_25790 = ~n_25776 & n_25777;
assign n_25791 = n_25778 ^ n_25164;
assign n_25792 = n_25779 ^ n_24568;
assign n_25793 = n_25781 ^ n_24083;
assign n_25794 = n_25782 ^ x114;
assign n_25795 = n_25783 ^ n_25782;
assign n_25796 = n_25309 ^ n_25785;
assign n_25797 = n_25786 ^ n_23858;
assign n_25798 = n_25787 ^ n_25785;
assign n_25799 = n_25787 ^ n_25309;
assign n_25800 = n_25788 ^ n_23858;
assign n_25801 = n_25786 ^ n_25788;
assign n_25802 = ~n_25741 & ~n_25789;
assign n_25803 = n_25789 ^ n_25741;
assign n_25804 = n_25790 ^ x197;
assign n_25805 = n_24990 ^ n_25791;
assign n_25806 = ~n_25791 & n_25173;
assign n_25807 = n_25792 ^ n_24132;
assign n_25808 = n_25793 ^ n_25792;
assign n_25809 = n_25793 ^ n_24132;
assign n_25810 = ~n_25795 & n_25794;
assign n_25811 = n_25795 ^ x114;
assign n_25812 = n_25797 ^ n_25788;
assign n_25813 = n_25796 & n_25798;
assign n_25814 = n_25799 ^ n_25785;
assign n_25815 = ~n_25800 & ~n_25801;
assign n_25816 = n_25805 ^ n_25164;
assign n_25817 = n_25478 ^ n_25805;
assign n_25818 = n_25806 ^ n_24990;
assign n_25819 = ~n_25807 & n_25808;
assign n_25820 = n_25809 ^ n_25792;
assign n_25821 = n_25810 ^ x114;
assign n_25822 = ~n_25784 & ~n_25811;
assign n_25823 = n_25811 ^ n_25784;
assign n_25824 = n_25804 ^ n_25812;
assign n_25825 = n_25812 ^ x196;
assign n_25826 = n_25813 ^ n_25309;
assign n_25827 = n_25814 ^ n_25298;
assign n_25828 = n_25815 ^ n_23858;
assign n_25829 = n_25816 ^ n_24585;
assign n_25830 = n_25818 ^ n_25194;
assign n_25831 = n_25818 ^ n_25184;
assign n_25832 = n_25819 ^ n_24132;
assign n_25833 = n_25820 ^ x113;
assign n_25834 = n_25821 ^ n_25820;
assign n_25835 = n_25348 ^ n_25823;
assign n_25836 = n_25824 ^ x196;
assign n_25837 = ~n_25824 & n_25825;
assign n_25838 = n_25826 ^ n_25823;
assign n_25839 = n_25826 ^ n_25348;
assign n_25840 = n_25827 ^ n_23897;
assign n_25841 = n_25828 ^ n_25827;
assign n_25842 = n_25828 ^ n_23897;
assign n_25843 = n_25829 ^ n_24171;
assign n_25844 = n_25830 ^ n_25184;
assign n_25845 = n_25502 ^ n_25830;
assign n_25846 = ~n_25194 & n_25831;
assign n_25847 = n_25832 ^ n_25829;
assign n_25848 = n_25832 ^ n_24171;
assign n_25849 = n_25834 & ~n_25833;
assign n_25850 = n_25834 ^ x113;
assign n_25851 = ~n_25802 & n_25836;
assign n_25852 = n_25836 ^ n_25802;
assign n_25853 = n_25837 ^ x196;
assign n_25854 = ~n_25835 & ~n_25838;
assign n_25855 = n_25839 ^ n_25823;
assign n_25856 = ~n_25840 & n_25841;
assign n_25857 = n_25842 ^ n_25827;
assign n_25858 = n_25844 ^ n_24604;
assign n_25859 = n_25846 ^ n_25009;
assign n_25860 = n_25843 & n_25847;
assign n_25861 = n_25848 ^ n_25829;
assign n_25862 = n_25849 ^ x113;
assign n_25863 = n_25822 & n_25850;
assign n_25864 = n_25850 ^ n_25822;
assign n_25865 = n_25854 ^ n_25348;
assign n_25866 = n_25855 ^ n_25337;
assign n_25867 = n_25856 ^ n_23897;
assign n_25868 = n_25853 ^ n_25857;
assign n_25869 = n_25857 ^ x195;
assign n_25870 = n_25858 ^ n_24211;
assign n_25871 = n_25859 ^ n_25029;
assign n_25872 = n_25859 ^ n_25218;
assign n_25873 = n_25860 ^ n_24171;
assign n_25874 = n_25861 ^ x112;
assign n_25875 = n_25862 ^ n_25861;
assign n_25876 = n_25387 ^ n_25864;
assign n_25877 = n_25865 ^ n_25864;
assign n_25878 = n_25865 ^ n_25387;
assign n_25879 = n_25866 ^ n_23934;
assign n_25880 = n_25867 ^ n_25866;
assign n_25881 = n_25867 ^ n_23934;
assign n_25882 = n_25868 ^ x195;
assign n_25883 = n_25868 & ~n_25869;
assign n_25884 = n_25871 ^ n_24624;
assign n_25885 = n_25871 ^ n_25218;
assign n_25886 = n_25231 & ~n_25872;
assign n_25887 = n_25873 ^ n_25858;
assign n_25888 = ~n_25875 & n_25874;
assign n_25889 = n_25875 ^ x112;
assign n_25890 = ~n_25876 & n_25877;
assign n_25891 = n_25878 ^ n_25864;
assign n_25892 = n_25879 & n_25880;
assign n_25893 = n_25881 ^ n_25866;
assign n_25894 = ~n_25882 & n_25851;
assign n_25895 = n_25851 ^ n_25882;
assign n_25896 = n_25883 ^ x195;
assign n_25897 = n_25884 ^ n_24251;
assign n_25898 = n_25521 ^ n_25885;
assign n_25899 = n_25886 ^ n_25029;
assign n_25900 = n_25887 ^ n_24211;
assign n_25901 = ~n_25887 & n_25870;
assign n_25902 = n_25888 ^ x112;
assign n_25903 = n_25863 & ~n_25889;
assign n_25904 = n_25889 ^ n_25863;
assign n_25905 = n_25890 ^ n_25387;
assign n_25906 = n_25891 ^ n_25376;
assign n_25907 = n_25892 ^ n_23934;
assign n_25908 = n_25893 ^ x194;
assign n_25909 = n_25896 ^ n_25893;
assign n_25910 = n_25899 ^ n_25047;
assign n_25911 = n_25899 ^ n_25255;
assign n_25912 = n_25900 ^ x127;
assign n_25913 = n_25901 ^ n_24211;
assign n_25914 = n_25902 ^ n_25900;
assign n_25915 = n_25902 ^ x127;
assign n_25916 = n_25426 ^ n_25904;
assign n_25917 = n_25905 ^ n_25904;
assign n_25918 = n_25905 ^ n_25426;
assign n_25919 = n_25906 ^ n_23974;
assign n_25920 = n_25907 ^ n_25906;
assign n_25921 = n_25907 ^ n_23974;
assign n_25922 = ~n_25909 & n_25908;
assign n_25923 = n_25909 ^ x194;
assign n_25924 = n_25910 ^ n_24643;
assign n_25925 = n_25910 ^ n_25255;
assign n_25926 = n_25266 & n_25911;
assign n_25927 = n_25913 ^ n_25884;
assign n_25928 = ~n_25912 & n_25914;
assign n_25929 = n_25915 ^ n_25900;
assign n_25930 = n_25916 & ~n_25917;
assign n_25931 = n_25918 ^ n_25904;
assign n_25932 = ~n_25919 & ~n_25920;
assign n_25933 = n_25921 ^ n_25906;
assign n_25934 = n_25922 ^ x194;
assign n_25935 = n_25894 & n_25923;
assign n_25936 = n_25923 ^ n_25894;
assign n_25937 = n_25924 ^ n_24292;
assign n_25938 = n_25537 ^ n_25925;
assign n_25939 = n_25926 ^ n_25047;
assign n_25940 = n_25927 ^ n_24251;
assign n_25941 = n_25927 & ~n_25897;
assign n_25942 = n_25928 ^ x127;
assign n_25943 = ~n_25903 & ~n_25929;
assign n_25944 = n_25929 ^ n_25903;
assign n_25945 = n_25930 ^ n_25426;
assign n_25946 = n_25931 ^ n_25415;
assign n_25947 = n_25932 ^ n_23974;
assign n_25948 = n_25933 ^ x193;
assign n_25949 = n_25934 ^ n_25933;
assign n_25950 = n_25939 ^ n_25290;
assign n_25951 = n_25940 ^ x126;
assign n_25952 = n_25941 ^ n_24251;
assign n_25953 = n_25942 ^ n_25940;
assign n_25954 = n_25462 ^ n_25944;
assign n_25955 = n_25945 ^ n_25944;
assign n_25956 = n_25945 ^ n_25462;
assign n_25957 = n_25946 ^ n_24012;
assign n_25958 = n_25947 ^ n_25946;
assign n_25959 = n_25947 ^ n_24012;
assign n_25960 = ~n_25949 & n_25948;
assign n_25961 = n_25949 ^ x193;
assign n_25962 = n_25066 ^ n_25950;
assign n_25963 = ~n_25950 & n_25304;
assign n_25964 = n_25952 ^ n_25924;
assign n_25965 = ~n_25953 & n_25951;
assign n_25966 = n_25953 ^ x126;
assign n_25967 = ~n_25954 & ~n_25955;
assign n_25968 = n_25956 ^ n_25944;
assign n_25969 = n_25957 & n_25958;
assign n_25970 = n_25959 ^ n_25946;
assign n_25971 = n_25960 ^ x193;
assign n_25972 = n_25935 & n_25961;
assign n_25973 = n_25961 ^ n_25935;
assign n_25974 = n_25962 ^ n_25290;
assign n_25975 = n_25962 ^ n_25561;
assign n_25976 = n_25963 ^ n_25066;
assign n_25977 = n_25964 ^ n_24292;
assign n_25978 = n_25964 & ~n_25937;
assign n_25979 = n_25965 ^ x126;
assign n_25980 = n_25943 & n_25966;
assign n_25981 = n_25966 ^ n_25943;
assign n_25982 = n_25967 ^ n_25462;
assign n_25983 = n_25968 ^ n_25453;
assign n_25984 = n_25969 ^ n_24012;
assign n_25985 = n_25970 ^ x192;
assign n_25986 = n_25971 ^ n_25970;
assign n_25987 = n_25974 ^ n_24654;
assign n_25988 = n_25976 ^ n_25329;
assign n_25989 = n_25977 ^ x125;
assign n_25990 = n_25978 ^ n_24292;
assign n_25991 = n_25979 ^ n_25977;
assign n_25992 = n_25490 ^ n_25981;
assign n_25993 = n_25982 ^ n_25981;
assign n_25994 = n_25982 ^ n_25490;
assign n_25995 = n_25983 ^ n_24051;
assign n_25996 = n_25984 ^ n_25983;
assign n_25997 = n_25984 ^ n_24051;
assign n_25998 = ~n_25986 & n_25985;
assign n_25999 = n_25986 ^ x192;
assign n_26000 = n_25987 ^ n_24331;
assign n_26001 = n_25084 ^ n_25988;
assign n_26002 = ~n_25988 & n_25343;
assign n_26003 = n_25990 ^ n_24331;
assign n_26004 = n_25990 ^ n_25987;
assign n_26005 = ~n_25991 & n_25989;
assign n_26006 = n_25991 ^ x125;
assign n_26007 = ~n_25992 & n_25993;
assign n_26008 = n_25994 ^ n_25981;
assign n_26009 = ~n_25995 & ~n_25996;
assign n_26010 = n_25997 ^ n_25983;
assign n_26011 = n_25998 ^ x192;
assign n_26012 = n_25972 & n_25999;
assign n_26013 = n_25999 ^ n_25972;
assign n_26014 = n_26001 ^ n_25329;
assign n_26015 = n_25582 ^ n_26001;
assign n_26016 = n_26002 ^ n_25084;
assign n_26017 = n_26003 ^ n_25987;
assign n_26018 = n_26000 & n_26004;
assign n_26019 = n_26005 ^ x125;
assign n_26020 = ~n_26006 & ~n_25980;
assign n_26021 = n_25980 ^ n_26006;
assign n_26022 = n_26007 ^ n_25490;
assign n_26023 = n_26008 ^ n_25484;
assign n_26024 = n_26009 ^ n_24051;
assign n_26025 = n_26010 ^ x207;
assign n_26026 = n_26011 ^ n_26010;
assign n_26027 = n_26014 ^ n_24677;
assign n_26028 = n_26016 ^ n_25368;
assign n_26029 = n_26017 ^ x124;
assign n_26030 = n_26018 ^ n_24331;
assign n_26031 = n_26019 ^ n_26017;
assign n_26032 = n_25513 ^ n_26021;
assign n_26033 = n_26022 ^ n_26021;
assign n_26034 = n_26022 ^ n_25513;
assign n_26035 = n_26023 ^ n_24091;
assign n_26036 = n_26024 ^ n_26023;
assign n_26037 = n_26024 ^ n_24091;
assign n_26038 = ~n_26026 & n_26025;
assign n_26039 = n_26026 ^ x207;
assign n_26040 = n_26027 ^ n_24371;
assign n_26041 = n_25103 ^ n_26028;
assign n_26042 = ~n_26028 & ~n_25382;
assign n_26043 = n_26030 ^ n_24371;
assign n_26044 = n_26030 ^ n_26027;
assign n_26045 = n_26031 & ~n_26029;
assign n_26046 = n_26031 ^ x124;
assign n_26047 = n_26032 & ~n_26033;
assign n_26048 = n_26034 ^ n_26021;
assign n_26049 = ~n_26035 & ~n_26036;
assign n_26050 = n_26037 ^ n_26023;
assign n_26051 = n_26038 ^ x207;
assign n_26052 = ~n_26012 & ~n_26039;
assign n_26053 = n_26041 ^ n_25368;
assign n_26054 = n_25604 ^ n_26041;
assign n_26055 = n_26042 ^ n_25103;
assign n_26056 = n_26043 ^ n_26027;
assign n_26057 = ~n_26040 & ~n_26044;
assign n_26058 = n_26045 ^ x124;
assign n_26059 = ~n_26046 & ~n_26020;
assign n_26060 = n_26020 ^ n_26046;
assign n_26061 = n_26047 ^ n_25513;
assign n_26062 = n_26048 ^ n_25506;
assign n_26063 = n_26049 ^ n_24091;
assign n_26064 = n_26050 ^ x206;
assign n_26065 = n_26051 ^ n_26050;
assign n_26066 = n_26053 ^ n_24697;
assign n_26067 = n_26055 ^ n_25407;
assign n_26068 = n_26056 ^ x123;
assign n_26069 = n_26057 ^ n_24371;
assign n_26070 = n_26058 ^ n_26056;
assign n_26071 = n_26060 ^ n_25529;
assign n_26072 = n_26061 ^ n_26060;
assign n_26073 = n_26061 ^ n_25529;
assign n_26074 = n_26062 ^ n_24128;
assign n_26075 = n_26063 ^ n_26062;
assign n_26076 = n_26063 ^ n_24128;
assign n_26077 = n_26065 & ~n_26064;
assign n_26078 = n_26065 ^ x206;
assign n_26079 = n_26066 ^ n_24411;
assign n_26080 = n_25122 ^ n_26067;
assign n_26081 = n_26067 & ~n_25421;
assign n_26082 = n_26069 ^ n_24411;
assign n_26083 = n_26069 ^ n_26066;
assign n_26084 = n_26070 & ~n_26068;
assign n_26085 = n_26070 ^ x123;
assign n_26086 = ~n_26071 & n_26072;
assign n_26087 = n_26073 ^ n_26060;
assign n_26088 = ~n_26074 & ~n_26075;
assign n_26089 = n_26076 ^ n_26062;
assign n_26090 = n_26077 ^ x206;
assign n_26091 = ~n_26078 & ~n_26052;
assign n_26092 = n_26052 ^ n_26078;
assign n_26093 = n_26080 ^ n_25407;
assign n_26094 = n_25625 ^ n_26080;
assign n_26095 = n_26081 ^ n_25122;
assign n_26096 = n_26082 ^ n_26066;
assign n_26097 = n_26079 & n_26083;
assign n_26098 = n_26084 ^ x123;
assign n_26099 = n_26085 & ~n_26059;
assign n_26100 = n_26059 ^ n_26085;
assign n_26101 = n_26086 ^ n_25529;
assign n_26102 = n_26087 ^ n_25534;
assign n_26103 = n_26088 ^ n_24128;
assign n_26104 = n_26089 ^ x205;
assign n_26105 = n_26090 ^ n_26089;
assign n_26106 = n_26092 & n_25680;
assign n_26107 = n_26092 ^ n_25159;
assign n_26108 = n_26093 ^ n_24719;
assign n_26109 = n_26095 ^ n_25446;
assign n_26110 = n_26096 ^ x122;
assign n_26111 = n_26097 ^ n_24411;
assign n_26112 = n_26098 ^ n_26096;
assign n_26113 = n_26100 ^ n_25542;
assign n_26114 = n_26101 ^ n_26100;
assign n_26115 = n_26101 ^ n_25542;
assign n_26116 = n_26102 ^ n_24167;
assign n_26117 = n_26103 ^ n_26102;
assign n_26118 = n_26103 ^ n_24167;
assign n_26119 = ~n_26105 & n_26104;
assign n_26120 = n_26105 ^ x205;
assign n_26121 = n_26106 ^ n_25699;
assign n_26122 = ~n_24732 & n_26107;
assign n_26123 = x295 & ~n_26107;
assign n_26124 = n_26107 ^ x295;
assign n_26125 = n_26107 ^ n_25670;
assign n_26126 = n_26108 ^ n_24450;
assign n_26127 = n_26109 ^ n_25141;
assign n_26128 = n_26111 ^ n_24450;
assign n_26129 = n_26111 ^ n_26108;
assign n_26130 = n_26112 & ~n_26110;
assign n_26131 = n_26112 ^ x122;
assign n_26132 = n_26113 & n_26114;
assign n_26133 = n_26115 ^ n_26100;
assign n_26134 = ~n_26116 & n_26117;
assign n_26135 = n_26118 ^ n_26102;
assign n_26136 = n_26119 ^ x205;
assign n_26137 = ~n_26091 & ~n_26120;
assign n_26138 = n_26120 ^ n_26091;
assign n_26139 = n_26122 ^ n_24754;
assign n_26140 = n_26123 ^ x294;
assign n_26141 = n_26127 ^ n_25446;
assign n_26142 = n_26128 ^ n_26108;
assign n_26143 = ~n_26126 & n_26129;
assign n_26144 = n_26130 ^ x122;
assign n_26145 = ~n_26099 & ~n_26131;
assign n_26146 = n_26131 ^ n_26099;
assign n_26147 = n_26132 ^ n_25542;
assign n_26148 = n_26133 ^ n_25547;
assign n_26149 = n_26134 ^ n_24167;
assign n_26150 = n_26135 ^ x204;
assign n_26151 = n_26136 ^ n_26135;
assign n_26152 = n_26138 ^ n_26106;
assign n_26153 = n_26121 ^ n_26138;
assign n_26154 = n_26141 ^ n_24736;
assign n_26155 = n_26142 ^ x121;
assign n_26156 = n_26143 ^ n_24450;
assign n_26157 = n_26144 ^ n_26142;
assign n_26158 = n_26146 ^ n_25557;
assign n_26159 = n_26147 ^ n_26146;
assign n_26160 = n_26147 ^ n_25557;
assign n_26161 = n_26148 ^ n_24207;
assign n_26162 = n_26149 ^ n_26148;
assign n_26163 = n_26149 ^ n_24207;
assign n_26164 = n_26151 & ~n_26150;
assign n_26165 = n_26151 ^ x204;
assign n_26166 = n_26152 & ~n_26121;
assign n_26167 = n_26152 ^ n_25197;
assign n_26168 = n_26154 ^ n_24478;
assign n_26169 = n_26156 ^ x120;
assign n_26170 = n_26157 & ~n_26155;
assign n_26171 = n_26157 ^ x121;
assign n_26172 = n_26158 & ~n_26159;
assign n_26173 = n_26160 ^ n_26146;
assign n_26174 = n_26161 & n_26162;
assign n_26175 = n_26163 ^ n_26148;
assign n_26176 = n_26164 ^ x204;
assign n_26177 = n_26165 & n_26137;
assign n_26178 = n_26137 ^ n_26165;
assign n_26179 = n_26166 ^ n_25699;
assign n_26180 = n_26167 ^ n_26122;
assign n_26181 = n_26167 ^ n_26139;
assign n_26182 = n_26169 ^ n_26168;
assign n_26183 = n_26170 ^ x121;
assign n_26184 = ~n_26145 & n_26171;
assign n_26185 = n_26171 ^ n_26145;
assign n_26186 = n_26172 ^ n_25557;
assign n_26187 = n_26173 ^ n_25564;
assign n_26188 = n_26174 ^ n_24207;
assign n_26189 = n_26175 ^ x203;
assign n_26190 = n_26176 ^ n_26175;
assign n_26191 = n_26178 ^ n_25737;
assign n_26192 = n_26179 ^ n_26178;
assign n_26193 = n_26179 ^ n_25737;
assign n_26194 = n_26139 & ~n_26180;
assign n_26195 = n_26181 ^ n_26123;
assign n_26196 = n_26181 ^ n_26140;
assign n_26197 = n_26183 ^ n_26184;
assign n_26198 = n_26185 ^ n_25573;
assign n_26199 = n_26186 ^ n_26185;
assign n_26200 = n_26186 ^ n_25573;
assign n_26201 = n_26187 ^ n_24247;
assign n_26202 = n_26188 ^ n_26187;
assign n_26203 = n_26188 ^ n_24247;
assign n_26204 = ~n_26190 & n_26189;
assign n_26205 = n_26190 ^ x203;
assign n_26206 = ~n_26192 & ~n_26191;
assign n_26207 = n_26192 ^ n_25237;
assign n_26208 = n_26193 ^ n_26178;
assign n_26209 = n_26194 ^ n_24754;
assign n_26210 = n_26140 & ~n_26195;
assign n_26211 = ~n_26124 & n_26196;
assign n_26212 = n_26196 ^ n_26124;
assign n_26213 = n_26197 ^ n_26182;
assign n_26214 = n_26198 & ~n_26199;
assign n_26215 = n_26200 ^ n_26185;
assign n_26216 = n_26201 & ~n_26202;
assign n_26217 = n_26203 ^ n_26187;
assign n_26218 = n_26204 ^ x203;
assign n_26219 = n_26177 & ~n_26205;
assign n_26220 = n_26205 ^ n_26177;
assign n_26221 = n_26206 ^ n_25737;
assign n_26222 = n_26207 ^ n_24780;
assign n_26223 = n_26209 ^ n_26207;
assign n_26224 = n_26209 ^ n_24780;
assign n_26225 = n_26210 ^ x294;
assign n_26226 = n_26213 ^ n_25592;
assign n_26227 = n_26214 ^ n_25573;
assign n_26228 = n_26215 ^ n_25580;
assign n_26229 = n_26216 ^ n_24247;
assign n_26230 = n_26217 ^ x202;
assign n_26231 = n_26218 ^ n_26217;
assign n_26232 = n_26220 ^ n_25775;
assign n_26233 = n_26221 ^ n_26220;
assign n_26234 = n_26221 ^ n_25775;
assign n_26235 = ~n_26222 & n_26223;
assign n_26236 = n_26224 ^ n_26207;
assign n_26237 = n_26227 ^ n_26213;
assign n_26238 = n_26227 ^ n_25592;
assign n_26239 = n_26228 ^ n_24288;
assign n_26240 = n_26229 ^ n_26228;
assign n_26241 = n_26229 ^ n_24288;
assign n_26242 = n_26231 & ~n_26230;
assign n_26243 = n_26231 ^ x202;
assign n_26244 = ~n_26233 & n_26232;
assign n_26245 = n_26233 ^ n_25271;
assign n_26246 = n_26234 ^ n_26220;
assign n_26247 = n_26235 ^ n_24780;
assign n_26248 = n_26225 ^ n_26236;
assign n_26249 = n_26236 ^ x293;
assign n_26250 = ~n_26226 & n_26237;
assign n_26251 = n_26238 ^ n_26213;
assign n_26252 = n_26239 & ~n_26240;
assign n_26253 = n_26241 ^ n_26228;
assign n_26254 = n_26242 ^ x202;
assign n_26255 = ~n_26243 & ~n_26219;
assign n_26256 = n_26219 ^ n_26243;
assign n_26257 = n_26244 ^ n_25775;
assign n_26258 = n_26245 ^ n_24797;
assign n_26259 = n_26247 ^ n_26245;
assign n_26260 = n_26247 ^ n_24797;
assign n_26261 = n_26248 ^ x293;
assign n_26262 = n_26248 & ~n_26249;
assign n_26263 = n_26250 ^ n_25592;
assign n_26264 = n_26251 ^ n_25599;
assign n_26265 = n_26252 ^ n_24288;
assign n_26266 = n_26253 ^ x201;
assign n_26267 = n_26254 ^ n_26253;
assign n_26268 = n_26256 ^ n_25814;
assign n_26269 = n_26257 ^ n_26256;
assign n_26270 = n_26257 ^ n_25814;
assign n_26271 = ~n_26258 & ~n_26259;
assign n_26272 = n_26260 ^ n_26245;
assign n_26273 = ~n_26261 & n_26211;
assign n_26274 = n_26211 ^ n_26261;
assign n_26275 = n_26262 ^ x293;
assign n_26276 = n_26263 ^ n_25606;
assign n_26277 = n_26263 ^ n_25177;
assign n_26278 = n_26264 ^ n_24327;
assign n_26279 = n_26265 ^ n_26264;
assign n_26280 = n_26265 ^ n_24327;
assign n_26281 = n_26267 & ~n_26266;
assign n_26282 = n_26267 ^ x201;
assign n_26283 = ~n_26269 & n_26268;
assign n_26284 = n_26269 ^ n_25309;
assign n_26285 = n_26270 ^ n_26256;
assign n_26286 = n_26271 ^ n_24797;
assign n_26287 = n_26272 ^ x292;
assign n_26288 = n_26275 ^ n_26272;
assign n_26289 = n_25612 & ~n_26276;
assign n_26290 = n_26277 ^ n_25606;
assign n_26291 = n_26278 & ~n_26279;
assign n_26292 = n_26280 ^ n_26264;
assign n_26293 = n_26281 ^ x201;
assign n_26294 = ~n_26282 & n_26255;
assign n_26295 = n_26255 ^ n_26282;
assign n_26296 = n_26283 ^ n_25814;
assign n_26297 = n_26284 ^ n_24812;
assign n_26298 = n_26285 ^ n_26124;
assign n_26299 = n_26286 ^ n_26284;
assign n_26300 = n_26286 ^ n_24812;
assign n_26301 = n_26288 & ~n_26287;
assign n_26302 = n_26288 ^ x292;
assign n_26303 = n_26289 ^ n_25177;
assign n_26304 = n_26290 ^ n_25613;
assign n_26305 = n_26291 ^ n_24327;
assign n_26306 = n_26292 ^ x200;
assign n_26307 = n_26293 ^ n_26292;
assign n_26308 = n_26295 ^ n_25855;
assign n_26309 = n_26296 ^ n_26295;
assign n_26310 = n_26296 ^ n_25855;
assign n_26311 = ~n_26297 & ~n_26299;
assign n_26312 = n_26300 ^ n_26284;
assign n_26313 = n_26301 ^ x292;
assign n_26314 = ~n_26273 & n_26302;
assign n_26315 = n_26302 ^ n_26273;
assign n_26316 = n_26303 ^ n_25633;
assign n_26317 = n_26303 ^ n_25235;
assign n_26318 = n_26304 ^ n_24367;
assign n_26319 = n_26305 ^ n_26304;
assign n_26320 = n_26307 & ~n_26306;
assign n_26321 = n_26307 ^ x200;
assign n_26322 = n_26309 & ~n_26308;
assign n_26323 = n_26309 ^ n_25348;
assign n_26324 = n_26310 ^ n_26295;
assign n_26325 = n_26311 ^ n_24812;
assign n_26326 = n_26312 ^ x291;
assign n_26327 = n_26313 ^ n_26312;
assign n_26328 = n_25639 & n_26316;
assign n_26329 = n_26317 ^ n_25633;
assign n_26330 = n_26319 & n_26318;
assign n_26331 = n_26319 ^ n_24367;
assign n_26332 = n_26320 ^ x200;
assign n_26333 = ~n_26321 & n_26294;
assign n_26334 = n_26294 ^ n_26321;
assign n_26335 = n_26322 ^ n_25855;
assign n_26336 = n_26323 ^ n_24824;
assign n_26337 = n_26212 ^ n_26324;
assign n_26338 = n_26325 ^ n_26323;
assign n_26339 = n_26325 ^ n_24824;
assign n_26340 = ~n_26327 & n_26326;
assign n_26341 = n_26327 ^ x291;
assign n_26342 = n_26328 ^ n_25235;
assign n_26343 = n_26329 ^ n_25627;
assign n_26344 = n_26330 ^ n_24367;
assign n_26345 = n_26331 ^ x215;
assign n_26346 = n_26332 ^ n_26331;
assign n_26347 = n_26332 ^ x215;
assign n_26348 = n_26334 ^ n_25891;
assign n_26349 = n_26334 ^ n_26335;
assign n_26350 = n_26335 ^ n_25891;
assign n_26351 = n_26336 & n_26338;
assign n_26352 = n_26339 ^ n_26323;
assign n_26353 = n_26340 ^ x291;
assign n_26354 = n_26314 & ~n_26341;
assign n_26355 = n_26341 ^ n_26314;
assign n_26356 = n_26342 ^ n_25652;
assign n_26357 = n_26343 ^ n_24406;
assign n_26358 = n_26344 ^ n_26343;
assign n_26359 = ~n_26345 & n_26346;
assign n_26360 = n_26347 ^ n_26331;
assign n_26361 = n_26349 & n_26348;
assign n_26362 = n_26349 ^ n_25387;
assign n_26363 = n_26350 ^ n_26334;
assign n_26364 = n_26351 ^ n_24824;
assign n_26365 = n_26352 ^ x290;
assign n_26366 = n_26353 ^ n_26352;
assign n_26367 = n_26356 & ~n_25658;
assign n_26368 = n_25293 ^ n_26356;
assign n_26369 = n_26358 & ~n_26357;
assign n_26370 = n_26358 ^ n_24406;
assign n_26371 = n_26359 ^ x215;
assign n_26372 = ~n_26360 & n_26333;
assign n_26373 = n_26333 ^ n_26360;
assign n_26374 = n_26361 ^ n_25891;
assign n_26375 = n_26362 ^ n_24847;
assign n_26376 = n_26274 ^ n_26363;
assign n_26377 = n_26364 ^ n_26362;
assign n_26378 = n_26364 ^ n_24847;
assign n_26379 = ~n_26366 & n_26365;
assign n_26380 = n_26366 ^ x290;
assign n_26381 = n_26367 ^ n_25293;
assign n_26382 = n_26368 ^ n_25657;
assign n_26383 = n_26369 ^ n_24406;
assign n_26384 = n_26370 ^ x214;
assign n_26385 = n_26371 ^ n_26370;
assign n_26386 = n_26373 ^ n_25931;
assign n_26387 = n_26373 ^ n_26374;
assign n_26388 = n_26374 ^ n_25931;
assign n_26389 = ~n_26375 & ~n_26377;
assign n_26390 = n_26378 ^ n_26362;
assign n_26391 = n_26379 ^ x290;
assign n_26392 = n_26354 & ~n_26380;
assign n_26393 = n_26380 ^ n_26354;
assign n_26394 = n_26381 ^ n_25673;
assign n_26395 = n_26383 ^ n_26382;
assign n_26396 = n_26383 ^ n_24446;
assign n_26397 = n_26385 & ~n_26384;
assign n_26398 = n_26385 ^ x214;
assign n_26399 = ~n_26387 & ~n_26386;
assign n_26400 = n_26387 ^ n_25426;
assign n_26401 = n_26388 ^ n_26373;
assign n_26402 = n_26389 ^ n_24847;
assign n_26403 = n_26390 ^ x289;
assign n_26404 = n_26391 ^ n_26390;
assign n_26405 = ~n_26394 & n_25685;
assign n_26406 = n_25332 ^ n_26394;
assign n_26407 = n_26395 ^ n_24446;
assign n_26408 = ~n_26395 & n_26396;
assign n_26409 = n_26397 ^ x214;
assign n_26410 = ~n_26398 & n_26372;
assign n_26411 = n_26372 ^ n_26398;
assign n_26412 = n_26399 ^ n_25931;
assign n_26413 = n_26400 ^ n_24865;
assign n_26414 = n_26315 ^ n_26401;
assign n_26415 = n_26402 ^ n_26400;
assign n_26416 = n_26402 ^ n_24865;
assign n_26417 = ~n_26404 & n_26403;
assign n_26418 = n_26404 ^ x289;
assign n_26419 = n_26405 ^ n_25332;
assign n_26420 = n_26406 ^ n_25684;
assign n_26421 = n_26407 ^ x213;
assign n_26422 = n_26408 ^ n_24446;
assign n_26423 = n_26409 ^ n_26407;
assign n_26424 = n_26411 ^ n_25968;
assign n_26425 = n_26412 ^ n_26411;
assign n_26426 = n_26412 ^ n_25968;
assign n_26427 = ~n_26413 & ~n_26415;
assign n_26428 = n_26416 ^ n_26400;
assign n_26429 = n_26417 ^ x289;
assign n_26430 = ~n_26392 & n_26418;
assign n_26431 = n_26418 ^ n_26392;
assign n_26432 = n_26419 ^ n_25701;
assign n_26433 = n_26420 ^ n_24485;
assign n_26434 = n_26422 ^ n_26420;
assign n_26435 = n_26422 ^ n_24485;
assign n_26436 = ~n_26423 & n_26421;
assign n_26437 = n_26423 ^ x213;
assign n_26438 = n_26425 & n_26424;
assign n_26439 = n_26425 ^ n_25462;
assign n_26440 = n_26426 ^ n_26411;
assign n_26441 = n_26427 ^ n_24865;
assign n_26442 = n_26428 ^ x288;
assign n_26443 = n_26429 ^ n_26428;
assign n_26444 = n_26432 & ~n_25711;
assign n_26445 = n_25371 ^ n_26432;
assign n_26446 = n_26433 & ~n_26434;
assign n_26447 = n_26435 ^ n_26420;
assign n_26448 = n_26436 ^ x213;
assign n_26449 = n_26437 & n_26410;
assign n_26450 = n_26410 ^ n_26437;
assign n_26451 = n_26438 ^ n_25968;
assign n_26452 = n_26439 ^ n_24883;
assign n_26453 = n_26355 ^ n_26440;
assign n_26454 = n_26441 ^ n_26439;
assign n_26455 = n_26441 ^ n_24883;
assign n_26456 = n_26443 & ~n_26442;
assign n_26457 = n_26443 ^ x288;
assign n_26458 = n_26444 ^ n_25371;
assign n_26459 = n_26445 ^ n_25710;
assign n_26460 = n_26446 ^ n_24485;
assign n_26461 = n_26447 ^ x212;
assign n_26462 = n_26448 ^ n_26447;
assign n_26463 = n_26450 ^ n_26008;
assign n_26464 = n_26450 ^ n_26451;
assign n_26465 = n_26451 ^ n_26008;
assign n_26466 = ~n_26452 & n_26454;
assign n_26467 = n_26455 ^ n_26439;
assign n_26468 = n_26456 ^ x288;
assign n_26469 = ~n_26457 & n_26430;
assign n_26470 = n_26430 ^ n_26457;
assign n_26471 = n_26458 ^ n_25730;
assign n_26472 = n_26458 ^ n_25410;
assign n_26473 = n_26459 ^ n_24520;
assign n_26474 = n_26460 ^ n_26459;
assign n_26475 = n_26460 ^ n_24520;
assign n_26476 = ~n_26462 & n_26461;
assign n_26477 = n_26462 ^ x212;
assign n_26478 = n_26464 & n_26463;
assign n_26479 = n_26464 ^ n_25490;
assign n_26480 = n_26465 ^ n_26450;
assign n_26481 = n_26466 ^ n_24883;
assign n_26482 = n_26467 ^ x303;
assign n_26483 = n_26468 ^ n_26467;
assign n_26484 = n_25743 & n_26471;
assign n_26485 = n_26472 ^ n_25730;
assign n_26486 = n_26473 & ~n_26474;
assign n_26487 = n_26475 ^ n_26459;
assign n_26488 = n_26476 ^ x212;
assign n_26489 = ~n_26477 & ~n_26449;
assign n_26490 = n_26449 ^ n_26477;
assign n_26491 = n_26478 ^ n_26008;
assign n_26492 = n_26479 ^ n_24901;
assign n_26493 = n_26393 ^ n_26480;
assign n_26494 = n_26481 ^ n_26479;
assign n_26495 = n_26481 ^ n_24901;
assign n_26496 = ~n_26483 & n_26482;
assign n_26497 = n_26483 ^ x303;
assign n_26498 = n_26484 ^ n_25410;
assign n_26499 = n_26485 ^ n_25744;
assign n_26500 = n_26486 ^ n_24520;
assign n_26501 = n_26487 ^ x211;
assign n_26502 = n_26488 ^ n_26487;
assign n_26503 = n_26490 ^ n_26048;
assign n_26504 = n_26490 ^ n_26491;
assign n_26505 = n_26491 ^ n_26048;
assign n_26506 = ~n_26492 & n_26494;
assign n_26507 = n_26495 ^ n_26479;
assign n_26508 = n_26496 ^ x303;
assign n_26509 = n_26469 & n_26497;
assign n_26510 = n_26497 ^ n_26469;
assign n_26511 = n_26498 ^ n_25768;
assign n_26512 = n_26499 ^ n_24547;
assign n_26513 = n_26500 ^ n_26499;
assign n_26514 = n_26500 ^ n_24547;
assign n_26515 = ~n_26502 & n_26501;
assign n_26516 = n_26502 ^ x211;
assign n_26517 = n_26504 & n_26503;
assign n_26518 = n_26504 ^ n_25513;
assign n_26519 = n_26505 ^ n_26490;
assign n_26520 = n_26506 ^ n_24901;
assign n_26521 = n_26507 ^ x302;
assign n_26522 = n_26508 ^ n_26507;
assign n_26523 = n_26511 & n_25780;
assign n_26524 = n_25448 ^ n_26511;
assign n_26525 = ~n_26512 & ~n_26513;
assign n_26526 = n_26514 ^ n_26499;
assign n_26527 = n_26515 ^ x211;
assign n_26528 = ~n_26489 & n_26516;
assign n_26529 = n_26516 ^ n_26489;
assign n_26530 = n_26517 ^ n_26048;
assign n_26531 = n_26518 ^ n_24919;
assign n_26532 = n_26431 ^ n_26519;
assign n_26533 = n_26520 ^ n_26518;
assign n_26534 = n_26520 ^ n_24919;
assign n_26535 = ~n_26522 & n_26521;
assign n_26536 = n_26522 ^ x302;
assign n_26537 = n_26523 ^ n_25448;
assign n_26538 = n_26524 ^ n_25779;
assign n_26539 = n_26525 ^ n_24547;
assign n_26540 = n_26526 ^ x210;
assign n_26541 = n_26527 ^ n_26526;
assign n_26542 = n_26529 ^ n_26087;
assign n_26543 = n_26530 ^ n_26529;
assign n_26544 = n_26530 ^ n_26087;
assign n_26545 = ~n_26531 & n_26533;
assign n_26546 = n_26534 ^ n_26518;
assign n_26547 = n_26535 ^ x302;
assign n_26548 = n_26509 & n_26536;
assign n_26549 = n_26536 ^ n_26509;
assign n_26550 = n_26537 ^ n_25805;
assign n_26551 = n_26538 ^ n_24568;
assign n_26552 = n_26539 ^ n_26538;
assign n_26553 = n_26539 ^ n_24568;
assign n_26554 = n_26541 & ~n_26540;
assign n_26555 = n_26541 ^ x210;
assign n_26556 = ~n_26543 & ~n_26542;
assign n_26557 = n_26543 ^ n_25529;
assign n_26558 = n_26544 ^ n_26529;
assign n_26559 = n_26545 ^ n_24919;
assign n_26560 = n_26546 ^ x301;
assign n_26561 = n_26547 ^ n_26546;
assign n_26562 = n_25478 ^ n_26550;
assign n_26563 = n_26550 & n_25817;
assign n_26564 = ~n_26551 & ~n_26552;
assign n_26565 = n_26553 ^ n_26538;
assign n_26566 = n_26554 ^ x210;
assign n_26567 = ~n_26555 & n_26528;
assign n_26568 = n_26528 ^ n_26555;
assign n_26569 = n_26556 ^ n_26087;
assign n_26570 = n_26557 ^ n_24937;
assign n_26571 = n_26470 ^ n_26558;
assign n_26572 = n_26559 ^ n_26557;
assign n_26573 = n_26559 ^ n_24937;
assign n_26574 = ~n_26561 & n_26560;
assign n_26575 = n_26561 ^ x301;
assign n_26576 = n_26562 ^ n_25816;
assign n_26577 = n_25682 ^ n_26562;
assign n_26578 = n_26563 ^ n_25478;
assign n_26579 = n_26564 ^ n_24568;
assign n_26580 = n_26565 ^ x209;
assign n_26581 = n_26566 ^ n_26565;
assign n_26582 = n_26568 ^ n_26133;
assign n_26583 = n_26569 ^ n_26568;
assign n_26584 = n_26569 ^ n_26133;
assign n_26585 = ~n_26570 & ~n_26572;
assign n_26586 = n_26573 ^ n_26557;
assign n_26587 = n_26574 ^ x301;
assign n_26588 = n_26575 & n_26548;
assign n_26589 = n_26548 ^ n_26575;
assign n_26590 = n_26576 ^ n_24585;
assign n_26591 = n_26578 ^ n_25830;
assign n_26592 = n_26579 ^ n_26576;
assign n_26593 = n_26579 ^ n_24585;
assign n_26594 = ~n_26581 & n_26580;
assign n_26595 = n_26581 ^ x209;
assign n_26596 = n_26583 & n_26582;
assign n_26597 = n_26583 ^ n_25542;
assign n_26598 = n_26584 ^ n_26568;
assign n_26599 = n_26585 ^ n_24937;
assign n_26600 = n_26586 ^ x300;
assign n_26601 = n_26587 ^ n_26586;
assign n_26602 = n_25502 ^ n_26591;
assign n_26603 = n_26591 & ~n_25845;
assign n_26604 = n_26590 & n_26592;
assign n_26605 = n_26593 ^ n_26576;
assign n_26606 = n_26594 ^ x209;
assign n_26607 = n_26595 & n_26567;
assign n_26608 = n_26567 ^ n_26595;
assign n_26609 = n_26596 ^ n_26133;
assign n_26610 = n_26597 ^ n_24956;
assign n_26611 = n_26510 ^ n_26598;
assign n_26612 = n_26599 ^ n_26597;
assign n_26613 = n_26599 ^ n_24956;
assign n_26614 = ~n_26601 & n_26600;
assign n_26615 = n_26601 ^ x300;
assign n_26616 = n_26602 ^ n_25844;
assign n_26617 = n_25742 ^ n_26602;
assign n_26618 = n_26603 ^ n_25502;
assign n_26619 = n_26604 ^ n_24585;
assign n_26620 = n_26605 ^ x208;
assign n_26621 = n_26606 ^ n_26605;
assign n_26622 = n_26608 ^ n_26173;
assign n_26623 = n_26609 ^ n_26608;
assign n_26624 = n_26609 ^ n_26173;
assign n_26625 = ~n_26610 & n_26612;
assign n_26626 = n_26613 ^ n_26597;
assign n_26627 = n_26614 ^ x300;
assign n_26628 = n_26588 & n_26615;
assign n_26629 = n_26615 ^ n_26588;
assign n_26630 = n_26616 ^ n_24604;
assign n_26631 = n_26618 ^ n_25521;
assign n_26632 = n_26618 ^ n_25885;
assign n_26633 = n_26619 ^ n_26616;
assign n_26634 = ~n_26621 & n_26620;
assign n_26635 = n_26621 ^ x208;
assign n_26636 = n_26623 & n_26622;
assign n_26637 = n_26623 ^ n_25557;
assign n_26638 = n_26624 ^ n_26608;
assign n_26639 = n_26625 ^ n_24956;
assign n_26640 = n_26626 ^ x299;
assign n_26641 = n_26627 ^ n_26626;
assign n_26642 = n_26631 ^ n_25885;
assign n_26643 = n_25898 & ~n_26632;
assign n_26644 = n_26633 ^ n_24604;
assign n_26645 = ~n_26633 & n_26630;
assign n_26646 = n_26634 ^ x208;
assign n_26647 = ~n_26635 & ~n_26607;
assign n_26648 = n_26607 ^ n_26635;
assign n_26649 = n_26636 ^ n_26173;
assign n_26650 = n_26637 ^ n_24975;
assign n_26651 = n_26638 ^ n_26549;
assign n_26652 = n_26639 ^ n_26637;
assign n_26653 = n_26639 ^ n_24975;
assign n_26654 = n_26641 & ~n_26640;
assign n_26655 = n_26641 ^ x299;
assign n_26656 = n_26642 ^ n_25871;
assign n_26657 = n_25803 ^ n_26642;
assign n_26658 = n_26643 ^ n_25521;
assign n_26659 = n_26644 ^ x223;
assign n_26660 = n_26645 ^ n_24604;
assign n_26661 = n_26646 ^ n_26644;
assign n_26662 = n_26646 ^ x223;
assign n_26663 = n_26648 ^ n_26215;
assign n_26664 = n_26649 ^ n_26648;
assign n_26665 = n_26649 ^ n_26215;
assign n_26666 = n_26650 & n_26652;
assign n_26667 = n_26653 ^ n_26637;
assign n_26668 = n_26654 ^ x299;
assign n_26669 = ~n_26628 & n_26655;
assign n_26670 = n_26655 ^ n_26628;
assign n_26671 = n_26656 ^ n_24624;
assign n_26672 = n_26658 ^ n_25925;
assign n_26673 = n_26660 ^ n_26656;
assign n_26674 = ~n_26659 & n_26661;
assign n_26675 = n_26662 ^ n_26644;
assign n_26676 = n_26664 & ~n_26663;
assign n_26677 = n_26664 ^ n_25573;
assign n_26678 = n_26665 ^ n_26648;
assign n_26679 = n_26666 ^ n_24975;
assign n_26680 = n_26667 ^ x298;
assign n_26681 = n_26668 ^ n_26667;
assign n_26682 = n_25537 ^ n_26672;
assign n_26683 = ~n_26672 & n_25938;
assign n_26684 = n_26673 ^ n_24624;
assign n_26685 = n_26673 & n_26671;
assign n_26686 = n_26674 ^ x223;
assign n_26687 = ~n_26675 & ~n_26647;
assign n_26688 = n_26647 ^ n_26675;
assign n_26689 = n_26676 ^ n_26215;
assign n_26690 = n_26677 ^ n_24994;
assign n_26691 = n_26589 ^ n_26678;
assign n_26692 = n_26679 ^ n_26677;
assign n_26693 = n_26679 ^ n_24994;
assign n_26694 = ~n_26681 & n_26680;
assign n_26695 = n_26681 ^ x298;
assign n_26696 = n_26682 ^ n_25910;
assign n_26697 = n_25852 ^ n_26682;
assign n_26698 = n_26683 ^ n_25537;
assign n_26699 = n_26684 ^ x222;
assign n_26700 = n_26685 ^ n_24624;
assign n_26701 = n_26686 ^ n_26684;
assign n_26702 = n_26688 ^ n_26251;
assign n_26703 = n_26689 ^ n_26688;
assign n_26704 = n_26689 ^ n_26251;
assign n_26705 = n_26690 & ~n_26692;
assign n_26706 = n_26693 ^ n_26677;
assign n_26707 = n_26694 ^ x298;
assign n_26708 = ~n_26669 & n_26695;
assign n_26709 = n_26695 ^ n_26669;
assign n_26710 = n_26696 ^ n_24643;
assign n_26711 = n_26698 ^ n_25561;
assign n_26712 = n_26698 ^ n_25962;
assign n_26713 = n_26700 ^ n_26696;
assign n_26714 = n_26701 & ~n_26699;
assign n_26715 = n_26701 ^ x222;
assign n_26716 = ~n_26703 & ~n_26702;
assign n_26717 = n_26703 ^ n_25592;
assign n_26718 = n_26704 ^ n_26688;
assign n_26719 = n_26705 ^ n_24994;
assign n_26720 = n_26706 ^ x297;
assign n_26721 = n_26707 ^ n_26706;
assign n_26722 = n_26711 ^ n_25962;
assign n_26723 = n_25975 & n_26712;
assign n_26724 = n_26713 ^ n_24643;
assign n_26725 = n_26713 & n_26710;
assign n_26726 = n_26714 ^ x222;
assign n_26727 = ~n_26715 & n_26687;
assign n_26728 = n_26687 ^ n_26715;
assign n_26729 = n_26716 ^ n_26251;
assign n_26730 = n_26717 ^ n_25013;
assign n_26731 = n_26718 ^ n_26629;
assign n_26732 = n_26719 ^ n_26717;
assign n_26733 = n_26719 ^ n_25013;
assign n_26734 = n_26721 & ~n_26720;
assign n_26735 = n_26721 ^ x297;
assign n_26736 = n_26722 ^ n_25974;
assign n_26737 = n_25895 ^ n_26722;
assign n_26738 = n_26723 ^ n_25561;
assign n_26739 = n_26724 ^ x221;
assign n_26740 = n_26725 ^ n_24643;
assign n_26741 = n_26726 ^ n_26724;
assign n_26742 = n_26728 ^ n_26290;
assign n_26743 = n_26729 ^ n_26728;
assign n_26744 = n_26730 & n_26732;
assign n_26745 = n_26733 ^ n_26717;
assign n_26746 = n_26734 ^ x297;
assign n_26747 = ~n_26708 & n_26735;
assign n_26748 = n_26735 ^ n_26708;
assign n_26749 = n_26736 ^ n_24654;
assign n_26750 = n_26738 ^ n_26001;
assign n_26751 = n_26740 ^ n_24654;
assign n_26752 = n_26740 ^ n_26736;
assign n_26753 = ~n_26741 & n_26739;
assign n_26754 = n_26741 ^ x221;
assign n_26755 = n_26742 ^ n_26729;
assign n_26756 = ~n_26743 & ~n_26742;
assign n_26757 = n_26743 ^ n_25606;
assign n_26758 = n_26744 ^ n_25013;
assign n_26759 = n_26745 ^ x296;
assign n_26760 = n_26746 ^ n_26745;
assign n_26761 = n_25582 ^ n_26750;
assign n_26762 = ~n_26750 & ~n_26015;
assign n_26763 = n_26751 ^ n_26736;
assign n_26764 = n_26749 & n_26752;
assign n_26765 = n_26753 ^ x221;
assign n_26766 = ~n_26754 & ~n_26727;
assign n_26767 = n_26727 ^ n_26754;
assign n_26768 = n_26670 ^ n_26755;
assign n_26769 = n_26756 ^ n_26290;
assign n_26770 = n_26757 ^ n_25026;
assign n_26771 = n_26758 ^ n_26757;
assign n_26772 = n_26760 & ~n_26759;
assign n_26773 = n_26760 ^ x296;
assign n_26774 = n_26761 ^ n_26014;
assign n_26775 = n_25936 ^ n_26761;
assign n_26776 = n_26762 ^ n_25582;
assign n_26777 = n_26763 ^ x220;
assign n_26778 = n_26764 ^ n_24654;
assign n_26779 = n_26765 ^ n_26763;
assign n_26780 = n_26767 ^ n_26329;
assign n_26781 = n_26769 ^ n_26767;
assign n_26782 = ~n_26771 & n_26770;
assign n_26783 = n_26771 ^ n_25026;
assign n_26784 = n_26772 ^ x296;
assign n_26785 = n_26747 & n_26773;
assign n_26786 = n_26773 ^ n_26747;
assign n_26787 = n_26774 ^ n_24677;
assign n_26788 = n_26776 ^ n_26041;
assign n_26789 = n_26778 ^ n_24677;
assign n_26790 = n_26778 ^ n_26774;
assign n_26791 = n_26779 & ~n_26777;
assign n_26792 = n_26779 ^ x220;
assign n_26793 = n_26781 & ~n_26780;
assign n_26794 = n_26781 ^ n_25633;
assign n_26795 = n_26781 ^ n_26329;
assign n_26796 = n_26782 ^ n_25026;
assign n_26797 = n_26783 ^ x311;
assign n_26798 = n_26784 ^ n_26783;
assign n_26799 = n_26784 ^ x311;
assign n_26800 = n_25604 ^ n_26788;
assign n_26801 = ~n_26788 & n_26054;
assign n_26802 = n_26789 ^ n_26774;
assign n_26803 = n_26787 & ~n_26790;
assign n_26804 = n_26791 ^ x220;
assign n_26805 = ~n_26792 & ~n_26766;
assign n_26806 = n_26766 ^ n_26792;
assign n_26807 = n_26793 ^ n_26329;
assign n_26808 = n_26794 ^ n_25051;
assign n_26809 = n_26795 ^ n_26709;
assign n_26810 = n_26796 ^ n_26794;
assign n_26811 = n_26797 & ~n_26798;
assign n_26812 = n_26799 ^ n_26783;
assign n_26813 = n_26800 ^ n_26053;
assign n_26814 = n_25973 ^ n_26800;
assign n_26815 = n_26801 ^ n_25604;
assign n_26816 = n_26802 ^ x219;
assign n_26817 = n_26803 ^ n_24677;
assign n_26818 = n_26804 ^ n_26802;
assign n_26819 = n_26806 ^ n_26368;
assign n_26820 = n_26807 ^ n_26806;
assign n_26821 = ~n_26810 & n_26808;
assign n_26822 = n_26810 ^ n_25051;
assign n_26823 = n_26811 ^ x311;
assign n_26824 = ~n_26785 & n_26812;
assign n_26825 = n_26812 ^ n_26785;
assign n_26826 = n_26813 ^ n_24697;
assign n_26827 = n_26815 ^ n_26080;
assign n_26828 = n_26817 ^ n_24697;
assign n_26829 = n_26817 ^ n_26813;
assign n_26830 = ~n_26818 & n_26816;
assign n_26831 = n_26818 ^ x219;
assign n_26832 = ~n_26820 & n_26819;
assign n_26833 = n_26820 ^ n_25652;
assign n_26834 = n_26820 ^ n_26368;
assign n_26835 = n_26821 ^ n_25051;
assign n_26836 = n_26822 ^ x310;
assign n_26837 = n_26823 ^ n_26822;
assign n_26838 = n_25625 ^ n_26827;
assign n_26839 = n_26827 & ~n_26094;
assign n_26840 = n_26828 ^ n_26813;
assign n_26841 = n_26826 & n_26829;
assign n_26842 = n_26830 ^ x219;
assign n_26843 = n_26831 & n_26805;
assign n_26844 = n_26805 ^ n_26831;
assign n_26845 = n_26832 ^ n_26368;
assign n_26846 = n_26833 ^ n_25070;
assign n_26847 = n_26748 ^ n_26834;
assign n_26848 = n_26835 ^ n_26833;
assign n_26849 = ~n_26837 & n_26836;
assign n_26850 = n_26837 ^ x310;
assign n_26851 = n_26838 ^ n_26093;
assign n_26852 = n_26013 ^ n_26838;
assign n_26853 = n_26839 ^ n_25625;
assign n_26854 = n_26840 ^ x218;
assign n_26855 = n_26841 ^ n_24697;
assign n_26856 = n_26842 ^ n_26840;
assign n_26857 = n_26844 ^ n_26406;
assign n_26858 = n_26845 ^ n_26844;
assign n_26859 = n_26845 ^ n_26406;
assign n_26860 = ~n_26848 & n_26846;
assign n_26861 = n_26848 ^ n_25070;
assign n_26862 = n_26849 ^ x310;
assign n_26863 = n_26824 & n_26850;
assign n_26864 = n_26850 ^ n_26824;
assign n_26865 = n_26851 ^ n_24719;
assign n_26866 = n_26853 ^ n_26127;
assign n_26867 = n_26855 ^ n_24719;
assign n_26868 = n_26855 ^ n_26851;
assign n_26869 = ~n_26856 & n_26854;
assign n_26870 = n_26856 ^ x218;
assign n_26871 = ~n_26858 & ~n_26857;
assign n_26872 = n_26858 ^ n_25673;
assign n_26873 = n_26859 ^ n_26844;
assign n_26874 = n_26860 ^ n_25070;
assign n_26875 = n_26861 ^ x309;
assign n_26876 = n_26862 ^ n_26861;
assign n_26877 = n_26866 ^ n_25645;
assign n_26878 = n_26867 ^ n_26851;
assign n_26879 = n_26865 & ~n_26868;
assign n_26880 = n_26869 ^ x218;
assign n_26881 = n_26843 & n_26870;
assign n_26882 = n_26870 ^ n_26843;
assign n_26883 = n_26871 ^ n_26406;
assign n_26884 = n_26872 ^ n_25088;
assign n_26885 = n_26786 ^ n_26873;
assign n_26886 = n_26872 ^ n_26874;
assign n_26887 = n_26874 ^ n_25088;
assign n_26888 = ~n_26876 & n_26875;
assign n_26889 = n_26876 ^ x309;
assign n_26890 = n_26877 ^ n_26154;
assign n_26891 = n_26877 ^ n_26012;
assign n_26892 = n_26878 ^ x217;
assign n_26893 = n_26879 ^ n_24719;
assign n_26894 = n_26880 ^ n_26878;
assign n_26895 = n_26882 ^ n_26445;
assign n_26896 = n_26883 ^ n_26882;
assign n_26897 = n_26883 ^ n_26445;
assign n_26898 = ~n_26884 & n_26886;
assign n_26899 = n_26872 ^ n_26887;
assign n_26900 = n_26888 ^ x309;
assign n_26901 = ~n_26863 & ~n_26889;
assign n_26902 = n_26889 ^ n_26863;
assign n_26903 = n_26891 ^ n_26039;
assign n_26904 = n_26893 ^ x216;
assign n_26905 = n_26894 & ~n_26892;
assign n_26906 = n_26894 ^ x217;
assign n_26907 = n_26896 & n_26895;
assign n_26908 = n_26896 ^ n_25701;
assign n_26909 = n_26897 ^ n_26882;
assign n_26910 = n_26898 ^ n_25088;
assign n_26911 = n_26899 ^ x308;
assign n_26912 = n_26900 ^ n_26899;
assign n_26913 = n_26904 ^ n_26890;
assign n_26914 = n_26905 ^ x217;
assign n_26915 = ~n_26906 & n_26881;
assign n_26916 = n_26881 ^ n_26906;
assign n_26917 = n_26907 ^ n_26445;
assign n_26918 = n_26908 ^ n_25107;
assign n_26919 = n_26825 ^ n_26909;
assign n_26920 = n_26910 ^ n_26908;
assign n_26921 = n_26910 ^ n_25107;
assign n_26922 = n_26912 & ~n_26911;
assign n_26923 = n_26912 ^ x308;
assign n_26924 = n_26914 ^ n_26913;
assign n_26925 = n_26916 ^ n_26485;
assign n_26926 = n_26917 ^ n_26916;
assign n_26927 = n_26917 ^ n_26485;
assign n_26928 = ~n_26918 & n_26920;
assign n_26929 = n_26921 ^ n_26908;
assign n_26930 = n_26922 ^ x308;
assign n_26931 = ~n_26923 & ~n_26901;
assign n_26932 = n_26901 ^ n_26923;
assign n_26933 = n_26924 ^ n_26915;
assign n_26934 = n_26926 & n_26925;
assign n_26935 = n_26926 ^ n_25730;
assign n_26936 = n_26927 ^ n_26916;
assign n_26937 = n_26928 ^ n_25107;
assign n_26938 = n_26929 ^ x307;
assign n_26939 = n_26930 ^ n_26929;
assign n_26940 = n_26933 ^ n_26524;
assign n_26941 = n_26934 ^ n_26485;
assign n_26942 = n_26935 ^ n_25126;
assign n_26943 = n_26864 ^ n_26936;
assign n_26944 = n_26937 ^ n_26935;
assign n_26945 = n_26937 ^ n_25126;
assign n_26946 = n_26939 & ~n_26938;
assign n_26947 = n_26939 ^ x307;
assign n_26948 = n_26933 ^ n_26941;
assign n_26949 = n_26941 ^ n_26524;
assign n_26950 = n_26942 & n_26944;
assign n_26951 = n_26945 ^ n_26935;
assign n_26952 = n_26946 ^ x307;
assign n_26953 = ~n_26931 & n_26947;
assign n_26954 = n_26947 ^ n_26931;
assign n_26955 = ~n_26948 & ~n_26940;
assign n_26956 = n_26948 ^ n_25768;
assign n_26957 = n_26949 ^ n_26933;
assign n_26958 = n_26950 ^ n_25126;
assign n_26959 = n_26951 ^ x306;
assign n_26960 = n_26952 ^ n_26951;
assign n_26961 = n_26955 ^ n_26524;
assign n_26962 = n_26956 ^ n_25145;
assign n_26963 = n_26957 ^ n_26902;
assign n_26964 = n_26958 ^ n_26956;
assign n_26965 = n_26958 ^ n_25145;
assign n_26966 = ~n_26960 & n_26959;
assign n_26967 = n_26960 ^ x306;
assign n_26968 = n_26961 ^ n_26577;
assign n_26969 = n_26961 ^ n_26562;
assign n_26970 = ~n_26962 & ~n_26964;
assign n_26971 = n_26965 ^ n_26956;
assign n_26972 = n_26966 ^ x306;
assign n_26973 = ~n_26953 & n_26967;
assign n_26974 = n_26967 ^ n_26953;
assign n_26975 = n_26968 ^ n_26562;
assign n_26976 = n_26968 ^ n_26932;
assign n_26977 = ~n_26577 & n_26969;
assign n_26978 = n_26970 ^ n_25145;
assign n_26979 = n_26971 ^ x305;
assign n_26980 = n_26972 ^ n_26971;
assign n_26981 = n_26975 ^ n_25805;
assign n_26982 = n_26977 ^ n_25682;
assign n_26983 = n_26978 ^ n_25164;
assign n_26984 = ~n_26980 & n_26979;
assign n_26985 = n_26980 ^ x305;
assign n_26986 = n_26981 ^ n_25164;
assign n_26987 = n_26978 ^ n_26981;
assign n_26988 = n_26982 ^ n_26617;
assign n_26989 = n_26982 ^ n_26602;
assign n_26990 = n_26983 ^ n_26981;
assign n_26991 = n_26984 ^ x305;
assign n_26992 = ~n_26973 & ~n_26985;
assign n_26993 = n_26985 ^ n_26973;
assign n_26994 = n_26986 & ~n_26987;
assign n_26995 = n_26988 ^ n_26602;
assign n_26996 = n_26954 ^ n_26988;
assign n_26997 = n_26617 & n_26989;
assign n_26998 = n_26990 ^ x304;
assign n_26999 = n_26991 ^ n_26990;
assign n_27000 = n_26994 ^ n_25164;
assign n_27001 = n_26995 ^ n_25830;
assign n_27002 = n_26997 ^ n_25742;
assign n_27003 = ~n_26999 & n_26998;
assign n_27004 = n_26999 ^ x304;
assign n_27005 = n_27000 ^ n_27001;
assign n_27006 = n_27001 ^ n_25184;
assign n_27007 = n_27002 ^ n_25803;
assign n_27008 = n_27002 ^ n_26642;
assign n_27009 = n_27003 ^ x304;
assign n_27010 = ~n_27004 & n_26992;
assign n_27011 = n_26992 ^ n_27004;
assign n_27012 = n_27005 ^ n_25184;
assign n_27013 = ~n_27005 & ~n_27006;
assign n_27014 = n_27007 ^ n_25885;
assign n_27015 = n_27007 ^ n_26642;
assign n_27016 = ~n_26657 & n_27008;
assign n_27017 = n_27009 ^ x319;
assign n_27018 = n_27012 ^ x319;
assign n_27019 = n_27012 ^ n_27009;
assign n_27020 = n_27013 ^ n_25184;
assign n_27021 = n_27014 ^ n_25218;
assign n_27022 = n_27015 ^ n_26974;
assign n_27023 = n_27016 ^ n_25803;
assign n_27024 = n_27012 ^ n_27017;
assign n_27025 = ~n_27018 & n_27019;
assign n_27026 = n_27020 ^ n_27014;
assign n_27027 = n_27023 ^ n_25852;
assign n_27028 = n_27023 ^ n_26682;
assign n_27029 = n_27024 & n_27010;
assign n_27030 = n_27010 ^ n_27024;
assign n_27031 = n_27025 ^ x319;
assign n_27032 = n_27026 ^ n_25218;
assign n_27033 = n_27026 & n_27021;
assign n_27034 = n_27027 ^ n_25925;
assign n_27035 = n_27027 ^ n_26682;
assign n_27036 = ~n_26697 & n_27028;
assign n_27037 = n_27031 ^ n_27032;
assign n_27038 = n_27032 ^ x318;
assign n_27039 = n_27033 ^ n_25218;
assign n_27040 = n_27034 ^ n_25255;
assign n_27041 = n_26993 ^ n_27035;
assign n_27042 = n_27036 ^ n_25852;
assign n_27043 = n_27037 ^ x318;
assign n_27044 = n_27037 & ~n_27038;
assign n_27045 = n_27039 ^ n_27034;
assign n_27046 = n_27042 ^ n_26722;
assign n_27047 = ~n_27029 & ~n_27043;
assign n_27048 = n_27043 ^ n_27029;
assign n_27049 = n_27044 ^ x318;
assign n_27050 = n_27045 ^ n_25255;
assign n_27051 = ~n_27045 & ~n_27040;
assign n_27052 = n_25895 ^ n_27046;
assign n_27053 = n_27046 & ~n_26737;
assign n_27054 = n_27049 ^ n_27050;
assign n_27055 = n_27050 ^ x317;
assign n_27056 = n_27051 ^ n_25255;
assign n_27057 = n_27052 ^ n_26722;
assign n_27058 = n_27011 ^ n_27052;
assign n_27059 = n_27053 ^ n_25895;
assign n_27060 = n_27054 ^ x317;
assign n_27061 = n_27054 & ~n_27055;
assign n_27062 = n_27056 ^ n_25290;
assign n_27063 = n_27057 ^ n_25962;
assign n_27064 = n_27059 ^ n_25936;
assign n_27065 = n_27059 ^ n_26761;
assign n_27066 = n_27047 & ~n_27060;
assign n_27067 = n_27060 ^ n_27047;
assign n_27068 = n_27061 ^ x317;
assign n_27069 = n_27062 ^ n_27063;
assign n_27070 = n_27063 ^ n_25290;
assign n_27071 = n_27056 ^ n_27063;
assign n_27072 = n_27064 ^ n_26001;
assign n_27073 = n_27064 ^ n_26761;
assign n_27074 = n_26775 & n_27065;
assign n_27075 = n_27068 ^ n_27069;
assign n_27076 = n_27069 ^ x316;
assign n_27077 = n_27070 & ~n_27071;
assign n_27078 = n_27072 ^ n_25329;
assign n_27079 = n_27030 ^ n_27073;
assign n_27080 = n_27074 ^ n_25936;
assign n_27081 = n_27075 ^ x316;
assign n_27082 = n_27075 & ~n_27076;
assign n_27083 = n_27077 ^ n_25290;
assign n_27084 = n_27080 ^ n_26800;
assign n_27085 = ~n_27066 & n_27081;
assign n_27086 = n_27082 ^ x316;
assign n_27087 = n_27083 ^ n_25329;
assign n_27088 = n_27083 ^ n_27072;
assign n_27089 = n_25973 ^ n_27084;
assign n_27090 = ~n_27084 & n_26814;
assign n_27091 = n_27087 ^ n_27072;
assign n_27092 = ~n_27078 & n_27088;
assign n_27093 = n_27089 ^ n_26800;
assign n_27094 = n_27048 ^ n_27089;
assign n_27095 = n_27090 ^ n_25973;
assign n_27096 = n_27086 ^ n_27091;
assign n_27097 = n_27091 ^ x315;
assign n_27098 = n_27092 ^ n_25329;
assign n_27099 = n_27093 ^ n_26041;
assign n_27100 = n_27095 ^ n_26013;
assign n_27101 = n_27095 ^ n_26838;
assign n_27102 = n_27096 ^ x315;
assign n_27103 = ~n_27096 & n_27097;
assign n_27104 = n_27098 ^ n_25368;
assign n_27105 = n_27099 ^ n_25368;
assign n_27106 = n_27098 ^ n_27099;
assign n_27107 = n_27100 ^ n_26080;
assign n_27108 = n_27100 ^ n_26838;
assign n_27109 = ~n_26852 & n_27101;
assign n_27110 = n_27085 & ~n_27102;
assign n_27111 = n_27102 ^ n_27085;
assign n_27112 = n_27103 ^ x315;
assign n_27113 = n_27104 ^ n_27099;
assign n_27114 = ~n_27105 & n_27106;
assign n_27115 = n_27107 ^ n_25407;
assign n_27116 = n_27108 ^ n_27067;
assign n_27117 = n_27109 ^ n_26013;
assign n_27118 = n_26125 & n_27111;
assign n_27119 = n_27111 ^ n_25680;
assign n_27120 = n_27111 ^ n_25663;
assign n_27121 = n_27111 ^ n_26125;
assign n_27122 = n_27112 ^ n_27113;
assign n_27123 = n_27113 ^ x314;
assign n_27124 = n_27114 ^ n_25368;
assign n_27125 = n_27117 ^ n_26903;
assign n_27126 = n_26153 ^ n_27118;
assign n_27127 = n_25168 & n_27119;
assign n_27128 = x391 & n_27120;
assign n_27129 = n_27120 ^ x391;
assign n_27130 = n_27122 ^ x314;
assign n_27131 = ~n_27122 & n_27123;
assign n_27132 = n_27124 ^ n_25407;
assign n_27133 = n_27124 ^ n_27107;
assign n_27134 = n_27125 ^ n_26877;
assign n_27135 = n_27066 ^ n_27125;
assign n_27136 = n_27127 ^ n_25197;
assign n_27137 = n_27128 ^ x390;
assign n_27138 = n_27130 ^ n_27110;
assign n_27139 = ~n_27110 & n_27130;
assign n_27140 = n_27131 ^ x314;
assign n_27141 = n_27132 ^ n_27107;
assign n_27142 = n_27115 & ~n_27133;
assign n_27143 = n_27134 ^ n_26127;
assign n_27144 = n_27135 ^ n_27081;
assign n_27145 = n_27138 ^ n_27126;
assign n_27146 = n_27138 ^ n_27118;
assign n_27147 = n_27140 ^ n_27141;
assign n_27148 = n_27141 ^ x313;
assign n_27149 = n_27142 ^ n_25407;
assign n_27150 = n_27143 ^ n_25446;
assign n_27151 = n_27145 ^ n_26152;
assign n_27152 = n_27126 & n_27146;
assign n_27153 = n_27147 ^ x313;
assign n_27154 = n_27147 & ~n_27148;
assign n_27155 = n_27149 ^ x312;
assign n_27156 = n_27151 ^ n_27127;
assign n_27157 = n_27152 ^ n_26153;
assign n_27158 = n_27153 ^ n_27139;
assign n_27159 = ~n_27139 & n_27153;
assign n_27160 = n_27154 ^ x313;
assign n_27161 = n_27155 ^ n_27150;
assign n_27162 = n_27156 ^ n_25197;
assign n_27163 = ~n_27156 & ~n_27136;
assign n_27164 = n_27157 ^ n_26208;
assign n_27165 = n_26208 ^ n_27158;
assign n_27166 = n_27157 ^ n_27158;
assign n_27167 = n_27160 ^ n_27159;
assign n_27168 = n_27162 ^ n_27128;
assign n_27169 = n_27163 ^ n_25197;
assign n_27170 = n_27164 ^ n_27158;
assign n_27171 = n_27165 & ~n_27166;
assign n_27172 = n_27167 ^ n_27161;
assign n_27173 = n_27168 & n_27137;
assign n_27174 = n_27168 ^ x390;
assign n_27175 = n_27169 ^ n_25237;
assign n_27176 = n_27170 ^ n_26192;
assign n_27177 = n_27171 ^ n_26208;
assign n_27178 = n_26246 ^ n_27172;
assign n_27179 = n_27173 ^ x390;
assign n_27180 = n_27129 & ~n_27174;
assign n_27181 = n_27174 ^ n_27129;
assign n_27182 = n_27175 ^ n_27176;
assign n_27183 = n_27176 ^ n_25237;
assign n_27184 = n_27169 ^ n_27176;
assign n_27185 = n_27177 ^ n_26246;
assign n_27186 = n_27177 ^ n_27172;
assign n_27187 = n_27179 ^ x389;
assign n_27188 = n_27179 ^ n_27182;
assign n_27189 = ~n_27183 & n_27184;
assign n_27190 = n_27185 ^ n_27172;
assign n_27191 = ~n_27178 & n_27186;
assign n_27192 = ~n_27188 & n_27187;
assign n_27193 = n_27188 ^ x389;
assign n_27194 = n_27189 ^ n_25237;
assign n_27195 = n_27190 ^ n_26233;
assign n_27196 = n_27191 ^ n_26246;
assign n_27197 = n_27192 ^ x389;
assign n_27198 = ~n_27180 & ~n_27193;
assign n_27199 = n_27193 ^ n_27180;
assign n_27200 = n_27194 ^ n_25271;
assign n_27201 = n_27195 ^ n_25271;
assign n_27202 = n_27194 ^ n_27195;
assign n_27203 = n_27196 ^ n_26298;
assign n_27204 = n_27196 ^ n_26124;
assign n_27205 = n_27197 ^ x388;
assign n_27206 = n_27200 ^ n_27195;
assign n_27207 = ~n_27201 & ~n_27202;
assign n_27208 = n_27203 ^ n_26269;
assign n_27209 = n_26298 & ~n_27204;
assign n_27210 = n_27197 ^ n_27206;
assign n_27211 = n_27207 ^ n_25271;
assign n_27212 = n_27209 ^ n_26285;
assign n_27213 = ~n_27210 & n_27205;
assign n_27214 = n_27210 ^ x388;
assign n_27215 = n_27211 ^ n_25309;
assign n_27216 = n_27208 ^ n_27211;
assign n_27217 = n_26324 ^ n_27212;
assign n_27218 = n_27213 ^ x388;
assign n_27219 = ~n_27198 & n_27214;
assign n_27220 = n_27214 ^ n_27198;
assign n_27221 = n_27208 ^ n_27215;
assign n_27222 = ~n_27215 & ~n_27216;
assign n_27223 = n_26212 ^ n_27217;
assign n_27224 = n_27217 & n_26337;
assign n_27225 = n_27218 ^ n_27221;
assign n_27226 = n_27221 ^ x387;
assign n_27227 = n_27222 ^ n_25309;
assign n_27228 = n_27223 ^ n_26309;
assign n_27229 = n_27224 ^ n_26212;
assign n_27230 = n_27225 ^ x387;
assign n_27231 = n_27225 & ~n_27226;
assign n_27232 = n_27227 ^ n_25348;
assign n_27233 = n_27228 ^ n_25348;
assign n_27234 = n_27227 ^ n_27228;
assign n_27235 = n_26363 ^ n_27229;
assign n_27236 = n_27219 & ~n_27230;
assign n_27237 = n_27230 ^ n_27219;
assign n_27238 = n_27231 ^ x387;
assign n_27239 = n_27232 ^ n_27228;
assign n_27240 = ~n_27233 & ~n_27234;
assign n_27241 = n_26274 ^ n_27235;
assign n_27242 = n_27235 & ~n_26376;
assign n_27243 = n_27238 ^ x386;
assign n_27244 = n_27238 ^ n_27239;
assign n_27245 = n_27240 ^ n_25348;
assign n_27246 = n_27241 ^ n_26349;
assign n_27247 = n_27242 ^ n_26274;
assign n_27248 = ~n_27244 & n_27243;
assign n_27249 = n_27244 ^ x386;
assign n_27250 = n_27245 ^ n_25387;
assign n_27251 = n_27246 ^ n_25387;
assign n_27252 = n_27245 ^ n_27246;
assign n_27253 = n_26401 ^ n_27247;
assign n_27254 = n_27248 ^ x386;
assign n_27255 = ~n_27236 & ~n_27249;
assign n_27256 = n_27249 ^ n_27236;
assign n_27257 = n_27250 ^ n_27246;
assign n_27258 = ~n_27251 & n_27252;
assign n_27259 = n_26315 ^ n_27253;
assign n_27260 = n_27253 & n_26414;
assign n_27261 = n_27254 ^ x385;
assign n_27262 = n_27254 ^ n_27257;
assign n_27263 = n_27258 ^ n_25387;
assign n_27264 = n_27259 ^ n_26387;
assign n_27265 = n_27260 ^ n_26315;
assign n_27266 = n_27262 & n_27261;
assign n_27267 = n_27262 ^ x385;
assign n_27268 = n_27263 ^ n_25426;
assign n_27269 = n_27264 ^ n_25426;
assign n_27270 = n_27263 ^ n_27264;
assign n_27271 = n_26440 ^ n_27265;
assign n_27272 = n_27266 ^ x385;
assign n_27273 = n_27255 & n_27267;
assign n_27274 = n_27267 ^ n_27255;
assign n_27275 = n_27268 ^ n_27264;
assign n_27276 = ~n_27269 & n_27270;
assign n_27277 = n_26355 ^ n_27271;
assign n_27278 = ~n_27271 & n_26453;
assign n_27279 = n_27272 ^ n_27275;
assign n_27280 = n_27275 ^ x384;
assign n_27281 = n_27276 ^ n_25426;
assign n_27282 = n_27277 ^ n_26425;
assign n_27283 = n_27278 ^ n_26355;
assign n_27284 = n_27279 ^ x384;
assign n_27285 = n_27279 & ~n_27280;
assign n_27286 = n_27281 ^ n_25462;
assign n_27287 = n_27282 ^ n_25462;
assign n_27288 = n_27281 ^ n_27282;
assign n_27289 = n_26480 ^ n_27283;
assign n_27290 = n_27284 & n_27273;
assign n_27291 = n_27273 ^ n_27284;
assign n_27292 = n_27285 ^ x384;
assign n_27293 = n_27286 ^ n_27282;
assign n_27294 = n_27287 & n_27288;
assign n_27295 = n_26393 ^ n_27289;
assign n_27296 = n_27289 & ~n_26493;
assign n_27297 = n_27292 ^ n_27293;
assign n_27298 = n_27293 ^ x399;
assign n_27299 = n_27294 ^ n_25462;
assign n_27300 = n_27295 ^ n_26464;
assign n_27301 = n_27296 ^ n_26393;
assign n_27302 = n_27297 ^ x399;
assign n_27303 = ~n_27297 & n_27298;
assign n_27304 = n_27299 ^ n_25490;
assign n_27305 = n_27300 ^ n_25490;
assign n_27306 = n_27299 ^ n_27300;
assign n_27307 = n_26519 ^ n_27301;
assign n_27308 = n_27290 & ~n_27302;
assign n_27309 = n_27302 ^ n_27290;
assign n_27310 = n_27303 ^ x399;
assign n_27311 = n_27304 ^ n_27300;
assign n_27312 = ~n_27305 & n_27306;
assign n_27313 = ~n_27307 & ~n_26532;
assign n_27314 = n_26431 ^ n_27307;
assign n_27315 = n_27310 ^ n_27311;
assign n_27316 = n_27311 ^ x398;
assign n_27317 = n_27312 ^ n_25490;
assign n_27318 = n_27313 ^ n_26431;
assign n_27319 = n_27314 ^ n_26504;
assign n_27320 = n_27315 ^ x398;
assign n_27321 = ~n_27315 & n_27316;
assign n_27322 = n_27317 ^ n_25513;
assign n_27323 = n_26558 ^ n_27318;
assign n_27324 = n_27319 ^ n_25513;
assign n_27325 = n_27317 ^ n_27319;
assign n_27326 = n_27320 ^ n_27308;
assign n_27327 = ~n_27308 & n_27320;
assign n_27328 = n_27321 ^ x398;
assign n_27329 = n_27322 ^ n_27319;
assign n_27330 = n_27323 & ~n_26571;
assign n_27331 = n_26470 ^ n_27323;
assign n_27332 = ~n_27324 & n_27325;
assign n_27333 = n_27328 ^ n_27329;
assign n_27334 = n_27329 ^ x397;
assign n_27335 = n_27330 ^ n_26470;
assign n_27336 = n_27129 ^ n_27331;
assign n_27337 = n_27331 ^ n_26543;
assign n_27338 = n_27332 ^ n_25513;
assign n_27339 = n_27333 ^ x397;
assign n_27340 = ~n_27333 & n_27334;
assign n_27341 = n_26598 ^ n_27335;
assign n_27342 = n_27337 ^ n_25529;
assign n_27343 = n_27338 ^ n_27337;
assign n_27344 = n_27338 ^ n_25529;
assign n_27345 = n_27327 & n_27339;
assign n_27346 = n_27339 ^ n_27327;
assign n_27347 = n_27340 ^ x397;
assign n_27348 = n_27341 & n_26611;
assign n_27349 = n_26510 ^ n_27341;
assign n_27350 = ~n_27342 & n_27343;
assign n_27351 = n_27344 ^ n_27337;
assign n_27352 = n_27348 ^ n_26510;
assign n_27353 = n_27349 ^ n_26583;
assign n_27354 = n_27181 ^ n_27349;
assign n_27355 = n_27350 ^ n_25529;
assign n_27356 = n_27347 ^ n_27351;
assign n_27357 = n_27351 ^ x396;
assign n_27358 = n_27352 ^ n_26638;
assign n_27359 = n_27352 ^ n_26549;
assign n_27360 = n_27353 ^ n_25542;
assign n_27361 = n_27355 ^ n_27353;
assign n_27362 = n_27355 ^ n_25542;
assign n_27363 = n_27356 ^ x396;
assign n_27364 = ~n_27356 & n_27357;
assign n_27365 = ~n_26651 & n_27358;
assign n_27366 = n_27359 ^ n_26638;
assign n_27367 = n_27360 & n_27361;
assign n_27368 = n_27362 ^ n_27353;
assign n_27369 = ~n_27345 & ~n_27363;
assign n_27370 = n_27363 ^ n_27345;
assign n_27371 = n_27364 ^ x396;
assign n_27372 = n_27365 ^ n_26549;
assign n_27373 = n_27199 ^ n_27366;
assign n_27374 = n_27366 ^ n_26623;
assign n_27375 = n_27367 ^ n_25542;
assign n_27376 = n_27368 ^ x395;
assign n_27377 = n_27371 ^ n_27368;
assign n_27378 = n_26678 ^ n_27372;
assign n_27379 = n_27374 ^ n_25557;
assign n_27380 = n_27375 ^ n_27374;
assign n_27381 = n_27375 ^ n_25557;
assign n_27382 = n_27377 & ~n_27376;
assign n_27383 = n_27377 ^ x395;
assign n_27384 = n_27378 & ~n_26691;
assign n_27385 = n_26589 ^ n_27378;
assign n_27386 = n_27379 & ~n_27380;
assign n_27387 = n_27381 ^ n_27374;
assign n_27388 = n_27382 ^ x395;
assign n_27389 = n_27383 & n_27369;
assign n_27390 = n_27369 ^ n_27383;
assign n_27391 = n_27384 ^ n_26589;
assign n_27392 = n_27220 ^ n_27385;
assign n_27393 = n_27385 ^ n_26664;
assign n_27394 = n_27386 ^ n_25557;
assign n_27395 = n_27387 ^ x394;
assign n_27396 = n_27388 ^ n_27387;
assign n_27397 = n_27391 ^ n_26718;
assign n_27398 = n_27391 ^ n_26629;
assign n_27399 = n_27393 ^ n_25573;
assign n_27400 = n_27394 ^ n_27393;
assign n_27401 = n_27394 ^ n_25573;
assign n_27402 = ~n_27396 & n_27395;
assign n_27403 = n_27396 ^ x394;
assign n_27404 = ~n_26731 & n_27397;
assign n_27405 = n_27398 ^ n_26718;
assign n_27406 = n_27399 & ~n_27400;
assign n_27407 = n_27401 ^ n_27393;
assign n_27408 = n_27402 ^ x394;
assign n_27409 = ~n_27389 & n_27403;
assign n_27410 = n_27403 ^ n_27389;
assign n_27411 = n_27404 ^ n_26629;
assign n_27412 = n_27237 ^ n_27405;
assign n_27413 = n_27405 ^ n_26703;
assign n_27414 = n_27406 ^ n_25573;
assign n_27415 = n_27407 ^ x393;
assign n_27416 = n_27408 ^ n_27407;
assign n_27417 = n_26755 ^ n_27411;
assign n_27418 = n_27413 ^ n_25592;
assign n_27419 = n_27414 ^ n_27413;
assign n_27420 = n_27414 ^ n_25592;
assign n_27421 = ~n_27416 & n_27415;
assign n_27422 = n_27416 ^ x393;
assign n_27423 = ~n_27417 & n_26768;
assign n_27424 = n_26670 ^ n_27417;
assign n_27425 = ~n_27418 & n_27419;
assign n_27426 = n_27420 ^ n_27413;
assign n_27427 = n_27421 ^ x393;
assign n_27428 = n_27409 & n_27422;
assign n_27429 = n_27422 ^ n_27409;
assign n_27430 = n_27423 ^ n_26670;
assign n_27431 = n_27256 ^ n_27424;
assign n_27432 = n_27424 ^ n_26743;
assign n_27433 = n_27425 ^ n_25592;
assign n_27434 = n_27426 ^ x392;
assign n_27435 = n_27427 ^ n_27426;
assign n_27436 = n_27430 ^ n_26795;
assign n_27437 = n_27430 ^ n_26709;
assign n_27438 = n_27432 ^ n_25606;
assign n_27439 = n_27433 ^ n_27432;
assign n_27440 = n_27435 & ~n_27434;
assign n_27441 = n_27435 ^ x392;
assign n_27442 = n_26809 & n_27436;
assign n_27443 = n_27437 ^ n_26795;
assign n_27444 = ~n_27439 & n_27438;
assign n_27445 = n_27439 ^ n_25606;
assign n_27446 = n_27440 ^ x392;
assign n_27447 = n_27441 & ~n_27428;
assign n_27448 = n_27428 ^ n_27441;
assign n_27449 = n_27442 ^ n_26709;
assign n_27450 = n_27443 ^ n_26781;
assign n_27451 = n_27274 ^ n_27443;
assign n_27452 = n_27444 ^ n_25606;
assign n_27453 = n_27445 ^ x407;
assign n_27454 = n_27446 ^ n_27445;
assign n_27455 = n_27446 ^ x407;
assign n_27456 = n_27449 ^ n_26834;
assign n_27457 = n_27450 ^ n_25633;
assign n_27458 = n_27452 ^ n_27450;
assign n_27459 = n_27453 & ~n_27454;
assign n_27460 = n_27455 ^ n_27445;
assign n_27461 = n_27456 & n_26847;
assign n_27462 = n_26748 ^ n_27456;
assign n_27463 = n_27458 & n_27457;
assign n_27464 = n_27458 ^ n_25633;
assign n_27465 = n_27459 ^ x407;
assign n_27466 = ~n_27460 & n_27447;
assign n_27467 = n_27447 ^ n_27460;
assign n_27468 = n_27461 ^ n_26748;
assign n_27469 = n_27291 ^ n_27462;
assign n_27470 = n_27462 ^ n_26820;
assign n_27471 = n_27463 ^ n_25633;
assign n_27472 = n_27464 ^ x406;
assign n_27473 = n_27465 ^ n_27464;
assign n_27474 = n_26873 ^ n_27468;
assign n_27475 = n_27470 ^ n_25652;
assign n_27476 = n_27471 ^ n_27470;
assign n_27477 = ~n_27473 & n_27472;
assign n_27478 = n_27473 ^ x406;
assign n_27479 = n_27474 & n_26885;
assign n_27480 = n_26786 ^ n_27474;
assign n_27481 = ~n_27476 & ~n_27475;
assign n_27482 = n_27476 ^ n_25652;
assign n_27483 = n_27477 ^ x406;
assign n_27484 = n_27466 & ~n_27478;
assign n_27485 = n_27478 ^ n_27466;
assign n_27486 = n_27479 ^ n_26786;
assign n_27487 = n_27309 ^ n_27480;
assign n_27488 = n_27480 ^ n_26858;
assign n_27489 = n_27481 ^ n_25652;
assign n_27490 = n_27482 ^ x405;
assign n_27491 = n_27483 ^ n_27482;
assign n_27492 = n_26909 ^ n_27486;
assign n_27493 = n_27488 ^ n_25673;
assign n_27494 = n_27489 ^ n_27488;
assign n_27495 = n_27489 ^ n_25673;
assign n_27496 = ~n_27491 & n_27490;
assign n_27497 = n_27491 ^ x405;
assign n_27498 = n_26825 ^ n_27492;
assign n_27499 = ~n_27492 & n_26919;
assign n_27500 = ~n_27493 & ~n_27494;
assign n_27501 = n_27495 ^ n_27488;
assign n_27502 = n_27496 ^ x405;
assign n_27503 = ~n_27484 & n_27497;
assign n_27504 = n_27497 ^ n_27484;
assign n_27505 = n_27326 ^ n_27498;
assign n_27506 = n_27498 ^ n_26896;
assign n_27507 = n_27499 ^ n_26825;
assign n_27508 = n_27500 ^ n_25673;
assign n_27509 = n_27501 ^ x404;
assign n_27510 = n_27502 ^ n_27501;
assign n_27511 = n_27502 ^ x404;
assign n_27512 = n_27506 ^ n_25701;
assign n_27513 = n_26936 ^ n_27507;
assign n_27514 = n_27508 ^ n_27506;
assign n_27515 = n_27508 ^ n_25701;
assign n_27516 = ~n_27509 & n_27510;
assign n_27517 = n_27511 ^ n_27501;
assign n_27518 = n_27513 & n_26943;
assign n_27519 = n_26864 ^ n_27513;
assign n_27520 = n_27512 & n_27514;
assign n_27521 = n_27515 ^ n_27506;
assign n_27522 = n_27516 ^ x404;
assign n_27523 = ~n_27503 & n_27517;
assign n_27524 = n_27517 ^ n_27503;
assign n_27525 = n_27518 ^ n_26864;
assign n_27526 = n_27519 ^ n_26926;
assign n_27527 = n_27346 ^ n_27519;
assign n_27528 = n_27520 ^ n_25701;
assign n_27529 = n_27521 ^ x403;
assign n_27530 = n_27522 ^ n_27521;
assign n_27531 = n_27525 ^ n_26957;
assign n_27532 = n_27525 ^ n_26963;
assign n_27533 = n_27526 ^ n_25730;
assign n_27534 = n_27528 ^ n_27526;
assign n_27535 = n_27522 ^ n_27529;
assign n_27536 = ~n_27529 & n_27530;
assign n_27537 = ~n_26963 & ~n_27531;
assign n_27538 = n_27532 ^ n_26948;
assign n_27539 = n_27370 ^ n_27532;
assign n_27540 = ~n_27534 & n_27533;
assign n_27541 = n_27534 ^ n_25730;
assign n_27542 = n_27523 & n_27535;
assign n_27543 = n_27535 ^ n_27523;
assign n_27544 = n_27536 ^ x403;
assign n_27545 = n_27537 ^ n_26902;
assign n_27546 = n_27538 ^ n_25768;
assign n_27547 = n_27540 ^ n_25730;
assign n_27548 = n_27541 ^ x402;
assign n_27549 = n_27544 ^ n_27541;
assign n_27550 = n_27545 ^ n_26968;
assign n_27551 = n_27545 ^ n_26976;
assign n_27552 = n_27547 ^ n_27538;
assign n_27553 = n_27547 ^ n_27546;
assign n_27554 = n_27544 ^ n_27548;
assign n_27555 = n_27548 & ~n_27549;
assign n_27556 = ~n_26976 & ~n_27550;
assign n_27557 = n_27551 ^ n_26975;
assign n_27558 = n_27390 ^ n_27551;
assign n_27559 = n_27546 & n_27552;
assign n_27560 = n_27553 ^ x401;
assign n_27561 = ~n_27542 & n_27554;
assign n_27562 = n_27554 ^ n_27542;
assign n_27563 = n_27555 ^ x402;
assign n_27564 = n_27556 ^ n_26932;
assign n_27565 = n_27557 ^ n_25805;
assign n_27566 = n_27559 ^ n_25768;
assign n_27567 = n_27121 & ~n_27562;
assign n_27568 = n_27562 ^ n_26125;
assign n_27569 = n_27562 ^ n_26092;
assign n_27570 = n_27563 ^ n_27553;
assign n_27571 = n_27564 ^ n_26988;
assign n_27572 = n_26954 ^ n_27564;
assign n_27573 = n_27566 ^ n_27557;
assign n_27574 = n_27566 ^ n_25805;
assign n_27575 = n_27567 ^ n_27145;
assign n_27576 = n_25680 & ~n_27568;
assign n_27577 = n_27568 ^ n_27111;
assign n_27578 = x487 & ~n_27569;
assign n_27579 = n_27569 ^ x487;
assign n_27580 = ~n_27570 & n_27560;
assign n_27581 = n_27570 ^ x401;
assign n_27582 = n_26996 & ~n_27571;
assign n_27583 = n_27572 ^ n_26988;
assign n_27584 = n_27565 & n_27573;
assign n_27585 = n_27574 ^ n_27557;
assign n_27586 = n_27576 ^ n_25699;
assign n_27587 = n_27578 ^ x486;
assign n_27588 = n_27580 ^ x401;
assign n_27589 = ~n_27561 & ~n_27581;
assign n_27590 = n_27581 ^ n_27561;
assign n_27591 = n_27582 ^ n_26954;
assign n_27592 = n_27583 ^ n_26995;
assign n_27593 = n_27410 ^ n_27583;
assign n_27594 = n_27584 ^ n_25805;
assign n_27595 = n_27585 ^ x400;
assign n_27596 = n_27588 ^ n_27585;
assign n_27597 = n_27590 ^ n_27567;
assign n_27598 = n_27590 ^ n_27575;
assign n_27599 = n_26974 ^ n_27591;
assign n_27600 = n_27015 ^ n_27591;
assign n_27601 = n_27592 ^ n_25830;
assign n_27602 = n_27594 ^ n_27592;
assign n_27603 = n_27596 & ~n_27595;
assign n_27604 = n_27596 ^ x400;
assign n_27605 = ~n_27575 & n_27597;
assign n_27606 = n_27597 ^ n_26153;
assign n_27607 = n_27015 ^ n_27599;
assign n_27608 = ~n_27022 & ~n_27600;
assign n_27609 = n_27602 & n_27601;
assign n_27610 = n_27602 ^ n_25830;
assign n_27611 = n_27603 ^ x400;
assign n_27612 = n_27604 & n_27589;
assign n_27613 = n_27589 ^ n_27604;
assign n_27614 = n_27605 ^ n_27145;
assign n_27615 = n_27606 ^ n_27576;
assign n_27616 = n_27606 ^ n_27586;
assign n_27617 = n_27607 ^ n_27007;
assign n_27618 = n_27429 ^ n_27607;
assign n_27619 = n_27608 ^ n_26974;
assign n_27620 = n_27609 ^ n_25830;
assign n_27621 = n_27610 ^ x415;
assign n_27622 = n_27611 ^ n_27610;
assign n_27623 = n_27613 ^ n_27170;
assign n_27624 = n_27614 ^ n_27613;
assign n_27625 = ~n_27586 & n_27615;
assign n_27626 = n_27616 ^ n_27578;
assign n_27627 = n_27616 ^ n_27587;
assign n_27628 = n_27617 ^ n_25885;
assign n_27629 = n_27619 ^ n_26993;
assign n_27630 = n_27619 ^ n_27035;
assign n_27631 = n_27617 ^ n_27620;
assign n_27632 = n_27611 ^ n_27621;
assign n_27633 = n_27621 & ~n_27622;
assign n_27634 = n_27614 ^ n_27623;
assign n_27635 = ~n_27623 & ~n_27624;
assign n_27636 = n_27624 ^ n_26208;
assign n_27637 = n_27625 ^ n_25699;
assign n_27638 = n_27587 & ~n_27626;
assign n_27639 = n_27628 ^ n_27620;
assign n_27640 = n_27629 ^ n_27035;
assign n_27641 = ~n_27041 & n_27630;
assign n_27642 = ~n_27628 & ~n_27631;
assign n_27643 = n_27632 & ~n_27612;
assign n_27644 = n_27612 ^ n_27632;
assign n_27645 = n_27633 ^ x415;
assign n_27646 = n_27635 ^ n_27170;
assign n_27647 = n_27636 ^ n_25737;
assign n_27648 = n_27637 ^ n_27636;
assign n_27649 = n_27638 ^ x486;
assign n_27650 = n_27639 ^ x414;
assign n_27651 = n_27640 ^ n_27027;
assign n_27652 = n_27448 ^ n_27640;
assign n_27653 = n_27641 ^ n_26993;
assign n_27654 = n_27642 ^ n_25885;
assign n_27655 = n_27645 ^ x414;
assign n_27656 = n_27639 ^ n_27645;
assign n_27657 = n_27646 ^ n_27190;
assign n_27658 = n_27644 ^ n_27646;
assign n_27659 = n_27637 ^ n_27647;
assign n_27660 = n_27647 & n_27648;
assign n_27661 = n_27649 ^ x485;
assign n_27662 = n_27651 ^ n_25925;
assign n_27663 = n_27653 ^ n_27058;
assign n_27664 = n_27653 ^ n_27052;
assign n_27665 = n_27651 ^ n_27654;
assign n_27666 = n_27639 ^ n_27655;
assign n_27667 = n_27650 & ~n_27656;
assign n_27668 = n_27644 ^ n_27657;
assign n_27669 = ~n_27657 & n_27658;
assign n_27670 = n_27658 ^ n_26246;
assign n_27671 = n_27659 ^ x485;
assign n_27672 = n_27649 ^ n_27659;
assign n_27673 = n_27660 ^ n_25737;
assign n_27674 = n_27661 ^ n_27659;
assign n_27675 = n_27662 ^ n_27654;
assign n_27676 = n_27663 ^ n_27057;
assign n_27677 = n_27467 ^ n_27663;
assign n_27678 = n_27058 & n_27664;
assign n_27679 = n_27662 & ~n_27665;
assign n_27680 = ~n_27666 & ~n_27643;
assign n_27681 = n_27643 ^ n_27666;
assign n_27682 = n_27667 ^ x414;
assign n_27683 = n_27669 ^ n_27190;
assign n_27684 = n_27670 ^ n_25775;
assign n_27685 = ~n_27671 & n_27672;
assign n_27686 = n_27673 ^ n_27670;
assign n_27687 = n_27675 ^ x413;
assign n_27688 = n_27676 ^ n_25962;
assign n_27689 = n_27678 ^ n_27011;
assign n_27690 = n_27679 ^ n_25925;
assign n_27691 = n_27681 ^ n_27203;
assign n_27692 = n_27682 ^ n_27675;
assign n_27693 = n_27681 ^ n_27683;
assign n_27694 = n_27683 ^ n_27203;
assign n_27695 = n_27673 ^ n_27684;
assign n_27696 = n_27685 ^ x485;
assign n_27697 = ~n_27684 & n_27686;
assign n_27698 = n_27689 ^ n_27079;
assign n_27699 = n_27689 ^ n_27073;
assign n_27700 = n_27690 ^ n_25962;
assign n_27701 = n_27690 ^ n_27676;
assign n_27702 = n_27692 ^ x413;
assign n_27703 = ~n_27692 & n_27687;
assign n_27704 = ~n_27693 & ~n_27691;
assign n_27705 = n_27693 ^ n_26285;
assign n_27706 = n_27694 ^ n_27681;
assign n_27707 = n_27695 ^ x484;
assign n_27708 = n_27696 ^ n_27695;
assign n_27709 = n_27697 ^ n_25775;
assign n_27710 = n_27698 ^ n_27064;
assign n_27711 = n_27485 ^ n_27698;
assign n_27712 = n_27079 & n_27699;
assign n_27713 = n_27700 ^ n_27676;
assign n_27714 = n_27688 & n_27701;
assign n_27715 = n_27680 & ~n_27702;
assign n_27716 = n_27702 ^ n_27680;
assign n_27717 = n_27703 ^ x413;
assign n_27718 = n_27704 ^ n_27203;
assign n_27719 = n_27705 ^ n_25814;
assign n_27720 = n_27708 & ~n_27707;
assign n_27721 = n_27708 ^ x484;
assign n_27722 = n_27709 ^ n_25814;
assign n_27723 = n_27709 ^ n_27705;
assign n_27724 = n_27710 ^ n_26001;
assign n_27725 = n_27712 ^ n_27030;
assign n_27726 = n_27713 ^ x412;
assign n_27727 = n_27714 ^ n_25962;
assign n_27728 = n_27716 ^ n_27223;
assign n_27729 = n_27713 ^ n_27717;
assign n_27730 = n_27718 ^ n_27716;
assign n_27731 = n_27718 ^ n_27223;
assign n_27732 = n_27720 ^ x484;
assign n_27733 = n_27722 ^ n_27705;
assign n_27734 = n_27719 & ~n_27723;
assign n_27735 = n_27725 ^ n_27089;
assign n_27736 = n_27726 ^ n_27717;
assign n_27737 = n_27727 ^ n_27724;
assign n_27738 = n_27727 ^ n_27710;
assign n_27739 = n_27726 & ~n_27729;
assign n_27740 = ~n_27730 & n_27728;
assign n_27741 = n_27730 ^ n_26324;
assign n_27742 = n_27731 ^ n_27716;
assign n_27743 = n_27732 ^ x483;
assign n_27744 = n_27733 ^ x483;
assign n_27745 = n_27732 ^ n_27733;
assign n_27746 = n_27734 ^ n_25814;
assign n_27747 = n_27048 ^ n_27735;
assign n_27748 = n_27735 & n_27094;
assign n_27749 = ~n_27715 & n_27736;
assign n_27750 = n_27736 ^ n_27715;
assign n_27751 = n_27737 ^ x411;
assign n_27752 = n_27724 & ~n_27738;
assign n_27753 = n_27739 ^ x412;
assign n_27754 = n_27740 ^ n_27223;
assign n_27755 = n_27741 ^ n_25855;
assign n_27756 = n_27743 ^ n_27733;
assign n_27757 = n_27744 & ~n_27745;
assign n_27758 = n_27746 ^ n_25855;
assign n_27759 = n_27746 ^ n_27741;
assign n_27760 = n_27747 ^ n_27093;
assign n_27761 = n_27504 ^ n_27747;
assign n_27762 = n_27748 ^ n_27048;
assign n_27763 = n_27750 ^ n_27241;
assign n_27764 = n_27752 ^ n_26001;
assign n_27765 = n_27753 ^ n_27737;
assign n_27766 = n_27754 ^ n_27750;
assign n_27767 = ~n_27756 & n_27721;
assign n_27768 = n_27721 ^ n_27756;
assign n_27769 = n_27757 ^ x483;
assign n_27770 = n_27758 ^ n_27741;
assign n_27771 = ~n_27755 & n_27759;
assign n_27772 = n_27760 ^ n_26041;
assign n_27773 = n_27116 ^ n_27762;
assign n_27774 = n_27108 ^ n_27762;
assign n_27775 = n_27763 ^ n_27754;
assign n_27776 = n_27764 ^ n_26041;
assign n_27777 = n_27764 ^ n_27760;
assign n_27778 = n_27765 ^ x411;
assign n_27779 = n_27765 & ~n_27751;
assign n_27780 = n_27766 & ~n_27763;
assign n_27781 = n_27766 ^ n_26363;
assign n_27782 = n_27770 ^ x482;
assign n_27783 = n_27769 ^ n_27770;
assign n_27784 = n_27771 ^ n_25855;
assign n_27785 = n_27773 ^ n_27100;
assign n_27786 = n_27524 ^ n_27773;
assign n_27787 = n_27116 & n_27774;
assign n_27788 = n_27776 ^ n_27760;
assign n_27789 = ~n_27772 & ~n_27777;
assign n_27790 = n_27749 & ~n_27778;
assign n_27791 = n_27778 ^ n_27749;
assign n_27792 = n_27779 ^ x411;
assign n_27793 = n_27780 ^ n_27241;
assign n_27794 = n_27781 ^ n_25891;
assign n_27795 = n_27769 ^ n_27782;
assign n_27796 = ~n_27782 & n_27783;
assign n_27797 = n_27784 ^ n_27781;
assign n_27798 = n_27785 ^ n_26080;
assign n_27799 = n_27787 ^ n_27067;
assign n_27800 = n_27788 ^ x410;
assign n_27801 = n_27789 ^ n_26041;
assign n_27802 = n_27791 ^ n_27259;
assign n_27803 = n_27792 ^ x410;
assign n_27804 = n_27792 ^ n_27788;
assign n_27805 = n_27793 ^ n_27791;
assign n_27806 = n_27793 ^ n_27259;
assign n_27807 = n_27784 ^ n_27794;
assign n_27808 = n_27795 ^ n_27767;
assign n_27809 = n_27767 & n_27795;
assign n_27810 = n_27796 ^ x482;
assign n_27811 = n_27794 & n_27797;
assign n_27812 = n_27799 ^ n_27144;
assign n_27813 = n_27801 ^ n_26080;
assign n_27814 = n_27801 ^ n_27785;
assign n_27815 = n_27803 ^ n_27788;
assign n_27816 = n_27800 & ~n_27804;
assign n_27817 = n_27802 & n_27805;
assign n_27818 = n_27805 ^ n_26401;
assign n_27819 = n_27806 ^ n_27791;
assign n_27820 = n_27807 ^ x481;
assign n_27821 = n_27810 ^ n_27807;
assign n_27822 = n_27811 ^ n_25891;
assign n_27823 = n_27812 ^ n_27143;
assign n_27824 = n_27543 ^ n_27812;
assign n_27825 = n_27813 ^ n_27785;
assign n_27826 = ~n_27798 & ~n_27814;
assign n_27827 = ~n_27790 & ~n_27815;
assign n_27828 = n_27815 ^ n_27790;
assign n_27829 = n_27816 ^ x410;
assign n_27830 = n_27817 ^ n_27259;
assign n_27831 = n_27818 ^ n_25931;
assign n_27832 = ~n_27821 & n_27820;
assign n_27833 = n_27821 ^ x481;
assign n_27834 = n_27822 ^ n_27818;
assign n_27835 = n_27823 ^ x408;
assign n_27836 = n_27824 ^ n_27524;
assign n_27837 = n_27825 ^ x409;
assign n_27838 = n_27826 ^ n_26080;
assign n_27839 = n_27828 ^ n_27277;
assign n_27840 = n_27829 ^ x409;
assign n_27841 = n_27829 ^ n_27825;
assign n_27842 = n_27828 ^ n_27830;
assign n_27843 = n_27832 ^ x481;
assign n_27844 = ~n_27833 & n_27809;
assign n_27845 = n_27809 ^ n_27833;
assign n_27846 = ~n_27834 & ~n_27831;
assign n_27847 = n_27834 ^ n_25931;
assign n_27848 = n_27838 ^ n_27835;
assign n_27849 = n_27839 ^ n_27830;
assign n_27850 = n_27840 ^ n_27825;
assign n_27851 = ~n_27837 & n_27841;
assign n_27852 = ~n_27842 & ~n_27839;
assign n_27853 = n_27842 ^ n_26440;
assign n_27854 = n_27846 ^ n_25931;
assign n_27855 = n_27847 ^ x480;
assign n_27856 = n_27843 ^ n_27847;
assign n_27857 = n_27827 ^ n_27850;
assign n_27858 = n_27850 & n_27827;
assign n_27859 = n_27851 ^ x409;
assign n_27860 = n_27852 ^ n_27277;
assign n_27861 = n_27853 ^ n_25968;
assign n_27862 = n_27854 ^ n_27853;
assign n_27863 = n_27843 ^ n_27855;
assign n_27864 = n_27855 & ~n_27856;
assign n_27865 = n_27857 ^ n_27295;
assign n_27866 = n_27859 ^ n_27848;
assign n_27867 = n_27857 ^ n_27860;
assign n_27868 = ~n_27862 & ~n_27861;
assign n_27869 = n_27862 ^ n_25968;
assign n_27870 = n_27844 & ~n_27863;
assign n_27871 = n_27863 ^ n_27844;
assign n_27872 = n_27864 ^ x480;
assign n_27873 = n_27865 ^ n_27860;
assign n_27874 = n_27866 ^ n_27858;
assign n_27875 = n_27867 & n_27865;
assign n_27876 = n_27867 ^ n_26480;
assign n_27877 = n_27868 ^ n_25968;
assign n_27878 = n_27869 ^ x495;
assign n_27879 = n_27872 ^ n_27869;
assign n_27880 = n_27874 ^ n_27314;
assign n_27881 = n_27875 ^ n_27295;
assign n_27882 = n_27876 ^ n_26008;
assign n_27883 = n_27876 ^ n_27877;
assign n_27884 = n_27877 ^ n_26008;
assign n_27885 = n_27872 ^ n_27878;
assign n_27886 = ~n_27878 & n_27879;
assign n_27887 = n_27881 ^ n_27874;
assign n_27888 = n_27882 & n_27883;
assign n_27889 = n_27876 ^ n_27884;
assign n_27890 = ~n_27885 & ~n_27870;
assign n_27891 = n_27870 ^ n_27885;
assign n_27892 = n_27886 ^ x495;
assign n_27893 = n_27887 & ~n_27880;
assign n_27894 = n_27887 ^ n_26519;
assign n_27895 = n_27887 ^ n_27314;
assign n_27896 = n_27888 ^ n_26008;
assign n_27897 = n_27889 ^ x494;
assign n_27898 = n_27889 ^ n_27892;
assign n_27899 = n_27893 ^ n_27314;
assign n_27900 = n_27894 ^ n_26048;
assign n_27901 = n_27894 ^ n_27896;
assign n_27902 = n_27896 ^ n_26048;
assign n_27903 = n_27897 ^ n_27892;
assign n_27904 = ~n_27897 & n_27898;
assign n_27905 = n_27899 ^ n_27331;
assign n_27906 = n_27899 ^ n_27129;
assign n_27907 = n_27900 & n_27901;
assign n_27908 = n_27894 ^ n_27902;
assign n_27909 = ~n_27903 & n_27890;
assign n_27910 = n_27890 ^ n_27903;
assign n_27911 = n_27904 ^ x494;
assign n_27912 = ~n_27336 & n_27905;
assign n_27913 = n_27906 ^ n_26558;
assign n_27914 = n_27906 ^ n_27331;
assign n_27915 = n_27907 ^ n_26048;
assign n_27916 = n_27908 ^ x493;
assign n_27917 = n_27908 ^ n_27911;
assign n_27918 = n_27912 ^ n_27129;
assign n_27919 = n_27913 ^ n_26087;
assign n_27920 = n_27913 ^ n_27915;
assign n_27921 = n_27915 ^ n_26087;
assign n_27922 = n_27916 ^ n_27911;
assign n_27923 = n_27916 & ~n_27917;
assign n_27924 = n_27918 ^ n_27349;
assign n_27925 = n_27919 & n_27920;
assign n_27926 = n_27913 ^ n_27921;
assign n_27927 = ~n_27909 & ~n_27922;
assign n_27928 = n_27922 ^ n_27909;
assign n_27929 = n_27923 ^ x493;
assign n_27930 = ~n_27924 & n_27354;
assign n_27931 = n_27924 ^ n_27181;
assign n_27932 = n_27925 ^ n_26087;
assign n_27933 = n_27926 ^ x492;
assign n_27934 = n_27929 ^ n_27926;
assign n_27935 = n_27930 ^ n_27181;
assign n_27936 = n_27931 ^ n_27349;
assign n_27937 = n_27932 ^ n_26133;
assign n_27938 = n_27934 & ~n_27933;
assign n_27939 = n_27934 ^ x492;
assign n_27940 = n_27935 ^ n_27366;
assign n_27941 = n_27373 ^ n_27935;
assign n_27942 = n_27936 ^ n_26598;
assign n_27943 = n_27938 ^ x492;
assign n_27944 = n_27927 & n_27939;
assign n_27945 = n_27939 ^ n_27927;
assign n_27946 = n_27373 & ~n_27940;
assign n_27947 = n_27941 ^ n_27366;
assign n_27948 = n_27942 ^ n_26133;
assign n_27949 = n_27942 ^ n_27932;
assign n_27950 = n_27942 ^ n_27937;
assign n_27951 = n_27943 ^ x491;
assign n_27952 = n_27946 ^ n_27199;
assign n_27953 = n_27947 ^ n_26638;
assign n_27954 = ~n_27948 & ~n_27949;
assign n_27955 = n_27950 ^ x491;
assign n_27956 = n_27950 ^ n_27943;
assign n_27957 = n_27950 ^ n_27951;
assign n_27958 = n_27952 ^ n_27385;
assign n_27959 = n_27392 ^ n_27952;
assign n_27960 = n_27953 ^ n_26173;
assign n_27961 = n_27954 ^ n_26133;
assign n_27962 = ~n_27955 & n_27956;
assign n_27963 = n_27944 & n_27957;
assign n_27964 = n_27957 ^ n_27944;
assign n_27965 = n_27392 & ~n_27958;
assign n_27966 = n_27959 ^ n_27385;
assign n_27967 = n_27953 ^ n_27961;
assign n_27968 = n_27961 ^ n_26173;
assign n_27969 = n_27962 ^ x491;
assign n_27970 = n_27965 ^ n_27220;
assign n_27971 = n_27966 ^ n_26678;
assign n_27972 = ~n_27960 & ~n_27967;
assign n_27973 = n_27953 ^ n_27968;
assign n_27974 = n_27969 ^ x490;
assign n_27975 = n_27970 ^ n_27405;
assign n_27976 = n_27237 ^ n_27970;
assign n_27977 = n_27971 ^ n_26215;
assign n_27978 = n_27972 ^ n_26173;
assign n_27979 = n_27973 ^ x490;
assign n_27980 = n_27973 ^ n_27969;
assign n_27981 = n_27973 ^ n_27974;
assign n_27982 = n_27412 & ~n_27975;
assign n_27983 = n_27976 ^ n_26718;
assign n_27984 = n_27976 ^ n_27405;
assign n_27985 = n_27971 ^ n_27978;
assign n_27986 = n_27977 ^ n_27978;
assign n_27987 = n_27979 & ~n_27980;
assign n_27988 = n_27963 & ~n_27981;
assign n_27989 = n_27981 ^ n_27963;
assign n_27990 = n_27982 ^ n_27237;
assign n_27991 = n_27983 ^ n_26251;
assign n_27992 = ~n_27977 & n_27985;
assign n_27993 = n_27986 ^ x489;
assign n_27994 = n_27987 ^ x490;
assign n_27995 = n_27990 ^ n_27424;
assign n_27996 = n_27990 ^ n_27431;
assign n_27997 = n_27992 ^ n_26215;
assign n_27998 = n_27986 ^ n_27994;
assign n_27999 = n_27993 ^ n_27994;
assign n_28000 = ~n_27431 & n_27995;
assign n_28001 = n_27579 ^ n_27996;
assign n_28002 = n_27996 ^ n_27424;
assign n_28003 = n_27983 ^ n_27997;
assign n_28004 = n_27991 ^ n_27997;
assign n_28005 = ~n_27993 & n_27998;
assign n_28006 = n_27988 & n_27999;
assign n_28007 = n_27999 ^ n_27988;
assign n_28008 = n_28000 ^ n_27256;
assign n_28009 = n_28002 ^ n_26755;
assign n_28010 = n_27991 & n_28003;
assign n_28011 = n_28004 ^ x488;
assign n_28012 = n_28005 ^ x489;
assign n_28013 = n_28008 ^ n_27443;
assign n_28014 = n_28009 ^ n_26290;
assign n_28015 = n_28010 ^ n_26251;
assign n_28016 = n_28012 ^ n_28004;
assign n_28017 = n_28013 & ~n_27451;
assign n_28018 = n_27274 ^ n_28013;
assign n_28019 = n_28009 ^ n_28015;
assign n_28020 = n_28014 ^ n_28015;
assign n_28021 = ~n_28016 & n_28011;
assign n_28022 = n_28016 ^ x488;
assign n_28023 = n_28017 ^ n_27274;
assign n_28024 = n_28018 ^ n_27443;
assign n_28025 = n_27627 ^ n_28018;
assign n_28026 = n_28014 & n_28019;
assign n_28027 = n_28020 ^ x503;
assign n_28028 = n_28021 ^ x488;
assign n_28029 = ~n_28006 & n_28022;
assign n_28030 = n_28022 ^ n_28006;
assign n_28031 = n_28023 ^ n_27462;
assign n_28032 = n_28023 ^ n_27469;
assign n_28033 = n_28024 ^ n_26795;
assign n_28034 = n_28026 ^ n_26290;
assign n_28035 = n_28020 ^ n_28028;
assign n_28036 = n_27469 & ~n_28031;
assign n_28037 = n_27674 ^ n_28032;
assign n_28038 = n_28032 ^ n_27462;
assign n_28039 = n_28033 ^ n_26329;
assign n_28040 = n_28034 ^ n_28033;
assign n_28041 = n_28035 & ~n_28027;
assign n_28042 = n_28035 ^ x503;
assign n_28043 = n_28036 ^ n_27291;
assign n_28044 = n_28038 ^ n_26834;
assign n_28045 = n_28040 & ~n_28039;
assign n_28046 = n_28040 ^ n_26329;
assign n_28047 = n_28041 ^ x503;
assign n_28048 = n_28029 & ~n_28042;
assign n_28049 = n_28042 ^ n_28029;
assign n_28050 = n_28043 ^ n_27480;
assign n_28051 = n_28043 ^ n_27487;
assign n_28052 = n_28044 ^ n_26368;
assign n_28053 = n_28045 ^ n_26329;
assign n_28054 = n_28046 ^ x502;
assign n_28055 = n_28047 ^ n_28046;
assign n_28056 = ~n_28049 & ~n_27577;
assign n_28057 = n_28049 ^ n_27111;
assign n_28058 = n_28049 ^ n_27562;
assign n_28059 = n_27487 & n_28050;
assign n_28060 = n_28051 ^ n_27721;
assign n_28061 = n_28051 ^ n_27480;
assign n_28062 = n_28053 ^ n_28044;
assign n_28063 = n_28047 ^ n_28054;
assign n_28064 = ~n_28054 & n_28055;
assign n_28065 = n_27598 ^ n_28056;
assign n_28066 = n_26125 & n_28057;
assign n_28067 = x71 & ~n_28057;
assign n_28068 = n_28057 ^ x71;
assign n_28069 = n_28057 ^ n_27568;
assign n_28070 = n_28059 ^ n_27309;
assign n_28071 = n_28061 ^ n_26873;
assign n_28072 = ~n_28062 & n_28052;
assign n_28073 = n_28062 ^ n_26368;
assign n_28074 = n_28063 & ~n_28048;
assign n_28075 = n_28048 ^ n_28063;
assign n_28076 = n_28064 ^ x502;
assign n_28077 = n_28066 ^ n_26153;
assign n_28078 = n_28067 ^ x70;
assign n_28079 = n_28070 ^ n_27498;
assign n_28080 = n_28070 ^ n_27505;
assign n_28081 = n_28071 ^ n_26406;
assign n_28082 = n_28072 ^ n_26368;
assign n_28083 = n_28073 ^ x501;
assign n_28084 = n_28056 ^ n_28075;
assign n_28085 = n_28065 ^ n_28075;
assign n_28086 = n_28076 ^ n_28073;
assign n_28087 = n_27505 & n_28079;
assign n_28088 = n_27768 ^ n_28080;
assign n_28089 = n_28080 ^ n_27498;
assign n_28090 = n_28082 ^ n_28071;
assign n_28091 = n_28076 ^ n_28083;
assign n_28092 = n_28065 & ~n_28084;
assign n_28093 = n_28085 ^ n_27597;
assign n_28094 = n_28083 & ~n_28086;
assign n_28095 = n_28087 ^ n_27326;
assign n_28096 = n_28089 ^ n_26909;
assign n_28097 = ~n_28090 & ~n_28081;
assign n_28098 = n_28090 ^ n_26406;
assign n_28099 = n_28091 & ~n_28074;
assign n_28100 = n_28074 ^ n_28091;
assign n_28101 = n_28092 ^ n_27598;
assign n_28102 = n_28066 ^ n_28093;
assign n_28103 = n_28077 ^ n_28093;
assign n_28104 = n_28094 ^ x501;
assign n_28105 = n_28095 ^ n_27346;
assign n_28106 = n_28095 ^ n_27519;
assign n_28107 = n_28096 ^ n_26445;
assign n_28108 = n_28097 ^ n_26406;
assign n_28109 = n_28098 ^ x500;
assign n_28110 = n_27634 ^ n_28100;
assign n_28111 = n_28101 ^ n_28100;
assign n_28112 = n_28077 & n_28102;
assign n_28113 = n_28067 ^ n_28103;
assign n_28114 = n_28078 ^ n_28103;
assign n_28115 = n_28104 ^ n_28098;
assign n_28116 = n_28105 ^ n_27519;
assign n_28117 = n_28105 ^ n_26936;
assign n_28118 = ~n_27527 & ~n_28106;
assign n_28119 = n_28108 ^ n_28096;
assign n_28120 = n_28104 ^ n_28109;
assign n_28121 = n_28111 & ~n_28110;
assign n_28122 = n_27634 ^ n_28111;
assign n_28123 = n_28112 ^ n_26153;
assign n_28124 = n_28078 & n_28113;
assign n_28125 = ~n_28068 & ~n_28114;
assign n_28126 = n_28114 ^ n_28068;
assign n_28127 = ~n_28109 & n_28115;
assign n_28128 = n_28116 ^ n_27808;
assign n_28129 = n_28117 ^ n_26485;
assign n_28130 = n_28118 ^ n_27346;
assign n_28131 = n_28119 & n_28107;
assign n_28132 = n_28119 ^ n_26445;
assign n_28133 = ~n_28120 & n_28099;
assign n_28134 = n_28099 ^ n_28120;
assign n_28135 = n_28121 ^ n_27634;
assign n_28136 = n_28122 ^ n_27624;
assign n_28137 = n_28123 ^ n_26208;
assign n_28138 = n_28124 ^ x70;
assign n_28139 = n_28127 ^ x500;
assign n_28140 = n_28130 ^ n_27532;
assign n_28141 = n_28130 ^ n_27370;
assign n_28142 = n_28131 ^ n_26445;
assign n_28143 = n_28132 ^ x499;
assign n_28144 = n_28134 ^ n_27668;
assign n_28145 = n_28134 ^ n_28135;
assign n_28146 = n_28136 ^ n_26208;
assign n_28147 = n_28136 ^ n_28123;
assign n_28148 = n_28136 ^ n_28137;
assign n_28149 = n_28139 ^ n_28132;
assign n_28150 = n_27539 & n_28140;
assign n_28151 = n_28141 ^ n_26957;
assign n_28152 = n_28141 ^ n_27532;
assign n_28153 = n_28142 ^ n_28117;
assign n_28154 = n_28142 ^ n_26485;
assign n_28155 = n_28139 ^ n_28143;
assign n_28156 = n_28144 ^ n_28135;
assign n_28157 = ~n_28144 & n_28145;
assign n_28158 = ~n_28146 & n_28147;
assign n_28159 = n_28148 ^ x69;
assign n_28160 = n_28148 ^ n_28138;
assign n_28161 = ~n_28143 & n_28149;
assign n_28162 = n_28150 ^ n_27370;
assign n_28163 = n_28151 ^ n_26524;
assign n_28164 = n_27845 ^ n_28152;
assign n_28165 = n_28129 & n_28153;
assign n_28166 = n_28154 ^ n_28117;
assign n_28167 = n_28133 & ~n_28155;
assign n_28168 = n_28155 ^ n_28133;
assign n_28169 = n_28156 ^ n_27658;
assign n_28170 = n_28157 ^ n_27668;
assign n_28171 = n_28158 ^ n_26208;
assign n_28172 = n_28159 ^ n_28138;
assign n_28173 = ~n_28159 & n_28160;
assign n_28174 = n_28161 ^ x499;
assign n_28175 = n_28162 ^ n_27551;
assign n_28176 = n_28162 ^ n_27558;
assign n_28177 = n_28165 ^ n_26485;
assign n_28178 = n_28166 ^ x498;
assign n_28179 = n_28168 ^ n_27706;
assign n_28180 = n_28169 ^ n_26246;
assign n_28181 = n_28170 ^ n_28168;
assign n_28182 = n_28171 ^ n_28169;
assign n_28183 = ~n_28125 & n_28172;
assign n_28184 = n_28172 ^ n_28125;
assign n_28185 = n_28173 ^ x69;
assign n_28186 = n_28174 ^ n_28166;
assign n_28187 = ~n_27558 & n_28175;
assign n_28188 = n_28176 ^ n_27551;
assign n_28189 = n_27871 ^ n_28176;
assign n_28190 = n_28177 ^ n_28151;
assign n_28191 = n_28174 ^ n_28178;
assign n_28192 = n_28181 & ~n_28179;
assign n_28193 = n_28181 ^ n_27706;
assign n_28194 = ~n_28182 & n_28180;
assign n_28195 = n_28182 ^ n_26246;
assign n_28196 = n_28178 & ~n_28186;
assign n_28197 = n_28187 ^ n_27390;
assign n_28198 = n_28188 ^ n_26968;
assign n_28199 = ~n_28190 & ~n_28163;
assign n_28200 = n_28190 ^ n_26524;
assign n_28201 = ~n_28167 & ~n_28191;
assign n_28202 = n_28191 ^ n_28167;
assign n_28203 = n_28192 ^ n_27706;
assign n_28204 = n_28193 ^ n_27693;
assign n_28205 = n_28194 ^ n_26246;
assign n_28206 = n_28185 ^ n_28195;
assign n_28207 = n_28195 ^ x68;
assign n_28208 = n_28196 ^ x498;
assign n_28209 = n_28197 ^ n_27583;
assign n_28210 = n_27593 ^ n_28197;
assign n_28211 = n_28198 ^ n_26562;
assign n_28212 = n_28199 ^ n_26524;
assign n_28213 = n_28200 ^ x497;
assign n_28214 = n_27742 ^ n_28202;
assign n_28215 = n_28203 ^ n_28202;
assign n_28216 = n_28204 ^ n_26285;
assign n_28217 = n_28204 ^ n_28205;
assign n_28218 = n_28205 ^ n_26285;
assign n_28219 = n_28206 ^ x68;
assign n_28220 = ~n_28206 & n_28207;
assign n_28221 = n_28208 ^ n_28200;
assign n_28222 = ~n_27593 & n_28209;
assign n_28223 = n_28210 ^ n_27583;
assign n_28224 = n_27891 ^ n_28210;
assign n_28225 = n_28212 ^ n_28198;
assign n_28226 = n_28212 ^ n_28211;
assign n_28227 = n_28208 ^ n_28213;
assign n_28228 = n_28203 ^ n_28214;
assign n_28229 = ~n_28214 & n_28215;
assign n_28230 = ~n_28216 & n_28217;
assign n_28231 = n_28204 ^ n_28218;
assign n_28232 = ~n_28183 & n_28219;
assign n_28233 = n_28219 ^ n_28183;
assign n_28234 = n_28220 ^ x68;
assign n_28235 = n_28213 & ~n_28221;
assign n_28236 = n_28222 ^ n_27410;
assign n_28237 = n_28223 ^ n_26988;
assign n_28238 = n_28211 & n_28225;
assign n_28239 = n_28226 ^ x496;
assign n_28240 = ~n_28201 & n_28227;
assign n_28241 = n_28227 ^ n_28201;
assign n_28242 = n_28228 ^ n_27730;
assign n_28243 = n_28229 ^ n_27742;
assign n_28244 = n_28230 ^ n_26285;
assign n_28245 = n_28231 ^ x67;
assign n_28246 = n_28234 ^ n_28231;
assign n_28247 = n_28235 ^ x497;
assign n_28248 = n_28236 ^ n_27607;
assign n_28249 = n_28236 ^ n_27618;
assign n_28250 = n_28237 ^ n_26602;
assign n_28251 = n_28238 ^ n_26562;
assign n_28252 = n_27775 ^ n_28241;
assign n_28253 = n_28242 ^ n_26324;
assign n_28254 = n_28241 ^ n_28243;
assign n_28255 = n_28242 ^ n_28244;
assign n_28256 = n_28246 & ~n_28245;
assign n_28257 = n_28246 ^ x67;
assign n_28258 = n_28247 ^ n_28226;
assign n_28259 = n_28247 ^ x496;
assign n_28260 = ~n_27618 & ~n_28248;
assign n_28261 = n_28249 ^ n_27607;
assign n_28262 = n_27910 ^ n_28249;
assign n_28263 = n_28251 ^ n_28237;
assign n_28264 = n_28252 ^ n_28243;
assign n_28265 = n_28253 ^ n_28244;
assign n_28266 = n_28252 & n_28254;
assign n_28267 = n_28253 & n_28255;
assign n_28268 = n_28256 ^ x67;
assign n_28269 = n_28232 & ~n_28257;
assign n_28270 = n_28257 ^ n_28232;
assign n_28271 = n_28239 & ~n_28258;
assign n_28272 = n_28259 ^ n_28226;
assign n_28273 = n_28260 ^ n_27429;
assign n_28274 = n_28261 ^ n_27015;
assign n_28275 = n_28263 & ~n_28250;
assign n_28276 = n_28263 ^ n_26602;
assign n_28277 = n_28264 ^ n_27766;
assign n_28278 = n_28265 ^ x66;
assign n_28279 = n_28266 ^ n_27775;
assign n_28280 = n_28267 ^ n_26324;
assign n_28281 = n_28268 ^ n_28265;
assign n_28282 = n_28271 ^ x496;
assign n_28283 = ~n_28240 & ~n_28272;
assign n_28284 = n_28272 ^ n_28240;
assign n_28285 = n_28273 ^ n_27640;
assign n_28286 = n_27448 ^ n_28273;
assign n_28287 = n_28274 ^ n_26642;
assign n_28288 = n_28275 ^ n_26602;
assign n_28289 = n_28276 ^ x511;
assign n_28290 = n_28277 ^ n_26363;
assign n_28291 = n_28280 ^ n_28277;
assign n_28292 = n_28280 ^ n_26363;
assign n_28293 = ~n_28281 & n_28278;
assign n_28294 = n_28281 ^ x66;
assign n_28295 = n_28282 ^ n_28276;
assign n_28296 = n_27819 ^ n_28284;
assign n_28297 = n_28279 ^ n_28284;
assign n_28298 = n_27652 & ~n_28285;
assign n_28299 = n_28286 ^ n_27035;
assign n_28300 = n_28286 ^ n_27640;
assign n_28301 = n_28288 ^ n_28274;
assign n_28302 = n_28282 ^ n_28289;
assign n_28303 = ~n_28290 & ~n_28291;
assign n_28304 = n_28292 ^ n_28277;
assign n_28305 = n_28293 ^ x66;
assign n_28306 = ~n_28269 & ~n_28294;
assign n_28307 = n_28294 ^ n_28269;
assign n_28308 = n_28289 & ~n_28295;
assign n_28309 = n_28279 ^ n_28296;
assign n_28310 = ~n_28296 & ~n_28297;
assign n_28311 = n_28298 ^ n_27448;
assign n_28312 = n_28299 ^ n_26682;
assign n_28313 = n_27928 ^ n_28300;
assign n_28314 = ~n_28301 & ~n_28287;
assign n_28315 = n_28301 ^ n_26642;
assign n_28316 = ~n_28302 & n_28283;
assign n_28317 = n_28283 ^ n_28302;
assign n_28318 = n_28303 ^ n_26363;
assign n_28319 = n_28304 ^ x65;
assign n_28320 = n_28304 ^ n_28305;
assign n_28321 = n_28308 ^ x511;
assign n_28322 = n_28309 ^ n_27805;
assign n_28323 = n_28310 ^ n_27819;
assign n_28324 = n_28311 ^ n_27663;
assign n_28325 = n_27677 ^ n_28311;
assign n_28326 = n_28314 ^ n_26642;
assign n_28327 = n_28315 ^ x510;
assign n_28328 = n_27849 ^ n_28317;
assign n_28329 = n_28318 ^ n_26401;
assign n_28330 = n_28319 ^ n_28305;
assign n_28331 = n_28319 & ~n_28320;
assign n_28332 = n_28321 ^ n_28315;
assign n_28333 = n_28321 ^ x510;
assign n_28334 = n_28322 ^ n_26401;
assign n_28335 = n_28318 ^ n_28322;
assign n_28336 = n_28323 ^ n_28317;
assign n_28337 = ~n_27677 & n_28324;
assign n_28338 = n_28325 ^ n_27663;
assign n_28339 = n_27945 ^ n_28325;
assign n_28340 = n_28299 ^ n_28326;
assign n_28341 = n_28312 ^ n_28326;
assign n_28342 = n_28329 ^ n_28322;
assign n_28343 = n_28306 & ~n_28330;
assign n_28344 = n_28330 ^ n_28306;
assign n_28345 = n_28331 ^ x65;
assign n_28346 = n_28327 & ~n_28332;
assign n_28347 = n_28333 ^ n_28315;
assign n_28348 = ~n_28334 & n_28335;
assign n_28349 = ~n_28336 & n_28328;
assign n_28350 = n_27849 ^ n_28336;
assign n_28351 = n_28337 ^ n_27467;
assign n_28352 = n_28338 ^ n_27052;
assign n_28353 = n_28312 & ~n_28340;
assign n_28354 = n_28341 ^ x509;
assign n_28355 = n_28342 ^ x64;
assign n_28356 = n_28345 ^ n_28342;
assign n_28357 = n_28346 ^ x510;
assign n_28358 = n_28316 & ~n_28347;
assign n_28359 = n_28347 ^ n_28316;
assign n_28360 = n_28348 ^ n_26401;
assign n_28361 = n_28349 ^ n_27849;
assign n_28362 = n_28350 ^ n_27842;
assign n_28363 = n_28351 ^ n_27698;
assign n_28364 = n_27711 ^ n_28351;
assign n_28365 = n_28352 ^ n_26722;
assign n_28366 = n_28353 ^ n_26682;
assign n_28367 = n_28356 & ~n_28355;
assign n_28368 = n_28356 ^ x64;
assign n_28369 = n_28341 ^ n_28357;
assign n_28370 = n_28357 ^ x509;
assign n_28371 = n_28359 ^ n_27873;
assign n_28372 = n_28361 ^ n_28359;
assign n_28373 = n_28360 ^ n_28362;
assign n_28374 = n_28362 ^ n_26440;
assign n_28375 = n_27711 & ~n_28363;
assign n_28376 = n_28364 ^ n_27698;
assign n_28377 = n_27964 ^ n_28364;
assign n_28378 = n_28352 ^ n_28366;
assign n_28379 = n_28366 ^ n_26722;
assign n_28380 = n_28367 ^ x64;
assign n_28381 = ~n_28343 & ~n_28368;
assign n_28382 = n_28368 ^ n_28343;
assign n_28383 = n_28354 & ~n_28369;
assign n_28384 = n_28341 ^ n_28370;
assign n_28385 = n_28361 ^ n_28371;
assign n_28386 = n_28371 & ~n_28372;
assign n_28387 = n_28373 ^ n_26440;
assign n_28388 = ~n_28373 & n_28374;
assign n_28389 = n_28375 ^ n_27485;
assign n_28390 = n_28376 ^ n_27073;
assign n_28391 = n_28365 & ~n_28378;
assign n_28392 = n_28352 ^ n_28379;
assign n_28393 = n_28383 ^ x509;
assign n_28394 = n_28358 & ~n_28384;
assign n_28395 = n_28384 ^ n_28358;
assign n_28396 = n_28385 ^ n_27867;
assign n_28397 = n_28386 ^ n_27873;
assign n_28398 = n_28380 ^ n_28387;
assign n_28399 = n_28387 ^ x79;
assign n_28400 = n_28388 ^ n_26440;
assign n_28401 = n_28389 ^ n_27747;
assign n_28402 = n_27504 ^ n_28389;
assign n_28403 = n_28390 ^ n_26761;
assign n_28404 = n_28391 ^ n_26722;
assign n_28405 = n_28392 ^ x508;
assign n_28406 = n_28392 ^ n_28393;
assign n_28407 = n_28393 ^ x508;
assign n_28408 = n_28395 ^ n_27895;
assign n_28409 = n_28396 ^ n_26480;
assign n_28410 = n_28395 ^ n_28397;
assign n_28411 = n_28398 ^ x79;
assign n_28412 = ~n_28398 & n_28399;
assign n_28413 = n_28400 ^ n_28396;
assign n_28414 = n_28400 ^ n_26480;
assign n_28415 = n_27761 & n_28401;
assign n_28416 = n_28402 ^ n_27089;
assign n_28417 = n_28402 ^ n_27747;
assign n_28418 = n_28390 ^ n_28404;
assign n_28419 = n_28404 ^ n_26761;
assign n_28420 = n_28405 & ~n_28406;
assign n_28421 = n_28392 ^ n_28407;
assign n_28422 = n_28408 ^ n_28397;
assign n_28423 = n_28408 & ~n_28410;
assign n_28424 = n_28381 & n_28411;
assign n_28425 = n_28412 ^ x79;
assign n_28426 = n_28409 & n_28413;
assign n_28427 = n_28414 ^ n_28396;
assign n_28428 = n_28415 ^ n_27504;
assign n_28429 = n_28416 ^ n_26800;
assign n_28430 = n_28417 ^ n_27989;
assign n_28431 = ~n_28403 & n_28418;
assign n_28432 = n_28390 ^ n_28419;
assign n_28433 = n_28420 ^ x508;
assign n_28434 = n_28394 & ~n_28421;
assign n_28435 = n_28421 ^ n_28394;
assign n_28436 = n_28422 ^ n_27887;
assign n_28437 = n_28423 ^ n_27895;
assign n_28438 = n_28426 ^ n_26480;
assign n_28439 = n_28427 ^ x78;
assign n_28440 = n_28425 ^ n_28427;
assign n_28441 = n_27524 ^ n_28428;
assign n_28442 = n_28428 ^ n_27773;
assign n_28443 = n_27786 ^ n_28428;
assign n_28444 = n_28431 ^ n_26761;
assign n_28445 = n_28432 ^ x507;
assign n_28446 = n_28432 ^ n_28433;
assign n_28447 = n_28435 ^ n_27914;
assign n_28448 = n_28436 ^ n_26519;
assign n_28449 = n_28437 ^ n_28435;
assign n_28450 = n_28436 ^ n_28438;
assign n_28451 = n_28425 ^ n_28439;
assign n_28452 = n_28439 & ~n_28440;
assign n_28453 = n_28441 ^ n_27108;
assign n_28454 = ~n_28441 & n_28442;
assign n_28455 = n_28007 ^ n_28443;
assign n_28456 = n_28444 ^ n_28416;
assign n_28457 = n_28445 ^ n_28433;
assign n_28458 = ~n_28445 & n_28446;
assign n_28459 = n_28448 ^ n_28438;
assign n_28460 = ~n_28449 & n_28447;
assign n_28461 = n_28449 ^ n_27914;
assign n_28462 = ~n_28448 & ~n_28450;
assign n_28463 = ~n_28424 & ~n_28451;
assign n_28464 = n_28451 ^ n_28424;
assign n_28465 = n_28452 ^ x78;
assign n_28466 = n_28453 ^ n_26838;
assign n_28467 = n_27836 ^ n_28454;
assign n_28468 = n_28456 & ~n_28429;
assign n_28469 = n_28456 ^ n_26800;
assign n_28470 = n_28434 & n_28457;
assign n_28471 = n_28457 ^ n_28434;
assign n_28472 = n_28458 ^ x507;
assign n_28473 = n_28459 ^ x77;
assign n_28474 = n_28460 ^ n_27914;
assign n_28475 = n_28461 ^ n_27906;
assign n_28476 = n_28462 ^ n_26519;
assign n_28477 = n_28069 & ~n_28464;
assign n_28478 = n_28464 ^ n_28069;
assign n_28479 = n_28464 ^ n_28049;
assign n_28480 = n_28459 ^ n_28465;
assign n_28481 = n_28465 ^ x77;
assign n_28482 = n_28467 ^ n_27812;
assign n_28483 = n_28030 ^ n_28467;
assign n_28484 = n_28468 ^ n_26800;
assign n_28485 = n_28469 ^ x506;
assign n_28486 = n_28471 ^ n_27931;
assign n_28487 = n_28472 ^ n_28469;
assign n_28488 = n_28471 ^ n_28474;
assign n_28489 = n_28475 ^ n_26558;
assign n_28490 = n_28475 ^ n_28476;
assign n_28491 = n_28476 ^ n_26558;
assign n_28492 = ~n_27577 & n_28478;
assign n_28493 = n_28473 & ~n_28480;
assign n_28494 = n_28459 ^ n_28481;
assign n_28495 = n_28482 ^ n_27125;
assign n_28496 = n_28483 ^ n_28007;
assign n_28497 = n_28453 ^ n_28484;
assign n_28498 = n_28484 ^ n_26838;
assign n_28499 = n_28472 ^ n_28485;
assign n_28500 = n_28486 ^ n_28474;
assign n_28501 = ~n_28485 & n_28487;
assign n_28502 = n_28486 & n_28488;
assign n_28503 = n_28489 & ~n_28490;
assign n_28504 = n_28475 ^ n_28491;
assign n_28505 = n_28492 ^ n_28069;
assign n_28506 = n_28492 ^ n_28058;
assign n_28507 = n_28493 ^ x77;
assign n_28508 = n_28463 & ~n_28494;
assign n_28509 = n_28494 ^ n_28463;
assign n_28510 = n_28495 ^ n_26877;
assign n_28511 = ~n_28466 & ~n_28497;
assign n_28512 = n_28453 ^ n_28498;
assign n_28513 = ~n_28470 & ~n_28499;
assign n_28514 = n_28499 ^ n_28470;
assign n_28515 = n_28500 ^ n_27936;
assign n_28516 = n_28501 ^ x506;
assign n_28517 = n_28502 ^ n_27931;
assign n_28518 = n_28503 ^ n_26558;
assign n_28519 = n_28504 ^ x76;
assign n_28520 = n_27121 & ~n_28505;
assign n_28521 = x7 & ~n_28506;
assign n_28522 = n_28506 ^ x7;
assign n_28523 = n_28504 ^ n_28507;
assign n_28524 = n_28477 ^ n_28509;
assign n_28525 = n_28509 ^ n_28085;
assign n_28526 = n_28511 ^ n_26838;
assign n_28527 = n_28512 ^ x505;
assign n_28528 = n_28514 ^ n_27941;
assign n_28529 = n_28515 ^ n_26598;
assign n_28530 = n_28516 ^ n_28512;
assign n_28531 = n_28516 ^ x505;
assign n_28532 = n_28517 ^ n_28514;
assign n_28533 = n_28515 ^ n_28518;
assign n_28534 = n_28519 ^ n_28507;
assign n_28535 = n_28521 ^ x6;
assign n_28536 = n_28519 & ~n_28523;
assign n_28537 = n_28524 ^ n_28085;
assign n_28538 = ~n_28524 & n_28525;
assign n_28539 = n_28526 ^ n_28510;
assign n_28540 = n_28516 ^ n_28527;
assign n_28541 = n_28529 ^ n_28518;
assign n_28542 = n_28530 & n_28531;
assign n_28543 = n_28532 & ~n_28528;
assign n_28544 = n_28532 ^ n_27941;
assign n_28545 = n_28529 & ~n_28533;
assign n_28546 = ~n_28508 & n_28534;
assign n_28547 = n_28534 ^ n_28508;
assign n_28548 = n_28536 ^ x76;
assign n_28549 = n_27598 & ~n_28537;
assign n_28550 = n_28538 ^ n_28085;
assign n_28551 = n_28539 ^ x504;
assign n_28552 = ~n_28540 & n_28513;
assign n_28553 = n_28513 ^ n_28540;
assign n_28554 = n_28541 ^ x75;
assign n_28555 = n_28543 ^ n_27941;
assign n_28556 = n_28544 ^ n_27947;
assign n_28557 = n_28545 ^ n_26598;
assign n_28558 = n_28547 ^ n_28122;
assign n_28559 = n_28541 ^ n_28548;
assign n_28560 = n_28549 ^ n_28085;
assign n_28561 = n_28547 ^ n_28550;
assign n_28562 = n_28550 ^ n_28122;
assign n_28563 = n_28551 ^ x505;
assign n_28564 = n_28553 ^ n_27959;
assign n_28565 = n_28554 ^ n_28548;
assign n_28566 = n_28555 ^ n_28553;
assign n_28567 = n_28555 ^ n_27959;
assign n_28568 = n_28556 ^ n_26638;
assign n_28569 = n_28557 ^ n_28556;
assign n_28570 = n_28557 ^ n_26638;
assign n_28571 = n_28554 & ~n_28559;
assign n_28572 = n_28560 ^ n_28520;
assign n_28573 = n_28560 ^ n_27145;
assign n_28574 = n_28558 & n_28561;
assign n_28575 = n_28547 ^ n_28562;
assign n_28576 = n_28563 ^ n_28542;
assign n_28577 = ~n_28565 & ~n_28546;
assign n_28578 = n_28546 ^ n_28565;
assign n_28579 = n_28564 & ~n_28566;
assign n_28580 = n_28567 ^ n_28553;
assign n_28581 = ~n_28568 & ~n_28569;
assign n_28582 = n_28570 ^ n_28556;
assign n_28583 = n_28571 ^ x75;
assign n_28584 = n_28572 ^ n_27145;
assign n_28585 = n_28572 & n_28573;
assign n_28586 = n_28574 ^ n_28122;
assign n_28587 = n_27634 & ~n_28575;
assign n_28588 = n_28576 ^ n_28552;
assign n_28589 = n_28578 ^ n_28156;
assign n_28590 = n_28579 ^ n_27959;
assign n_28591 = n_28580 ^ n_27966;
assign n_28592 = n_28581 ^ n_26638;
assign n_28593 = n_28582 ^ x74;
assign n_28594 = n_28583 ^ n_28582;
assign n_28595 = n_28583 ^ x74;
assign n_28596 = n_28584 ^ n_28521;
assign n_28597 = n_28584 ^ n_28535;
assign n_28598 = n_28585 ^ n_27145;
assign n_28599 = n_28578 ^ n_28586;
assign n_28600 = n_28586 ^ n_28156;
assign n_28601 = n_28587 ^ n_28122;
assign n_28602 = n_28588 ^ n_27984;
assign n_28603 = n_28588 ^ n_28590;
assign n_28604 = n_27984 ^ n_28590;
assign n_28605 = n_28591 ^ n_26678;
assign n_28606 = n_28592 ^ n_28591;
assign n_28607 = ~n_28593 & n_28594;
assign n_28608 = n_28595 ^ n_28582;
assign n_28609 = n_28535 & ~n_28596;
assign n_28610 = n_28598 ^ n_27170;
assign n_28611 = n_28589 & ~n_28599;
assign n_28612 = n_28578 ^ n_28600;
assign n_28613 = n_28598 ^ n_28601;
assign n_28614 = n_28602 & ~n_28603;
assign n_28615 = n_28588 ^ n_28604;
assign n_28616 = n_28592 ^ n_28605;
assign n_28617 = n_28605 & ~n_28606;
assign n_28618 = n_28607 ^ x74;
assign n_28619 = ~n_28608 & ~n_28577;
assign n_28620 = n_28577 ^ n_28608;
assign n_28621 = n_28609 ^ x6;
assign n_28622 = n_28610 ^ n_28601;
assign n_28623 = n_28611 ^ n_28156;
assign n_28624 = n_27668 & n_28612;
assign n_28625 = ~n_28610 & n_28613;
assign n_28626 = n_28614 ^ n_27984;
assign n_28627 = n_28615 ^ n_27976;
assign n_28628 = n_28616 ^ x73;
assign n_28629 = n_28617 ^ n_26678;
assign n_28630 = n_28618 ^ n_28616;
assign n_28631 = n_28620 ^ n_28193;
assign n_28632 = n_28621 ^ x5;
assign n_28633 = n_28622 ^ x5;
assign n_28634 = n_28622 ^ n_28621;
assign n_28635 = n_28623 ^ n_28620;
assign n_28636 = n_28624 ^ n_28156;
assign n_28637 = n_28625 ^ n_27170;
assign n_28638 = n_28626 ^ n_27996;
assign n_28639 = n_28001 ^ n_28626;
assign n_28640 = n_28618 ^ n_28628;
assign n_28641 = n_28629 ^ n_26718;
assign n_28642 = n_28629 ^ n_28627;
assign n_28643 = ~n_28628 & n_28630;
assign n_28644 = n_28622 ^ n_28632;
assign n_28645 = ~n_28633 & n_28634;
assign n_28646 = n_28635 & ~n_28631;
assign n_28647 = n_28635 ^ n_28193;
assign n_28648 = n_28636 ^ n_27190;
assign n_28649 = n_28636 ^ n_28637;
assign n_28650 = n_28637 ^ n_27190;
assign n_28651 = ~n_28001 & n_28638;
assign n_28652 = n_28639 ^ n_28002;
assign n_28653 = ~n_28619 & n_28640;
assign n_28654 = n_28640 ^ n_28619;
assign n_28655 = n_28641 ^ n_28627;
assign n_28656 = n_28641 & ~n_28642;
assign n_28657 = n_28643 ^ x73;
assign n_28658 = n_28645 ^ x5;
assign n_28659 = n_28646 ^ n_28193;
assign n_28660 = n_27706 & ~n_28647;
assign n_28661 = ~n_28648 & ~n_28649;
assign n_28662 = n_28636 ^ n_28650;
assign n_28663 = n_28651 ^ n_27579;
assign n_28664 = n_28652 ^ n_26755;
assign n_28665 = n_28654 ^ n_28228;
assign n_28666 = n_28655 ^ x72;
assign n_28667 = n_28656 ^ n_26718;
assign n_28668 = n_28657 ^ n_28655;
assign n_28669 = n_28658 ^ x4;
assign n_28670 = n_28659 ^ n_28654;
assign n_28671 = n_28660 ^ n_28193;
assign n_28672 = n_28661 ^ n_27190;
assign n_28673 = n_28658 ^ n_28662;
assign n_28674 = n_28663 ^ n_28018;
assign n_28675 = n_28659 ^ n_28665;
assign n_28676 = n_28657 ^ n_28666;
assign n_28677 = n_28652 ^ n_28667;
assign n_28678 = n_28664 ^ n_28667;
assign n_28679 = ~n_28666 & n_28668;
assign n_28680 = n_28669 ^ n_28662;
assign n_28681 = ~n_28665 & n_28670;
assign n_28682 = n_28671 ^ n_27203;
assign n_28683 = n_28672 ^ n_28671;
assign n_28684 = n_28672 ^ n_27203;
assign n_28685 = n_28669 & n_28673;
assign n_28686 = n_28674 & n_28025;
assign n_28687 = n_28674 ^ n_27627;
assign n_28688 = n_27742 & ~n_28675;
assign n_28689 = ~n_28676 & ~n_28653;
assign n_28690 = n_28653 ^ n_28676;
assign n_28691 = n_28664 & n_28677;
assign n_28692 = n_28678 ^ x87;
assign n_28693 = n_28679 ^ x72;
assign n_28694 = ~n_28644 & ~n_28680;
assign n_28695 = n_28680 ^ n_28644;
assign n_28696 = n_28681 ^ n_28228;
assign n_28697 = n_28682 & n_28683;
assign n_28698 = n_28684 ^ n_28671;
assign n_28699 = n_28685 ^ x4;
assign n_28700 = n_28686 ^ n_27627;
assign n_28701 = n_28687 ^ n_28024;
assign n_28702 = n_28688 ^ n_28228;
assign n_28703 = n_28690 ^ n_28264;
assign n_28704 = n_28691 ^ n_26755;
assign n_28705 = n_28678 ^ n_28693;
assign n_28706 = n_28692 ^ n_28693;
assign n_28707 = n_28696 ^ n_28690;
assign n_28708 = n_28697 ^ n_27203;
assign n_28709 = n_28698 ^ x3;
assign n_28710 = n_28699 ^ n_28698;
assign n_28711 = n_28699 ^ x3;
assign n_28712 = n_28700 ^ n_28032;
assign n_28713 = n_28037 ^ n_28700;
assign n_28714 = n_28701 ^ n_26795;
assign n_28715 = n_28702 ^ n_27223;
assign n_28716 = n_28704 ^ n_28701;
assign n_28717 = ~n_28692 & n_28705;
assign n_28718 = ~n_28706 & n_28689;
assign n_28719 = n_28689 ^ n_28706;
assign n_28720 = n_28707 & n_28703;
assign n_28721 = n_28707 ^ n_28264;
assign n_28722 = n_28708 ^ n_28702;
assign n_28723 = ~n_28709 & n_28710;
assign n_28724 = n_28711 ^ n_28698;
assign n_28725 = n_28037 & n_28712;
assign n_28726 = n_28713 ^ n_28038;
assign n_28727 = n_28708 ^ n_28715;
assign n_28728 = n_28716 & n_28714;
assign n_28729 = n_28716 ^ n_26795;
assign n_28730 = n_28717 ^ x87;
assign n_28731 = n_28719 ^ n_28309;
assign n_28732 = n_28720 ^ n_28264;
assign n_28733 = ~n_27775 & n_28721;
assign n_28734 = n_28721 ^ n_28522;
assign n_28735 = n_28715 & ~n_28722;
assign n_28736 = n_28723 ^ x3;
assign n_28737 = n_28694 & ~n_28724;
assign n_28738 = n_28724 ^ n_28694;
assign n_28739 = n_28725 ^ n_27674;
assign n_28740 = n_28726 ^ n_26834;
assign n_28741 = n_28727 ^ x2;
assign n_28742 = n_28728 ^ n_26795;
assign n_28743 = n_28729 ^ x86;
assign n_28744 = n_28730 ^ x86;
assign n_28745 = n_28730 ^ n_28729;
assign n_28746 = n_28732 ^ n_28719;
assign n_28747 = n_28733 ^ n_28264;
assign n_28748 = n_28735 ^ n_27223;
assign n_28749 = n_28736 ^ n_28727;
assign n_28750 = n_28736 ^ x2;
assign n_28751 = n_28739 ^ n_28051;
assign n_28752 = n_28739 ^ n_28060;
assign n_28753 = n_28726 ^ n_28742;
assign n_28754 = n_28742 ^ n_26834;
assign n_28755 = n_28730 ^ n_28743;
assign n_28756 = n_28744 & ~n_28745;
assign n_28757 = n_28746 & ~n_28731;
assign n_28758 = n_28746 ^ n_28309;
assign n_28759 = n_28747 ^ n_27241;
assign n_28760 = n_28748 ^ n_28747;
assign n_28761 = n_28748 ^ n_27241;
assign n_28762 = n_28741 & ~n_28749;
assign n_28763 = n_28750 ^ n_28727;
assign n_28764 = ~n_28060 & ~n_28751;
assign n_28765 = n_28752 ^ n_28061;
assign n_28766 = n_28740 & n_28753;
assign n_28767 = n_28726 ^ n_28754;
assign n_28768 = n_28718 & n_28755;
assign n_28769 = n_28755 ^ n_28718;
assign n_28770 = n_28756 ^ x86;
assign n_28771 = n_28757 ^ n_28309;
assign n_28772 = n_27819 & n_28758;
assign n_28773 = n_28758 ^ n_28597;
assign n_28774 = ~n_28759 & n_28760;
assign n_28775 = n_28761 ^ n_28747;
assign n_28776 = n_28762 ^ x2;
assign n_28777 = n_28763 & n_28737;
assign n_28778 = n_28737 ^ n_28763;
assign n_28779 = n_28764 ^ n_27721;
assign n_28780 = n_28765 ^ n_26873;
assign n_28781 = n_28766 ^ n_26834;
assign n_28782 = n_28767 ^ x85;
assign n_28783 = n_28769 ^ n_28350;
assign n_28784 = n_28770 ^ n_28767;
assign n_28785 = n_28771 ^ n_28769;
assign n_28786 = n_28772 ^ n_28309;
assign n_28787 = n_28774 ^ n_27241;
assign n_28788 = n_28775 ^ x1;
assign n_28789 = n_28776 ^ n_28775;
assign n_28790 = n_28779 ^ n_28080;
assign n_28791 = n_28779 ^ n_28088;
assign n_28792 = n_28781 ^ n_28765;
assign n_28793 = n_28781 ^ n_28780;
assign n_28794 = n_28771 ^ n_28783;
assign n_28795 = n_28784 & ~n_28782;
assign n_28796 = n_28784 ^ x85;
assign n_28797 = n_28783 & ~n_28785;
assign n_28798 = n_28786 ^ n_27259;
assign n_28799 = n_28787 ^ n_28786;
assign n_28800 = n_28776 ^ n_28788;
assign n_28801 = ~n_28788 & n_28789;
assign n_28802 = n_28088 & ~n_28790;
assign n_28803 = n_28791 ^ n_28089;
assign n_28804 = n_28780 & n_28792;
assign n_28805 = n_28793 ^ x84;
assign n_28806 = n_27849 & ~n_28794;
assign n_28807 = n_28794 ^ n_28644;
assign n_28808 = n_28795 ^ x85;
assign n_28809 = ~n_28768 & n_28796;
assign n_28810 = n_28796 ^ n_28768;
assign n_28811 = n_28797 ^ n_28350;
assign n_28812 = n_28799 & n_28798;
assign n_28813 = n_28799 ^ n_27259;
assign n_28814 = ~n_28777 & n_28800;
assign n_28815 = n_28800 ^ n_28777;
assign n_28816 = n_28801 ^ x1;
assign n_28817 = n_28802 ^ n_27768;
assign n_28818 = n_28803 ^ n_26909;
assign n_28819 = n_28804 ^ n_26873;
assign n_28820 = n_28806 ^ n_28350;
assign n_28821 = n_28808 ^ n_28793;
assign n_28822 = n_28808 ^ n_28805;
assign n_28823 = n_28810 ^ n_28385;
assign n_28824 = n_28810 ^ n_28811;
assign n_28825 = n_28812 ^ n_27259;
assign n_28826 = n_28813 ^ x0;
assign n_28827 = n_28816 ^ n_28813;
assign n_28828 = n_28816 ^ x0;
assign n_28829 = n_28817 ^ n_28116;
assign n_28830 = n_28817 ^ n_28128;
assign n_28831 = n_28819 ^ n_28803;
assign n_28832 = n_28819 ^ n_28818;
assign n_28833 = n_28820 ^ n_27277;
assign n_28834 = n_28805 & ~n_28821;
assign n_28835 = ~n_28822 & n_28809;
assign n_28836 = n_28809 ^ n_28822;
assign n_28837 = n_28823 ^ n_28811;
assign n_28838 = n_28823 & ~n_28824;
assign n_28839 = n_28825 ^ n_28820;
assign n_28840 = n_28825 ^ n_27277;
assign n_28841 = n_28826 & ~n_28827;
assign n_28842 = n_28828 ^ n_28813;
assign n_28843 = ~n_28128 & ~n_28829;
assign n_28844 = n_28830 ^ n_28105;
assign n_28845 = n_28818 & ~n_28831;
assign n_28846 = n_28832 ^ x83;
assign n_28847 = n_28834 ^ x84;
assign n_28848 = n_28836 ^ n_28422;
assign n_28849 = n_27873 & ~n_28837;
assign n_28850 = n_28837 ^ n_28695;
assign n_28851 = n_28838 ^ n_28385;
assign n_28852 = ~n_28833 & ~n_28839;
assign n_28853 = n_28840 ^ n_28820;
assign n_28854 = n_28841 ^ x0;
assign n_28855 = ~n_28814 & n_28842;
assign n_28856 = n_28842 ^ n_28814;
assign n_28857 = n_28843 ^ n_27808;
assign n_28858 = n_28844 ^ n_26936;
assign n_28859 = n_28845 ^ n_26909;
assign n_28860 = n_28847 ^ n_28832;
assign n_28861 = n_28849 ^ n_28385;
assign n_28862 = n_28851 ^ n_28836;
assign n_28863 = n_28851 ^ n_28422;
assign n_28864 = n_28852 ^ n_27277;
assign n_28865 = n_28853 ^ x15;
assign n_28866 = n_28854 ^ n_28853;
assign n_28867 = n_28857 ^ n_28152;
assign n_28868 = n_28859 ^ n_28844;
assign n_28869 = n_28859 ^ n_28858;
assign n_28870 = n_28860 & ~n_28846;
assign n_28871 = n_28860 ^ x83;
assign n_28872 = n_28861 ^ n_27295;
assign n_28873 = n_28848 & ~n_28862;
assign n_28874 = n_28863 ^ n_28836;
assign n_28875 = n_28864 ^ n_28861;
assign n_28876 = n_28864 ^ n_27295;
assign n_28877 = ~n_28866 & n_28865;
assign n_28878 = n_28866 ^ x15;
assign n_28879 = n_28867 & n_28164;
assign n_28880 = n_27845 ^ n_28867;
assign n_28881 = n_28858 & n_28868;
assign n_28882 = n_28869 ^ x82;
assign n_28883 = n_28870 ^ x83;
assign n_28884 = ~n_28871 & ~n_28835;
assign n_28885 = n_28835 ^ n_28871;
assign n_28886 = n_28873 ^ n_28422;
assign n_28887 = n_27895 & ~n_28874;
assign n_28888 = n_28738 ^ n_28874;
assign n_28889 = n_28872 & n_28875;
assign n_28890 = n_28876 ^ n_28861;
assign n_28891 = n_28877 ^ x15;
assign n_28892 = n_28855 & n_28878;
assign n_28893 = n_28878 ^ n_28855;
assign n_28894 = n_28879 ^ n_27845;
assign n_28895 = n_28880 ^ n_28141;
assign n_28896 = n_28881 ^ n_26936;
assign n_28897 = n_28883 ^ n_28869;
assign n_28898 = n_28885 ^ n_28461;
assign n_28899 = n_28886 ^ n_28885;
assign n_28900 = n_28887 ^ n_28422;
assign n_28901 = n_28889 ^ n_27295;
assign n_28902 = n_28890 ^ x14;
assign n_28903 = n_28891 ^ n_28890;
assign n_28904 = n_28891 ^ x14;
assign n_28905 = n_28894 ^ n_27871;
assign n_28906 = n_28894 ^ n_28176;
assign n_28907 = n_28895 ^ n_26957;
assign n_28908 = n_28896 ^ n_28895;
assign n_28909 = n_28896 ^ n_26957;
assign n_28910 = n_28897 & ~n_28882;
assign n_28911 = n_28897 ^ x82;
assign n_28912 = n_28886 ^ n_28898;
assign n_28913 = n_28898 & ~n_28899;
assign n_28914 = n_28900 ^ n_27314;
assign n_28915 = n_28901 ^ n_28900;
assign n_28916 = n_28901 ^ n_27314;
assign n_28917 = n_28902 & ~n_28903;
assign n_28918 = n_28904 ^ n_28890;
assign n_28919 = n_28905 ^ n_28176;
assign n_28920 = n_28189 & ~n_28906;
assign n_28921 = n_28907 & ~n_28908;
assign n_28922 = n_28909 ^ n_28895;
assign n_28923 = n_28910 ^ x82;
assign n_28924 = ~n_28884 & n_28911;
assign n_28925 = n_28911 ^ n_28884;
assign n_28926 = n_27914 & ~n_28912;
assign n_28927 = n_28778 ^ n_28912;
assign n_28928 = n_28913 ^ n_28461;
assign n_28929 = n_28914 & ~n_28915;
assign n_28930 = n_28916 ^ n_28900;
assign n_28931 = n_28917 ^ x14;
assign n_28932 = ~n_28892 & ~n_28918;
assign n_28933 = n_28918 ^ n_28892;
assign n_28934 = n_28919 ^ n_28188;
assign n_28935 = n_28919 ^ n_28068;
assign n_28936 = n_28920 ^ n_27871;
assign n_28937 = n_28921 ^ n_26957;
assign n_28938 = n_28922 ^ x81;
assign n_28939 = n_28923 ^ n_28922;
assign n_28940 = n_28925 ^ n_28500;
assign n_28941 = n_28926 ^ n_28461;
assign n_28942 = n_28928 ^ n_28925;
assign n_28943 = n_28929 ^ n_27314;
assign n_28944 = n_28930 ^ x13;
assign n_28945 = n_28931 ^ n_28930;
assign n_28946 = n_28934 ^ n_26968;
assign n_28947 = n_28936 ^ n_28224;
assign n_28948 = n_28936 ^ n_28210;
assign n_28949 = n_28937 ^ n_28934;
assign n_28950 = n_28937 ^ n_26968;
assign n_28951 = ~n_28939 & n_28938;
assign n_28952 = n_28939 ^ x81;
assign n_28953 = n_28928 ^ n_28940;
assign n_28954 = n_28941 ^ n_27331;
assign n_28955 = n_28940 & ~n_28942;
assign n_28956 = n_28941 ^ n_28943;
assign n_28957 = n_28931 ^ n_28944;
assign n_28958 = ~n_28944 & n_28945;
assign n_28959 = n_28947 ^ n_28223;
assign n_28960 = n_28947 ^ n_28126;
assign n_28961 = n_28224 & ~n_28948;
assign n_28962 = ~n_28946 & ~n_28949;
assign n_28963 = n_28950 ^ n_28934;
assign n_28964 = n_28951 ^ x81;
assign n_28965 = n_28952 & ~n_28924;
assign n_28966 = n_28924 ^ n_28952;
assign n_28967 = ~n_27931 & ~n_28953;
assign n_28968 = n_28815 ^ n_28953;
assign n_28969 = n_28955 ^ n_28500;
assign n_28970 = ~n_28956 & ~n_28954;
assign n_28971 = n_28956 ^ n_27331;
assign n_28972 = ~n_28957 & ~n_28932;
assign n_28973 = n_28932 ^ n_28957;
assign n_28974 = n_28958 ^ x13;
assign n_28975 = n_28959 ^ n_26988;
assign n_28976 = n_28961 ^ n_27891;
assign n_28977 = n_28962 ^ n_26968;
assign n_28978 = n_28963 ^ x80;
assign n_28979 = n_28964 ^ n_28963;
assign n_28980 = n_28966 ^ n_28544;
assign n_28981 = n_28967 ^ n_28500;
assign n_28982 = n_28969 ^ n_28966;
assign n_28983 = n_28970 ^ n_27331;
assign n_28984 = n_28971 ^ x12;
assign n_28985 = n_28974 ^ n_28971;
assign n_28986 = n_28976 ^ n_28262;
assign n_28987 = n_28976 ^ n_28249;
assign n_28988 = n_28977 ^ n_28959;
assign n_28989 = n_28964 ^ n_28978;
assign n_28990 = ~n_28978 & n_28979;
assign n_28991 = n_28969 ^ n_28980;
assign n_28992 = n_28981 ^ n_27349;
assign n_28993 = ~n_28980 & n_28982;
assign n_28994 = n_28983 ^ n_28981;
assign n_28995 = n_28974 ^ n_28984;
assign n_28996 = n_28984 & ~n_28985;
assign n_28997 = n_28986 ^ n_28261;
assign n_28998 = n_28184 ^ n_28986;
assign n_28999 = ~n_28262 & ~n_28987;
assign n_29000 = n_28988 & n_28975;
assign n_29001 = n_28988 ^ n_26988;
assign n_29002 = n_28989 & ~n_28965;
assign n_29003 = n_28965 ^ n_28989;
assign n_29004 = n_28990 ^ x80;
assign n_29005 = ~n_27941 & n_28991;
assign n_29006 = n_28856 ^ n_28991;
assign n_29007 = n_28983 ^ n_28992;
assign n_29008 = n_28993 ^ n_28544;
assign n_29009 = n_28992 & n_28994;
assign n_29010 = n_28995 & n_28972;
assign n_29011 = n_28972 ^ n_28995;
assign n_29012 = n_28996 ^ x12;
assign n_29013 = n_28997 ^ n_27015;
assign n_29014 = n_28999 ^ n_27910;
assign n_29015 = n_29000 ^ n_26988;
assign n_29016 = n_29001 ^ x95;
assign n_29017 = n_29003 ^ n_28580;
assign n_29018 = n_29004 ^ n_29001;
assign n_29019 = n_29005 ^ n_28544;
assign n_29020 = n_29007 ^ x11;
assign n_29021 = n_29008 ^ n_29003;
assign n_29022 = n_29009 ^ n_27349;
assign n_29023 = n_29012 ^ n_29007;
assign n_29024 = n_29014 ^ n_28313;
assign n_29025 = n_29014 ^ n_28300;
assign n_29026 = n_29015 ^ n_28997;
assign n_29027 = n_29004 ^ n_29016;
assign n_29028 = ~n_29016 & n_29018;
assign n_29029 = n_29019 ^ n_27366;
assign n_29030 = n_29012 ^ n_29020;
assign n_29031 = ~n_29021 & ~n_29017;
assign n_29032 = n_29021 ^ n_28580;
assign n_29033 = n_29022 ^ n_29019;
assign n_29034 = n_29020 & ~n_29023;
assign n_29035 = n_29024 ^ n_28286;
assign n_29036 = n_29024 ^ n_28233;
assign n_29037 = ~n_28313 & n_29025;
assign n_29038 = ~n_29026 & n_29013;
assign n_29039 = n_29026 ^ n_27015;
assign n_29040 = ~n_29027 & ~n_29002;
assign n_29041 = n_29002 ^ n_29027;
assign n_29042 = n_29028 ^ x95;
assign n_29043 = n_29022 ^ n_29029;
assign n_29044 = n_29010 & n_29030;
assign n_29045 = n_29030 ^ n_29010;
assign n_29046 = n_29031 ^ n_28580;
assign n_29047 = ~n_27959 & n_29032;
assign n_29048 = n_28893 ^ n_29032;
assign n_29049 = n_29029 & ~n_29033;
assign n_29050 = n_29034 ^ x11;
assign n_29051 = n_29035 ^ n_27035;
assign n_29052 = n_29037 ^ n_27928;
assign n_29053 = n_29038 ^ n_27015;
assign n_29054 = n_29039 ^ x94;
assign n_29055 = n_29041 ^ n_28615;
assign n_29056 = n_29042 ^ n_29039;
assign n_29057 = n_29043 ^ x10;
assign n_29058 = n_29046 ^ n_29041;
assign n_29059 = n_29047 ^ n_28580;
assign n_29060 = n_29049 ^ n_27366;
assign n_29061 = n_29050 ^ n_29043;
assign n_29062 = n_29052 ^ n_28339;
assign n_29063 = n_29052 ^ n_28325;
assign n_29064 = n_29053 ^ n_29035;
assign n_29065 = n_29042 ^ n_29054;
assign n_29066 = n_29046 ^ n_29055;
assign n_29067 = n_29054 & ~n_29056;
assign n_29068 = ~n_29055 & n_29058;
assign n_29069 = n_29059 ^ n_27385;
assign n_29070 = n_29060 ^ n_29059;
assign n_29071 = n_29061 & ~n_29057;
assign n_29072 = n_29061 ^ x10;
assign n_29073 = n_29062 ^ n_28338;
assign n_29074 = n_29062 ^ n_28270;
assign n_29075 = n_28339 & ~n_29063;
assign n_29076 = n_29064 ^ n_27035;
assign n_29077 = ~n_29064 & n_29051;
assign n_29078 = n_29040 & n_29065;
assign n_29079 = n_29065 ^ n_29040;
assign n_29080 = ~n_27984 & ~n_29066;
assign n_29081 = n_28933 ^ n_29066;
assign n_29082 = n_29067 ^ x94;
assign n_29083 = n_29068 ^ n_28615;
assign n_29084 = n_29060 ^ n_29069;
assign n_29085 = ~n_29069 & n_29070;
assign n_29086 = n_29071 ^ x10;
assign n_29087 = ~n_29044 & n_29072;
assign n_29088 = n_29072 ^ n_29044;
assign n_29089 = n_29073 ^ n_27052;
assign n_29090 = n_29075 ^ n_27945;
assign n_29091 = n_29076 ^ x93;
assign n_29092 = n_29077 ^ n_27035;
assign n_29093 = n_29079 ^ n_28639;
assign n_29094 = n_29080 ^ n_28615;
assign n_29095 = n_29082 ^ n_29076;
assign n_29096 = n_29082 ^ x93;
assign n_29097 = n_29083 ^ n_29079;
assign n_29098 = n_29084 ^ x9;
assign n_29099 = n_29085 ^ n_27385;
assign n_29100 = n_29086 ^ n_29084;
assign n_29101 = n_29090 ^ n_28377;
assign n_29102 = n_29090 ^ n_28364;
assign n_29103 = n_29092 ^ n_27052;
assign n_29104 = n_29092 ^ n_29073;
assign n_29105 = n_29083 ^ n_29093;
assign n_29106 = n_29094 ^ n_27405;
assign n_29107 = n_29091 & ~n_29095;
assign n_29108 = n_29096 ^ n_29076;
assign n_29109 = n_29093 & n_29097;
assign n_29110 = n_29099 ^ n_29094;
assign n_29111 = ~n_29100 & n_29098;
assign n_29112 = n_29100 ^ x9;
assign n_29113 = n_29101 ^ n_28376;
assign n_29114 = n_28307 ^ n_29101;
assign n_29115 = ~n_28377 & n_29102;
assign n_29116 = n_29103 ^ n_29073;
assign n_29117 = ~n_29089 & n_29104;
assign n_29118 = n_27996 & n_29105;
assign n_29119 = n_28973 ^ n_29105;
assign n_29120 = n_29107 ^ x93;
assign n_29121 = ~n_29108 & ~n_29078;
assign n_29122 = n_29078 ^ n_29108;
assign n_29123 = n_29109 ^ n_28639;
assign n_29124 = n_29110 & ~n_29106;
assign n_29125 = n_29110 ^ n_27405;
assign n_29126 = n_29111 ^ x9;
assign n_29127 = ~n_29087 & n_29112;
assign n_29128 = n_29112 ^ n_29087;
assign n_29129 = n_29113 ^ n_27073;
assign n_29130 = n_29115 ^ n_27964;
assign n_29131 = n_29116 ^ x92;
assign n_29132 = n_29117 ^ n_27052;
assign n_29133 = n_29118 ^ n_28639;
assign n_29134 = n_29120 ^ n_29116;
assign n_29135 = n_29122 ^ n_28687;
assign n_29136 = n_29123 ^ n_29122;
assign n_29137 = n_29124 ^ n_27405;
assign n_29138 = n_29125 ^ x8;
assign n_29139 = n_29126 ^ n_29125;
assign n_29140 = n_29130 ^ n_28430;
assign n_29141 = n_29130 ^ n_28417;
assign n_29142 = n_29132 ^ n_27073;
assign n_29143 = n_29132 ^ n_29113;
assign n_29144 = n_29133 ^ n_27424;
assign n_29145 = n_29134 ^ x92;
assign n_29146 = n_29134 & ~n_29131;
assign n_29147 = n_29123 ^ n_29135;
assign n_29148 = n_29135 & n_29136;
assign n_29149 = n_29137 ^ n_29133;
assign n_29150 = ~n_29139 & n_29138;
assign n_29151 = n_29139 ^ x8;
assign n_29152 = n_29140 ^ n_28402;
assign n_29153 = n_28344 ^ n_29140;
assign n_29154 = n_28430 & n_29141;
assign n_29155 = n_29142 ^ n_29113;
assign n_29156 = ~n_29129 & ~n_29143;
assign n_29157 = n_29137 ^ n_29144;
assign n_29158 = ~n_29145 & ~n_29121;
assign n_29159 = n_29121 ^ n_29145;
assign n_29160 = n_29146 ^ x92;
assign n_29161 = n_28018 & ~n_29147;
assign n_29162 = n_29011 ^ n_29147;
assign n_29163 = n_29148 ^ n_28687;
assign n_29164 = ~n_29144 & ~n_29149;
assign n_29165 = n_29150 ^ x8;
assign n_29166 = n_29151 & n_29127;
assign n_29167 = n_29127 ^ n_29151;
assign n_29168 = n_29152 ^ n_27089;
assign n_29169 = n_29154 ^ n_27989;
assign n_29170 = n_29155 ^ x91;
assign n_29171 = n_29156 ^ n_27073;
assign n_29172 = n_29157 ^ x23;
assign n_29173 = n_29159 ^ n_28713;
assign n_29174 = n_29160 ^ x91;
assign n_29175 = n_29160 ^ n_29155;
assign n_29176 = n_29161 ^ n_28687;
assign n_29177 = n_29163 ^ n_29159;
assign n_29178 = n_29164 ^ n_27424;
assign n_29179 = n_29165 ^ n_29157;
assign n_29180 = n_28455 ^ n_29169;
assign n_29181 = n_28443 ^ n_29169;
assign n_29182 = n_28007 ^ n_29169;
assign n_29183 = n_29171 ^ n_27089;
assign n_29184 = n_29171 ^ n_29152;
assign n_29185 = n_29174 ^ n_29155;
assign n_29186 = ~n_29170 & n_29175;
assign n_29187 = n_29176 ^ n_27443;
assign n_29188 = n_29177 & n_29173;
assign n_29189 = n_29177 ^ n_28713;
assign n_29190 = n_29178 ^ n_29176;
assign n_29191 = ~n_29179 & n_29172;
assign n_29192 = n_29179 ^ x23;
assign n_29193 = n_29180 ^ n_28441;
assign n_29194 = n_28382 ^ n_29180;
assign n_29195 = n_29181 & ~n_29182;
assign n_29196 = n_29183 ^ n_29152;
assign n_29197 = n_29168 & n_29184;
assign n_29198 = n_29158 ^ n_29185;
assign n_29199 = ~n_29185 & n_29158;
assign n_29200 = n_29186 ^ x91;
assign n_29201 = n_29178 ^ n_29187;
assign n_29202 = n_29188 ^ n_28713;
assign n_29203 = ~n_28032 & n_29189;
assign n_29204 = n_29045 ^ n_29189;
assign n_29205 = n_29187 & ~n_29190;
assign n_29206 = n_29191 ^ x23;
assign n_29207 = ~n_29166 & ~n_29192;
assign n_29208 = n_29192 ^ n_29166;
assign n_29209 = n_29193 ^ n_27108;
assign n_29210 = n_28496 ^ n_29195;
assign n_29211 = n_29196 ^ x90;
assign n_29212 = n_29197 ^ n_27089;
assign n_29213 = n_29198 ^ n_28752;
assign n_29214 = n_29200 ^ x90;
assign n_29215 = n_29196 ^ n_29200;
assign n_29216 = n_29201 ^ x22;
assign n_29217 = n_29202 ^ n_29198;
assign n_29218 = n_29203 ^ n_28713;
assign n_29219 = n_29205 ^ n_27443;
assign n_29220 = n_29206 ^ n_29201;
assign n_29221 = n_29206 ^ x22;
assign n_29222 = n_29210 ^ n_28495;
assign n_29223 = n_29210 ^ n_28411;
assign n_29224 = n_29211 ^ n_29200;
assign n_29225 = n_29212 ^ n_27108;
assign n_29226 = n_29212 ^ n_29193;
assign n_29227 = n_29202 ^ n_29213;
assign n_29228 = n_29214 & n_29215;
assign n_29229 = ~n_29213 & n_29217;
assign n_29230 = n_29218 ^ n_27462;
assign n_29231 = n_29219 ^ n_29218;
assign n_29232 = n_29219 ^ n_27462;
assign n_29233 = n_29216 & ~n_29220;
assign n_29234 = n_29221 ^ n_29201;
assign n_29235 = n_29223 ^ n_28381;
assign n_29236 = n_29224 ^ n_29199;
assign n_29237 = n_29199 & ~n_29224;
assign n_29238 = n_29225 ^ n_29193;
assign n_29239 = n_29209 & n_29226;
assign n_29240 = ~n_28051 & n_29227;
assign n_29241 = n_29088 ^ n_29227;
assign n_29242 = n_29228 ^ x90;
assign n_29243 = n_29229 ^ n_28752;
assign n_29244 = n_29230 & n_29231;
assign n_29245 = n_29232 ^ n_29218;
assign n_29246 = n_29233 ^ x22;
assign n_29247 = n_29234 & ~n_29207;
assign n_29248 = n_29207 ^ n_29234;
assign n_29249 = n_29235 ^ n_28382;
assign n_29250 = n_29236 ^ n_28791;
assign n_29251 = n_29238 ^ x89;
assign n_29252 = n_29239 ^ n_27108;
assign n_29253 = n_29240 ^ n_28752;
assign n_29254 = n_29242 ^ n_29238;
assign n_29255 = n_29243 ^ n_29236;
assign n_29256 = n_29244 ^ n_27462;
assign n_29257 = n_29245 ^ x21;
assign n_29258 = n_29246 ^ n_29245;
assign n_29259 = n_29243 ^ n_29250;
assign n_29260 = n_29252 ^ n_29222;
assign n_29261 = n_29253 ^ n_27480;
assign n_29262 = n_29254 ^ x89;
assign n_29263 = ~n_29254 & n_29251;
assign n_29264 = ~n_29250 & n_29255;
assign n_29265 = n_29256 ^ n_29253;
assign n_29266 = n_29246 ^ n_29257;
assign n_29267 = n_29257 & ~n_29258;
assign n_29268 = n_28080 & n_29259;
assign n_29269 = n_29128 ^ n_29259;
assign n_29270 = n_29260 ^ x88;
assign n_29271 = n_29256 ^ n_29261;
assign n_29272 = n_29237 ^ n_29262;
assign n_29273 = ~n_29262 & ~n_29237;
assign n_29274 = n_29263 ^ x89;
assign n_29275 = n_29264 ^ n_28791;
assign n_29276 = ~n_29261 & ~n_29265;
assign n_29277 = n_29247 & n_29266;
assign n_29278 = n_29266 ^ n_29247;
assign n_29279 = n_29267 ^ x21;
assign n_29280 = n_29268 ^ n_28791;
assign n_29281 = n_29271 ^ x20;
assign n_29282 = n_29272 ^ n_28830;
assign n_29283 = n_29274 ^ n_29273;
assign n_29284 = n_29275 ^ n_29272;
assign n_29285 = n_29276 ^ n_27480;
assign n_29286 = n_29279 ^ n_29271;
assign n_29287 = n_29280 ^ n_27498;
assign n_29288 = n_29279 ^ n_29281;
assign n_29289 = n_29283 ^ n_29270;
assign n_29290 = n_29284 & n_29282;
assign n_29291 = n_29284 ^ n_28830;
assign n_29292 = n_29285 ^ n_29280;
assign n_29293 = n_29285 ^ n_27498;
assign n_29294 = n_29281 & ~n_29286;
assign n_29295 = ~n_29288 & ~n_29277;
assign n_29296 = n_29277 ^ n_29288;
assign n_29297 = n_29289 ^ n_28880;
assign n_29298 = n_29290 ^ n_28830;
assign n_29299 = n_28116 & ~n_29291;
assign n_29300 = n_29167 ^ n_29291;
assign n_29301 = n_29287 & n_29292;
assign n_29302 = n_29293 ^ n_29280;
assign n_29303 = n_29294 ^ x20;
assign n_29304 = n_29298 ^ n_29289;
assign n_29305 = n_29299 ^ n_28830;
assign n_29306 = n_29301 ^ n_27498;
assign n_29307 = n_29302 ^ x19;
assign n_29308 = n_29303 ^ n_29302;
assign n_29309 = n_29303 ^ x19;
assign n_29310 = n_29304 & ~n_29297;
assign n_29311 = n_29304 ^ n_28880;
assign n_29312 = n_29305 ^ n_27519;
assign n_29313 = n_29306 ^ n_29305;
assign n_29314 = n_29307 & ~n_29308;
assign n_29315 = n_29309 ^ n_29302;
assign n_29316 = n_29310 ^ n_28880;
assign n_29317 = n_28152 & ~n_29311;
assign n_29318 = n_29208 ^ n_29311;
assign n_29319 = n_29306 ^ n_29312;
assign n_29320 = ~n_29312 & n_29313;
assign n_29321 = n_29314 ^ x19;
assign n_29322 = ~n_29295 & n_29315;
assign n_29323 = n_29315 ^ n_29295;
assign n_29324 = n_29316 ^ n_28919;
assign n_29325 = n_29316 ^ n_28935;
assign n_29326 = n_29317 ^ n_28880;
assign n_29327 = n_29319 ^ x18;
assign n_29328 = n_29320 ^ n_27519;
assign n_29329 = n_29321 ^ n_29319;
assign n_29330 = n_29321 ^ x18;
assign n_29331 = n_28935 & n_29324;
assign n_29332 = n_28176 & n_29325;
assign n_29333 = n_29248 ^ n_29325;
assign n_29334 = n_29326 ^ n_27532;
assign n_29335 = n_29328 ^ n_29326;
assign n_29336 = n_29328 ^ n_27532;
assign n_29337 = n_29327 & ~n_29329;
assign n_29338 = n_29330 ^ n_29319;
assign n_29339 = n_29331 ^ n_28068;
assign n_29340 = n_29332 ^ n_28919;
assign n_29341 = ~n_29334 & n_29335;
assign n_29342 = n_29336 ^ n_29326;
assign n_29343 = n_29337 ^ x18;
assign n_29344 = ~n_29322 & ~n_29338;
assign n_29345 = n_29338 ^ n_29322;
assign n_29346 = n_29339 ^ n_28960;
assign n_29347 = n_29339 ^ n_28947;
assign n_29348 = n_29340 ^ n_27551;
assign n_29349 = n_29341 ^ n_27532;
assign n_29350 = n_29342 ^ x17;
assign n_29351 = n_29343 ^ n_29342;
assign n_29352 = n_28210 & ~n_29346;
assign n_29353 = n_29278 ^ n_29346;
assign n_29354 = n_28960 & ~n_29347;
assign n_29355 = n_29349 ^ n_29340;
assign n_29356 = n_29349 ^ n_29348;
assign n_29357 = n_29343 ^ n_29350;
assign n_29358 = n_29350 & ~n_29351;
assign n_29359 = n_29352 ^ n_28947;
assign n_29360 = n_29354 ^ n_28126;
assign n_29361 = ~n_29348 & ~n_29355;
assign n_29362 = n_29356 ^ x16;
assign n_29363 = ~n_29344 & n_29357;
assign n_29364 = n_29357 ^ n_29344;
assign n_29365 = n_29358 ^ x17;
assign n_29366 = n_29359 ^ n_27583;
assign n_29367 = n_29360 ^ n_28986;
assign n_29368 = n_29361 ^ n_27551;
assign n_29369 = n_29365 ^ n_29356;
assign n_29370 = n_29365 ^ x16;
assign n_29371 = n_28184 ^ n_29367;
assign n_29372 = n_29367 & ~n_28998;
assign n_29373 = n_29368 ^ n_29359;
assign n_29374 = n_29368 ^ n_27583;
assign n_29375 = n_29362 & ~n_29369;
assign n_29376 = n_29370 ^ n_29356;
assign n_29377 = n_28249 & n_29371;
assign n_29378 = n_29296 ^ n_29371;
assign n_29379 = n_29372 ^ n_28184;
assign n_29380 = ~n_29366 & n_29373;
assign n_29381 = n_29374 ^ n_29359;
assign n_29382 = n_29375 ^ x16;
assign n_29383 = n_29376 & n_29363;
assign n_29384 = n_29363 ^ n_29376;
assign n_29385 = n_29377 ^ n_28986;
assign n_29386 = n_29379 ^ n_29036;
assign n_29387 = n_29379 ^ n_29024;
assign n_29388 = n_29380 ^ n_27583;
assign n_29389 = n_29381 ^ x31;
assign n_29390 = n_29382 ^ n_29381;
assign n_29391 = n_29385 ^ n_27607;
assign n_29392 = n_28300 & n_29386;
assign n_29393 = n_29323 ^ n_29386;
assign n_29394 = ~n_29036 & ~n_29387;
assign n_29395 = n_29388 ^ n_29385;
assign n_29396 = n_29390 & ~n_29389;
assign n_29397 = n_29390 ^ x31;
assign n_29398 = n_29388 ^ n_29391;
assign n_29399 = n_29392 ^ n_29024;
assign n_29400 = n_29394 ^ n_28233;
assign n_29401 = ~n_29391 & ~n_29395;
assign n_29402 = n_29396 ^ x31;
assign n_29403 = n_29383 & ~n_29397;
assign n_29404 = n_29397 ^ n_29383;
assign n_29405 = n_29398 ^ x30;
assign n_29406 = n_29399 ^ n_27640;
assign n_29407 = n_29400 ^ n_29074;
assign n_29408 = n_29400 ^ n_29062;
assign n_29409 = n_29401 ^ n_27607;
assign n_29410 = n_29402 ^ n_29398;
assign n_29411 = n_29402 ^ n_29405;
assign n_29412 = ~n_28325 & n_29407;
assign n_29413 = n_29345 ^ n_29407;
assign n_29414 = n_29074 & ~n_29408;
assign n_29415 = n_29409 ^ n_27640;
assign n_29416 = n_29409 ^ n_29399;
assign n_29417 = ~n_29405 & n_29410;
assign n_29418 = n_29403 & ~n_29411;
assign n_29419 = n_29411 ^ n_29403;
assign n_29420 = n_29412 ^ n_29062;
assign n_29421 = n_29414 ^ n_28270;
assign n_29422 = n_29415 ^ n_29399;
assign n_29423 = ~n_29406 & ~n_29416;
assign n_29424 = n_29417 ^ x30;
assign n_29425 = n_29420 ^ n_27663;
assign n_29426 = n_29421 ^ n_29101;
assign n_29427 = n_29422 ^ x29;
assign n_29428 = n_29423 ^ n_27640;
assign n_29429 = n_29424 ^ n_29422;
assign n_29430 = n_28307 ^ n_29426;
assign n_29431 = n_29426 & ~n_29114;
assign n_29432 = n_29424 ^ n_29427;
assign n_29433 = n_29428 ^ n_29420;
assign n_29434 = n_29427 & ~n_29429;
assign n_29435 = n_28364 & ~n_29430;
assign n_29436 = n_29364 ^ n_29430;
assign n_29437 = n_29431 ^ n_28307;
assign n_29438 = n_29432 ^ n_29418;
assign n_29439 = ~n_29418 & ~n_29432;
assign n_29440 = n_29433 ^ n_27663;
assign n_29441 = ~n_29433 & ~n_29425;
assign n_29442 = n_29434 ^ x29;
assign n_29443 = n_29435 ^ n_29101;
assign n_29444 = n_29437 ^ n_29140;
assign n_29445 = ~n_28478 & ~n_29438;
assign n_29446 = n_29438 ^ n_28478;
assign n_29447 = n_29438 ^ n_28464;
assign n_29448 = n_29440 ^ x28;
assign n_29449 = n_29441 ^ n_27663;
assign n_29450 = n_29442 ^ n_29440;
assign n_29451 = n_29443 ^ n_27698;
assign n_29452 = n_28344 ^ n_29444;
assign n_29453 = ~n_29444 & ~n_29153;
assign n_29454 = n_29445 ^ n_28537;
assign n_29455 = n_28069 & ~n_29446;
assign n_29456 = n_29442 ^ n_29448;
assign n_29457 = n_29449 ^ n_27698;
assign n_29458 = n_29449 ^ n_29443;
assign n_29459 = ~n_29448 & n_29450;
assign n_29460 = n_28417 & ~n_29452;
assign n_29461 = n_29384 ^ n_29452;
assign n_29462 = n_29453 ^ n_28344;
assign n_29463 = n_29455 ^ n_28478;
assign n_29464 = n_28479 ^ n_29455;
assign n_29465 = n_29456 ^ n_29439;
assign n_29466 = ~n_29439 & ~n_29456;
assign n_29467 = n_29457 ^ n_29443;
assign n_29468 = ~n_29451 & ~n_29458;
assign n_29469 = n_29459 ^ x28;
assign n_29470 = n_29460 ^ n_29140;
assign n_29471 = n_29194 ^ n_29462;
assign n_29472 = n_29462 ^ n_29180;
assign n_29473 = n_28382 ^ n_29462;
assign n_29474 = ~n_27577 & n_29463;
assign n_29475 = x231 & ~n_29464;
assign n_29476 = n_29464 ^ x231;
assign n_29477 = n_29465 ^ n_29445;
assign n_29478 = n_29465 ^ n_29454;
assign n_29479 = n_29467 ^ x27;
assign n_29480 = n_29468 ^ n_27698;
assign n_29481 = n_29469 ^ n_29467;
assign n_29482 = n_29470 ^ n_27747;
assign n_29483 = ~n_28443 & ~n_29471;
assign n_29484 = n_29404 ^ n_29471;
assign n_29485 = ~n_29472 & n_29473;
assign n_29486 = n_29474 ^ n_27598;
assign n_29487 = n_29454 & ~n_29477;
assign n_29488 = n_28085 & ~n_29478;
assign n_29489 = n_29480 ^ n_29470;
assign n_29490 = n_29481 ^ x27;
assign n_29491 = ~n_29481 & n_29479;
assign n_29492 = n_29480 ^ n_29482;
assign n_29493 = n_29483 ^ n_29180;
assign n_29494 = n_29249 ^ n_29485;
assign n_29495 = n_29487 ^ n_28537;
assign n_29496 = n_29488 ^ n_28537;
assign n_29497 = ~n_29482 & ~n_29489;
assign n_29498 = n_29490 ^ n_29466;
assign n_29499 = ~n_29466 & ~n_29490;
assign n_29500 = n_29491 ^ x27;
assign n_29501 = n_29492 ^ x26;
assign n_29502 = n_29493 ^ n_27773;
assign n_29503 = ~n_28467 & n_29494;
assign n_29504 = n_29419 ^ n_29494;
assign n_29505 = n_29495 ^ n_28575;
assign n_29506 = n_29496 ^ n_29474;
assign n_29507 = n_29496 ^ n_29486;
assign n_29508 = n_29497 ^ n_27747;
assign n_29509 = n_29498 ^ n_28575;
assign n_29510 = n_29495 ^ n_29498;
assign n_29511 = n_29500 ^ n_29492;
assign n_29512 = n_29500 ^ n_29501;
assign n_29513 = n_29503 ^ n_29210;
assign n_29514 = n_29505 ^ n_29498;
assign n_29515 = n_29486 & n_29506;
assign n_29516 = n_29507 ^ x230;
assign n_29517 = n_29475 ^ n_29507;
assign n_29518 = n_29508 ^ n_27773;
assign n_29519 = n_29508 ^ n_29493;
assign n_29520 = ~n_29509 & n_29510;
assign n_29521 = ~n_29501 & n_29511;
assign n_29522 = n_29512 ^ n_29499;
assign n_29523 = n_29499 & n_29512;
assign n_29524 = n_29513 ^ n_27812;
assign n_29525 = ~n_28122 & n_29514;
assign n_29526 = n_29515 ^ n_27598;
assign n_29527 = n_29475 ^ n_29516;
assign n_29528 = ~n_29516 & n_29517;
assign n_29529 = n_29518 ^ n_29493;
assign n_29530 = ~n_29502 & ~n_29519;
assign n_29531 = n_29520 ^ n_28575;
assign n_29532 = n_29521 ^ x26;
assign n_29533 = n_29522 ^ n_28612;
assign n_29534 = n_29525 ^ n_28575;
assign n_29535 = n_29526 ^ n_27634;
assign n_29536 = n_29527 & n_29476;
assign n_29537 = n_29476 ^ n_29527;
assign n_29538 = n_29528 ^ x230;
assign n_29539 = n_29529 ^ x25;
assign n_29540 = n_29530 ^ n_27773;
assign n_29541 = n_29531 ^ n_29522;
assign n_29542 = n_29532 ^ n_29529;
assign n_29543 = n_29531 ^ n_29533;
assign n_29544 = n_29534 ^ n_27634;
assign n_29545 = n_29526 ^ n_29534;
assign n_29546 = n_29535 ^ n_29534;
assign n_29547 = n_29538 ^ x229;
assign n_29548 = n_29532 ^ n_29539;
assign n_29549 = n_29540 ^ n_29524;
assign n_29550 = n_29533 & n_29541;
assign n_29551 = n_29539 & ~n_29542;
assign n_29552 = ~n_28156 & ~n_29543;
assign n_29553 = ~n_29544 & n_29545;
assign n_29554 = n_29546 ^ n_29538;
assign n_29555 = n_29546 ^ n_29547;
assign n_29556 = n_29523 ^ n_29548;
assign n_29557 = ~n_29548 & n_29523;
assign n_29558 = n_29550 ^ n_28612;
assign n_29559 = n_29551 ^ x25;
assign n_29560 = n_29552 ^ n_28612;
assign n_29561 = n_29553 ^ n_27634;
assign n_29562 = n_29547 & n_29554;
assign n_29563 = n_29536 & n_29555;
assign n_29564 = n_29555 ^ n_29536;
assign n_29565 = n_29556 ^ n_28647;
assign n_29566 = n_29558 ^ n_29556;
assign n_29567 = n_29559 ^ n_29549;
assign n_29568 = n_29560 ^ n_27668;
assign n_29569 = n_29561 ^ n_27668;
assign n_29570 = n_29561 ^ n_29560;
assign n_29571 = n_29562 ^ x229;
assign n_29572 = n_29558 ^ n_29565;
assign n_29573 = n_29565 & n_29566;
assign n_29574 = n_29567 ^ x24;
assign n_29575 = n_29569 ^ n_29560;
assign n_29576 = n_29568 & ~n_29570;
assign n_29577 = ~n_28193 & n_29572;
assign n_29578 = n_29573 ^ n_28647;
assign n_29579 = n_29557 ^ n_29574;
assign n_29580 = n_29575 ^ x228;
assign n_29581 = n_29571 ^ n_29575;
assign n_29582 = n_29576 ^ n_27668;
assign n_29583 = n_29577 ^ n_28647;
assign n_29584 = n_29578 ^ n_28675;
assign n_29585 = n_29579 ^ n_28675;
assign n_29586 = n_29578 ^ n_29579;
assign n_29587 = n_29571 ^ n_29580;
assign n_29588 = n_29580 & ~n_29581;
assign n_29589 = n_29583 ^ n_27706;
assign n_29590 = n_29582 ^ n_29583;
assign n_29591 = n_29584 ^ n_29579;
assign n_29592 = n_29585 & ~n_29586;
assign n_29593 = n_29587 & ~n_29563;
assign n_29594 = n_29563 ^ n_29587;
assign n_29595 = n_29588 ^ x228;
assign n_29596 = n_29582 ^ n_29589;
assign n_29597 = ~n_29589 & n_29590;
assign n_29598 = ~n_28228 & ~n_29591;
assign n_29599 = n_29592 ^ n_28675;
assign n_29600 = n_29595 ^ n_29596;
assign n_29601 = n_29596 ^ x227;
assign n_29602 = n_29597 ^ n_27706;
assign n_29603 = n_29598 ^ n_28675;
assign n_29604 = n_29599 ^ n_28522;
assign n_29605 = n_29599 ^ n_28721;
assign n_29606 = n_29600 ^ x227;
assign n_29607 = n_29600 & ~n_29601;
assign n_29608 = n_29603 ^ n_27742;
assign n_29609 = n_29602 ^ n_29603;
assign n_29610 = n_29604 ^ n_28721;
assign n_29611 = n_28734 & n_29605;
assign n_29612 = ~n_29593 & n_29606;
assign n_29613 = n_29606 ^ n_29593;
assign n_29614 = n_29607 ^ x227;
assign n_29615 = n_29602 ^ n_29608;
assign n_29616 = ~n_29608 & n_29609;
assign n_29617 = n_28264 & ~n_29610;
assign n_29618 = n_29611 ^ n_28522;
assign n_29619 = n_29614 ^ n_29615;
assign n_29620 = n_29615 ^ x226;
assign n_29621 = n_29616 ^ n_27742;
assign n_29622 = n_29617 ^ n_28721;
assign n_29623 = n_29618 ^ n_28773;
assign n_29624 = n_29618 ^ n_28758;
assign n_29625 = n_29619 ^ x226;
assign n_29626 = n_29619 & ~n_29620;
assign n_29627 = n_29622 ^ n_27775;
assign n_29628 = n_29621 ^ n_29622;
assign n_29629 = n_28309 & ~n_29623;
assign n_29630 = ~n_28773 & ~n_29624;
assign n_29631 = ~n_29625 & ~n_29612;
assign n_29632 = n_29612 ^ n_29625;
assign n_29633 = n_29626 ^ x226;
assign n_29634 = n_29621 ^ n_29627;
assign n_29635 = ~n_29627 & ~n_29628;
assign n_29636 = n_29629 ^ n_28758;
assign n_29637 = n_29630 ^ n_28597;
assign n_29638 = n_29634 ^ x225;
assign n_29639 = n_29633 ^ n_29634;
assign n_29640 = n_29635 ^ n_27775;
assign n_29641 = n_29636 ^ n_27819;
assign n_29642 = n_29637 ^ n_28794;
assign n_29643 = n_29633 ^ n_29638;
assign n_29644 = ~n_29638 & n_29639;
assign n_29645 = n_29640 ^ n_27819;
assign n_29646 = n_29640 ^ n_29636;
assign n_29647 = n_29642 ^ n_28644;
assign n_29648 = ~n_29642 & n_28807;
assign n_29649 = ~n_29643 & n_29631;
assign n_29650 = n_29631 ^ n_29643;
assign n_29651 = n_29644 ^ x225;
assign n_29652 = n_29645 ^ n_29636;
assign n_29653 = n_29641 & n_29646;
assign n_29654 = n_28350 & ~n_29647;
assign n_29655 = n_29648 ^ n_28644;
assign n_29656 = n_29651 ^ n_29652;
assign n_29657 = n_29652 ^ x224;
assign n_29658 = n_29653 ^ n_27819;
assign n_29659 = n_29654 ^ n_28794;
assign n_29660 = n_29655 ^ n_28695;
assign n_29661 = n_29655 ^ n_28837;
assign n_29662 = n_29656 ^ x224;
assign n_29663 = n_29656 & ~n_29657;
assign n_29664 = n_29658 ^ n_29659;
assign n_29665 = n_29659 ^ n_27849;
assign n_29666 = n_29660 ^ n_28837;
assign n_29667 = n_28850 & ~n_29661;
assign n_29668 = ~n_29649 & n_29662;
assign n_29669 = n_29662 ^ n_29649;
assign n_29670 = n_29663 ^ x224;
assign n_29671 = n_29664 ^ n_27849;
assign n_29672 = n_29664 & ~n_29665;
assign n_29673 = n_28385 & ~n_29666;
assign n_29674 = n_29667 ^ n_28695;
assign n_29675 = n_29671 ^ x239;
assign n_29676 = n_29670 ^ n_29671;
assign n_29677 = n_29672 ^ n_27849;
assign n_29678 = n_29673 ^ n_28837;
assign n_29679 = n_28738 ^ n_29674;
assign n_29680 = n_29674 ^ n_28874;
assign n_29681 = n_29670 ^ n_29675;
assign n_29682 = ~n_29675 & n_29676;
assign n_29683 = n_29677 ^ n_27873;
assign n_29684 = n_29678 ^ n_27873;
assign n_29685 = n_29677 ^ n_29678;
assign n_29686 = n_29679 ^ n_28874;
assign n_29687 = ~n_28888 & ~n_29680;
assign n_29688 = n_29668 & n_29681;
assign n_29689 = n_29681 ^ n_29668;
assign n_29690 = n_29682 ^ x239;
assign n_29691 = n_29683 ^ n_29678;
assign n_29692 = ~n_29684 & n_29685;
assign n_29693 = n_28422 & n_29686;
assign n_29694 = n_29476 ^ n_29686;
assign n_29695 = n_29687 ^ n_28738;
assign n_29696 = n_29691 ^ x238;
assign n_29697 = n_29690 ^ n_29691;
assign n_29698 = n_29692 ^ n_27873;
assign n_29699 = n_29693 ^ n_28874;
assign n_29700 = n_29695 ^ n_28912;
assign n_29701 = n_28927 ^ n_29695;
assign n_29702 = n_29690 ^ n_29696;
assign n_29703 = ~n_29696 & n_29697;
assign n_29704 = n_29698 ^ n_29699;
assign n_29705 = n_29699 ^ n_27895;
assign n_29706 = n_28927 & n_29700;
assign n_29707 = n_29537 ^ n_29701;
assign n_29708 = n_28461 & n_29701;
assign n_29709 = n_29688 & n_29702;
assign n_29710 = n_29702 ^ n_29688;
assign n_29711 = n_29703 ^ x238;
assign n_29712 = n_29704 ^ n_27895;
assign n_29713 = n_29704 & ~n_29705;
assign n_29714 = n_29706 ^ n_28778;
assign n_29715 = n_29708 ^ n_28912;
assign n_29716 = n_29712 ^ x237;
assign n_29717 = n_29711 ^ n_29712;
assign n_29718 = n_29713 ^ n_27895;
assign n_29719 = n_29714 ^ n_28953;
assign n_29720 = n_29715 ^ n_27914;
assign n_29721 = n_29711 ^ n_29716;
assign n_29722 = ~n_29716 & n_29717;
assign n_29723 = n_29715 ^ n_29718;
assign n_29724 = ~n_29719 & n_28968;
assign n_29725 = n_28815 ^ n_29719;
assign n_29726 = n_29720 ^ n_29718;
assign n_29727 = n_29709 ^ n_29721;
assign n_29728 = n_29721 & n_29709;
assign n_29729 = n_29722 ^ x237;
assign n_29730 = ~n_29720 & n_29723;
assign n_29731 = n_29724 ^ n_28815;
assign n_29732 = n_29564 ^ n_29725;
assign n_29733 = n_28500 & ~n_29725;
assign n_29734 = n_29726 ^ x236;
assign n_29735 = n_29729 ^ n_29726;
assign n_29736 = n_29730 ^ n_27914;
assign n_29737 = n_29731 ^ n_28991;
assign n_29738 = n_29731 ^ n_29006;
assign n_29739 = n_29733 ^ n_28953;
assign n_29740 = n_29735 & ~n_29734;
assign n_29741 = n_29735 ^ x236;
assign n_29742 = n_29736 ^ n_27931;
assign n_29743 = n_29006 & n_29737;
assign n_29744 = n_29594 ^ n_29738;
assign n_29745 = n_28544 & ~n_29738;
assign n_29746 = n_29739 ^ n_27931;
assign n_29747 = n_29739 ^ n_29736;
assign n_29748 = n_29740 ^ x236;
assign n_29749 = n_29741 & n_29728;
assign n_29750 = n_29728 ^ n_29741;
assign n_29751 = n_29739 ^ n_29742;
assign n_29752 = n_29743 ^ n_28856;
assign n_29753 = n_29745 ^ n_28991;
assign n_29754 = n_29746 & n_29747;
assign n_29755 = n_29748 ^ n_29751;
assign n_29756 = n_29751 ^ x235;
assign n_29757 = n_29752 ^ n_29032;
assign n_29758 = n_29753 ^ n_27941;
assign n_29759 = n_29754 ^ n_27931;
assign n_29760 = n_29755 ^ x235;
assign n_29761 = ~n_29755 & n_29756;
assign n_29762 = ~n_29757 & ~n_29048;
assign n_29763 = n_28893 ^ n_29757;
assign n_29764 = n_29759 ^ n_29753;
assign n_29765 = n_29749 & ~n_29760;
assign n_29766 = n_29760 ^ n_29749;
assign n_29767 = n_29761 ^ x235;
assign n_29768 = n_29762 ^ n_28893;
assign n_29769 = n_29613 ^ n_29763;
assign n_29770 = ~n_28580 & ~n_29763;
assign n_29771 = n_29764 & ~n_29758;
assign n_29772 = n_29764 ^ n_27941;
assign n_29773 = n_29767 ^ x234;
assign n_29774 = n_29768 ^ n_29066;
assign n_29775 = n_29768 ^ n_29081;
assign n_29776 = n_29770 ^ n_29032;
assign n_29777 = n_29771 ^ n_27941;
assign n_29778 = n_29772 ^ n_29767;
assign n_29779 = n_29772 ^ x234;
assign n_29780 = ~n_29081 & ~n_29774;
assign n_29781 = n_29632 ^ n_29775;
assign n_29782 = ~n_28615 & n_29775;
assign n_29783 = n_29776 ^ n_27959;
assign n_29784 = n_29777 ^ n_29776;
assign n_29785 = n_29773 & ~n_29778;
assign n_29786 = n_29779 ^ n_29767;
assign n_29787 = n_29780 ^ n_28933;
assign n_29788 = n_29782 ^ n_29066;
assign n_29789 = n_29777 ^ n_29783;
assign n_29790 = ~n_29783 & n_29784;
assign n_29791 = n_29785 ^ x234;
assign n_29792 = ~n_29786 & n_29765;
assign n_29793 = n_29765 ^ n_29786;
assign n_29794 = n_29787 ^ n_29105;
assign n_29795 = n_29787 ^ n_28973;
assign n_29796 = n_29788 ^ n_27984;
assign n_29797 = n_29789 ^ x233;
assign n_29798 = n_29790 ^ n_27959;
assign n_29799 = n_29791 ^ n_29789;
assign n_29800 = n_29791 ^ x233;
assign n_29801 = ~n_29119 & ~n_29794;
assign n_29802 = n_29795 ^ n_29105;
assign n_29803 = n_29798 ^ n_29788;
assign n_29804 = n_29798 ^ n_29796;
assign n_29805 = n_29797 & ~n_29799;
assign n_29806 = n_29800 ^ n_29789;
assign n_29807 = n_29801 ^ n_28973;
assign n_29808 = n_28639 & ~n_29802;
assign n_29809 = n_29650 ^ n_29802;
assign n_29810 = n_29796 & ~n_29803;
assign n_29811 = n_29804 ^ x232;
assign n_29812 = n_29805 ^ x233;
assign n_29813 = n_29792 & ~n_29806;
assign n_29814 = n_29806 ^ n_29792;
assign n_29815 = n_29807 ^ n_29147;
assign n_29816 = n_29807 ^ n_29162;
assign n_29817 = n_29808 ^ n_29105;
assign n_29818 = n_29810 ^ n_27984;
assign n_29819 = n_29812 ^ n_29804;
assign n_29820 = n_29812 ^ x232;
assign n_29821 = n_29162 & ~n_29815;
assign n_29822 = n_29669 ^ n_29816;
assign n_29823 = ~n_28687 & ~n_29816;
assign n_29824 = n_29817 ^ n_27996;
assign n_29825 = n_29818 ^ n_29817;
assign n_29826 = n_29818 ^ n_27996;
assign n_29827 = ~n_29811 & n_29819;
assign n_29828 = n_29820 ^ n_29804;
assign n_29829 = n_29821 ^ n_29011;
assign n_29830 = n_29823 ^ n_29147;
assign n_29831 = n_29824 & n_29825;
assign n_29832 = n_29826 ^ n_29817;
assign n_29833 = n_29827 ^ x232;
assign n_29834 = n_29813 & n_29828;
assign n_29835 = n_29828 ^ n_29813;
assign n_29836 = n_29829 ^ n_29189;
assign n_29837 = n_29829 ^ n_29204;
assign n_29838 = n_29830 ^ n_28018;
assign n_29839 = n_29831 ^ n_27996;
assign n_29840 = n_29832 ^ x247;
assign n_29841 = n_29833 ^ n_29832;
assign n_29842 = ~n_29204 & n_29836;
assign n_29843 = n_29837 ^ n_29689;
assign n_29844 = n_28713 & n_29837;
assign n_29845 = n_29839 ^ n_29830;
assign n_29846 = n_29839 ^ n_29838;
assign n_29847 = n_29841 & ~n_29840;
assign n_29848 = n_29841 ^ x247;
assign n_29849 = n_29842 ^ n_29045;
assign n_29850 = n_29844 ^ n_29189;
assign n_29851 = ~n_29838 & n_29845;
assign n_29852 = n_29846 ^ x246;
assign n_29853 = n_29847 ^ x247;
assign n_29854 = ~n_29834 & ~n_29848;
assign n_29855 = n_29848 ^ n_29834;
assign n_29856 = n_29849 ^ n_29241;
assign n_29857 = n_29849 ^ n_29227;
assign n_29858 = n_29850 ^ n_28032;
assign n_29859 = n_29851 ^ n_28018;
assign n_29860 = n_29853 ^ n_29846;
assign n_29861 = n_29853 ^ n_29852;
assign n_29862 = n_29856 ^ n_29710;
assign n_29863 = n_28752 & n_29856;
assign n_29864 = ~n_29241 & n_29857;
assign n_29865 = n_29859 ^ n_29850;
assign n_29866 = ~n_29852 & n_29860;
assign n_29867 = ~n_29854 & n_29861;
assign n_29868 = n_29861 ^ n_29854;
assign n_29869 = n_29863 ^ n_29227;
assign n_29870 = n_29864 ^ n_29088;
assign n_29871 = ~n_29865 & ~n_29858;
assign n_29872 = n_29865 ^ n_28032;
assign n_29873 = n_29866 ^ x246;
assign n_29874 = n_29869 ^ n_28051;
assign n_29875 = n_29870 ^ n_29259;
assign n_29876 = n_29870 ^ n_29269;
assign n_29877 = n_29871 ^ n_28032;
assign n_29878 = n_29872 ^ x245;
assign n_29879 = n_29873 ^ n_29872;
assign n_29880 = n_29269 & n_29875;
assign n_29881 = n_28791 & ~n_29876;
assign n_29882 = n_29727 ^ n_29876;
assign n_29883 = n_29877 ^ n_29869;
assign n_29884 = n_29877 ^ n_28051;
assign n_29885 = n_29879 & ~n_29878;
assign n_29886 = n_29879 ^ x245;
assign n_29887 = n_29880 ^ n_29128;
assign n_29888 = n_29881 ^ n_29259;
assign n_29889 = ~n_29874 & n_29883;
assign n_29890 = n_29884 ^ n_29869;
assign n_29891 = n_29885 ^ x245;
assign n_29892 = ~n_29867 & ~n_29886;
assign n_29893 = n_29886 ^ n_29867;
assign n_29894 = n_29887 ^ n_29291;
assign n_29895 = n_29888 ^ n_28080;
assign n_29896 = n_29889 ^ n_28051;
assign n_29897 = n_29890 ^ x244;
assign n_29898 = n_29891 ^ n_29890;
assign n_29899 = n_29894 & n_29300;
assign n_29900 = n_29167 ^ n_29894;
assign n_29901 = n_29896 ^ n_29888;
assign n_29902 = n_29891 ^ n_29897;
assign n_29903 = n_29897 & ~n_29898;
assign n_29904 = n_29899 ^ n_29167;
assign n_29905 = ~n_28830 & n_29900;
assign n_29906 = n_29900 ^ n_29750;
assign n_29907 = n_29901 & n_29895;
assign n_29908 = n_29901 ^ n_28080;
assign n_29909 = ~n_29892 & ~n_29902;
assign n_29910 = n_29902 ^ n_29892;
assign n_29911 = n_29903 ^ x244;
assign n_29912 = n_29904 ^ n_29311;
assign n_29913 = n_29208 ^ n_29904;
assign n_29914 = n_29905 ^ n_29291;
assign n_29915 = n_29907 ^ n_28080;
assign n_29916 = n_29908 ^ x243;
assign n_29917 = n_29911 ^ n_29908;
assign n_29918 = ~n_29318 & ~n_29912;
assign n_29919 = n_29913 ^ n_29311;
assign n_29920 = n_29914 ^ n_28116;
assign n_29921 = n_29915 ^ n_29914;
assign n_29922 = n_29915 ^ n_28116;
assign n_29923 = n_29911 ^ n_29916;
assign n_29924 = ~n_29916 & n_29917;
assign n_29925 = n_29918 ^ n_29208;
assign n_29926 = ~n_28880 & n_29919;
assign n_29927 = n_29919 ^ n_29766;
assign n_29928 = ~n_29920 & n_29921;
assign n_29929 = n_29922 ^ n_29914;
assign n_29930 = ~n_29909 & ~n_29923;
assign n_29931 = n_29923 ^ n_29909;
assign n_29932 = n_29924 ^ x243;
assign n_29933 = n_29925 ^ n_29325;
assign n_29934 = n_29925 ^ n_29248;
assign n_29935 = n_29926 ^ n_29311;
assign n_29936 = n_29928 ^ n_28116;
assign n_29937 = n_29929 ^ x242;
assign n_29938 = n_29932 ^ n_29929;
assign n_29939 = n_29932 ^ x242;
assign n_29940 = n_29333 & ~n_29933;
assign n_29941 = n_29934 ^ n_29325;
assign n_29942 = n_29935 ^ n_28152;
assign n_29943 = n_29936 ^ n_29935;
assign n_29944 = ~n_29937 & n_29938;
assign n_29945 = n_29939 ^ n_29929;
assign n_29946 = n_29940 ^ n_29248;
assign n_29947 = n_28919 & n_29941;
assign n_29948 = n_29793 ^ n_29941;
assign n_29949 = n_29936 ^ n_29942;
assign n_29950 = ~n_29942 & n_29943;
assign n_29951 = n_29944 ^ x242;
assign n_29952 = ~n_29930 & n_29945;
assign n_29953 = n_29945 ^ n_29930;
assign n_29954 = n_29946 ^ n_29346;
assign n_29955 = n_29946 ^ n_29353;
assign n_29956 = n_29947 ^ n_29325;
assign n_29957 = n_29949 ^ x241;
assign n_29958 = n_29950 ^ n_28152;
assign n_29959 = n_29951 ^ n_29949;
assign n_29960 = n_29353 & n_29954;
assign n_29961 = n_28947 & n_29955;
assign n_29962 = n_29814 ^ n_29955;
assign n_29963 = n_29956 ^ n_28176;
assign n_29964 = n_29951 ^ n_29957;
assign n_29965 = n_29958 ^ n_29956;
assign n_29966 = ~n_29957 & n_29959;
assign n_29967 = n_29960 ^ n_29278;
assign n_29968 = n_29961 ^ n_29346;
assign n_29969 = ~n_29952 & ~n_29964;
assign n_29970 = n_29964 ^ n_29952;
assign n_29971 = ~n_29965 & n_29963;
assign n_29972 = n_29965 ^ n_28176;
assign n_29973 = n_29966 ^ x241;
assign n_29974 = n_29967 ^ n_29371;
assign n_29975 = n_29968 ^ n_28210;
assign n_29976 = n_29446 & n_29970;
assign n_29977 = n_29970 ^ n_29438;
assign n_29978 = n_29971 ^ n_28176;
assign n_29979 = n_29972 ^ x240;
assign n_29980 = n_29973 ^ n_29972;
assign n_29981 = n_29974 & n_29378;
assign n_29982 = n_29296 ^ n_29974;
assign n_29983 = n_29976 ^ n_29478;
assign n_29984 = n_29977 ^ n_28478;
assign n_29985 = n_29978 ^ n_29968;
assign n_29986 = n_29978 ^ n_29975;
assign n_29987 = n_29973 ^ n_29979;
assign n_29988 = n_29979 & ~n_29980;
assign n_29989 = n_29981 ^ n_29296;
assign n_29990 = ~n_28986 & ~n_29982;
assign n_29991 = n_29835 ^ n_29982;
assign n_29992 = ~n_28478 & ~n_29984;
assign n_29993 = ~n_29975 & n_29985;
assign n_29994 = n_29986 ^ x255;
assign n_29995 = n_29987 & n_29969;
assign n_29996 = n_29969 ^ n_29987;
assign n_29997 = n_29988 ^ x240;
assign n_29998 = n_29989 ^ n_29386;
assign n_29999 = n_29989 ^ n_29393;
assign n_30000 = n_29990 ^ n_29371;
assign n_30001 = n_29992 ^ n_29446;
assign n_30002 = n_29447 ^ n_29992;
assign n_30003 = n_29993 ^ n_28210;
assign n_30004 = n_29996 ^ n_29976;
assign n_30005 = n_29996 ^ n_29983;
assign n_30006 = n_29997 ^ n_29986;
assign n_30007 = n_29997 ^ x255;
assign n_30008 = n_29393 & ~n_29998;
assign n_30009 = n_29024 & n_29999;
assign n_30010 = n_29855 ^ n_29999;
assign n_30011 = n_30000 ^ n_28249;
assign n_30012 = n_28069 & ~n_30001;
assign n_30013 = x455 & ~n_30002;
assign n_30014 = n_30002 ^ x455;
assign n_30015 = n_30003 ^ n_30000;
assign n_30016 = n_29983 & ~n_30004;
assign n_30017 = n_28537 & ~n_30005;
assign n_30018 = ~n_29994 & n_30006;
assign n_30019 = n_30007 ^ n_29986;
assign n_30020 = n_30008 ^ n_29323;
assign n_30021 = n_30009 ^ n_29386;
assign n_30022 = n_30003 ^ n_30011;
assign n_30023 = n_30012 ^ n_28085;
assign n_30024 = n_30013 ^ x454;
assign n_30025 = n_30011 & ~n_30015;
assign n_30026 = n_30016 ^ n_29478;
assign n_30027 = n_30017 ^ n_29478;
assign n_30028 = n_30018 ^ x255;
assign n_30029 = n_30019 & ~n_29995;
assign n_30030 = n_29995 ^ n_30019;
assign n_30031 = n_30020 ^ n_29407;
assign n_30032 = n_30021 ^ n_28300;
assign n_30033 = n_30022 ^ x254;
assign n_30034 = n_30025 ^ n_28249;
assign n_30035 = n_30026 ^ n_29514;
assign n_30036 = n_30027 ^ n_30012;
assign n_30037 = n_30027 ^ n_30023;
assign n_30038 = n_30028 ^ n_30022;
assign n_30039 = n_30030 ^ n_29514;
assign n_30040 = n_30026 ^ n_30030;
assign n_30041 = n_29345 ^ n_30031;
assign n_30042 = ~n_30031 & n_29413;
assign n_30043 = n_30028 ^ n_30033;
assign n_30044 = n_30034 ^ n_30021;
assign n_30045 = n_30034 ^ n_30032;
assign n_30046 = n_30035 ^ n_30030;
assign n_30047 = n_30023 & n_30036;
assign n_30048 = n_30037 ^ n_30013;
assign n_30049 = n_30037 ^ n_30024;
assign n_30050 = n_30033 & ~n_30038;
assign n_30051 = ~n_30039 & ~n_30040;
assign n_30052 = ~n_29062 & n_30041;
assign n_30053 = n_29868 ^ n_30041;
assign n_30054 = n_30042 ^ n_29345;
assign n_30055 = n_30029 & ~n_30043;
assign n_30056 = n_30043 ^ n_30029;
assign n_30057 = n_30032 & ~n_30044;
assign n_30058 = n_30045 ^ x253;
assign n_30059 = n_28575 & n_30046;
assign n_30060 = n_30047 ^ n_28085;
assign n_30061 = n_30024 & n_30048;
assign n_30062 = n_30049 & n_30014;
assign n_30063 = n_30014 ^ n_30049;
assign n_30064 = n_30050 ^ x254;
assign n_30065 = n_30051 ^ n_29514;
assign n_30066 = n_30052 ^ n_29407;
assign n_30067 = n_30054 ^ n_29436;
assign n_30068 = n_30054 ^ n_29430;
assign n_30069 = n_30056 ^ n_29543;
assign n_30070 = n_30057 ^ n_28300;
assign n_30071 = n_30059 ^ n_29514;
assign n_30072 = n_30061 ^ x454;
assign n_30073 = n_30064 ^ n_30045;
assign n_30074 = n_30065 ^ n_30056;
assign n_30075 = n_30066 ^ n_28325;
assign n_30076 = n_29101 & ~n_30067;
assign n_30077 = n_29893 ^ n_30067;
assign n_30078 = ~n_29436 & n_30068;
assign n_30079 = n_30070 ^ n_30066;
assign n_30080 = n_30070 ^ n_28325;
assign n_30081 = n_30071 ^ n_28122;
assign n_30082 = n_30060 ^ n_30071;
assign n_30083 = n_30072 ^ x453;
assign n_30084 = ~n_30073 & n_30058;
assign n_30085 = n_30073 ^ x253;
assign n_30086 = n_30074 & n_30069;
assign n_30087 = n_30074 ^ n_29543;
assign n_30088 = n_30076 ^ n_29430;
assign n_30089 = n_30078 ^ n_29364;
assign n_30090 = ~n_30075 & ~n_30079;
assign n_30091 = n_30080 ^ n_30066;
assign n_30092 = n_30060 ^ n_30081;
assign n_30093 = ~n_30081 & ~n_30082;
assign n_30094 = n_30084 ^ x253;
assign n_30095 = n_30085 & ~n_30055;
assign n_30096 = n_30055 ^ n_30085;
assign n_30097 = n_30086 ^ n_29543;
assign n_30098 = ~n_28612 & n_30087;
assign n_30099 = n_30088 ^ n_28364;
assign n_30100 = n_30089 ^ n_29452;
assign n_30101 = n_30090 ^ n_28325;
assign n_30102 = n_30091 ^ x252;
assign n_30103 = n_30092 ^ x453;
assign n_30104 = n_30072 ^ n_30092;
assign n_30105 = n_30083 ^ n_30092;
assign n_30106 = n_30093 ^ n_28122;
assign n_30107 = n_30094 ^ n_30091;
assign n_30108 = n_30094 ^ x252;
assign n_30109 = n_30096 ^ n_29572;
assign n_30110 = n_30097 ^ n_30096;
assign n_30111 = n_30097 ^ n_29572;
assign n_30112 = n_30098 ^ n_29543;
assign n_30113 = n_29384 ^ n_30100;
assign n_30114 = n_30100 & n_29461;
assign n_30115 = n_30101 ^ n_30099;
assign n_30116 = n_30101 ^ n_30088;
assign n_30117 = ~n_30103 & n_30104;
assign n_30118 = n_30062 & n_30105;
assign n_30119 = n_30105 ^ n_30062;
assign n_30120 = ~n_30102 & n_30107;
assign n_30121 = n_30108 ^ n_30091;
assign n_30122 = n_30109 & n_30110;
assign n_30123 = n_30111 ^ n_30096;
assign n_30124 = n_30106 ^ n_30112;
assign n_30125 = n_30112 ^ n_28156;
assign n_30126 = ~n_29140 & n_30113;
assign n_30127 = n_29910 ^ n_30113;
assign n_30128 = n_30114 ^ n_29384;
assign n_30129 = n_30115 ^ x251;
assign n_30130 = ~n_30099 & ~n_30116;
assign n_30131 = n_30117 ^ x453;
assign n_30132 = n_30120 ^ x252;
assign n_30133 = ~n_30121 & n_30095;
assign n_30134 = n_30095 ^ n_30121;
assign n_30135 = n_30122 ^ n_29572;
assign n_30136 = n_28647 & ~n_30123;
assign n_30137 = n_30124 ^ n_28156;
assign n_30138 = ~n_30124 & n_30125;
assign n_30139 = n_30126 ^ n_29452;
assign n_30140 = n_30128 ^ n_29404;
assign n_30141 = n_30128 ^ n_29471;
assign n_30142 = n_30130 ^ n_28364;
assign n_30143 = n_30132 ^ n_30115;
assign n_30144 = n_30132 ^ n_30129;
assign n_30145 = n_30134 ^ n_29591;
assign n_30146 = n_30135 ^ n_30134;
assign n_30147 = n_30136 ^ n_29572;
assign n_30148 = n_30137 ^ x452;
assign n_30149 = n_30131 ^ n_30137;
assign n_30150 = n_30138 ^ n_28156;
assign n_30151 = n_30139 ^ n_28417;
assign n_30152 = n_30140 ^ n_29471;
assign n_30153 = ~n_29484 & ~n_30141;
assign n_30154 = n_30142 ^ n_28417;
assign n_30155 = n_30142 ^ n_30139;
assign n_30156 = n_30129 & ~n_30143;
assign n_30157 = n_30144 & n_30133;
assign n_30158 = n_30133 ^ n_30144;
assign n_30159 = ~n_30146 & ~n_30145;
assign n_30160 = n_30146 ^ n_29591;
assign n_30161 = n_30147 ^ n_28193;
assign n_30162 = n_30131 ^ n_30148;
assign n_30163 = ~n_30148 & n_30149;
assign n_30164 = n_30150 ^ n_30147;
assign n_30165 = n_29180 & n_30152;
assign n_30166 = n_30153 ^ n_29404;
assign n_30167 = n_30154 ^ n_30139;
assign n_30168 = ~n_30151 & n_30155;
assign n_30169 = n_30156 ^ x251;
assign n_30170 = n_30158 ^ n_29610;
assign n_30171 = n_30159 ^ n_29591;
assign n_30172 = n_28675 & ~n_30160;
assign n_30173 = n_30150 ^ n_30161;
assign n_30174 = ~n_30118 & ~n_30162;
assign n_30175 = n_30162 ^ n_30118;
assign n_30176 = n_30163 ^ x452;
assign n_30177 = ~n_30161 & n_30164;
assign n_30178 = n_30165 ^ n_29471;
assign n_30179 = n_30166 ^ n_29504;
assign n_30180 = n_30167 ^ x250;
assign n_30181 = n_30168 ^ n_28417;
assign n_30182 = n_30169 ^ n_30167;
assign n_30183 = n_30171 ^ n_30158;
assign n_30184 = n_30171 ^ n_30170;
assign n_30185 = n_30172 ^ n_29591;
assign n_30186 = n_30173 ^ x451;
assign n_30187 = n_30176 ^ n_30173;
assign n_30188 = n_30177 ^ n_28193;
assign n_30189 = n_30178 ^ n_28443;
assign n_30190 = ~n_29210 & n_30179;
assign n_30191 = n_29953 ^ n_30179;
assign n_30192 = n_30181 ^ n_28443;
assign n_30193 = n_30181 ^ n_30178;
assign n_30194 = n_30182 & ~n_30180;
assign n_30195 = n_30182 ^ x250;
assign n_30196 = n_30170 & ~n_30183;
assign n_30197 = ~n_28721 & ~n_30184;
assign n_30198 = n_30185 ^ n_28228;
assign n_30199 = ~n_30187 & n_30186;
assign n_30200 = n_30187 ^ x451;
assign n_30201 = n_30188 ^ n_30185;
assign n_30202 = n_30188 ^ n_28228;
assign n_30203 = n_30190 ^ n_29494;
assign n_30204 = n_30191 ^ n_29931;
assign n_30205 = n_30192 ^ n_30178;
assign n_30206 = n_30189 & n_30193;
assign n_30207 = n_30194 ^ x250;
assign n_30208 = ~n_30195 & n_30157;
assign n_30209 = n_30157 ^ n_30195;
assign n_30210 = n_30196 ^ n_29610;
assign n_30211 = n_30197 ^ n_29610;
assign n_30212 = n_30199 ^ x451;
assign n_30213 = n_30174 & n_30200;
assign n_30214 = n_30200 ^ n_30174;
assign n_30215 = n_30198 & ~n_30201;
assign n_30216 = n_30202 ^ n_30185;
assign n_30217 = n_30203 ^ n_28467;
assign n_30218 = n_30205 ^ x249;
assign n_30219 = n_30206 ^ n_28443;
assign n_30220 = n_30207 ^ n_30205;
assign n_30221 = n_30209 ^ n_29623;
assign n_30222 = n_30210 ^ n_30209;
assign n_30223 = n_30211 ^ n_28264;
assign n_30224 = n_30215 ^ n_28228;
assign n_30225 = n_30216 ^ x450;
assign n_30226 = n_30212 ^ n_30216;
assign n_30227 = n_30219 ^ n_30217;
assign n_30228 = ~n_30220 & n_30218;
assign n_30229 = n_30220 ^ x249;
assign n_30230 = n_30222 & ~n_30221;
assign n_30231 = n_30222 ^ n_29623;
assign n_30232 = n_30224 ^ n_30211;
assign n_30233 = n_30224 ^ n_30223;
assign n_30234 = n_30212 ^ n_30225;
assign n_30235 = ~n_30225 & n_30226;
assign n_30236 = n_30228 ^ x249;
assign n_30237 = ~n_30208 & ~n_30229;
assign n_30238 = n_30229 ^ n_30208;
assign n_30239 = n_30230 ^ n_29623;
assign n_30240 = ~n_28758 & n_30231;
assign n_30241 = ~n_30223 & ~n_30232;
assign n_30242 = n_30233 ^ x449;
assign n_30243 = ~n_30213 & n_30234;
assign n_30244 = n_30234 ^ n_30213;
assign n_30245 = n_30235 ^ x450;
assign n_30246 = n_30236 ^ n_30227;
assign n_30247 = n_30238 ^ n_29647;
assign n_30248 = n_30239 ^ n_30238;
assign n_30249 = n_30240 ^ n_29623;
assign n_30250 = n_30241 ^ n_28264;
assign n_30251 = n_30245 ^ n_30233;
assign n_30252 = n_30245 ^ n_30242;
assign n_30253 = n_30246 ^ x248;
assign n_30254 = n_30248 & ~n_30247;
assign n_30255 = n_30248 ^ n_29647;
assign n_30256 = n_30249 ^ n_28309;
assign n_30257 = n_30250 ^ n_30249;
assign n_30258 = n_30242 & ~n_30251;
assign n_30259 = ~n_30243 & n_30252;
assign n_30260 = n_30252 ^ n_30243;
assign n_30261 = n_30253 ^ n_30237;
assign n_30262 = n_30254 ^ n_29647;
assign n_30263 = n_28794 & n_30255;
assign n_30264 = n_30250 ^ n_30256;
assign n_30265 = ~n_30256 & n_30257;
assign n_30266 = n_30258 ^ x449;
assign n_30267 = n_30261 ^ n_29666;
assign n_30268 = n_30262 ^ n_30261;
assign n_30269 = n_30263 ^ n_29647;
assign n_30270 = n_30264 ^ x448;
assign n_30271 = n_30265 ^ n_28309;
assign n_30272 = n_30266 ^ n_30264;
assign n_30273 = n_30262 ^ n_30267;
assign n_30274 = ~n_30267 & n_30268;
assign n_30275 = n_30269 ^ n_28350;
assign n_30276 = n_30266 ^ n_30270;
assign n_30277 = n_30271 ^ n_30269;
assign n_30278 = ~n_30270 & n_30272;
assign n_30279 = n_28837 & n_30273;
assign n_30280 = n_30274 ^ n_29666;
assign n_30281 = n_30271 ^ n_30275;
assign n_30282 = ~n_30259 & n_30276;
assign n_30283 = n_30276 ^ n_30259;
assign n_30284 = ~n_30275 & n_30277;
assign n_30285 = n_30278 ^ x448;
assign n_30286 = n_30279 ^ n_29666;
assign n_30287 = n_30280 ^ n_29476;
assign n_30288 = n_30280 ^ n_29694;
assign n_30289 = n_30281 ^ x463;
assign n_30290 = n_30284 ^ n_28350;
assign n_30291 = n_30285 ^ n_30281;
assign n_30292 = n_30286 ^ n_28385;
assign n_30293 = ~n_29694 & ~n_30287;
assign n_30294 = n_28874 & n_30288;
assign n_30295 = n_30290 ^ n_30286;
assign n_30296 = n_30291 & ~n_30289;
assign n_30297 = n_30291 ^ x463;
assign n_30298 = n_30290 ^ n_30292;
assign n_30299 = n_30293 ^ n_29686;
assign n_30300 = n_30294 ^ n_29686;
assign n_30301 = ~n_30292 & n_30295;
assign n_30302 = n_30296 ^ x463;
assign n_30303 = n_30297 & n_30282;
assign n_30304 = n_30282 ^ n_30297;
assign n_30305 = n_30298 ^ x462;
assign n_30306 = n_30299 ^ n_29701;
assign n_30307 = n_30299 ^ n_29707;
assign n_30308 = n_30301 ^ n_28385;
assign n_30309 = n_30302 ^ n_30298;
assign n_30310 = n_29707 & ~n_30306;
assign n_30311 = n_28912 & n_30307;
assign n_30312 = n_30308 ^ n_30300;
assign n_30313 = n_30308 ^ n_28422;
assign n_30314 = n_30309 & ~n_30305;
assign n_30315 = n_30309 ^ x462;
assign n_30316 = n_30310 ^ n_29537;
assign n_30317 = n_30311 ^ n_29701;
assign n_30318 = n_30312 ^ n_28422;
assign n_30319 = ~n_30312 & n_30313;
assign n_30320 = n_30314 ^ x462;
assign n_30321 = n_30303 & n_30315;
assign n_30322 = n_30315 ^ n_30303;
assign n_30323 = n_30316 ^ n_29725;
assign n_30324 = n_30316 ^ n_29564;
assign n_30325 = n_30317 ^ n_28461;
assign n_30326 = n_30318 ^ x461;
assign n_30327 = n_30319 ^ n_28422;
assign n_30328 = n_30320 ^ n_30318;
assign n_30329 = ~n_29732 & n_30323;
assign n_30330 = n_30324 ^ n_29725;
assign n_30331 = n_30320 ^ n_30326;
assign n_30332 = n_30327 ^ n_30317;
assign n_30333 = n_30327 ^ n_30325;
assign n_30334 = n_30326 & ~n_30328;
assign n_30335 = n_30329 ^ n_29564;
assign n_30336 = n_28953 & ~n_30330;
assign n_30337 = n_30331 & ~n_30321;
assign n_30338 = n_30321 ^ n_30331;
assign n_30339 = n_30325 & ~n_30332;
assign n_30340 = n_30333 ^ x460;
assign n_30341 = n_30334 ^ x461;
assign n_30342 = n_30335 ^ n_29738;
assign n_30343 = n_30335 ^ n_29744;
assign n_30344 = n_30336 ^ n_29725;
assign n_30345 = n_30339 ^ n_28461;
assign n_30346 = n_30341 ^ n_30333;
assign n_30347 = n_30341 ^ x460;
assign n_30348 = ~n_29744 & n_30342;
assign n_30349 = ~n_28991 & ~n_30343;
assign n_30350 = n_30344 ^ n_28500;
assign n_30351 = n_30345 ^ n_30344;
assign n_30352 = n_30345 ^ n_28500;
assign n_30353 = n_30340 & ~n_30346;
assign n_30354 = n_30347 ^ n_30333;
assign n_30355 = n_30348 ^ n_29594;
assign n_30356 = n_30349 ^ n_29738;
assign n_30357 = ~n_30350 & n_30351;
assign n_30358 = n_30352 ^ n_30344;
assign n_30359 = n_30353 ^ x460;
assign n_30360 = n_30337 & n_30354;
assign n_30361 = n_30354 ^ n_30337;
assign n_30362 = n_30355 ^ n_29763;
assign n_30363 = n_30355 ^ n_29769;
assign n_30364 = n_30356 ^ n_28544;
assign n_30365 = n_30357 ^ n_28500;
assign n_30366 = n_30358 ^ x459;
assign n_30367 = n_30359 ^ n_30358;
assign n_30368 = n_30359 ^ x459;
assign n_30369 = n_29769 & n_30362;
assign n_30370 = ~n_29032 & n_30363;
assign n_30371 = n_30365 ^ n_30356;
assign n_30372 = n_30365 ^ n_30364;
assign n_30373 = ~n_30366 & n_30367;
assign n_30374 = n_30368 ^ n_30358;
assign n_30375 = n_30369 ^ n_29613;
assign n_30376 = n_30370 ^ n_29763;
assign n_30377 = ~n_30364 & n_30371;
assign n_30378 = n_30372 ^ x458;
assign n_30379 = n_30373 ^ x459;
assign n_30380 = n_30360 & ~n_30374;
assign n_30381 = n_30374 ^ n_30360;
assign n_30382 = n_30375 ^ n_29775;
assign n_30383 = n_30375 ^ n_29781;
assign n_30384 = n_30376 ^ n_28580;
assign n_30385 = n_30377 ^ n_28544;
assign n_30386 = n_30379 ^ n_30372;
assign n_30387 = ~n_29781 & n_30382;
assign n_30388 = n_29066 & n_30383;
assign n_30389 = n_30014 ^ n_30383;
assign n_30390 = n_30385 ^ n_30376;
assign n_30391 = n_30386 & ~n_30378;
assign n_30392 = n_30386 ^ x458;
assign n_30393 = n_30387 ^ n_29632;
assign n_30394 = n_30388 ^ n_29775;
assign n_30395 = n_30390 & n_30384;
assign n_30396 = n_30390 ^ n_28580;
assign n_30397 = n_30391 ^ x458;
assign n_30398 = n_30392 & ~n_30380;
assign n_30399 = n_30380 ^ n_30392;
assign n_30400 = n_30393 ^ n_29802;
assign n_30401 = n_30394 ^ n_28615;
assign n_30402 = n_30395 ^ n_28580;
assign n_30403 = n_30396 ^ x457;
assign n_30404 = n_30397 ^ n_30396;
assign n_30405 = ~n_30400 & ~n_29809;
assign n_30406 = n_29650 ^ n_30400;
assign n_30407 = n_30402 ^ n_30394;
assign n_30408 = n_30402 ^ n_30401;
assign n_30409 = n_30397 ^ n_30403;
assign n_30410 = n_30403 & ~n_30404;
assign n_30411 = n_30405 ^ n_29650;
assign n_30412 = ~n_29105 & n_30406;
assign n_30413 = n_30063 ^ n_30406;
assign n_30414 = ~n_30401 & n_30407;
assign n_30415 = n_30408 ^ x456;
assign n_30416 = ~n_30398 & n_30409;
assign n_30417 = n_30409 ^ n_30398;
assign n_30418 = n_30410 ^ x457;
assign n_30419 = n_30411 ^ n_29816;
assign n_30420 = n_30411 ^ n_29822;
assign n_30421 = n_30412 ^ n_29802;
assign n_30422 = n_30414 ^ n_28615;
assign n_30423 = n_30418 ^ n_30408;
assign n_30424 = n_29822 & n_30419;
assign n_30425 = n_29147 & n_30420;
assign n_30426 = n_30119 ^ n_30420;
assign n_30427 = n_30421 ^ n_28639;
assign n_30428 = n_30422 ^ n_30421;
assign n_30429 = n_30422 ^ n_28639;
assign n_30430 = ~n_30423 & n_30415;
assign n_30431 = n_30423 ^ x456;
assign n_30432 = n_30424 ^ n_29669;
assign n_30433 = n_30425 ^ n_29816;
assign n_30434 = ~n_30427 & ~n_30428;
assign n_30435 = n_30429 ^ n_30421;
assign n_30436 = n_30430 ^ x456;
assign n_30437 = n_30416 & n_30431;
assign n_30438 = n_30431 ^ n_30416;
assign n_30439 = n_30432 ^ n_29837;
assign n_30440 = n_30432 ^ n_29689;
assign n_30441 = n_30433 ^ n_28687;
assign n_30442 = n_30434 ^ n_28639;
assign n_30443 = n_30435 ^ x471;
assign n_30444 = n_30436 ^ n_30435;
assign n_30445 = n_29843 & n_30439;
assign n_30446 = n_30440 ^ n_29837;
assign n_30447 = n_30442 ^ n_30433;
assign n_30448 = n_30442 ^ n_30441;
assign n_30449 = n_30436 ^ n_30443;
assign n_30450 = n_30443 & ~n_30444;
assign n_30451 = n_30445 ^ n_29689;
assign n_30452 = ~n_29189 & ~n_30446;
assign n_30453 = n_30175 ^ n_30446;
assign n_30454 = n_30441 & n_30447;
assign n_30455 = n_30448 ^ x470;
assign n_30456 = n_30437 & n_30449;
assign n_30457 = n_30449 ^ n_30437;
assign n_30458 = n_30450 ^ x471;
assign n_30459 = n_30451 ^ n_29856;
assign n_30460 = n_30451 ^ n_29710;
assign n_30461 = n_30452 ^ n_29837;
assign n_30462 = n_30454 ^ n_28687;
assign n_30463 = n_30458 ^ n_30448;
assign n_30464 = n_30458 ^ x470;
assign n_30465 = n_29862 & ~n_30459;
assign n_30466 = n_30460 ^ n_29856;
assign n_30467 = n_30461 ^ n_28713;
assign n_30468 = n_30462 ^ n_30461;
assign n_30469 = n_30462 ^ n_28713;
assign n_30470 = n_30455 & ~n_30463;
assign n_30471 = n_30464 ^ n_30448;
assign n_30472 = n_30465 ^ n_29710;
assign n_30473 = ~n_29227 & n_30466;
assign n_30474 = n_30214 ^ n_30466;
assign n_30475 = n_30467 & n_30468;
assign n_30476 = n_30469 ^ n_30461;
assign n_30477 = n_30470 ^ x470;
assign n_30478 = n_30456 & n_30471;
assign n_30479 = n_30471 ^ n_30456;
assign n_30480 = n_30472 ^ n_29876;
assign n_30481 = n_30473 ^ n_29856;
assign n_30482 = n_30475 ^ n_28713;
assign n_30483 = n_30476 ^ x469;
assign n_30484 = n_30477 ^ n_30476;
assign n_30485 = n_29984 & n_30479;
assign n_30486 = n_30479 ^ n_29970;
assign n_30487 = n_30479 ^ n_29984;
assign n_30488 = n_29727 ^ n_30480;
assign n_30489 = n_30480 & ~n_29882;
assign n_30490 = n_30481 ^ n_28752;
assign n_30491 = n_30482 ^ n_30481;
assign n_30492 = n_30477 ^ n_30483;
assign n_30493 = ~n_30483 & n_30484;
assign n_30494 = n_30485 ^ n_30005;
assign n_30495 = n_29446 & ~n_30487;
assign n_30496 = ~n_29259 & ~n_30488;
assign n_30497 = n_30244 ^ n_30488;
assign n_30498 = n_30489 ^ n_29727;
assign n_30499 = ~n_30491 & n_30490;
assign n_30500 = n_30491 ^ n_28752;
assign n_30501 = ~n_30478 & n_30492;
assign n_30502 = n_30492 ^ n_30478;
assign n_30503 = n_30493 ^ x469;
assign n_30504 = n_30495 ^ n_29977;
assign n_30505 = n_30496 ^ n_29876;
assign n_30506 = n_30498 ^ n_29906;
assign n_30507 = n_30498 ^ n_29900;
assign n_30508 = n_30499 ^ n_28752;
assign n_30509 = n_30500 ^ x468;
assign n_30510 = n_30502 ^ n_30485;
assign n_30511 = n_30502 ^ n_30494;
assign n_30512 = n_30503 ^ n_30500;
assign n_30513 = ~n_28478 & ~n_30504;
assign n_30514 = x167 & n_30504;
assign n_30515 = n_30504 ^ x167;
assign n_30516 = n_30505 ^ n_28791;
assign n_30517 = n_29291 & n_30506;
assign n_30518 = n_30260 ^ n_30506;
assign n_30519 = n_29906 & ~n_30507;
assign n_30520 = n_30508 ^ n_30505;
assign n_30521 = n_30508 ^ n_28791;
assign n_30522 = n_30503 ^ n_30509;
assign n_30523 = n_30494 & ~n_30510;
assign n_30524 = n_29478 & ~n_30511;
assign n_30525 = n_30509 & ~n_30512;
assign n_30526 = n_30513 ^ n_28537;
assign n_30527 = n_30514 ^ x166;
assign n_30528 = n_30517 ^ n_29900;
assign n_30529 = n_30519 ^ n_29750;
assign n_30530 = ~n_30516 & n_30520;
assign n_30531 = n_30521 ^ n_30505;
assign n_30532 = ~n_30501 & n_30522;
assign n_30533 = n_30522 ^ n_30501;
assign n_30534 = n_30523 ^ n_30005;
assign n_30535 = n_30524 ^ n_30005;
assign n_30536 = n_30525 ^ x468;
assign n_30537 = n_30528 ^ n_28830;
assign n_30538 = n_30529 ^ n_29927;
assign n_30539 = n_30529 ^ n_29919;
assign n_30540 = n_30530 ^ n_28791;
assign n_30541 = n_30531 ^ x467;
assign n_30542 = n_30533 ^ n_30046;
assign n_30543 = n_30534 ^ n_30533;
assign n_30544 = n_30535 ^ n_30513;
assign n_30545 = n_30535 ^ n_30526;
assign n_30546 = n_30536 ^ n_30531;
assign n_30547 = n_29311 & ~n_30538;
assign n_30548 = n_30283 ^ n_30538;
assign n_30549 = ~n_29927 & ~n_30539;
assign n_30550 = n_30540 ^ n_30528;
assign n_30551 = n_30536 ^ n_30541;
assign n_30552 = n_30534 ^ n_30542;
assign n_30553 = n_30542 & n_30543;
assign n_30554 = n_30526 & n_30544;
assign n_30555 = n_30545 ^ n_30514;
assign n_30556 = n_30545 ^ n_30527;
assign n_30557 = ~n_30541 & n_30546;
assign n_30558 = n_30547 ^ n_29919;
assign n_30559 = n_30549 ^ n_29766;
assign n_30560 = ~n_30550 & ~n_30537;
assign n_30561 = n_30550 ^ n_28830;
assign n_30562 = ~n_30532 & n_30551;
assign n_30563 = n_30551 ^ n_30532;
assign n_30564 = ~n_29514 & ~n_30552;
assign n_30565 = n_30553 ^ n_30046;
assign n_30566 = n_30554 ^ n_28537;
assign n_30567 = n_30527 & n_30555;
assign n_30568 = n_30515 & ~n_30556;
assign n_30569 = n_30556 ^ n_30515;
assign n_30570 = n_30557 ^ x467;
assign n_30571 = n_30558 ^ n_28880;
assign n_30572 = n_29948 ^ n_30559;
assign n_30573 = n_30559 ^ n_29941;
assign n_30574 = n_30560 ^ n_28830;
assign n_30575 = n_30561 ^ x466;
assign n_30576 = n_30563 ^ n_30087;
assign n_30577 = n_30564 ^ n_30046;
assign n_30578 = n_30565 ^ n_30563;
assign n_30579 = n_30567 ^ x166;
assign n_30580 = n_30570 ^ n_30561;
assign n_30581 = n_30570 ^ x466;
assign n_30582 = ~n_29325 & n_30572;
assign n_30583 = n_30304 ^ n_30572;
assign n_30584 = ~n_29948 & n_30573;
assign n_30585 = n_30574 ^ n_28880;
assign n_30586 = n_30574 ^ n_30558;
assign n_30587 = n_30565 ^ n_30576;
assign n_30588 = n_30577 ^ n_28575;
assign n_30589 = n_30566 ^ n_30577;
assign n_30590 = ~n_30576 & n_30578;
assign n_30591 = ~n_30575 & n_30580;
assign n_30592 = n_30581 ^ n_30561;
assign n_30593 = n_30582 ^ n_29941;
assign n_30594 = n_30584 ^ n_29793;
assign n_30595 = n_30585 ^ n_30558;
assign n_30596 = ~n_30571 & n_30586;
assign n_30597 = n_29543 & ~n_30587;
assign n_30598 = n_30566 ^ n_30588;
assign n_30599 = n_30588 & ~n_30589;
assign n_30600 = n_30590 ^ n_30087;
assign n_30601 = n_30591 ^ x466;
assign n_30602 = ~n_30592 & ~n_30562;
assign n_30603 = n_30562 ^ n_30592;
assign n_30604 = n_30593 ^ n_28919;
assign n_30605 = n_29962 ^ n_30594;
assign n_30606 = n_30594 ^ n_29955;
assign n_30607 = n_30595 ^ x465;
assign n_30608 = n_30596 ^ n_28880;
assign n_30609 = n_30597 ^ n_30087;
assign n_30610 = n_30598 ^ x165;
assign n_30611 = n_30579 ^ n_30598;
assign n_30612 = n_30599 ^ n_28575;
assign n_30613 = n_30600 ^ n_30123;
assign n_30614 = n_30601 ^ n_30595;
assign n_30615 = n_30603 ^ n_30123;
assign n_30616 = n_30600 ^ n_30603;
assign n_30617 = n_29346 & n_30605;
assign n_30618 = n_30322 ^ n_30605;
assign n_30619 = ~n_29962 & n_30606;
assign n_30620 = n_30601 ^ n_30607;
assign n_30621 = n_30608 ^ n_30604;
assign n_30622 = n_30608 ^ n_30593;
assign n_30623 = n_30609 ^ n_28612;
assign n_30624 = n_30579 ^ n_30610;
assign n_30625 = n_30610 & ~n_30611;
assign n_30626 = n_30612 ^ n_30609;
assign n_30627 = n_30613 ^ n_30603;
assign n_30628 = n_30607 & ~n_30614;
assign n_30629 = n_30615 & n_30616;
assign n_30630 = n_30617 ^ n_29955;
assign n_30631 = n_30619 ^ n_29814;
assign n_30632 = n_30620 & n_30602;
assign n_30633 = n_30602 ^ n_30620;
assign n_30634 = n_30621 ^ x464;
assign n_30635 = n_30604 & n_30622;
assign n_30636 = n_30568 & n_30624;
assign n_30637 = n_30624 ^ n_30568;
assign n_30638 = n_30625 ^ x165;
assign n_30639 = ~n_30626 & ~n_30623;
assign n_30640 = n_30626 ^ n_28612;
assign n_30641 = ~n_29572 & n_30627;
assign n_30642 = n_30628 ^ x465;
assign n_30643 = n_30629 ^ n_30123;
assign n_30644 = n_30630 ^ n_28947;
assign n_30645 = n_30631 ^ n_29982;
assign n_30646 = n_30633 ^ n_30160;
assign n_30647 = n_30635 ^ n_28919;
assign n_30648 = n_30639 ^ n_28612;
assign n_30649 = n_30640 ^ x164;
assign n_30650 = n_30638 ^ n_30640;
assign n_30651 = n_30641 ^ n_30123;
assign n_30652 = n_30642 ^ n_30634;
assign n_30653 = n_30642 ^ n_30621;
assign n_30654 = n_30643 ^ n_30633;
assign n_30655 = n_30643 ^ n_30160;
assign n_30656 = n_29835 ^ n_30645;
assign n_30657 = ~n_30645 & ~n_29991;
assign n_30658 = n_30647 ^ n_28947;
assign n_30659 = n_30630 ^ n_30647;
assign n_30660 = n_30638 ^ n_30649;
assign n_30661 = ~n_30649 & n_30650;
assign n_30662 = n_30648 ^ n_30651;
assign n_30663 = n_30651 ^ n_28647;
assign n_30664 = n_30652 ^ n_30632;
assign n_30665 = ~n_30632 & n_30652;
assign n_30666 = ~n_30634 & n_30653;
assign n_30667 = n_30646 & ~n_30654;
assign n_30668 = n_30655 ^ n_30633;
assign n_30669 = ~n_29371 & n_30656;
assign n_30670 = n_30338 ^ n_30656;
assign n_30671 = n_30657 ^ n_29835;
assign n_30672 = n_30630 ^ n_30658;
assign n_30673 = n_30644 & ~n_30659;
assign n_30674 = ~n_30636 & n_30660;
assign n_30675 = n_30660 ^ n_30636;
assign n_30676 = n_30661 ^ x164;
assign n_30677 = n_30662 ^ n_28647;
assign n_30678 = ~n_30662 & ~n_30663;
assign n_30679 = n_30664 ^ n_30184;
assign n_30680 = n_30666 ^ x464;
assign n_30681 = n_30667 ^ n_30160;
assign n_30682 = n_29591 & ~n_30668;
assign n_30683 = n_30669 ^ n_29982;
assign n_30684 = n_30671 ^ n_29999;
assign n_30685 = n_30672 ^ x479;
assign n_30686 = n_30673 ^ n_28947;
assign n_30687 = n_30677 ^ x163;
assign n_30688 = n_30676 ^ n_30677;
assign n_30689 = n_30678 ^ n_28647;
assign n_30690 = n_30680 ^ n_30672;
assign n_30691 = n_30681 ^ n_30664;
assign n_30692 = n_30681 ^ n_30184;
assign n_30693 = n_30682 ^ n_30160;
assign n_30694 = n_30683 ^ n_28986;
assign n_30695 = n_30684 ^ n_29855;
assign n_30696 = ~n_30684 & ~n_30010;
assign n_30697 = n_30680 ^ n_30685;
assign n_30698 = n_30686 ^ n_30683;
assign n_30699 = n_30676 ^ n_30687;
assign n_30700 = n_30687 & ~n_30688;
assign n_30701 = n_30685 & ~n_30690;
assign n_30702 = n_30679 & ~n_30691;
assign n_30703 = n_30692 ^ n_30664;
assign n_30704 = n_30689 ^ n_30693;
assign n_30705 = n_30693 ^ n_28675;
assign n_30706 = ~n_29386 & ~n_30695;
assign n_30707 = n_30361 ^ n_30695;
assign n_30708 = n_30696 ^ n_29855;
assign n_30709 = n_30665 ^ n_30697;
assign n_30710 = ~n_30697 & n_30665;
assign n_30711 = n_30698 ^ n_28986;
assign n_30712 = n_30698 & n_30694;
assign n_30713 = n_30674 & ~n_30699;
assign n_30714 = n_30699 ^ n_30674;
assign n_30715 = n_30700 ^ x163;
assign n_30716 = n_30701 ^ x479;
assign n_30717 = n_30702 ^ n_30184;
assign n_30718 = n_29610 & ~n_30703;
assign n_30719 = n_30704 ^ n_28675;
assign n_30720 = n_30704 & ~n_30705;
assign n_30721 = n_30706 ^ n_29999;
assign n_30722 = n_30708 ^ n_30053;
assign n_30723 = n_30708 ^ n_30041;
assign n_30724 = n_30709 ^ n_30231;
assign n_30725 = n_30711 ^ x478;
assign n_30726 = n_30712 ^ n_28986;
assign n_30727 = n_30716 ^ x478;
assign n_30728 = n_30711 ^ n_30716;
assign n_30729 = n_30717 ^ n_30709;
assign n_30730 = n_30718 ^ n_30184;
assign n_30731 = n_30719 ^ x162;
assign n_30732 = n_30715 ^ n_30719;
assign n_30733 = n_30720 ^ n_28675;
assign n_30734 = n_30721 ^ n_29024;
assign n_30735 = ~n_29407 & n_30722;
assign n_30736 = n_30381 ^ n_30722;
assign n_30737 = ~n_30053 & n_30723;
assign n_30738 = n_30717 ^ n_30724;
assign n_30739 = n_30725 ^ n_30716;
assign n_30740 = n_30721 ^ n_30726;
assign n_30741 = n_30727 & ~n_30728;
assign n_30742 = ~n_30724 & ~n_30729;
assign n_30743 = n_30730 ^ n_28721;
assign n_30744 = n_30715 ^ n_30731;
assign n_30745 = ~n_30731 & n_30732;
assign n_30746 = n_30730 ^ n_30733;
assign n_30747 = n_30734 ^ n_30726;
assign n_30748 = n_30735 ^ n_30041;
assign n_30749 = n_30737 ^ n_29868;
assign n_30750 = n_29623 & n_30738;
assign n_30751 = n_30710 ^ n_30739;
assign n_30752 = ~n_30739 & n_30710;
assign n_30753 = n_30734 & n_30740;
assign n_30754 = n_30741 ^ x478;
assign n_30755 = n_30742 ^ n_30231;
assign n_30756 = n_30713 & n_30744;
assign n_30757 = n_30744 ^ n_30713;
assign n_30758 = n_30745 ^ x162;
assign n_30759 = n_30746 ^ n_28721;
assign n_30760 = n_30746 & n_30743;
assign n_30761 = n_30747 ^ x477;
assign n_30762 = n_30748 ^ n_29062;
assign n_30763 = n_30749 ^ n_30067;
assign n_30764 = n_30750 ^ n_30231;
assign n_30765 = n_30751 ^ n_30255;
assign n_30766 = n_30753 ^ n_29024;
assign n_30767 = n_30747 ^ n_30754;
assign n_30768 = n_30755 ^ n_30255;
assign n_30769 = n_30755 ^ n_30751;
assign n_30770 = n_30759 ^ x161;
assign n_30771 = n_30758 ^ n_30759;
assign n_30772 = n_30760 ^ n_28721;
assign n_30773 = n_30761 ^ n_30754;
assign n_30774 = n_30763 ^ n_29893;
assign n_30775 = ~n_30763 & n_30077;
assign n_30776 = n_30764 ^ n_28758;
assign n_30777 = n_30762 ^ n_30766;
assign n_30778 = n_30748 ^ n_30766;
assign n_30779 = ~n_30761 & n_30767;
assign n_30780 = n_30768 ^ n_30751;
assign n_30781 = ~n_30765 & n_30769;
assign n_30782 = n_30758 ^ n_30770;
assign n_30783 = n_30770 & ~n_30771;
assign n_30784 = n_30772 ^ n_30764;
assign n_30785 = n_30752 ^ n_30773;
assign n_30786 = ~n_30773 & ~n_30752;
assign n_30787 = n_29430 & ~n_30774;
assign n_30788 = n_30399 ^ n_30774;
assign n_30789 = n_30775 ^ n_29893;
assign n_30790 = n_30777 ^ x476;
assign n_30791 = ~n_30762 & ~n_30778;
assign n_30792 = n_30779 ^ x477;
assign n_30793 = n_29647 & ~n_30780;
assign n_30794 = n_30781 ^ n_30255;
assign n_30795 = ~n_30756 & n_30782;
assign n_30796 = n_30782 ^ n_30756;
assign n_30797 = n_30783 ^ x161;
assign n_30798 = n_30784 ^ n_28758;
assign n_30799 = n_30784 & ~n_30776;
assign n_30800 = n_30785 ^ n_30273;
assign n_30801 = n_30787 ^ n_30067;
assign n_30802 = n_30789 ^ n_30127;
assign n_30803 = n_30789 ^ n_30113;
assign n_30804 = n_30791 ^ n_29062;
assign n_30805 = n_30790 ^ n_30792;
assign n_30806 = n_30777 ^ n_30792;
assign n_30807 = n_30793 ^ n_30255;
assign n_30808 = n_30794 ^ n_30785;
assign n_30809 = n_30797 ^ x160;
assign n_30810 = n_30798 ^ x160;
assign n_30811 = n_30797 ^ n_30798;
assign n_30812 = n_30799 ^ n_28758;
assign n_30813 = n_30794 ^ n_30800;
assign n_30814 = n_30801 ^ n_29101;
assign n_30815 = n_29452 & ~n_30802;
assign n_30816 = n_30417 ^ n_30802;
assign n_30817 = n_30127 & n_30803;
assign n_30818 = n_30804 ^ n_30801;
assign n_30819 = n_30786 ^ n_30805;
assign n_30820 = n_30805 & ~n_30786;
assign n_30821 = ~n_30790 & n_30806;
assign n_30822 = n_30807 ^ n_28794;
assign n_30823 = ~n_30800 & n_30808;
assign n_30824 = n_30809 ^ n_30798;
assign n_30825 = n_30810 & ~n_30811;
assign n_30826 = n_30812 ^ n_28794;
assign n_30827 = n_30812 ^ n_30807;
assign n_30828 = n_29666 & ~n_30813;
assign n_30829 = n_30815 ^ n_30113;
assign n_30830 = n_30817 ^ n_29910;
assign n_30831 = n_30818 ^ n_29101;
assign n_30832 = ~n_30818 & ~n_30814;
assign n_30833 = n_30819 ^ n_30288;
assign n_30834 = n_30821 ^ x476;
assign n_30835 = n_30823 ^ n_30273;
assign n_30836 = n_30824 & n_30795;
assign n_30837 = n_30795 ^ n_30824;
assign n_30838 = n_30825 ^ x160;
assign n_30839 = n_30826 ^ n_30807;
assign n_30840 = n_30822 & n_30827;
assign n_30841 = n_30828 ^ n_30273;
assign n_30842 = n_30829 ^ n_29140;
assign n_30843 = n_30830 ^ n_30152;
assign n_30844 = n_29931 ^ n_30830;
assign n_30845 = n_30831 ^ x475;
assign n_30846 = n_30832 ^ n_29101;
assign n_30847 = n_30831 ^ n_30834;
assign n_30848 = n_30833 ^ n_30835;
assign n_30849 = n_30819 ^ n_30835;
assign n_30850 = n_30839 ^ x175;
assign n_30851 = n_30838 ^ n_30839;
assign n_30852 = n_30840 ^ n_28794;
assign n_30853 = n_30841 ^ n_28837;
assign n_30854 = n_29931 ^ n_30843;
assign n_30855 = ~n_30843 & ~n_30844;
assign n_30856 = n_30845 ^ n_30834;
assign n_30857 = n_30846 ^ n_29140;
assign n_30858 = n_30846 ^ n_30829;
assign n_30859 = n_30845 & ~n_30847;
assign n_30860 = ~n_29686 & ~n_30848;
assign n_30861 = ~n_30833 & n_30849;
assign n_30862 = n_30838 ^ n_30850;
assign n_30863 = ~n_30850 & n_30851;
assign n_30864 = n_30841 ^ n_30852;
assign n_30865 = n_29471 & ~n_30854;
assign n_30866 = n_30438 ^ n_30854;
assign n_30867 = n_30204 ^ n_30855;
assign n_30868 = n_30856 ^ n_30820;
assign n_30869 = ~n_30820 & n_30856;
assign n_30870 = n_30857 ^ n_30829;
assign n_30871 = ~n_30842 & ~n_30858;
assign n_30872 = n_30859 ^ x475;
assign n_30873 = n_30860 ^ n_30288;
assign n_30874 = n_30861 ^ n_30288;
assign n_30875 = n_30836 & ~n_30862;
assign n_30876 = n_30862 ^ n_30836;
assign n_30877 = n_30863 ^ x175;
assign n_30878 = n_30864 ^ n_28837;
assign n_30879 = ~n_30864 & n_30853;
assign n_30880 = n_30865 ^ n_30152;
assign n_30881 = ~n_29494 & n_30867;
assign n_30882 = n_30457 ^ n_30867;
assign n_30883 = n_30868 ^ n_30307;
assign n_30884 = n_30870 ^ x474;
assign n_30885 = n_30871 ^ n_29140;
assign n_30886 = n_30870 ^ n_30872;
assign n_30887 = n_30873 ^ n_28874;
assign n_30888 = n_30868 ^ n_30874;
assign n_30889 = n_30878 ^ x174;
assign n_30890 = n_30877 ^ n_30878;
assign n_30891 = n_30879 ^ n_28837;
assign n_30892 = n_30880 ^ n_29180;
assign n_30893 = n_30881 ^ n_30179;
assign n_30894 = n_30882 ^ n_30854;
assign n_30895 = n_30883 ^ n_30874;
assign n_30896 = n_30884 ^ n_30872;
assign n_30897 = n_30885 ^ n_30880;
assign n_30898 = ~n_30884 & n_30886;
assign n_30899 = n_30883 & ~n_30888;
assign n_30900 = n_30877 ^ n_30889;
assign n_30901 = n_30889 & ~n_30890;
assign n_30902 = n_30891 ^ n_30873;
assign n_30903 = n_30885 ^ n_30892;
assign n_30904 = ~n_29701 & n_30895;
assign n_30905 = ~n_30869 & n_30896;
assign n_30906 = n_30896 ^ n_30869;
assign n_30907 = n_30892 & n_30897;
assign n_30908 = n_30898 ^ x474;
assign n_30909 = n_30899 ^ n_30307;
assign n_30910 = n_30875 & n_30900;
assign n_30911 = n_30900 ^ n_30875;
assign n_30912 = n_30901 ^ x174;
assign n_30913 = n_30902 ^ n_28874;
assign n_30914 = ~n_30902 & n_30887;
assign n_30915 = n_30903 ^ x473;
assign n_30916 = n_30904 ^ n_30307;
assign n_30917 = n_30906 ^ n_30330;
assign n_30918 = n_30907 ^ n_29180;
assign n_30919 = n_30908 ^ n_30903;
assign n_30920 = n_30906 ^ n_30909;
assign n_30921 = n_30909 ^ n_30330;
assign n_30922 = n_30912 ^ x173;
assign n_30923 = n_30913 ^ x173;
assign n_30924 = n_30913 ^ n_30912;
assign n_30925 = n_30914 ^ n_28874;
assign n_30926 = n_30916 ^ n_28912;
assign n_30927 = n_30918 ^ n_29210;
assign n_30928 = n_30919 & ~n_30915;
assign n_30929 = n_30919 ^ x473;
assign n_30930 = n_30917 & n_30920;
assign n_30931 = n_30906 ^ n_30921;
assign n_30932 = n_30923 ^ n_30912;
assign n_30933 = n_30922 & ~n_30924;
assign n_30934 = n_30925 ^ n_28912;
assign n_30935 = n_30916 ^ n_30925;
assign n_30936 = n_30927 ^ n_30893;
assign n_30937 = n_30928 ^ x473;
assign n_30938 = ~n_30929 & ~n_30905;
assign n_30939 = n_30905 ^ n_30929;
assign n_30940 = n_30930 ^ n_30330;
assign n_30941 = n_29725 & n_30931;
assign n_30942 = n_30910 & n_30932;
assign n_30943 = n_30933 ^ x173;
assign n_30944 = n_30916 ^ n_30934;
assign n_30945 = n_30926 & ~n_30935;
assign n_30946 = n_30936 ^ x472;
assign n_30947 = n_30939 ^ n_30343;
assign n_30948 = n_30939 ^ n_30940;
assign n_30949 = n_30940 ^ n_30343;
assign n_30950 = n_30941 ^ n_30330;
assign n_30951 = n_30944 ^ x172;
assign n_30952 = n_30943 ^ n_30944;
assign n_30953 = n_30945 ^ n_28912;
assign n_30954 = n_30937 ^ n_30946;
assign n_30955 = n_30947 & ~n_30948;
assign n_30956 = n_30939 ^ n_30949;
assign n_30957 = n_30950 ^ n_28953;
assign n_30958 = n_30943 ^ n_30951;
assign n_30959 = n_30951 & ~n_30952;
assign n_30960 = n_30950 ^ n_30953;
assign n_30961 = n_30954 ^ n_30938;
assign n_30962 = n_30955 ^ n_30343;
assign n_30963 = n_29738 & ~n_30956;
assign n_30964 = n_30957 ^ n_30953;
assign n_30965 = n_30942 ^ n_30958;
assign n_30966 = n_30958 & n_30942;
assign n_30967 = n_30959 ^ x172;
assign n_30968 = ~n_30957 & n_30960;
assign n_30969 = n_30961 ^ n_30363;
assign n_30970 = n_30961 ^ n_30962;
assign n_30971 = n_30963 ^ n_30343;
assign n_30972 = n_30964 ^ x171;
assign n_30973 = n_30965 ^ n_30487;
assign n_30974 = n_30487 & n_30965;
assign n_30975 = n_30965 ^ n_30479;
assign n_30976 = n_30964 ^ n_30967;
assign n_30977 = n_30968 ^ n_28953;
assign n_30978 = n_30969 ^ n_30962;
assign n_30979 = ~n_30969 & ~n_30970;
assign n_30980 = n_30971 ^ n_28991;
assign n_30981 = n_30972 ^ n_30967;
assign n_30982 = n_29984 & ~n_30973;
assign n_30983 = n_30974 ^ n_30511;
assign n_30984 = ~n_30972 & n_30976;
assign n_30985 = n_30971 ^ n_30977;
assign n_30986 = n_29763 & n_30978;
assign n_30987 = n_30979 ^ n_30363;
assign n_30988 = n_30980 ^ n_30977;
assign n_30989 = ~n_30981 & n_30966;
assign n_30990 = n_30966 ^ n_30981;
assign n_30991 = n_30486 ^ n_30982;
assign n_30992 = n_30982 ^ n_30487;
assign n_30993 = n_30984 ^ x171;
assign n_30994 = n_30980 & n_30985;
assign n_30995 = n_30986 ^ n_30363;
assign n_30996 = n_30987 ^ n_30383;
assign n_30997 = n_30389 ^ n_30987;
assign n_30998 = n_30988 ^ x170;
assign n_30999 = n_30990 ^ n_30974;
assign n_31000 = n_30990 ^ n_30983;
assign n_31001 = n_30991 ^ x391;
assign n_31002 = x391 & ~n_30991;
assign n_31003 = n_29446 & ~n_30992;
assign n_31004 = n_30993 ^ n_30988;
assign n_31005 = n_30994 ^ n_28991;
assign n_31006 = n_30995 ^ n_29032;
assign n_31007 = ~n_30389 & ~n_30996;
assign n_31008 = ~n_29775 & ~n_30997;
assign n_31009 = n_30983 & n_30999;
assign n_31010 = n_30005 & n_31000;
assign n_31011 = n_31002 ^ x390;
assign n_31012 = n_31003 ^ n_29478;
assign n_31013 = ~n_31004 & n_30998;
assign n_31014 = n_31004 ^ x170;
assign n_31015 = n_30995 ^ n_31005;
assign n_31016 = n_31005 ^ n_29032;
assign n_31017 = n_31007 ^ n_30014;
assign n_31018 = n_31008 ^ n_30383;
assign n_31019 = n_31009 ^ n_30511;
assign n_31020 = n_31010 ^ n_30511;
assign n_31021 = n_31013 ^ x170;
assign n_31022 = ~n_30989 & ~n_31014;
assign n_31023 = n_31014 ^ n_30989;
assign n_31024 = ~n_31006 & n_31015;
assign n_31025 = n_30995 ^ n_31016;
assign n_31026 = n_30063 ^ n_31017;
assign n_31027 = n_31017 ^ n_30406;
assign n_31028 = n_31018 ^ n_29066;
assign n_31029 = n_31020 ^ n_31003;
assign n_31030 = n_31020 ^ n_31012;
assign n_31031 = n_31019 ^ n_31023;
assign n_31032 = n_31023 ^ n_30552;
assign n_31033 = n_31024 ^ n_29032;
assign n_31034 = n_31025 ^ x169;
assign n_31035 = n_31025 ^ n_31021;
assign n_31036 = n_31026 ^ n_30406;
assign n_31037 = n_30413 & n_31027;
assign n_31038 = n_31012 & n_31029;
assign n_31039 = n_31030 ^ n_31002;
assign n_31040 = n_31030 ^ n_31011;
assign n_31041 = n_31031 ^ n_30552;
assign n_31042 = n_31031 & ~n_31032;
assign n_31043 = n_31018 ^ n_31033;
assign n_31044 = n_31033 ^ n_29066;
assign n_31045 = n_31034 ^ n_31021;
assign n_31046 = n_31034 & ~n_31035;
assign n_31047 = n_29802 & ~n_31036;
assign n_31048 = n_31037 ^ n_30063;
assign n_31049 = n_31038 ^ n_29478;
assign n_31050 = n_31011 & n_31039;
assign n_31051 = n_31001 & n_31040;
assign n_31052 = n_31040 ^ n_31001;
assign n_31053 = ~n_30046 & n_31041;
assign n_31054 = n_31042 ^ n_30552;
assign n_31055 = n_31028 & n_31043;
assign n_31056 = n_31018 ^ n_31044;
assign n_31057 = ~n_31022 & n_31045;
assign n_31058 = n_31045 ^ n_31022;
assign n_31059 = n_31046 ^ x169;
assign n_31060 = n_31047 ^ n_30406;
assign n_31061 = n_30119 ^ n_31048;
assign n_31062 = n_31048 ^ n_30420;
assign n_31063 = n_31050 ^ x390;
assign n_31064 = n_31053 ^ n_30552;
assign n_31065 = n_31055 ^ n_29066;
assign n_31066 = n_31056 ^ x168;
assign n_31067 = n_31058 ^ n_30587;
assign n_31068 = n_31054 ^ n_31058;
assign n_31069 = n_31056 ^ n_31059;
assign n_31070 = n_31060 ^ n_29105;
assign n_31071 = n_31061 ^ n_30420;
assign n_31072 = n_30426 & ~n_31062;
assign n_31073 = n_31064 ^ n_31049;
assign n_31074 = n_31064 ^ n_29514;
assign n_31075 = n_31060 ^ n_31065;
assign n_31076 = n_31066 ^ n_31059;
assign n_31077 = n_31054 ^ n_31067;
assign n_31078 = ~n_31067 & n_31068;
assign n_31079 = ~n_31066 & n_31069;
assign n_31080 = n_31070 ^ n_31065;
assign n_31081 = n_29816 & n_31071;
assign n_31082 = n_31072 ^ n_30119;
assign n_31083 = n_31073 ^ n_29514;
assign n_31084 = n_31073 & n_31074;
assign n_31085 = ~n_31070 & ~n_31075;
assign n_31086 = ~n_31057 & n_31076;
assign n_31087 = n_31076 ^ n_31057;
assign n_31088 = ~n_30087 & n_31077;
assign n_31089 = n_31078 ^ n_30587;
assign n_31090 = n_31079 ^ x168;
assign n_31091 = n_31080 ^ x183;
assign n_31092 = n_31081 ^ n_30420;
assign n_31093 = n_31082 ^ n_30446;
assign n_31094 = n_31083 ^ x389;
assign n_31095 = n_31063 ^ n_31083;
assign n_31096 = n_31084 ^ n_29514;
assign n_31097 = n_31085 ^ n_29105;
assign n_31098 = n_31087 ^ n_30627;
assign n_31099 = n_31088 ^ n_30587;
assign n_31100 = n_31089 ^ n_31087;
assign n_31101 = n_31080 ^ n_31090;
assign n_31102 = n_31091 ^ n_31090;
assign n_31103 = n_31092 ^ n_29147;
assign n_31104 = n_31093 & n_30453;
assign n_31105 = n_31093 ^ n_30175;
assign n_31106 = n_31063 ^ n_31094;
assign n_31107 = n_31094 & ~n_31095;
assign n_31108 = n_31097 ^ n_31092;
assign n_31109 = n_31099 ^ n_29543;
assign n_31110 = n_31096 ^ n_31099;
assign n_31111 = ~n_31100 & ~n_31098;
assign n_31112 = n_31100 ^ n_30627;
assign n_31113 = ~n_31091 & n_31101;
assign n_31114 = n_31102 ^ n_31086;
assign n_31115 = n_31086 & n_31102;
assign n_31116 = n_31104 ^ n_30175;
assign n_31117 = ~n_29837 & n_31105;
assign n_31118 = ~n_31051 & n_31106;
assign n_31119 = n_31106 ^ n_31051;
assign n_31120 = n_31107 ^ x389;
assign n_31121 = n_31108 ^ n_29147;
assign n_31122 = n_31108 & n_31103;
assign n_31123 = n_31096 ^ n_31109;
assign n_31124 = ~n_31109 & ~n_31110;
assign n_31125 = n_31111 ^ n_30627;
assign n_31126 = n_30123 & n_31112;
assign n_31127 = n_31113 ^ x183;
assign n_31128 = n_31114 ^ n_30668;
assign n_31129 = n_31116 ^ n_30466;
assign n_31130 = n_31117 ^ n_30446;
assign n_31131 = n_31120 ^ x388;
assign n_31132 = n_31121 ^ x182;
assign n_31133 = n_31122 ^ n_29147;
assign n_31134 = n_31120 ^ n_31123;
assign n_31135 = n_31124 ^ n_29543;
assign n_31136 = n_31125 ^ n_31114;
assign n_31137 = n_31126 ^ n_30627;
assign n_31138 = n_31127 ^ n_31121;
assign n_31139 = n_31125 ^ n_31128;
assign n_31140 = n_31129 & ~n_30474;
assign n_31141 = n_31129 ^ n_30214;
assign n_31142 = n_31130 ^ n_29189;
assign n_31143 = n_31130 ^ n_31133;
assign n_31144 = n_31133 ^ n_29189;
assign n_31145 = ~n_31134 & n_31131;
assign n_31146 = n_31134 ^ x388;
assign n_31147 = ~n_31128 & ~n_31136;
assign n_31148 = n_31137 ^ n_29572;
assign n_31149 = n_31135 ^ n_31137;
assign n_31150 = n_31138 ^ x182;
assign n_31151 = n_31138 & ~n_31132;
assign n_31152 = n_30160 & ~n_31139;
assign n_31153 = n_31140 ^ n_30214;
assign n_31154 = ~n_29856 & n_31141;
assign n_31155 = n_31142 & n_31143;
assign n_31156 = n_31130 ^ n_31144;
assign n_31157 = n_31145 ^ x388;
assign n_31158 = n_31146 & n_31118;
assign n_31159 = n_31118 ^ n_31146;
assign n_31160 = n_31147 ^ n_30668;
assign n_31161 = n_31135 ^ n_31148;
assign n_31162 = ~n_31148 & ~n_31149;
assign n_31163 = n_31150 ^ n_31115;
assign n_31164 = n_31115 & n_31150;
assign n_31165 = n_31151 ^ x182;
assign n_31166 = n_31152 ^ n_30668;
assign n_31167 = n_31153 ^ n_30488;
assign n_31168 = n_30497 ^ n_31153;
assign n_31169 = n_31154 ^ n_30466;
assign n_31170 = n_31155 ^ n_29189;
assign n_31171 = n_31156 ^ x181;
assign n_31172 = n_31161 ^ x387;
assign n_31173 = n_31157 ^ n_31161;
assign n_31174 = n_31162 ^ n_29572;
assign n_31175 = n_31160 ^ n_31163;
assign n_31176 = n_31163 ^ n_30703;
assign n_31177 = n_31156 ^ n_31165;
assign n_31178 = n_31166 ^ n_29591;
assign n_31179 = n_30497 & ~n_31167;
assign n_31180 = n_29876 & ~n_31168;
assign n_31181 = n_31169 ^ n_29227;
assign n_31182 = n_31169 ^ n_31170;
assign n_31183 = n_31170 ^ n_29227;
assign n_31184 = n_31171 ^ n_31165;
assign n_31185 = n_31157 ^ n_31172;
assign n_31186 = ~n_31172 & n_31173;
assign n_31187 = n_31174 ^ n_31166;
assign n_31188 = n_31175 ^ n_30703;
assign n_31189 = n_31175 & ~n_31176;
assign n_31190 = n_31171 & ~n_31177;
assign n_31191 = n_31174 ^ n_31178;
assign n_31192 = n_31179 ^ n_30244;
assign n_31193 = n_31180 ^ n_30488;
assign n_31194 = ~n_31181 & n_31182;
assign n_31195 = n_31169 ^ n_31183;
assign n_31196 = ~n_31164 & n_31184;
assign n_31197 = n_31184 ^ n_31164;
assign n_31198 = ~n_31185 & n_31158;
assign n_31199 = n_31158 ^ n_31185;
assign n_31200 = n_31186 ^ x387;
assign n_31201 = ~n_31178 & ~n_31187;
assign n_31202 = n_31001 ^ n_31188;
assign n_31203 = n_30184 & n_31188;
assign n_31204 = n_31189 ^ n_30703;
assign n_31205 = n_31190 ^ x181;
assign n_31206 = n_31191 ^ x386;
assign n_31207 = n_31192 ^ n_30506;
assign n_31208 = n_30518 ^ n_31192;
assign n_31209 = n_31193 ^ n_29259;
assign n_31210 = n_31194 ^ n_29227;
assign n_31211 = n_31195 ^ x180;
assign n_31212 = n_31197 ^ n_30738;
assign n_31213 = n_31200 ^ n_31191;
assign n_31214 = n_31201 ^ n_29591;
assign n_31215 = n_31203 ^ n_30703;
assign n_31216 = n_31204 ^ n_31197;
assign n_31217 = n_31195 ^ n_31205;
assign n_31218 = n_31205 ^ x180;
assign n_31219 = n_31200 ^ n_31206;
assign n_31220 = n_30518 & n_31207;
assign n_31221 = n_31208 ^ n_30515;
assign n_31222 = ~n_29900 & ~n_31208;
assign n_31223 = n_31193 ^ n_31210;
assign n_31224 = n_31210 ^ n_29259;
assign n_31225 = n_31204 ^ n_31212;
assign n_31226 = n_31206 & ~n_31213;
assign n_31227 = n_31214 ^ n_31215;
assign n_31228 = n_31215 ^ n_29610;
assign n_31229 = n_31212 & n_31216;
assign n_31230 = n_31211 & ~n_31217;
assign n_31231 = n_31195 ^ n_31218;
assign n_31232 = n_31198 & n_31219;
assign n_31233 = n_31219 ^ n_31198;
assign n_31234 = n_31220 ^ n_30260;
assign n_31235 = n_31222 ^ n_30506;
assign n_31236 = n_31209 & ~n_31223;
assign n_31237 = n_31193 ^ n_31224;
assign n_31238 = ~n_30231 & ~n_31225;
assign n_31239 = n_31052 ^ n_31225;
assign n_31240 = n_31226 ^ x386;
assign n_31241 = n_31227 ^ n_29610;
assign n_31242 = n_31227 & ~n_31228;
assign n_31243 = n_31229 ^ n_30738;
assign n_31244 = n_31230 ^ x180;
assign n_31245 = n_31196 & n_31231;
assign n_31246 = n_31231 ^ n_31196;
assign n_31247 = n_31234 ^ n_30538;
assign n_31248 = n_30548 ^ n_31234;
assign n_31249 = n_31235 ^ n_29291;
assign n_31250 = n_31236 ^ n_29259;
assign n_31251 = n_31237 ^ x179;
assign n_31252 = n_31238 ^ n_30738;
assign n_31253 = n_31240 ^ n_31241;
assign n_31254 = n_31241 ^ x385;
assign n_31255 = n_31242 ^ n_29610;
assign n_31256 = n_31237 ^ n_31244;
assign n_31257 = n_31244 ^ x179;
assign n_31258 = n_31243 ^ n_31246;
assign n_31259 = n_31246 ^ n_30780;
assign n_31260 = n_30548 & n_31247;
assign n_31261 = ~n_29919 & n_31248;
assign n_31262 = n_30569 ^ n_31248;
assign n_31263 = n_31235 ^ n_31250;
assign n_31264 = n_31249 ^ n_31250;
assign n_31265 = n_31252 ^ n_29623;
assign n_31266 = n_31253 ^ x385;
assign n_31267 = n_31253 & ~n_31254;
assign n_31268 = n_31252 ^ n_31255;
assign n_31269 = ~n_31251 & n_31256;
assign n_31270 = n_31237 ^ n_31257;
assign n_31271 = n_31258 ^ n_30780;
assign n_31272 = n_31258 & n_31259;
assign n_31273 = n_31260 ^ n_30283;
assign n_31274 = n_31261 ^ n_30538;
assign n_31275 = n_31249 & n_31263;
assign n_31276 = n_31264 ^ x178;
assign n_31277 = n_31265 ^ n_31255;
assign n_31278 = ~n_31232 & n_31266;
assign n_31279 = n_31266 ^ n_31232;
assign n_31280 = n_31267 ^ x385;
assign n_31281 = ~n_31268 & n_31265;
assign n_31282 = n_31269 ^ x179;
assign n_31283 = ~n_31245 & n_31270;
assign n_31284 = n_31270 ^ n_31245;
assign n_31285 = ~n_30255 & n_31271;
assign n_31286 = n_31119 ^ n_31271;
assign n_31287 = n_31272 ^ n_30780;
assign n_31288 = n_31273 ^ n_30572;
assign n_31289 = n_31274 ^ n_29311;
assign n_31290 = n_31275 ^ n_29291;
assign n_31291 = n_31277 ^ x384;
assign n_31292 = n_31280 ^ n_31277;
assign n_31293 = n_31281 ^ n_29623;
assign n_31294 = n_31264 ^ n_31282;
assign n_31295 = n_31276 ^ n_31282;
assign n_31296 = n_31284 ^ n_30813;
assign n_31297 = n_31285 ^ n_30780;
assign n_31298 = n_31287 ^ n_31284;
assign n_31299 = n_31288 & n_30583;
assign n_31300 = n_30304 ^ n_31288;
assign n_31301 = n_31290 ^ n_31274;
assign n_31302 = n_31280 ^ n_31291;
assign n_31303 = n_31291 & ~n_31292;
assign n_31304 = ~n_31276 & n_31294;
assign n_31305 = ~n_31283 & ~n_31295;
assign n_31306 = n_31295 ^ n_31283;
assign n_31307 = n_31287 ^ n_31296;
assign n_31308 = n_31297 ^ n_29647;
assign n_31309 = n_31293 ^ n_31297;
assign n_31310 = n_31296 & ~n_31298;
assign n_31311 = n_31299 ^ n_30304;
assign n_31312 = ~n_29941 & ~n_31300;
assign n_31313 = n_30637 ^ n_31300;
assign n_31314 = n_31301 & ~n_31289;
assign n_31315 = n_31301 ^ n_29311;
assign n_31316 = n_31278 & ~n_31302;
assign n_31317 = n_31302 ^ n_31278;
assign n_31318 = n_31303 ^ x384;
assign n_31319 = n_31304 ^ x178;
assign n_31320 = n_31306 ^ n_30848;
assign n_31321 = ~n_30273 & ~n_31307;
assign n_31322 = n_31159 ^ n_31307;
assign n_31323 = n_31293 ^ n_31308;
assign n_31324 = ~n_31308 & n_31309;
assign n_31325 = n_31310 ^ n_30813;
assign n_31326 = n_31311 ^ n_30605;
assign n_31327 = n_30618 ^ n_31311;
assign n_31328 = n_31312 ^ n_30572;
assign n_31329 = n_31314 ^ n_29311;
assign n_31330 = n_31315 ^ x177;
assign n_31331 = n_31319 ^ n_31315;
assign n_31332 = n_31321 ^ n_30813;
assign n_31333 = n_31323 ^ x399;
assign n_31334 = n_31318 ^ n_31323;
assign n_31335 = n_31324 ^ n_29647;
assign n_31336 = n_31325 ^ n_31306;
assign n_31337 = n_31325 ^ n_31320;
assign n_31338 = n_30618 & ~n_31326;
assign n_31339 = n_31327 ^ n_30675;
assign n_31340 = ~n_29955 & n_31327;
assign n_31341 = n_31328 ^ n_29325;
assign n_31342 = n_31329 ^ n_31328;
assign n_31343 = n_31331 & ~n_31330;
assign n_31344 = n_31331 ^ x177;
assign n_31345 = n_31332 ^ n_29666;
assign n_31346 = n_31318 ^ n_31333;
assign n_31347 = ~n_31333 & n_31334;
assign n_31348 = n_31335 ^ n_31332;
assign n_31349 = n_31320 & ~n_31336;
assign n_31350 = ~n_30288 & ~n_31337;
assign n_31351 = n_31199 ^ n_31337;
assign n_31352 = n_31338 ^ n_30322;
assign n_31353 = n_31340 ^ n_30605;
assign n_31354 = n_31329 ^ n_31341;
assign n_31355 = ~n_31341 & ~n_31342;
assign n_31356 = n_31343 ^ x177;
assign n_31357 = ~n_31344 & n_31305;
assign n_31358 = n_31305 ^ n_31344;
assign n_31359 = n_31335 ^ n_31345;
assign n_31360 = n_31316 & n_31346;
assign n_31361 = n_31346 ^ n_31316;
assign n_31362 = n_31347 ^ x399;
assign n_31363 = ~n_31345 & n_31348;
assign n_31364 = n_31349 ^ n_30848;
assign n_31365 = n_31350 ^ n_30848;
assign n_31366 = n_31352 ^ n_30656;
assign n_31367 = n_31352 ^ n_30338;
assign n_31368 = n_31353 ^ n_29346;
assign n_31369 = n_31354 ^ x176;
assign n_31370 = n_31355 ^ n_29325;
assign n_31371 = n_31356 ^ n_31354;
assign n_31372 = n_31356 ^ x176;
assign n_31373 = n_31358 ^ n_30895;
assign n_31374 = n_31359 ^ x398;
assign n_31375 = n_31362 ^ x398;
assign n_31376 = n_31359 ^ n_31362;
assign n_31377 = n_31363 ^ n_29666;
assign n_31378 = n_31358 ^ n_31364;
assign n_31379 = n_31365 ^ n_29686;
assign n_31380 = n_30670 & ~n_31366;
assign n_31381 = n_31367 ^ n_30656;
assign n_31382 = n_31370 ^ n_31353;
assign n_31383 = n_31370 ^ n_29346;
assign n_31384 = ~n_31369 & n_31371;
assign n_31385 = n_31372 ^ n_31354;
assign n_31386 = n_31373 ^ n_31364;
assign n_31387 = n_31374 ^ n_31362;
assign n_31388 = n_31375 & n_31376;
assign n_31389 = n_31377 ^ n_31365;
assign n_31390 = n_31373 & n_31378;
assign n_31391 = n_31377 ^ n_31379;
assign n_31392 = n_31380 ^ n_30338;
assign n_31393 = n_29982 & n_31381;
assign n_31394 = n_31381 ^ n_30714;
assign n_31395 = n_31368 & n_31382;
assign n_31396 = n_31383 ^ n_31353;
assign n_31397 = n_31384 ^ x176;
assign n_31398 = ~n_31357 & n_31385;
assign n_31399 = n_31385 ^ n_31357;
assign n_31400 = ~n_30307 & ~n_31386;
assign n_31401 = n_31233 ^ n_31386;
assign n_31402 = ~n_31387 & ~n_31360;
assign n_31403 = n_31360 ^ n_31387;
assign n_31404 = n_31388 ^ x398;
assign n_31405 = n_31379 & n_31389;
assign n_31406 = n_31390 ^ n_30895;
assign n_31407 = n_31391 ^ x397;
assign n_31408 = n_31392 ^ n_30695;
assign n_31409 = n_31392 ^ n_30707;
assign n_31410 = n_31393 ^ n_30656;
assign n_31411 = n_31395 ^ n_29346;
assign n_31412 = n_31396 ^ x191;
assign n_31413 = n_31397 ^ n_31396;
assign n_31414 = n_31399 ^ n_30931;
assign n_31415 = n_31400 ^ n_30895;
assign n_31416 = n_31404 ^ n_31391;
assign n_31417 = n_31405 ^ n_29686;
assign n_31418 = n_31406 ^ n_31399;
assign n_31419 = n_31404 ^ n_31407;
assign n_31420 = n_30707 & n_31408;
assign n_31421 = n_30757 ^ n_31409;
assign n_31422 = ~n_29999 & n_31409;
assign n_31423 = n_31410 ^ n_29371;
assign n_31424 = n_31411 ^ n_29371;
assign n_31425 = n_31410 ^ n_31411;
assign n_31426 = n_31397 ^ n_31412;
assign n_31427 = ~n_31412 & n_31413;
assign n_31428 = n_31406 ^ n_31414;
assign n_31429 = n_31415 ^ n_29701;
assign n_31430 = n_31407 & ~n_31416;
assign n_31431 = n_31415 ^ n_31417;
assign n_31432 = ~n_31414 & n_31418;
assign n_31433 = n_31419 & n_31402;
assign n_31434 = n_31402 ^ n_31419;
assign n_31435 = n_31420 ^ n_30361;
assign n_31436 = n_31422 ^ n_30695;
assign n_31437 = n_31423 ^ n_31411;
assign n_31438 = ~n_31424 & ~n_31425;
assign n_31439 = ~n_31398 & ~n_31426;
assign n_31440 = n_31426 ^ n_31398;
assign n_31441 = n_31427 ^ x191;
assign n_31442 = n_30330 & ~n_31428;
assign n_31443 = n_31279 ^ n_31428;
assign n_31444 = n_31430 ^ x397;
assign n_31445 = n_31431 & ~n_31429;
assign n_31446 = n_31431 ^ n_29701;
assign n_31447 = n_31432 ^ n_30931;
assign n_31448 = n_31435 ^ n_30722;
assign n_31449 = n_31435 ^ n_30736;
assign n_31450 = n_31436 ^ n_29386;
assign n_31451 = n_31437 ^ x190;
assign n_31452 = n_31438 ^ n_29371;
assign n_31453 = n_31440 ^ n_30956;
assign n_31454 = n_31441 ^ n_31437;
assign n_31455 = n_31441 ^ x190;
assign n_31456 = n_31442 ^ n_30931;
assign n_31457 = n_31444 ^ x396;
assign n_31458 = n_31445 ^ n_29701;
assign n_31459 = n_31446 ^ x396;
assign n_31460 = n_31444 ^ n_31446;
assign n_31461 = n_31447 ^ n_31440;
assign n_31462 = n_31447 ^ n_30956;
assign n_31463 = n_30736 & n_31448;
assign n_31464 = n_30796 ^ n_31449;
assign n_31465 = ~n_30041 & ~n_31449;
assign n_31466 = n_31452 ^ n_31436;
assign n_31467 = n_31452 ^ n_31450;
assign n_31468 = ~n_31451 & n_31454;
assign n_31469 = n_31455 ^ n_31437;
assign n_31470 = n_31456 ^ n_29725;
assign n_31471 = n_31457 ^ n_31446;
assign n_31472 = n_31458 ^ n_31456;
assign n_31473 = n_31459 & ~n_31460;
assign n_31474 = n_31453 & n_31461;
assign n_31475 = n_31462 ^ n_31440;
assign n_31476 = n_31463 ^ n_30381;
assign n_31477 = n_31465 ^ n_30722;
assign n_31478 = n_31450 & ~n_31466;
assign n_31479 = n_31467 ^ x189;
assign n_31480 = n_31468 ^ x190;
assign n_31481 = n_31439 & ~n_31469;
assign n_31482 = n_31469 ^ n_31439;
assign n_31483 = n_31458 ^ n_31470;
assign n_31484 = ~n_31433 & ~n_31471;
assign n_31485 = n_31471 ^ n_31433;
assign n_31486 = n_31470 & n_31472;
assign n_31487 = n_31473 ^ x396;
assign n_31488 = n_31474 ^ n_30956;
assign n_31489 = n_30343 & n_31475;
assign n_31490 = n_31317 ^ n_31475;
assign n_31491 = n_31476 ^ n_30788;
assign n_31492 = n_31476 ^ n_30774;
assign n_31493 = n_31477 ^ n_29407;
assign n_31494 = n_31478 ^ n_29386;
assign n_31495 = n_31480 ^ x189;
assign n_31496 = n_31467 ^ n_31480;
assign n_31497 = n_31479 ^ n_31480;
assign n_31498 = n_31482 ^ n_30978;
assign n_31499 = n_31483 ^ x395;
assign n_31500 = n_31486 ^ n_29725;
assign n_31501 = n_31487 ^ n_31483;
assign n_31502 = n_31487 ^ x395;
assign n_31503 = n_31488 ^ n_31482;
assign n_31504 = n_31489 ^ n_30956;
assign n_31505 = n_30837 ^ n_31491;
assign n_31506 = n_30067 & n_31491;
assign n_31507 = n_30788 & n_31492;
assign n_31508 = n_31494 ^ n_31477;
assign n_31509 = n_31494 ^ n_31493;
assign n_31510 = n_31495 & n_31496;
assign n_31511 = n_31497 & ~n_31481;
assign n_31512 = n_31481 ^ n_31497;
assign n_31513 = n_31488 ^ n_31498;
assign n_31514 = ~n_31499 & n_31501;
assign n_31515 = n_31502 ^ n_31483;
assign n_31516 = n_31498 & n_31503;
assign n_31517 = n_31504 ^ n_29738;
assign n_31518 = n_31500 ^ n_31504;
assign n_31519 = n_31506 ^ n_30774;
assign n_31520 = n_31507 ^ n_30399;
assign n_31521 = ~n_31493 & n_31508;
assign n_31522 = n_31509 ^ x188;
assign n_31523 = n_31510 ^ x189;
assign n_31524 = n_31512 ^ n_30997;
assign n_31525 = ~n_30363 & ~n_31513;
assign n_31526 = n_31361 ^ n_31513;
assign n_31527 = n_31514 ^ x395;
assign n_31528 = n_31484 & n_31515;
assign n_31529 = n_31515 ^ n_31484;
assign n_31530 = n_31516 ^ n_30978;
assign n_31531 = n_31500 ^ n_31517;
assign n_31532 = ~n_31517 & n_31518;
assign n_31533 = n_31519 ^ n_29430;
assign n_31534 = n_31520 ^ n_30816;
assign n_31535 = n_31520 ^ n_30802;
assign n_31536 = n_31521 ^ n_29407;
assign n_31537 = n_31523 ^ x188;
assign n_31538 = n_31509 ^ n_31523;
assign n_31539 = n_31522 ^ n_31523;
assign n_31540 = n_31525 ^ n_30978;
assign n_31541 = n_31530 ^ n_31512;
assign n_31542 = n_31530 ^ n_31524;
assign n_31543 = n_31527 ^ n_31531;
assign n_31544 = n_31531 ^ x394;
assign n_31545 = n_31532 ^ n_29738;
assign n_31546 = ~n_30113 & n_31534;
assign n_31547 = n_30876 ^ n_31534;
assign n_31548 = ~n_30816 & ~n_31535;
assign n_31549 = n_31536 ^ n_31519;
assign n_31550 = n_31536 ^ n_31533;
assign n_31551 = n_31537 & ~n_31538;
assign n_31552 = ~n_31539 & n_31511;
assign n_31553 = n_31511 ^ n_31539;
assign n_31554 = n_31540 ^ n_29763;
assign n_31555 = n_31524 & n_31541;
assign n_31556 = ~n_30383 & n_31542;
assign n_31557 = n_31403 ^ n_31542;
assign n_31558 = n_31543 ^ x394;
assign n_31559 = n_31543 & ~n_31544;
assign n_31560 = n_31545 ^ n_31540;
assign n_31561 = n_31545 ^ n_29763;
assign n_31562 = n_31546 ^ n_30802;
assign n_31563 = n_31548 ^ n_30417;
assign n_31564 = ~n_31533 & ~n_31549;
assign n_31565 = n_31550 ^ x187;
assign n_31566 = n_31551 ^ x188;
assign n_31567 = n_31553 ^ n_31036;
assign n_31568 = n_31555 ^ n_30997;
assign n_31569 = n_31556 ^ n_30997;
assign n_31570 = ~n_31528 & ~n_31558;
assign n_31571 = n_31558 ^ n_31528;
assign n_31572 = n_31559 ^ x394;
assign n_31573 = n_31554 & ~n_31560;
assign n_31574 = n_31561 ^ n_31540;
assign n_31575 = n_31562 ^ n_29452;
assign n_31576 = n_30866 ^ n_31563;
assign n_31577 = n_31563 ^ n_30854;
assign n_31578 = n_30438 ^ n_31563;
assign n_31579 = n_31564 ^ n_29430;
assign n_31580 = n_31566 ^ x187;
assign n_31581 = n_31550 ^ n_31566;
assign n_31582 = n_31565 ^ n_31566;
assign n_31583 = n_31568 ^ n_31553;
assign n_31584 = n_31568 ^ n_31567;
assign n_31585 = n_31569 ^ n_29775;
assign n_31586 = n_31573 ^ n_29763;
assign n_31587 = n_31574 ^ x393;
assign n_31588 = n_31572 ^ n_31574;
assign n_31589 = ~n_30152 & n_31576;
assign n_31590 = n_30911 ^ n_31576;
assign n_31591 = ~n_31577 & n_31578;
assign n_31592 = n_31579 ^ n_29452;
assign n_31593 = n_31579 ^ n_31562;
assign n_31594 = n_31580 & ~n_31581;
assign n_31595 = ~n_31582 & n_31552;
assign n_31596 = n_31552 ^ n_31582;
assign n_31597 = n_31567 & ~n_31583;
assign n_31598 = ~n_30406 & ~n_31584;
assign n_31599 = n_31434 ^ n_31584;
assign n_31600 = n_31586 ^ n_31569;
assign n_31601 = n_31572 ^ n_31587;
assign n_31602 = n_31587 & ~n_31588;
assign n_31603 = n_31589 ^ n_30854;
assign n_31604 = n_30894 ^ n_31591;
assign n_31605 = n_31592 ^ n_31562;
assign n_31606 = ~n_31575 & n_31593;
assign n_31607 = n_31594 ^ x187;
assign n_31608 = n_31596 ^ n_31071;
assign n_31609 = n_31597 ^ n_31036;
assign n_31610 = n_31598 ^ n_31036;
assign n_31611 = n_31600 & n_31585;
assign n_31612 = n_31600 ^ n_29775;
assign n_31613 = ~n_31570 & ~n_31601;
assign n_31614 = n_31601 ^ n_31570;
assign n_31615 = n_31602 ^ x393;
assign n_31616 = n_31603 ^ n_29471;
assign n_31617 = ~n_30179 & n_31604;
assign n_31618 = n_31604 ^ n_30910;
assign n_31619 = n_31605 ^ x186;
assign n_31620 = n_31606 ^ n_29452;
assign n_31621 = n_31607 ^ x186;
assign n_31622 = n_31605 ^ n_31607;
assign n_31623 = n_31609 ^ n_31596;
assign n_31624 = n_31610 ^ n_29802;
assign n_31625 = n_31611 ^ n_29775;
assign n_31626 = n_31612 ^ x392;
assign n_31627 = n_31615 ^ n_31612;
assign n_31628 = n_31615 ^ x392;
assign n_31629 = n_31617 ^ n_30867;
assign n_31630 = n_31618 ^ n_30932;
assign n_31631 = n_31619 ^ n_31607;
assign n_31632 = n_31620 ^ n_31616;
assign n_31633 = n_31620 ^ n_31603;
assign n_31634 = n_31621 & n_31622;
assign n_31635 = ~n_31623 & ~n_31608;
assign n_31636 = n_31623 ^ n_31071;
assign n_31637 = n_31625 ^ n_31610;
assign n_31638 = n_31625 ^ n_31624;
assign n_31639 = n_31626 & ~n_31627;
assign n_31640 = n_31628 ^ n_31612;
assign n_31641 = n_31630 ^ n_30911;
assign n_31642 = n_31631 & n_31595;
assign n_31643 = n_31595 ^ n_31631;
assign n_31644 = n_31632 ^ x185;
assign n_31645 = ~n_31616 & n_31633;
assign n_31646 = n_31634 ^ x186;
assign n_31647 = n_31635 ^ n_31071;
assign n_31648 = ~n_30420 & n_31636;
assign n_31649 = n_31485 ^ n_31636;
assign n_31650 = ~n_31624 & ~n_31637;
assign n_31651 = n_31638 ^ x407;
assign n_31652 = n_31639 ^ x392;
assign n_31653 = ~n_31613 & n_31640;
assign n_31654 = n_31640 ^ n_31613;
assign n_31655 = n_31643 ^ n_31105;
assign n_31656 = n_31645 ^ n_29471;
assign n_31657 = n_31644 ^ n_31646;
assign n_31658 = n_31646 ^ x185;
assign n_31659 = n_31632 ^ n_31646;
assign n_31660 = n_31647 ^ n_31643;
assign n_31661 = n_31648 ^ n_31071;
assign n_31662 = n_31650 ^ n_29802;
assign n_31663 = n_31652 ^ n_31638;
assign n_31664 = n_31652 ^ x407;
assign n_31665 = n_31647 ^ n_31655;
assign n_31666 = n_31656 ^ n_29494;
assign n_31667 = n_31642 & n_31657;
assign n_31668 = n_31657 ^ n_31642;
assign n_31669 = n_31658 & n_31659;
assign n_31670 = n_31655 & ~n_31660;
assign n_31671 = n_31661 ^ n_29816;
assign n_31672 = n_31662 ^ n_31661;
assign n_31673 = n_31662 ^ n_29816;
assign n_31674 = n_31651 & ~n_31663;
assign n_31675 = n_31664 ^ n_31638;
assign n_31676 = n_30446 & n_31665;
assign n_31677 = n_31529 ^ n_31665;
assign n_31678 = n_31666 ^ n_31629;
assign n_31679 = n_31668 ^ n_31141;
assign n_31680 = n_31669 ^ x185;
assign n_31681 = n_31670 ^ n_31105;
assign n_31682 = n_31671 & ~n_31672;
assign n_31683 = n_31673 ^ n_31661;
assign n_31684 = n_31674 ^ x407;
assign n_31685 = ~n_31653 & ~n_31675;
assign n_31686 = n_31675 ^ n_31653;
assign n_31687 = n_31676 ^ n_31105;
assign n_31688 = n_31678 ^ x184;
assign n_31689 = n_31681 ^ n_31668;
assign n_31690 = n_31681 ^ n_31141;
assign n_31691 = n_31682 ^ n_29816;
assign n_31692 = n_31683 ^ x406;
assign n_31693 = n_31684 ^ n_31683;
assign n_31694 = n_31687 ^ n_29837;
assign n_31695 = n_31680 ^ n_31688;
assign n_31696 = n_31679 & ~n_31689;
assign n_31697 = n_31690 ^ n_31668;
assign n_31698 = n_31691 ^ n_31687;
assign n_31699 = n_31691 ^ n_29837;
assign n_31700 = n_31684 ^ n_31692;
assign n_31701 = n_31692 & ~n_31693;
assign n_31702 = n_31667 ^ n_31695;
assign n_31703 = n_31696 ^ n_31141;
assign n_31704 = ~n_30466 & n_31697;
assign n_31705 = n_31571 ^ n_31697;
assign n_31706 = ~n_31694 & ~n_31698;
assign n_31707 = n_31699 ^ n_31687;
assign n_31708 = n_31685 & ~n_31700;
assign n_31709 = n_31700 ^ n_31685;
assign n_31710 = n_31701 ^ x406;
assign n_31711 = n_31702 ^ n_31168;
assign n_31712 = n_31703 ^ n_31702;
assign n_31713 = n_31704 ^ n_31141;
assign n_31714 = n_31706 ^ n_29837;
assign n_31715 = n_31707 ^ x405;
assign n_31716 = n_31710 ^ n_31707;
assign n_31717 = n_31703 ^ n_31711;
assign n_31718 = ~n_31711 & ~n_31712;
assign n_31719 = n_31713 ^ n_29856;
assign n_31720 = n_31714 ^ n_31713;
assign n_31721 = n_31710 ^ n_31715;
assign n_31722 = ~n_31715 & n_31716;
assign n_31723 = n_30488 & ~n_31717;
assign n_31724 = n_31614 ^ n_31717;
assign n_31725 = n_31718 ^ n_31168;
assign n_31726 = n_31714 ^ n_31719;
assign n_31727 = ~n_31719 & n_31720;
assign n_31728 = ~n_31721 & ~n_31708;
assign n_31729 = n_31708 ^ n_31721;
assign n_31730 = n_31722 ^ x405;
assign n_31731 = n_31723 ^ n_31168;
assign n_31732 = n_31725 ^ n_31208;
assign n_31733 = n_31725 ^ n_31221;
assign n_31734 = n_31726 ^ x404;
assign n_31735 = n_31727 ^ n_29856;
assign n_31736 = n_31730 ^ n_31726;
assign n_31737 = n_31730 ^ x404;
assign n_31738 = n_31731 ^ n_29876;
assign n_31739 = ~n_31221 & ~n_31732;
assign n_31740 = ~n_30506 & n_31733;
assign n_31741 = n_31654 ^ n_31733;
assign n_31742 = n_31735 ^ n_31731;
assign n_31743 = n_31734 & ~n_31736;
assign n_31744 = n_31737 ^ n_31726;
assign n_31745 = n_31735 ^ n_31738;
assign n_31746 = n_31739 ^ n_30515;
assign n_31747 = n_31740 ^ n_31208;
assign n_31748 = ~n_31738 & ~n_31742;
assign n_31749 = n_31743 ^ x404;
assign n_31750 = ~n_31728 & ~n_31744;
assign n_31751 = n_31744 ^ n_31728;
assign n_31752 = n_31745 ^ x403;
assign n_31753 = n_31746 ^ n_31248;
assign n_31754 = n_31747 ^ n_29900;
assign n_31755 = n_31748 ^ n_29876;
assign n_31756 = n_31749 ^ n_31745;
assign n_31757 = ~n_31753 & n_31262;
assign n_31758 = n_30569 ^ n_31753;
assign n_31759 = n_31755 ^ n_31747;
assign n_31760 = n_31755 ^ n_31754;
assign n_31761 = ~n_31756 & n_31752;
assign n_31762 = n_31756 ^ x403;
assign n_31763 = n_31757 ^ n_30569;
assign n_31764 = n_30538 & n_31758;
assign n_31765 = n_31686 ^ n_31758;
assign n_31766 = n_31754 & n_31759;
assign n_31767 = n_31760 ^ x402;
assign n_31768 = n_31761 ^ x403;
assign n_31769 = ~n_31762 & n_31750;
assign n_31770 = n_31750 ^ n_31762;
assign n_31771 = n_31763 ^ n_31300;
assign n_31772 = n_31764 ^ n_31248;
assign n_31773 = n_31766 ^ n_29900;
assign n_31774 = n_31768 ^ n_31760;
assign n_31775 = n_31768 ^ n_31767;
assign n_31776 = n_31771 & n_31313;
assign n_31777 = n_30637 ^ n_31771;
assign n_31778 = n_31772 ^ n_29919;
assign n_31779 = n_31773 ^ n_31772;
assign n_31780 = n_31773 ^ n_29919;
assign n_31781 = n_31767 & ~n_31774;
assign n_31782 = ~n_31769 & n_31775;
assign n_31783 = n_31775 ^ n_31769;
assign n_31784 = n_31776 ^ n_30637;
assign n_31785 = ~n_30572 & n_31777;
assign n_31786 = n_31709 ^ n_31777;
assign n_31787 = ~n_31778 & n_31779;
assign n_31788 = n_31780 ^ n_31772;
assign n_31789 = n_31781 ^ x402;
assign n_31790 = n_31784 ^ n_31327;
assign n_31791 = n_31784 ^ n_31339;
assign n_31792 = n_31785 ^ n_31300;
assign n_31793 = n_31787 ^ n_29919;
assign n_31794 = n_31788 ^ x401;
assign n_31795 = n_31789 ^ n_31788;
assign n_31796 = ~n_31339 & n_31790;
assign n_31797 = ~n_30605 & n_31791;
assign n_31798 = n_31729 ^ n_31791;
assign n_31799 = n_31792 ^ n_29941;
assign n_31800 = n_31793 ^ n_31792;
assign n_31801 = n_31793 ^ n_29941;
assign n_31802 = ~n_31795 & n_31794;
assign n_31803 = n_31795 ^ x401;
assign n_31804 = n_31796 ^ n_30675;
assign n_31805 = n_31797 ^ n_31327;
assign n_31806 = n_31799 & ~n_31800;
assign n_31807 = n_31801 ^ n_31792;
assign n_31808 = n_31802 ^ x401;
assign n_31809 = ~n_31782 & ~n_31803;
assign n_31810 = n_31803 ^ n_31782;
assign n_31811 = n_31804 ^ n_31381;
assign n_31812 = n_31805 ^ n_29955;
assign n_31813 = n_31806 ^ n_29941;
assign n_31814 = n_31807 ^ x400;
assign n_31815 = n_31808 ^ n_31807;
assign n_31816 = n_31811 & ~n_31394;
assign n_31817 = n_31811 ^ n_30714;
assign n_31818 = n_31813 ^ n_31805;
assign n_31819 = n_31813 ^ n_29955;
assign n_31820 = n_31815 & ~n_31814;
assign n_31821 = n_31815 ^ x400;
assign n_31822 = n_31816 ^ n_30714;
assign n_31823 = ~n_30656 & n_31817;
assign n_31824 = n_31751 ^ n_31817;
assign n_31825 = ~n_31812 & n_31818;
assign n_31826 = n_31819 ^ n_31805;
assign n_31827 = n_31820 ^ x400;
assign n_31828 = ~n_31809 & ~n_31821;
assign n_31829 = n_31821 ^ n_31809;
assign n_31830 = n_31822 ^ n_31409;
assign n_31831 = n_31421 ^ n_31822;
assign n_31832 = n_31823 ^ n_31381;
assign n_31833 = n_31825 ^ n_29955;
assign n_31834 = n_31826 ^ x415;
assign n_31835 = n_31827 ^ n_31826;
assign n_31836 = n_31421 & n_31830;
assign n_31837 = n_30695 & ~n_31831;
assign n_31838 = n_31770 ^ n_31831;
assign n_31839 = n_31832 ^ n_29982;
assign n_31840 = n_31833 ^ n_31832;
assign n_31841 = n_31833 ^ n_29982;
assign n_31842 = n_31827 ^ n_31834;
assign n_31843 = n_31834 & ~n_31835;
assign n_31844 = n_31836 ^ n_30757;
assign n_31845 = n_31837 ^ n_31409;
assign n_31846 = n_31839 & n_31840;
assign n_31847 = n_31841 ^ n_31832;
assign n_31848 = ~n_31828 & ~n_31842;
assign n_31849 = n_31842 ^ n_31828;
assign n_31850 = n_31843 ^ x415;
assign n_31851 = n_31844 ^ n_31449;
assign n_31852 = n_31464 ^ n_31844;
assign n_31853 = n_31845 ^ n_29999;
assign n_31854 = n_31846 ^ n_29982;
assign n_31855 = n_31847 ^ x414;
assign n_31856 = n_31850 ^ n_31847;
assign n_31857 = ~n_31464 & n_31851;
assign n_31858 = ~n_30722 & ~n_31852;
assign n_31859 = n_31783 ^ n_31852;
assign n_31860 = n_31845 ^ n_31854;
assign n_31861 = n_31853 ^ n_31854;
assign n_31862 = n_31850 ^ n_31855;
assign n_31863 = ~n_31855 & n_31856;
assign n_31864 = n_31857 ^ n_30796;
assign n_31865 = n_31858 ^ n_31449;
assign n_31866 = ~n_31853 & ~n_31860;
assign n_31867 = n_31861 ^ x413;
assign n_31868 = ~n_31848 & ~n_31862;
assign n_31869 = n_31863 ^ x414;
assign n_31870 = n_31864 ^ n_31491;
assign n_31871 = n_31505 ^ n_31864;
assign n_31872 = n_31865 ^ n_30041;
assign n_31873 = n_31866 ^ n_29999;
assign n_31874 = n_31869 ^ n_31861;
assign n_31875 = ~n_31505 & ~n_31870;
assign n_31876 = n_30774 & ~n_31871;
assign n_31877 = n_31810 ^ n_31871;
assign n_31878 = n_31865 ^ n_31873;
assign n_31879 = n_31873 ^ n_30041;
assign n_31880 = n_31874 & ~n_31867;
assign n_31881 = n_31874 ^ x413;
assign n_31882 = n_31875 ^ n_30837;
assign n_31883 = n_31876 ^ n_31491;
assign n_31884 = n_31872 & ~n_31878;
assign n_31885 = n_31865 ^ n_31879;
assign n_31886 = n_31880 ^ x413;
assign n_31887 = n_31881 & ~n_31868;
assign n_31888 = n_31868 ^ n_31881;
assign n_31889 = n_31882 ^ n_30876;
assign n_31890 = n_31882 ^ n_31534;
assign n_31891 = n_31883 ^ n_30067;
assign n_31892 = n_31884 ^ n_30041;
assign n_31893 = n_31885 ^ x412;
assign n_31894 = n_31885 ^ n_31886;
assign n_31895 = n_30973 & n_31888;
assign n_31896 = n_31888 ^ n_30973;
assign n_31897 = n_31888 ^ n_30965;
assign n_31898 = n_31889 ^ n_31534;
assign n_31899 = n_31547 & n_31890;
assign n_31900 = n_31883 ^ n_31892;
assign n_31901 = n_31892 ^ n_30067;
assign n_31902 = n_31893 ^ n_31886;
assign n_31903 = ~n_31893 & n_31894;
assign n_31904 = n_31895 ^ n_31000;
assign n_31905 = n_30487 & ~n_31896;
assign n_31906 = n_30802 & ~n_31898;
assign n_31907 = n_31829 ^ n_31898;
assign n_31908 = n_31899 ^ n_30876;
assign n_31909 = n_31891 & n_31900;
assign n_31910 = n_31883 ^ n_31901;
assign n_31911 = ~n_31887 & ~n_31902;
assign n_31912 = n_31902 ^ n_31887;
assign n_31913 = n_31903 ^ x412;
assign n_31914 = n_31905 ^ n_30973;
assign n_31915 = n_31905 ^ n_30975;
assign n_31916 = n_31906 ^ n_31534;
assign n_31917 = n_31590 ^ n_31908;
assign n_31918 = n_31908 ^ n_31576;
assign n_31919 = n_30911 ^ n_31908;
assign n_31920 = n_31909 ^ n_30067;
assign n_31921 = n_31910 ^ x411;
assign n_31922 = n_31912 ^ n_31895;
assign n_31923 = n_31912 ^ n_31904;
assign n_31924 = n_31910 ^ n_31913;
assign n_31925 = n_29984 & ~n_31914;
assign n_31926 = x103 & ~n_31915;
assign n_31927 = n_31915 ^ x103;
assign n_31928 = n_31916 ^ n_30113;
assign n_31929 = n_30854 & ~n_31917;
assign n_31930 = n_31849 ^ n_31917;
assign n_31931 = ~n_31918 & ~n_31919;
assign n_31932 = n_31916 ^ n_31920;
assign n_31933 = n_31921 ^ n_31913;
assign n_31934 = ~n_31904 & ~n_31922;
assign n_31935 = n_30511 & n_31923;
assign n_31936 = ~n_31921 & n_31924;
assign n_31937 = n_31925 ^ n_30005;
assign n_31938 = n_31926 ^ x102;
assign n_31939 = n_31929 ^ n_31576;
assign n_31940 = n_31641 ^ n_31931;
assign n_31941 = ~n_31932 & ~n_31928;
assign n_31942 = n_31932 ^ n_30113;
assign n_31943 = n_31911 & ~n_31933;
assign n_31944 = n_31933 ^ n_31911;
assign n_31945 = n_31934 ^ n_31000;
assign n_31946 = n_31935 ^ n_31000;
assign n_31947 = n_31936 ^ x411;
assign n_31948 = n_31939 ^ n_30152;
assign n_31949 = ~n_30867 & n_31940;
assign n_31950 = n_31940 ^ n_31862;
assign n_31951 = n_31941 ^ n_30113;
assign n_31952 = n_31942 ^ x410;
assign n_31953 = n_31944 ^ n_31041;
assign n_31954 = n_31945 ^ n_31944;
assign n_31955 = n_31945 ^ n_31041;
assign n_31956 = n_31946 ^ n_31925;
assign n_31957 = n_31946 ^ n_31937;
assign n_31958 = n_31942 ^ n_31947;
assign n_31959 = n_31949 ^ n_31604;
assign n_31960 = n_31950 ^ n_31848;
assign n_31961 = n_31951 ^ n_30152;
assign n_31962 = n_31951 ^ n_31939;
assign n_31963 = n_31952 ^ n_31947;
assign n_31964 = n_31953 & ~n_31954;
assign n_31965 = n_31955 ^ n_31944;
assign n_31966 = n_31937 & ~n_31956;
assign n_31967 = n_31957 ^ n_31926;
assign n_31968 = n_31957 ^ n_31938;
assign n_31969 = ~n_31952 & n_31958;
assign n_31970 = n_31959 ^ n_30179;
assign n_31971 = n_31960 ^ n_31917;
assign n_31972 = n_31961 ^ n_31939;
assign n_31973 = ~n_31948 & n_31962;
assign n_31974 = ~n_31943 & n_31963;
assign n_31975 = n_31963 ^ n_31943;
assign n_31976 = n_31964 ^ n_31041;
assign n_31977 = n_30552 & n_31965;
assign n_31978 = n_31966 ^ n_30005;
assign n_31979 = n_31938 & ~n_31967;
assign n_31980 = n_31969 ^ x410;
assign n_31981 = n_31972 ^ x409;
assign n_31982 = n_31973 ^ n_30152;
assign n_31983 = n_31975 ^ n_31077;
assign n_31984 = n_31976 ^ n_31975;
assign n_31985 = n_31977 ^ n_31041;
assign n_31986 = n_31979 ^ x102;
assign n_31987 = n_31972 ^ n_31980;
assign n_31988 = n_31980 ^ x409;
assign n_31989 = n_31982 ^ n_31970;
assign n_31990 = n_31983 ^ n_31976;
assign n_31991 = n_31984 & ~n_31983;
assign n_31992 = n_31985 ^ n_30046;
assign n_31993 = n_31978 ^ n_31985;
assign n_31994 = n_31986 ^ x101;
assign n_31995 = n_31981 & ~n_31987;
assign n_31996 = n_31972 ^ n_31988;
assign n_31997 = n_30587 & ~n_31990;
assign n_31998 = n_31991 ^ n_31077;
assign n_31999 = n_31978 ^ n_31992;
assign n_32000 = ~n_31992 & ~n_31993;
assign n_32001 = n_31995 ^ x409;
assign n_32002 = n_31974 & ~n_31996;
assign n_32003 = n_31996 ^ n_31974;
assign n_32004 = n_31997 ^ n_31077;
assign n_32005 = n_31999 ^ x101;
assign n_32006 = n_31986 ^ n_31999;
assign n_32007 = n_31994 ^ n_31999;
assign n_32008 = n_32000 ^ n_30046;
assign n_32009 = n_32001 ^ n_31989;
assign n_32010 = n_31998 ^ n_32003;
assign n_32011 = n_32003 ^ n_31112;
assign n_32012 = n_32004 ^ n_30087;
assign n_32013 = ~n_32005 & n_32006;
assign n_32014 = n_31968 & ~n_32007;
assign n_32015 = n_32007 ^ n_31968;
assign n_32016 = n_32008 ^ n_32004;
assign n_32017 = n_32008 ^ n_30087;
assign n_32018 = n_32009 ^ x408;
assign n_32019 = n_32010 ^ n_31112;
assign n_32020 = n_32010 & ~n_32011;
assign n_32021 = n_32013 ^ x101;
assign n_32022 = ~n_32012 & n_32016;
assign n_32023 = n_32017 ^ n_32004;
assign n_32024 = n_32018 ^ n_32002;
assign n_32025 = ~n_30627 & ~n_32019;
assign n_32026 = n_32020 ^ n_31112;
assign n_32027 = n_32021 ^ x100;
assign n_32028 = n_32022 ^ n_30087;
assign n_32029 = n_32023 ^ x100;
assign n_32030 = n_32021 ^ n_32023;
assign n_32031 = n_32024 ^ n_31139;
assign n_32032 = n_32025 ^ n_31112;
assign n_32033 = n_32026 ^ n_32024;
assign n_32034 = n_32027 ^ n_32023;
assign n_32035 = n_32029 & ~n_32030;
assign n_32036 = n_32026 ^ n_32031;
assign n_32037 = n_32028 ^ n_32032;
assign n_32038 = n_32032 ^ n_30123;
assign n_32039 = ~n_32031 & ~n_32033;
assign n_32040 = n_32014 & n_32034;
assign n_32041 = n_32034 ^ n_32014;
assign n_32042 = n_32035 ^ x100;
assign n_32043 = n_30668 & ~n_32036;
assign n_32044 = n_32037 ^ n_30123;
assign n_32045 = n_32037 & n_32038;
assign n_32046 = n_32039 ^ n_31139;
assign n_32047 = n_32043 ^ n_31139;
assign n_32048 = n_32044 ^ x99;
assign n_32049 = n_32042 ^ n_32044;
assign n_32050 = n_32045 ^ n_30123;
assign n_32051 = n_32046 ^ n_31188;
assign n_32052 = n_32046 ^ n_31001;
assign n_32053 = n_32047 ^ n_30160;
assign n_32054 = n_32042 ^ n_32048;
assign n_32055 = ~n_32048 & n_32049;
assign n_32056 = n_32050 ^ n_32047;
assign n_32057 = ~n_31202 & n_32051;
assign n_32058 = n_32052 ^ n_31188;
assign n_32059 = n_32050 ^ n_32053;
assign n_32060 = ~n_32040 & n_32054;
assign n_32061 = n_32054 ^ n_32040;
assign n_32062 = n_32055 ^ x99;
assign n_32063 = ~n_32053 & n_32056;
assign n_32064 = n_32057 ^ n_31001;
assign n_32065 = n_30703 & n_32058;
assign n_32066 = n_32059 ^ x98;
assign n_32067 = n_32062 ^ n_32059;
assign n_32068 = n_32062 ^ x98;
assign n_32069 = n_32063 ^ n_30160;
assign n_32070 = n_32064 ^ n_31239;
assign n_32071 = n_32064 ^ n_31225;
assign n_32072 = n_32065 ^ n_31188;
assign n_32073 = ~n_32066 & n_32067;
assign n_32074 = n_32068 ^ n_32059;
assign n_32075 = ~n_30738 & n_32070;
assign n_32076 = ~n_31239 & ~n_32071;
assign n_32077 = n_32072 ^ n_30184;
assign n_32078 = n_32069 ^ n_32072;
assign n_32079 = n_32073 ^ x98;
assign n_32080 = ~n_32060 & ~n_32074;
assign n_32081 = n_32074 ^ n_32060;
assign n_32082 = n_32075 ^ n_31225;
assign n_32083 = n_32076 ^ n_31052;
assign n_32084 = n_32069 ^ n_32077;
assign n_32085 = n_32077 & ~n_32078;
assign n_32086 = n_32082 ^ n_30231;
assign n_32087 = n_32083 ^ n_31286;
assign n_32088 = n_32083 ^ n_31271;
assign n_32089 = n_32084 ^ x97;
assign n_32090 = n_32079 ^ n_32084;
assign n_32091 = n_32085 ^ n_30184;
assign n_32092 = n_30780 & n_32087;
assign n_32093 = n_31286 & ~n_32088;
assign n_32094 = n_32079 ^ n_32089;
assign n_32095 = n_32089 & ~n_32090;
assign n_32096 = n_32091 ^ n_32082;
assign n_32097 = n_32091 ^ n_30231;
assign n_32098 = n_32092 ^ n_31271;
assign n_32099 = n_32093 ^ n_31119;
assign n_32100 = n_32094 & n_32080;
assign n_32101 = n_32080 ^ n_32094;
assign n_32102 = n_32095 ^ x97;
assign n_32103 = n_32086 & n_32096;
assign n_32104 = n_32097 ^ n_32082;
assign n_32105 = n_32098 ^ n_30255;
assign n_32106 = n_32099 ^ n_31159;
assign n_32107 = n_32099 ^ n_31307;
assign n_32108 = n_32103 ^ n_30231;
assign n_32109 = n_32102 ^ n_32104;
assign n_32110 = n_32104 ^ x96;
assign n_32111 = n_32106 ^ n_31307;
assign n_32112 = n_31322 & n_32107;
assign n_32113 = n_32108 ^ n_30255;
assign n_32114 = n_32108 ^ n_32098;
assign n_32115 = n_32109 ^ x96;
assign n_32116 = ~n_32109 & n_32110;
assign n_32117 = n_30813 & n_32111;
assign n_32118 = n_32112 ^ n_31159;
assign n_32119 = n_32113 ^ n_32098;
assign n_32120 = ~n_32105 & n_32114;
assign n_32121 = ~n_32115 & ~n_32100;
assign n_32122 = n_32100 ^ n_32115;
assign n_32123 = n_32116 ^ x96;
assign n_32124 = n_32117 ^ n_31307;
assign n_32125 = n_32118 ^ n_31337;
assign n_32126 = n_31351 ^ n_32118;
assign n_32127 = n_32119 ^ x111;
assign n_32128 = n_32120 ^ n_30255;
assign n_32129 = n_32123 ^ n_32119;
assign n_32130 = n_32124 ^ n_30273;
assign n_32131 = ~n_31351 & ~n_32125;
assign n_32132 = n_32126 ^ n_31927;
assign n_32133 = n_30848 & n_32126;
assign n_32134 = n_32123 ^ n_32127;
assign n_32135 = n_32128 ^ n_32124;
assign n_32136 = n_32127 & ~n_32129;
assign n_32137 = n_32128 ^ n_32130;
assign n_32138 = n_32131 ^ n_31199;
assign n_32139 = n_32133 ^ n_31337;
assign n_32140 = n_32134 & ~n_32121;
assign n_32141 = n_32121 ^ n_32134;
assign n_32142 = n_32130 & ~n_32135;
assign n_32143 = n_32136 ^ x111;
assign n_32144 = n_32137 ^ x110;
assign n_32145 = n_32138 ^ n_31386;
assign n_32146 = n_32138 ^ n_31401;
assign n_32147 = n_32139 ^ n_30288;
assign n_32148 = n_32142 ^ n_30273;
assign n_32149 = n_32143 ^ n_32137;
assign n_32150 = n_31401 & n_32145;
assign n_32151 = n_31968 ^ n_32146;
assign n_32152 = ~n_30895 & n_32146;
assign n_32153 = n_32148 ^ n_32139;
assign n_32154 = n_32148 ^ n_30288;
assign n_32155 = n_32149 ^ x110;
assign n_32156 = n_32149 & ~n_32144;
assign n_32157 = n_32150 ^ n_31233;
assign n_32158 = n_32152 ^ n_31386;
assign n_32159 = n_32147 & ~n_32153;
assign n_32160 = n_32154 ^ n_32139;
assign n_32161 = n_32155 ^ n_32140;
assign n_32162 = n_32140 & ~n_32155;
assign n_32163 = n_32156 ^ x110;
assign n_32164 = n_32157 ^ n_31428;
assign n_32165 = n_32157 ^ n_31443;
assign n_32166 = n_32158 ^ n_30307;
assign n_32167 = n_32159 ^ n_30288;
assign n_32168 = n_32160 ^ x109;
assign n_32169 = n_32163 ^ n_32160;
assign n_32170 = n_31443 & ~n_32164;
assign n_32171 = n_32015 ^ n_32165;
assign n_32172 = ~n_30931 & ~n_32165;
assign n_32173 = n_32167 ^ n_32158;
assign n_32174 = n_32167 ^ n_30307;
assign n_32175 = n_32169 & ~n_32168;
assign n_32176 = n_32169 ^ x109;
assign n_32177 = n_32170 ^ n_31279;
assign n_32178 = n_32172 ^ n_31428;
assign n_32179 = n_32166 & ~n_32173;
assign n_32180 = n_32174 ^ n_32158;
assign n_32181 = n_32175 ^ x109;
assign n_32182 = ~n_32162 & n_32176;
assign n_32183 = n_32176 ^ n_32162;
assign n_32184 = n_32177 ^ n_31475;
assign n_32185 = n_32177 ^ n_31317;
assign n_32186 = n_32178 ^ n_30330;
assign n_32187 = n_32179 ^ n_30307;
assign n_32188 = n_32180 ^ x108;
assign n_32189 = n_32181 ^ n_32180;
assign n_32190 = n_32181 ^ x108;
assign n_32191 = ~n_31490 & n_32184;
assign n_32192 = n_32185 ^ n_31475;
assign n_32193 = n_32187 ^ n_32178;
assign n_32194 = n_32187 ^ n_32186;
assign n_32195 = ~n_32188 & n_32189;
assign n_32196 = n_32190 ^ n_32180;
assign n_32197 = n_32191 ^ n_31317;
assign n_32198 = n_30956 & n_32192;
assign n_32199 = n_32041 ^ n_32192;
assign n_32200 = ~n_32186 & ~n_32193;
assign n_32201 = n_32194 ^ x107;
assign n_32202 = n_32195 ^ x108;
assign n_32203 = n_32196 & n_32182;
assign n_32204 = n_32182 ^ n_32196;
assign n_32205 = n_32197 ^ n_31513;
assign n_32206 = n_32197 ^ n_31526;
assign n_32207 = n_32198 ^ n_31475;
assign n_32208 = n_32200 ^ n_30330;
assign n_32209 = n_32202 ^ n_32194;
assign n_32210 = ~n_31526 & ~n_32205;
assign n_32211 = n_32061 ^ n_32206;
assign n_32212 = ~n_30978 & n_32206;
assign n_32213 = n_32207 ^ n_30343;
assign n_32214 = n_32208 ^ n_32207;
assign n_32215 = ~n_32209 & n_32201;
assign n_32216 = n_32209 ^ x107;
assign n_32217 = n_32210 ^ n_31361;
assign n_32218 = n_32212 ^ n_31513;
assign n_32219 = ~n_32214 & n_32213;
assign n_32220 = n_32214 ^ n_30343;
assign n_32221 = n_32215 ^ x107;
assign n_32222 = ~n_32203 & n_32216;
assign n_32223 = n_32216 ^ n_32203;
assign n_32224 = n_32217 ^ n_31542;
assign n_32225 = n_32217 ^ n_31557;
assign n_32226 = n_32218 ^ n_30363;
assign n_32227 = n_32219 ^ n_30343;
assign n_32228 = n_32220 ^ x106;
assign n_32229 = n_32221 ^ n_32220;
assign n_32230 = ~n_31557 & ~n_32224;
assign n_32231 = n_30997 & ~n_32225;
assign n_32232 = n_32081 ^ n_32225;
assign n_32233 = n_32227 ^ n_32218;
assign n_32234 = n_32227 ^ n_30363;
assign n_32235 = n_32221 ^ n_32228;
assign n_32236 = n_32228 & ~n_32229;
assign n_32237 = n_32230 ^ n_31403;
assign n_32238 = n_32231 ^ n_31542;
assign n_32239 = n_32226 & n_32233;
assign n_32240 = n_32234 ^ n_32218;
assign n_32241 = n_32222 & n_32235;
assign n_32242 = n_32235 ^ n_32222;
assign n_32243 = n_32236 ^ x106;
assign n_32244 = n_32237 ^ n_31584;
assign n_32245 = n_32238 ^ n_30383;
assign n_32246 = n_32239 ^ n_30363;
assign n_32247 = n_32240 ^ x105;
assign n_32248 = n_32243 ^ n_32240;
assign n_32249 = ~n_32244 & n_31599;
assign n_32250 = n_31434 ^ n_32244;
assign n_32251 = n_32246 ^ n_32238;
assign n_32252 = n_32246 ^ n_30383;
assign n_32253 = ~n_32248 & n_32247;
assign n_32254 = n_32248 ^ x105;
assign n_32255 = n_32249 ^ n_31434;
assign n_32256 = n_32101 ^ n_32250;
assign n_32257 = n_31036 & ~n_32250;
assign n_32258 = ~n_32245 & n_32251;
assign n_32259 = n_32252 ^ n_32238;
assign n_32260 = n_32253 ^ x105;
assign n_32261 = ~n_32241 & ~n_32254;
assign n_32262 = n_32254 ^ n_32241;
assign n_32263 = n_32255 ^ n_31636;
assign n_32264 = n_32257 ^ n_31584;
assign n_32265 = n_32258 ^ n_30383;
assign n_32266 = n_32259 ^ x104;
assign n_32267 = n_32260 ^ n_32259;
assign n_32268 = n_32263 & n_31649;
assign n_32269 = n_31485 ^ n_32263;
assign n_32270 = n_32264 ^ n_30406;
assign n_32271 = n_32265 ^ n_32264;
assign n_32272 = n_32260 ^ n_32266;
assign n_32273 = n_32266 & ~n_32267;
assign n_32274 = n_32268 ^ n_31485;
assign n_32275 = ~n_31071 & ~n_32269;
assign n_32276 = n_32122 ^ n_32269;
assign n_32277 = ~n_32271 & n_32270;
assign n_32278 = n_32271 ^ n_30406;
assign n_32279 = n_32261 & ~n_32272;
assign n_32280 = n_32272 ^ n_32261;
assign n_32281 = n_32273 ^ x104;
assign n_32282 = n_32274 ^ n_31529;
assign n_32283 = n_32274 ^ n_31665;
assign n_32284 = n_32275 ^ n_31636;
assign n_32285 = n_32277 ^ n_30406;
assign n_32286 = n_32278 ^ x119;
assign n_32287 = n_32281 ^ n_32278;
assign n_32288 = n_32282 ^ n_31665;
assign n_32289 = n_31677 & ~n_32283;
assign n_32290 = n_32284 ^ n_30420;
assign n_32291 = n_32285 ^ n_32284;
assign n_32292 = n_32287 & ~n_32286;
assign n_32293 = n_32287 ^ x119;
assign n_32294 = n_32141 ^ n_32288;
assign n_32295 = ~n_31105 & n_32288;
assign n_32296 = n_32289 ^ n_31529;
assign n_32297 = n_32285 ^ n_32290;
assign n_32298 = ~n_32290 & n_32291;
assign n_32299 = n_32292 ^ x119;
assign n_32300 = ~n_32279 & ~n_32293;
assign n_32301 = n_32293 ^ n_32279;
assign n_32302 = n_32295 ^ n_31665;
assign n_32303 = n_32296 ^ n_31697;
assign n_32304 = n_32296 ^ n_31705;
assign n_32305 = n_32297 ^ x118;
assign n_32306 = n_32298 ^ n_30420;
assign n_32307 = n_32299 ^ n_32297;
assign n_32308 = n_32299 ^ x118;
assign n_32309 = n_32302 ^ n_30446;
assign n_32310 = ~n_31705 & ~n_32303;
assign n_32311 = ~n_31141 & ~n_32304;
assign n_32312 = n_32161 ^ n_32304;
assign n_32313 = n_32306 ^ n_32302;
assign n_32314 = n_32306 ^ n_30446;
assign n_32315 = n_32305 & ~n_32307;
assign n_32316 = n_32308 ^ n_32297;
assign n_32317 = n_32310 ^ n_31571;
assign n_32318 = n_32311 ^ n_31697;
assign n_32319 = n_32309 & n_32313;
assign n_32320 = n_32314 ^ n_32302;
assign n_32321 = n_32315 ^ x118;
assign n_32322 = n_32300 & n_32316;
assign n_32323 = n_32316 ^ n_32300;
assign n_32324 = n_32317 ^ n_31717;
assign n_32325 = n_32317 ^ n_31724;
assign n_32326 = n_32318 ^ n_30466;
assign n_32327 = n_32319 ^ n_30446;
assign n_32328 = n_32320 ^ x117;
assign n_32329 = n_32321 ^ n_32320;
assign n_32330 = ~n_31724 & ~n_32324;
assign n_32331 = n_31168 & n_32325;
assign n_32332 = n_32183 ^ n_32325;
assign n_32333 = n_32327 ^ n_32318;
assign n_32334 = n_32321 ^ n_32328;
assign n_32335 = ~n_32328 & n_32329;
assign n_32336 = n_32330 ^ n_31614;
assign n_32337 = n_32331 ^ n_31717;
assign n_32338 = ~n_32333 & ~n_32326;
assign n_32339 = n_32333 ^ n_30466;
assign n_32340 = ~n_32322 & n_32334;
assign n_32341 = n_32334 ^ n_32322;
assign n_32342 = n_32335 ^ x117;
assign n_32343 = n_32336 ^ n_31733;
assign n_32344 = n_32336 ^ n_31741;
assign n_32345 = n_32337 ^ n_30488;
assign n_32346 = n_32338 ^ n_30466;
assign n_32347 = n_32339 ^ x116;
assign n_32348 = n_32342 ^ n_32339;
assign n_32349 = n_31741 & ~n_32343;
assign n_32350 = n_31208 & n_32344;
assign n_32351 = n_32204 ^ n_32344;
assign n_32352 = n_32346 ^ n_32337;
assign n_32353 = n_32346 ^ n_32345;
assign n_32354 = n_32342 ^ n_32347;
assign n_32355 = ~n_32347 & n_32348;
assign n_32356 = n_32349 ^ n_31654;
assign n_32357 = n_32350 ^ n_31733;
assign n_32358 = ~n_32345 & ~n_32352;
assign n_32359 = n_32353 ^ x115;
assign n_32360 = n_32340 & n_32354;
assign n_32361 = n_32354 ^ n_32340;
assign n_32362 = n_32355 ^ x116;
assign n_32363 = n_32356 ^ n_31758;
assign n_32364 = n_32356 ^ n_31765;
assign n_32365 = n_32357 ^ n_30506;
assign n_32366 = n_32358 ^ n_30488;
assign n_32367 = n_32362 ^ n_32353;
assign n_32368 = n_31765 & ~n_32363;
assign n_32369 = ~n_31248 & n_32364;
assign n_32370 = n_32223 ^ n_32364;
assign n_32371 = n_32366 ^ n_32357;
assign n_32372 = ~n_32367 & n_32359;
assign n_32373 = n_32367 ^ x115;
assign n_32374 = n_32368 ^ n_31686;
assign n_32375 = n_32369 ^ n_31758;
assign n_32376 = ~n_32371 & ~n_32365;
assign n_32377 = n_32371 ^ n_30506;
assign n_32378 = n_32372 ^ x115;
assign n_32379 = ~n_32360 & n_32373;
assign n_32380 = n_32373 ^ n_32360;
assign n_32381 = n_32374 ^ n_31777;
assign n_32382 = n_32374 ^ n_31709;
assign n_32383 = n_32375 ^ n_30538;
assign n_32384 = n_32376 ^ n_30506;
assign n_32385 = n_32377 ^ x114;
assign n_32386 = n_32378 ^ n_32377;
assign n_32387 = ~n_31786 & ~n_32381;
assign n_32388 = n_32382 ^ n_31777;
assign n_32389 = n_32384 ^ n_32375;
assign n_32390 = n_32384 ^ n_30538;
assign n_32391 = n_32386 & ~n_32385;
assign n_32392 = n_32386 ^ x114;
assign n_32393 = n_32387 ^ n_31709;
assign n_32394 = n_31300 & ~n_32388;
assign n_32395 = n_32242 ^ n_32388;
assign n_32396 = n_32383 & n_32389;
assign n_32397 = n_32390 ^ n_32375;
assign n_32398 = n_32391 ^ x114;
assign n_32399 = n_32379 & ~n_32392;
assign n_32400 = n_32393 ^ n_31791;
assign n_32401 = n_32393 ^ n_31729;
assign n_32402 = n_32394 ^ n_31777;
assign n_32403 = n_32396 ^ n_30538;
assign n_32404 = n_32397 ^ x113;
assign n_32405 = n_32398 ^ n_32397;
assign n_32406 = n_32398 ^ x113;
assign n_32407 = ~n_31798 & n_32400;
assign n_32408 = n_32401 ^ n_31791;
assign n_32409 = n_32402 ^ n_30572;
assign n_32410 = n_32403 ^ n_32402;
assign n_32411 = n_32403 ^ n_30572;
assign n_32412 = ~n_32404 & n_32405;
assign n_32413 = n_32406 ^ n_32397;
assign n_32414 = n_32407 ^ n_31729;
assign n_32415 = ~n_31327 & n_32408;
assign n_32416 = n_32262 ^ n_32408;
assign n_32417 = ~n_32409 & ~n_32410;
assign n_32418 = n_32411 ^ n_32402;
assign n_32419 = n_32412 ^ x113;
assign n_32420 = n_32399 & ~n_32413;
assign n_32421 = n_32413 ^ n_32399;
assign n_32422 = n_32414 ^ n_31817;
assign n_32423 = n_32414 ^ n_31751;
assign n_32424 = n_32415 ^ n_31791;
assign n_32425 = n_32417 ^ n_30572;
assign n_32426 = n_32418 ^ x112;
assign n_32427 = n_32419 ^ n_32418;
assign n_32428 = n_31896 & ~n_32421;
assign n_32429 = n_32421 ^ n_31888;
assign n_32430 = n_31824 & n_32422;
assign n_32431 = n_32423 ^ n_31817;
assign n_32432 = n_32424 ^ n_30605;
assign n_32433 = n_32425 ^ n_32424;
assign n_32434 = n_32419 ^ n_32426;
assign n_32435 = ~n_32426 & n_32427;
assign n_32436 = n_32428 ^ n_31923;
assign n_32437 = n_32429 ^ n_30973;
assign n_32438 = n_32430 ^ n_31751;
assign n_32439 = ~n_31381 & ~n_32431;
assign n_32440 = n_32280 ^ n_32431;
assign n_32441 = n_32425 ^ n_32432;
assign n_32442 = ~n_32432 & n_32433;
assign n_32443 = n_32420 & ~n_32434;
assign n_32444 = n_32434 ^ n_32420;
assign n_32445 = n_32435 ^ x112;
assign n_32446 = n_30973 & n_32437;
assign n_32447 = n_32438 ^ n_31770;
assign n_32448 = n_32438 ^ n_31831;
assign n_32449 = n_32439 ^ n_31817;
assign n_32450 = n_32441 ^ x127;
assign n_32451 = n_32442 ^ n_30605;
assign n_32452 = n_32444 ^ n_32428;
assign n_32453 = n_32444 ^ n_32436;
assign n_32454 = n_32445 ^ n_32441;
assign n_32455 = n_31897 ^ n_32446;
assign n_32456 = n_32446 ^ n_31896;
assign n_32457 = n_32447 ^ n_31831;
assign n_32458 = n_31838 & n_32448;
assign n_32459 = n_32449 ^ n_30656;
assign n_32460 = n_32451 ^ n_32449;
assign n_32461 = ~n_32436 & n_32452;
assign n_32462 = ~n_31000 & ~n_32453;
assign n_32463 = ~n_32454 & n_32450;
assign n_32464 = n_32454 ^ x127;
assign n_32465 = n_32455 ^ x327;
assign n_32466 = x327 & ~n_32455;
assign n_32467 = n_30487 & ~n_32456;
assign n_32468 = ~n_31409 & n_32457;
assign n_32469 = n_32301 ^ n_32457;
assign n_32470 = n_32458 ^ n_31770;
assign n_32471 = n_32460 & ~n_32459;
assign n_32472 = n_32460 ^ n_30656;
assign n_32473 = n_32461 ^ n_31923;
assign n_32474 = n_32462 ^ n_31923;
assign n_32475 = n_32463 ^ x127;
assign n_32476 = ~n_32443 & ~n_32464;
assign n_32477 = n_32464 ^ n_32443;
assign n_32478 = n_32466 ^ x326;
assign n_32479 = n_32467 ^ n_30511;
assign n_32480 = n_32468 ^ n_31831;
assign n_32481 = n_32470 ^ n_31859;
assign n_32482 = n_32470 ^ n_31852;
assign n_32483 = n_32471 ^ n_30656;
assign n_32484 = n_32472 ^ x126;
assign n_32485 = n_32473 ^ n_31965;
assign n_32486 = n_32474 ^ n_32467;
assign n_32487 = n_32475 ^ n_32472;
assign n_32488 = n_32475 ^ x126;
assign n_32489 = n_32477 ^ n_31965;
assign n_32490 = n_32473 ^ n_32477;
assign n_32491 = n_32474 ^ n_32479;
assign n_32492 = n_32480 ^ n_30695;
assign n_32493 = n_31449 & n_32481;
assign n_32494 = n_32323 ^ n_32481;
assign n_32495 = ~n_31859 & ~n_32482;
assign n_32496 = n_32483 ^ n_32480;
assign n_32497 = n_32483 ^ n_30695;
assign n_32498 = n_32485 ^ n_32477;
assign n_32499 = n_32479 & ~n_32486;
assign n_32500 = n_32484 & ~n_32487;
assign n_32501 = n_32488 ^ n_32472;
assign n_32502 = n_32489 & ~n_32490;
assign n_32503 = n_32491 ^ n_32478;
assign n_32504 = n_32491 ^ n_32466;
assign n_32505 = n_32493 ^ n_31852;
assign n_32506 = n_32495 ^ n_31783;
assign n_32507 = ~n_32492 & ~n_32496;
assign n_32508 = n_32497 ^ n_32480;
assign n_32509 = ~n_31041 & n_32498;
assign n_32510 = n_32499 ^ n_30511;
assign n_32511 = n_32500 ^ x126;
assign n_32512 = n_32476 & ~n_32501;
assign n_32513 = n_32501 ^ n_32476;
assign n_32514 = n_32502 ^ n_31965;
assign n_32515 = ~n_32465 & n_32503;
assign n_32516 = n_32503 ^ n_32465;
assign n_32517 = n_32478 & ~n_32504;
assign n_32518 = n_32505 ^ n_30722;
assign n_32519 = n_32506 ^ n_31877;
assign n_32520 = n_32506 ^ n_31871;
assign n_32521 = n_32507 ^ n_30695;
assign n_32522 = n_32508 ^ x125;
assign n_32523 = n_32509 ^ n_31965;
assign n_32524 = n_32511 ^ n_32508;
assign n_32525 = n_32513 ^ n_31990;
assign n_32526 = n_32514 ^ n_32513;
assign n_32527 = n_32517 ^ x326;
assign n_32528 = ~n_31491 & ~n_32519;
assign n_32529 = n_32341 ^ n_32519;
assign n_32530 = ~n_31877 & n_32520;
assign n_32531 = n_32521 ^ n_32518;
assign n_32532 = n_32521 ^ n_32505;
assign n_32533 = n_32511 ^ n_32522;
assign n_32534 = n_32523 ^ n_30552;
assign n_32535 = n_32510 ^ n_32523;
assign n_32536 = n_32522 & ~n_32524;
assign n_32537 = n_32525 ^ n_32514;
assign n_32538 = n_32526 & n_32525;
assign n_32539 = n_32527 ^ x325;
assign n_32540 = n_32528 ^ n_31871;
assign n_32541 = n_32530 ^ n_31810;
assign n_32542 = n_32531 ^ x124;
assign n_32543 = n_32518 & n_32532;
assign n_32544 = ~n_32533 & n_32512;
assign n_32545 = n_32512 ^ n_32533;
assign n_32546 = n_32510 ^ n_32534;
assign n_32547 = n_32534 & ~n_32535;
assign n_32548 = n_32536 ^ x125;
assign n_32549 = ~n_31077 & n_32537;
assign n_32550 = n_32538 ^ n_31990;
assign n_32551 = n_32540 ^ n_30774;
assign n_32552 = n_32541 ^ n_31907;
assign n_32553 = n_32541 ^ n_31898;
assign n_32554 = n_32543 ^ n_30722;
assign n_32555 = n_32545 ^ n_32019;
assign n_32556 = n_32539 ^ n_32546;
assign n_32557 = n_32546 ^ x325;
assign n_32558 = n_32527 ^ n_32546;
assign n_32559 = n_32547 ^ n_30552;
assign n_32560 = n_32548 ^ n_32531;
assign n_32561 = n_32548 ^ n_32542;
assign n_32562 = n_32549 ^ n_31990;
assign n_32563 = n_32550 ^ n_32545;
assign n_32564 = ~n_31534 & n_32552;
assign n_32565 = n_32361 ^ n_32552;
assign n_32566 = n_31907 & n_32553;
assign n_32567 = n_32554 ^ n_32551;
assign n_32568 = n_32554 ^ n_32540;
assign n_32569 = n_32550 ^ n_32555;
assign n_32570 = ~n_32515 & ~n_32556;
assign n_32571 = n_32556 ^ n_32515;
assign n_32572 = n_32557 & ~n_32558;
assign n_32573 = n_32559 ^ n_30587;
assign n_32574 = n_32542 & ~n_32560;
assign n_32575 = ~n_32561 & n_32544;
assign n_32576 = n_32544 ^ n_32561;
assign n_32577 = n_32562 ^ n_30587;
assign n_32578 = n_32559 ^ n_32562;
assign n_32579 = n_32555 & ~n_32563;
assign n_32580 = n_32564 ^ n_31898;
assign n_32581 = n_32566 ^ n_31829;
assign n_32582 = n_32567 ^ x123;
assign n_32583 = ~n_32551 & ~n_32568;
assign n_32584 = ~n_31112 & ~n_32569;
assign n_32585 = n_32572 ^ x325;
assign n_32586 = n_32573 ^ n_32562;
assign n_32587 = n_32574 ^ x124;
assign n_32588 = n_32576 ^ n_32036;
assign n_32589 = ~n_32577 & n_32578;
assign n_32590 = n_32579 ^ n_32019;
assign n_32591 = n_32580 ^ n_30802;
assign n_32592 = n_31930 ^ n_32581;
assign n_32593 = n_32581 ^ n_31917;
assign n_32594 = n_31849 ^ n_32581;
assign n_32595 = n_32583 ^ n_30774;
assign n_32596 = n_32584 ^ n_32019;
assign n_32597 = n_32586 ^ x324;
assign n_32598 = n_32585 ^ n_32586;
assign n_32599 = n_32587 ^ n_32582;
assign n_32600 = n_32587 ^ n_32567;
assign n_32601 = n_32589 ^ n_30587;
assign n_32602 = n_32590 ^ n_32576;
assign n_32603 = n_32590 ^ n_32588;
assign n_32604 = ~n_31576 & n_32592;
assign n_32605 = n_32593 & n_32594;
assign n_32606 = n_32595 ^ n_30802;
assign n_32607 = n_32595 ^ n_32580;
assign n_32608 = n_32596 ^ n_30627;
assign n_32609 = n_32585 ^ n_32597;
assign n_32610 = ~n_32597 & n_32598;
assign n_32611 = n_32599 & ~n_32575;
assign n_32612 = n_32575 ^ n_32599;
assign n_32613 = n_32582 & ~n_32600;
assign n_32614 = n_32601 ^ n_32596;
assign n_32615 = n_32588 & ~n_32602;
assign n_32616 = n_31139 & ~n_32603;
assign n_32617 = n_32604 ^ n_31917;
assign n_32618 = n_31971 ^ n_32605;
assign n_32619 = n_32606 ^ n_32580;
assign n_32620 = ~n_32591 & n_32607;
assign n_32621 = n_32601 ^ n_32608;
assign n_32622 = n_32570 & n_32609;
assign n_32623 = n_32609 ^ n_32570;
assign n_32624 = n_32610 ^ x324;
assign n_32625 = n_32612 ^ n_32058;
assign n_32626 = n_32613 ^ x123;
assign n_32627 = n_32608 & n_32614;
assign n_32628 = n_32615 ^ n_32036;
assign n_32629 = n_32616 ^ n_32036;
assign n_32630 = n_32617 ^ n_30854;
assign n_32631 = ~n_31604 & n_32618;
assign n_32632 = n_32618 ^ n_32379;
assign n_32633 = n_32619 ^ x122;
assign n_32634 = n_32620 ^ n_30802;
assign n_32635 = n_32621 ^ x323;
assign n_32636 = n_32624 ^ x323;
assign n_32637 = n_32621 ^ n_32624;
assign n_32638 = n_32626 ^ x122;
assign n_32639 = n_32626 ^ n_32619;
assign n_32640 = n_32627 ^ n_30627;
assign n_32641 = n_32628 ^ n_32612;
assign n_32642 = n_32628 ^ n_32625;
assign n_32643 = n_32629 ^ n_30668;
assign n_32644 = n_32631 ^ n_31940;
assign n_32645 = n_32632 ^ n_32392;
assign n_32646 = n_32630 ^ n_32634;
assign n_32647 = n_32617 ^ n_32634;
assign n_32648 = n_32635 ^ n_32624;
assign n_32649 = n_32636 & ~n_32637;
assign n_32650 = n_32638 ^ n_32619;
assign n_32651 = ~n_32633 & n_32639;
assign n_32652 = n_32640 ^ n_32629;
assign n_32653 = n_32625 & n_32641;
assign n_32654 = ~n_31188 & ~n_32642;
assign n_32655 = n_32640 ^ n_32643;
assign n_32656 = n_32645 ^ n_32380;
assign n_32657 = n_32646 ^ x121;
assign n_32658 = ~n_32630 & n_32647;
assign n_32659 = n_32622 ^ n_32648;
assign n_32660 = ~n_32648 & n_32622;
assign n_32661 = n_32649 ^ x323;
assign n_32662 = n_32611 ^ n_32650;
assign n_32663 = ~n_32650 & n_32611;
assign n_32664 = n_32651 ^ x122;
assign n_32665 = ~n_32643 & ~n_32652;
assign n_32666 = n_32653 ^ n_32058;
assign n_32667 = n_32654 ^ n_32058;
assign n_32668 = n_32655 ^ x322;
assign n_32669 = n_32658 ^ n_30854;
assign n_32670 = n_32661 ^ n_32655;
assign n_32671 = n_32662 ^ n_32070;
assign n_32672 = n_32646 ^ n_32664;
assign n_32673 = n_32665 ^ n_30668;
assign n_32674 = n_32666 ^ n_32662;
assign n_32675 = n_32666 ^ n_32070;
assign n_32676 = n_32667 ^ n_30703;
assign n_32677 = n_32661 ^ n_32668;
assign n_32678 = n_32669 ^ n_30867;
assign n_32679 = n_32668 & ~n_32670;
assign n_32680 = n_32672 ^ x121;
assign n_32681 = n_32672 & ~n_32657;
assign n_32682 = n_32673 ^ n_32667;
assign n_32683 = n_32673 ^ n_30703;
assign n_32684 = n_32671 & ~n_32674;
assign n_32685 = n_32675 ^ n_32662;
assign n_32686 = n_32660 & ~n_32677;
assign n_32687 = n_32677 ^ n_32660;
assign n_32688 = n_32678 ^ n_32644;
assign n_32689 = n_32679 ^ x322;
assign n_32690 = n_32663 ^ n_32680;
assign n_32691 = ~n_32680 & n_32663;
assign n_32692 = n_32681 ^ x121;
assign n_32693 = n_32676 & ~n_32682;
assign n_32694 = n_32683 ^ n_32667;
assign n_32695 = n_32684 ^ n_32070;
assign n_32696 = n_31225 & n_32685;
assign n_32697 = n_32688 ^ x120;
assign n_32698 = n_32689 ^ x321;
assign n_32699 = n_32690 ^ n_32087;
assign n_32700 = n_32693 ^ n_30703;
assign n_32701 = n_32694 ^ x321;
assign n_32702 = n_32689 ^ n_32694;
assign n_32703 = n_32695 ^ n_32690;
assign n_32704 = n_32696 ^ n_32070;
assign n_32705 = n_32692 ^ n_32697;
assign n_32706 = n_32698 ^ n_32694;
assign n_32707 = n_32701 & ~n_32702;
assign n_32708 = ~n_32703 & n_32699;
assign n_32709 = n_32703 ^ n_32087;
assign n_32710 = n_32704 ^ n_30738;
assign n_32711 = n_32700 ^ n_32704;
assign n_32712 = n_32705 ^ n_32691;
assign n_32713 = n_32686 & ~n_32706;
assign n_32714 = n_32706 ^ n_32686;
assign n_32715 = n_32707 ^ x321;
assign n_32716 = n_32708 ^ n_32087;
assign n_32717 = ~n_31271 & n_32709;
assign n_32718 = n_32700 ^ n_32710;
assign n_32719 = ~n_32710 & ~n_32711;
assign n_32720 = n_32712 ^ n_32111;
assign n_32721 = n_32715 ^ x320;
assign n_32722 = n_32716 ^ n_32712;
assign n_32723 = n_32717 ^ n_32087;
assign n_32724 = n_32718 ^ x320;
assign n_32725 = n_32715 ^ n_32718;
assign n_32726 = n_32719 ^ n_30738;
assign n_32727 = n_32721 ^ n_32718;
assign n_32728 = n_32722 & ~n_32720;
assign n_32729 = n_32722 ^ n_32111;
assign n_32730 = n_32723 ^ n_30780;
assign n_32731 = ~n_32724 & n_32725;
assign n_32732 = n_32726 ^ n_32723;
assign n_32733 = ~n_32727 & ~n_32713;
assign n_32734 = n_32713 ^ n_32727;
assign n_32735 = n_32728 ^ n_32111;
assign n_32736 = n_31307 & ~n_32729;
assign n_32737 = n_32726 ^ n_32730;
assign n_32738 = n_32731 ^ x320;
assign n_32739 = n_32730 & n_32732;
assign n_32740 = n_32735 ^ n_32126;
assign n_32741 = n_32735 ^ n_32132;
assign n_32742 = n_32736 ^ n_32111;
assign n_32743 = n_32737 ^ x335;
assign n_32744 = n_32738 ^ n_32737;
assign n_32745 = n_32738 ^ x335;
assign n_32746 = n_32739 ^ n_30780;
assign n_32747 = n_32132 & ~n_32740;
assign n_32748 = n_31337 & n_32741;
assign n_32749 = n_32742 ^ n_30813;
assign n_32750 = ~n_32743 & n_32744;
assign n_32751 = n_32745 ^ n_32737;
assign n_32752 = n_32746 ^ n_32742;
assign n_32753 = n_32746 ^ n_30813;
assign n_32754 = n_32747 ^ n_31927;
assign n_32755 = n_32748 ^ n_32126;
assign n_32756 = n_32750 ^ x335;
assign n_32757 = n_32733 & ~n_32751;
assign n_32758 = n_32751 ^ n_32733;
assign n_32759 = n_32749 & ~n_32752;
assign n_32760 = n_32753 ^ n_32742;
assign n_32761 = n_32754 ^ n_32146;
assign n_32762 = n_32151 ^ n_32754;
assign n_32763 = n_32755 ^ n_30848;
assign n_32764 = n_32759 ^ n_30813;
assign n_32765 = n_32760 ^ x334;
assign n_32766 = n_32756 ^ n_32760;
assign n_32767 = n_32151 & ~n_32761;
assign n_32768 = n_31386 & n_32762;
assign n_32769 = n_32764 ^ n_32755;
assign n_32770 = n_32756 ^ n_32765;
assign n_32771 = n_32765 & ~n_32766;
assign n_32772 = n_32767 ^ n_31968;
assign n_32773 = n_32768 ^ n_32146;
assign n_32774 = ~n_32769 & n_32763;
assign n_32775 = n_32769 ^ n_30848;
assign n_32776 = n_32757 & n_32770;
assign n_32777 = n_32770 ^ n_32757;
assign n_32778 = n_32771 ^ x334;
assign n_32779 = n_32772 ^ n_32165;
assign n_32780 = n_32171 ^ n_32772;
assign n_32781 = n_32773 ^ n_30895;
assign n_32782 = n_32774 ^ n_30848;
assign n_32783 = n_32775 ^ x333;
assign n_32784 = n_32778 ^ n_32775;
assign n_32785 = n_32778 ^ x333;
assign n_32786 = ~n_32171 & n_32779;
assign n_32787 = n_31428 & ~n_32780;
assign n_32788 = n_32782 ^ n_32773;
assign n_32789 = n_32782 ^ n_32781;
assign n_32790 = n_32783 & ~n_32784;
assign n_32791 = n_32785 ^ n_32775;
assign n_32792 = n_32786 ^ n_32015;
assign n_32793 = n_32787 ^ n_32165;
assign n_32794 = ~n_32781 & ~n_32788;
assign n_32795 = n_32789 ^ x332;
assign n_32796 = n_32790 ^ x333;
assign n_32797 = ~n_32776 & ~n_32791;
assign n_32798 = n_32791 ^ n_32776;
assign n_32799 = n_32792 ^ n_32192;
assign n_32800 = n_32793 ^ n_30931;
assign n_32801 = n_32794 ^ n_30895;
assign n_32802 = n_32796 ^ n_32789;
assign n_32803 = n_32796 ^ n_32795;
assign n_32804 = ~n_32799 & ~n_32199;
assign n_32805 = n_32799 ^ n_32041;
assign n_32806 = n_32793 ^ n_32801;
assign n_32807 = n_32800 ^ n_32801;
assign n_32808 = ~n_32795 & n_32802;
assign n_32809 = ~n_32797 & ~n_32803;
assign n_32810 = n_32803 ^ n_32797;
assign n_32811 = n_32804 ^ n_32041;
assign n_32812 = ~n_31475 & ~n_32805;
assign n_32813 = n_32800 & ~n_32806;
assign n_32814 = n_32807 ^ x331;
assign n_32815 = n_32808 ^ x332;
assign n_32816 = n_32811 ^ n_32206;
assign n_32817 = n_32811 ^ n_32211;
assign n_32818 = n_32812 ^ n_32192;
assign n_32819 = n_32813 ^ n_30931;
assign n_32820 = n_32815 ^ n_32807;
assign n_32821 = ~n_32211 & n_32816;
assign n_32822 = n_31513 & n_32817;
assign n_32823 = n_32818 ^ n_30956;
assign n_32824 = n_32818 ^ n_32819;
assign n_32825 = n_32819 ^ n_30956;
assign n_32826 = n_32820 & ~n_32814;
assign n_32827 = n_32820 ^ x331;
assign n_32828 = n_32821 ^ n_32061;
assign n_32829 = n_32822 ^ n_32206;
assign n_32830 = n_32823 & n_32824;
assign n_32831 = n_32818 ^ n_32825;
assign n_32832 = n_32826 ^ x331;
assign n_32833 = n_32827 & ~n_32809;
assign n_32834 = n_32809 ^ n_32827;
assign n_32835 = n_32828 ^ n_32225;
assign n_32836 = n_32829 ^ n_30978;
assign n_32837 = n_32830 ^ n_30956;
assign n_32838 = n_32831 ^ x330;
assign n_32839 = n_32831 ^ n_32832;
assign n_32840 = ~n_32835 & n_32232;
assign n_32841 = n_32081 ^ n_32835;
assign n_32842 = n_32837 ^ n_32829;
assign n_32843 = n_32837 ^ n_32836;
assign n_32844 = n_32838 ^ n_32832;
assign n_32845 = ~n_32838 & n_32839;
assign n_32846 = n_32840 ^ n_32081;
assign n_32847 = n_32841 ^ n_32465;
assign n_32848 = ~n_31542 & ~n_32841;
assign n_32849 = ~n_32836 & ~n_32842;
assign n_32850 = n_32843 ^ x329;
assign n_32851 = n_32844 & n_32833;
assign n_32852 = n_32833 ^ n_32844;
assign n_32853 = n_32845 ^ x330;
assign n_32854 = n_32846 ^ n_32250;
assign n_32855 = n_32846 ^ n_32256;
assign n_32856 = n_32848 ^ n_32225;
assign n_32857 = n_32849 ^ n_30978;
assign n_32858 = n_32853 ^ n_32843;
assign n_32859 = n_32853 ^ x329;
assign n_32860 = n_32256 & ~n_32854;
assign n_32861 = n_32855 ^ n_32516;
assign n_32862 = n_31584 & ~n_32855;
assign n_32863 = n_32856 ^ n_30997;
assign n_32864 = n_32857 ^ n_32856;
assign n_32865 = ~n_32850 & n_32858;
assign n_32866 = n_32859 ^ n_32843;
assign n_32867 = n_32860 ^ n_32101;
assign n_32868 = n_32862 ^ n_32250;
assign n_32869 = n_32857 ^ n_32863;
assign n_32870 = ~n_32863 & ~n_32864;
assign n_32871 = n_32865 ^ x329;
assign n_32872 = n_32851 & n_32866;
assign n_32873 = n_32866 ^ n_32851;
assign n_32874 = n_32867 ^ n_32269;
assign n_32875 = n_32868 ^ n_31036;
assign n_32876 = n_32869 ^ x328;
assign n_32877 = n_32870 ^ n_30997;
assign n_32878 = n_32871 ^ n_32869;
assign n_32879 = ~n_32874 & ~n_32276;
assign n_32880 = n_32122 ^ n_32874;
assign n_32881 = n_32871 ^ n_32876;
assign n_32882 = n_32877 ^ n_32868;
assign n_32883 = n_32877 ^ n_32875;
assign n_32884 = n_32876 & ~n_32878;
assign n_32885 = n_32879 ^ n_32122;
assign n_32886 = n_32880 ^ n_32571;
assign n_32887 = ~n_31636 & n_32880;
assign n_32888 = n_32872 & ~n_32881;
assign n_32889 = n_32881 ^ n_32872;
assign n_32890 = ~n_32875 & n_32882;
assign n_32891 = n_32883 ^ x343;
assign n_32892 = n_32884 ^ x328;
assign n_32893 = n_32885 ^ n_32288;
assign n_32894 = n_32885 ^ n_32294;
assign n_32895 = n_32887 ^ n_32269;
assign n_32896 = n_32890 ^ n_31036;
assign n_32897 = n_32892 ^ n_32883;
assign n_32898 = n_32892 ^ n_32891;
assign n_32899 = n_32294 & ~n_32893;
assign n_32900 = n_32894 ^ n_32623;
assign n_32901 = ~n_31665 & n_32894;
assign n_32902 = n_32895 ^ n_31071;
assign n_32903 = n_32896 ^ n_32895;
assign n_32904 = n_32896 ^ n_31071;
assign n_32905 = ~n_32891 & n_32897;
assign n_32906 = n_32888 & n_32898;
assign n_32907 = n_32898 ^ n_32888;
assign n_32908 = n_32899 ^ n_32141;
assign n_32909 = n_32901 ^ n_32288;
assign n_32910 = n_32902 & n_32903;
assign n_32911 = n_32904 ^ n_32895;
assign n_32912 = n_32905 ^ x343;
assign n_32913 = n_32908 ^ n_32304;
assign n_32914 = n_32909 ^ n_31105;
assign n_32915 = n_32910 ^ n_31071;
assign n_32916 = n_32911 ^ x342;
assign n_32917 = n_32912 ^ n_32911;
assign n_32918 = n_32161 ^ n_32913;
assign n_32919 = n_32913 & ~n_32312;
assign n_32920 = n_32915 ^ n_32909;
assign n_32921 = n_32915 ^ n_31105;
assign n_32922 = n_32912 ^ n_32916;
assign n_32923 = n_32916 & ~n_32917;
assign n_32924 = n_32918 ^ n_32659;
assign n_32925 = ~n_31697 & ~n_32918;
assign n_32926 = n_32919 ^ n_32161;
assign n_32927 = ~n_32914 & n_32920;
assign n_32928 = n_32921 ^ n_32909;
assign n_32929 = n_32906 & ~n_32922;
assign n_32930 = n_32922 ^ n_32906;
assign n_32931 = n_32923 ^ x342;
assign n_32932 = n_32925 ^ n_32304;
assign n_32933 = n_32926 ^ n_32325;
assign n_32934 = n_32926 ^ n_32183;
assign n_32935 = n_32927 ^ n_31105;
assign n_32936 = n_32928 ^ x341;
assign n_32937 = ~n_32437 & n_32930;
assign n_32938 = n_32930 ^ n_32437;
assign n_32939 = n_32930 ^ n_32421;
assign n_32940 = n_32931 ^ n_32928;
assign n_32941 = n_32932 ^ n_31141;
assign n_32942 = ~n_32332 & ~n_32933;
assign n_32943 = n_32934 ^ n_32325;
assign n_32944 = n_32935 ^ n_32932;
assign n_32945 = n_32935 ^ n_31141;
assign n_32946 = n_32931 ^ n_32936;
assign n_32947 = n_32937 ^ n_32453;
assign n_32948 = n_31896 & n_32938;
assign n_32949 = n_32936 & ~n_32940;
assign n_32950 = n_32942 ^ n_32183;
assign n_32951 = n_31717 & ~n_32943;
assign n_32952 = n_32943 ^ n_32687;
assign n_32953 = n_32941 & ~n_32944;
assign n_32954 = n_32945 ^ n_32932;
assign n_32955 = n_32929 & ~n_32946;
assign n_32956 = n_32946 ^ n_32929;
assign n_32957 = n_32948 ^ n_32429;
assign n_32958 = n_32949 ^ x341;
assign n_32959 = n_32950 ^ n_32344;
assign n_32960 = n_32950 ^ n_32204;
assign n_32961 = n_32951 ^ n_32325;
assign n_32962 = n_32953 ^ n_31141;
assign n_32963 = n_32954 ^ x340;
assign n_32964 = n_32956 ^ n_32937;
assign n_32965 = n_30973 & ~n_32957;
assign n_32966 = x39 & n_32957;
assign n_32967 = n_32957 ^ x39;
assign n_32968 = n_32958 ^ n_32954;
assign n_32969 = n_32351 & n_32959;
assign n_32970 = n_32960 ^ n_32344;
assign n_32971 = n_32961 ^ n_31168;
assign n_32972 = n_32962 ^ n_32961;
assign n_32973 = n_32958 ^ n_32963;
assign n_32974 = ~n_32964 & n_32947;
assign n_32975 = n_32964 ^ n_32453;
assign n_32976 = n_32965 ^ n_31000;
assign n_32977 = n_32966 ^ x38;
assign n_32978 = ~n_32963 & n_32968;
assign n_32979 = n_32969 ^ n_32204;
assign n_32980 = ~n_31733 & ~n_32970;
assign n_32981 = n_32970 ^ n_32714;
assign n_32982 = n_32962 ^ n_32971;
assign n_32983 = n_32971 & n_32972;
assign n_32984 = n_32955 & n_32973;
assign n_32985 = n_32973 ^ n_32955;
assign n_32986 = n_32974 ^ n_32453;
assign n_32987 = ~n_31923 & ~n_32975;
assign n_32988 = n_32978 ^ x340;
assign n_32989 = n_32979 ^ n_32364;
assign n_32990 = n_32979 ^ n_32370;
assign n_32991 = n_32980 ^ n_32344;
assign n_32992 = n_32982 ^ x339;
assign n_32993 = n_32983 ^ n_31168;
assign n_32994 = n_32985 ^ n_32498;
assign n_32995 = n_32986 ^ n_32985;
assign n_32996 = n_32986 ^ n_32498;
assign n_32997 = n_32987 ^ n_32453;
assign n_32998 = n_32988 ^ n_32982;
assign n_32999 = n_32370 & ~n_32989;
assign n_33000 = ~n_31758 & n_32990;
assign n_33001 = n_32734 ^ n_32990;
assign n_33002 = n_32991 ^ n_31208;
assign n_33003 = n_32988 ^ n_32992;
assign n_33004 = n_32991 ^ n_32993;
assign n_33005 = n_32994 & n_32995;
assign n_33006 = n_32996 ^ n_32985;
assign n_33007 = n_32997 ^ n_32965;
assign n_33008 = n_32997 ^ n_32976;
assign n_33009 = ~n_32992 & n_32998;
assign n_33010 = n_32999 ^ n_32223;
assign n_33011 = n_33000 ^ n_32364;
assign n_33012 = ~n_32984 & ~n_33003;
assign n_33013 = n_33003 ^ n_32984;
assign n_33014 = ~n_33004 & n_33002;
assign n_33015 = n_33004 ^ n_31208;
assign n_33016 = n_33005 ^ n_32498;
assign n_33017 = ~n_31965 & ~n_33006;
assign n_33018 = ~n_32976 & n_33007;
assign n_33019 = n_33008 ^ n_32966;
assign n_33020 = n_33008 ^ n_32977;
assign n_33021 = n_33009 ^ x339;
assign n_33022 = n_33010 ^ n_32388;
assign n_33023 = n_33010 ^ n_32395;
assign n_33024 = n_33011 ^ n_31248;
assign n_33025 = n_33013 ^ n_32537;
assign n_33026 = n_33014 ^ n_31208;
assign n_33027 = n_33015 ^ x338;
assign n_33028 = n_33016 ^ n_33013;
assign n_33029 = n_33017 ^ n_32498;
assign n_33030 = n_33018 ^ n_31000;
assign n_33031 = n_32977 & ~n_33019;
assign n_33032 = n_32967 & n_33020;
assign n_33033 = n_33020 ^ n_32967;
assign n_33034 = n_33021 ^ n_33015;
assign n_33035 = n_33021 ^ x338;
assign n_33036 = n_32395 & n_33022;
assign n_33037 = ~n_31777 & n_33023;
assign n_33038 = n_33023 ^ n_32758;
assign n_33039 = n_33026 ^ n_33011;
assign n_33040 = n_33026 ^ n_33024;
assign n_33041 = n_33028 & ~n_33025;
assign n_33042 = n_33028 ^ n_32537;
assign n_33043 = n_33030 ^ n_33029;
assign n_33044 = n_33030 ^ n_31041;
assign n_33045 = n_33031 ^ x38;
assign n_33046 = n_33027 & ~n_33034;
assign n_33047 = n_33035 ^ n_33015;
assign n_33048 = n_33036 ^ n_32242;
assign n_33049 = n_33037 ^ n_32388;
assign n_33050 = ~n_33024 & ~n_33039;
assign n_33051 = n_33040 ^ x337;
assign n_33052 = n_33041 ^ n_32537;
assign n_33053 = n_31990 & ~n_33042;
assign n_33054 = n_33043 ^ n_31041;
assign n_33055 = n_33043 & n_33044;
assign n_33056 = n_33045 ^ x37;
assign n_33057 = n_33046 ^ x338;
assign n_33058 = ~n_33047 & ~n_33012;
assign n_33059 = n_33012 ^ n_33047;
assign n_33060 = n_33048 ^ n_32408;
assign n_33061 = n_33048 ^ n_32416;
assign n_33062 = n_33049 ^ n_31300;
assign n_33063 = n_33050 ^ n_31248;
assign n_33064 = n_33052 ^ n_32569;
assign n_33065 = n_33053 ^ n_32537;
assign n_33066 = n_33054 ^ x37;
assign n_33067 = n_33045 ^ n_33054;
assign n_33068 = n_33055 ^ n_31041;
assign n_33069 = n_33056 ^ n_33054;
assign n_33070 = n_33057 ^ n_33040;
assign n_33071 = n_33057 ^ x337;
assign n_33072 = n_33059 ^ n_32569;
assign n_33073 = n_33052 ^ n_33059;
assign n_33074 = n_32416 & n_33060;
assign n_33075 = ~n_31791 & ~n_33061;
assign n_33076 = n_33061 ^ n_32777;
assign n_33077 = n_33063 ^ n_33049;
assign n_33078 = n_33063 ^ n_31300;
assign n_33079 = n_33064 ^ n_33059;
assign n_33080 = n_33065 ^ n_31077;
assign n_33081 = n_33066 & ~n_33067;
assign n_33082 = n_33068 ^ n_33065;
assign n_33083 = n_33032 & n_33069;
assign n_33084 = n_33069 ^ n_33032;
assign n_33085 = ~n_33051 & n_33070;
assign n_33086 = n_33071 ^ n_33040;
assign n_33087 = ~n_33072 & ~n_33073;
assign n_33088 = n_33074 ^ n_32262;
assign n_33089 = n_33075 ^ n_32408;
assign n_33090 = ~n_33062 & ~n_33077;
assign n_33091 = n_33078 ^ n_33049;
assign n_33092 = n_32019 & ~n_33079;
assign n_33093 = n_33068 ^ n_33080;
assign n_33094 = n_33081 ^ x37;
assign n_33095 = ~n_33080 & n_33082;
assign n_33096 = n_33085 ^ x337;
assign n_33097 = n_33086 & n_33058;
assign n_33098 = n_33058 ^ n_33086;
assign n_33099 = n_33087 ^ n_32569;
assign n_33100 = n_33088 ^ n_32431;
assign n_33101 = n_33088 ^ n_32440;
assign n_33102 = n_33089 ^ n_31327;
assign n_33103 = n_33090 ^ n_31300;
assign n_33104 = n_33091 ^ x336;
assign n_33105 = n_33092 ^ n_32569;
assign n_33106 = n_33093 ^ x36;
assign n_33107 = n_33094 ^ n_33093;
assign n_33108 = n_33094 ^ x36;
assign n_33109 = n_33095 ^ n_31077;
assign n_33110 = n_33096 ^ n_33091;
assign n_33111 = n_33098 ^ n_32603;
assign n_33112 = n_33099 ^ n_33098;
assign n_33113 = n_33099 ^ n_32603;
assign n_33114 = n_32440 & n_33100;
assign n_33115 = ~n_31817 & n_33101;
assign n_33116 = n_33101 ^ n_32798;
assign n_33117 = n_33089 ^ n_33103;
assign n_33118 = n_33102 ^ n_33103;
assign n_33119 = n_33106 & ~n_33107;
assign n_33120 = n_33108 ^ n_33093;
assign n_33121 = n_33109 ^ n_33105;
assign n_33122 = n_33109 ^ n_31112;
assign n_33123 = ~n_33110 & n_33104;
assign n_33124 = n_33110 ^ x336;
assign n_33125 = ~n_33111 & n_33112;
assign n_33126 = n_33113 ^ n_33098;
assign n_33127 = n_33114 ^ n_32280;
assign n_33128 = n_33115 ^ n_32431;
assign n_33129 = ~n_33102 & ~n_33117;
assign n_33130 = n_33118 ^ x351;
assign n_33131 = n_33119 ^ x36;
assign n_33132 = n_33083 & n_33120;
assign n_33133 = n_33120 ^ n_33083;
assign n_33134 = n_33121 ^ n_31112;
assign n_33135 = ~n_33121 & n_33122;
assign n_33136 = n_33123 ^ x336;
assign n_33137 = n_33097 & ~n_33124;
assign n_33138 = n_33124 ^ n_33097;
assign n_33139 = n_33125 ^ n_32603;
assign n_33140 = n_32036 & n_33126;
assign n_33141 = n_33127 ^ n_32457;
assign n_33142 = n_33127 ^ n_32301;
assign n_33143 = n_33128 ^ n_31381;
assign n_33144 = n_33129 ^ n_31327;
assign n_33145 = n_33131 ^ n_33134;
assign n_33146 = n_33134 ^ x35;
assign n_33147 = n_33135 ^ n_31112;
assign n_33148 = n_33136 ^ n_33118;
assign n_33149 = n_33136 ^ n_33130;
assign n_33150 = n_33138 ^ n_32642;
assign n_33151 = n_33139 ^ n_33138;
assign n_33152 = n_33139 ^ n_32642;
assign n_33153 = n_33140 ^ n_32603;
assign n_33154 = ~n_32469 & n_33141;
assign n_33155 = n_33142 ^ n_32457;
assign n_33156 = n_33144 ^ n_33128;
assign n_33157 = n_33145 ^ x35;
assign n_33158 = n_33145 & ~n_33146;
assign n_33159 = ~n_33130 & n_33148;
assign n_33160 = n_33149 & n_33137;
assign n_33161 = n_33137 ^ n_33149;
assign n_33162 = n_33150 & ~n_33151;
assign n_33163 = n_33152 ^ n_33138;
assign n_33164 = n_33147 ^ n_33153;
assign n_33165 = n_33153 ^ n_31139;
assign n_33166 = n_33154 ^ n_32301;
assign n_33167 = n_31831 & n_33155;
assign n_33168 = n_33155 ^ n_32810;
assign n_33169 = ~n_33156 & n_33143;
assign n_33170 = n_33156 ^ n_31381;
assign n_33171 = ~n_33132 & n_33157;
assign n_33172 = n_33157 ^ n_33132;
assign n_33173 = n_33158 ^ x35;
assign n_33174 = n_33159 ^ x351;
assign n_33175 = n_33161 ^ n_32685;
assign n_33176 = n_33162 ^ n_32642;
assign n_33177 = ~n_32058 & ~n_33163;
assign n_33178 = n_33164 ^ n_31139;
assign n_33179 = ~n_33164 & ~n_33165;
assign n_33180 = n_33166 ^ n_32481;
assign n_33181 = n_33166 ^ n_32323;
assign n_33182 = n_33167 ^ n_32457;
assign n_33183 = n_33169 ^ n_31381;
assign n_33184 = n_33170 ^ x350;
assign n_33185 = n_33173 ^ x34;
assign n_33186 = n_33170 ^ n_33174;
assign n_33187 = n_33176 ^ n_33161;
assign n_33188 = n_33176 ^ n_33175;
assign n_33189 = n_33177 ^ n_32642;
assign n_33190 = n_33178 ^ x34;
assign n_33191 = n_33173 ^ n_33178;
assign n_33192 = n_33179 ^ n_31139;
assign n_33193 = ~n_32494 & n_33180;
assign n_33194 = n_33181 ^ n_32481;
assign n_33195 = n_33182 ^ n_31409;
assign n_33196 = n_33182 ^ n_33183;
assign n_33197 = n_33184 ^ n_33174;
assign n_33198 = n_33185 ^ n_33178;
assign n_33199 = ~n_33184 & n_33186;
assign n_33200 = n_33175 & n_33187;
assign n_33201 = ~n_32070 & ~n_33188;
assign n_33202 = n_33189 ^ n_31188;
assign n_33203 = n_33190 & ~n_33191;
assign n_33204 = n_33192 ^ n_33189;
assign n_33205 = n_33193 ^ n_32323;
assign n_33206 = n_31852 & n_33194;
assign n_33207 = n_33194 ^ n_32834;
assign n_33208 = n_33195 ^ n_33183;
assign n_33209 = ~n_33195 & n_33196;
assign n_33210 = n_33197 & n_33160;
assign n_33211 = n_33160 ^ n_33197;
assign n_33212 = ~n_33171 & n_33198;
assign n_33213 = n_33198 ^ n_33171;
assign n_33214 = n_33199 ^ x350;
assign n_33215 = n_33200 ^ n_32685;
assign n_33216 = n_33201 ^ n_32685;
assign n_33217 = n_33192 ^ n_33202;
assign n_33218 = n_33203 ^ x34;
assign n_33219 = n_33202 & n_33204;
assign n_33220 = n_33205 ^ n_32529;
assign n_33221 = n_33205 ^ n_32519;
assign n_33222 = n_33206 ^ n_32481;
assign n_33223 = n_33208 ^ x349;
assign n_33224 = n_33209 ^ n_31409;
assign n_33225 = n_33211 ^ n_32709;
assign n_33226 = n_33208 ^ n_33214;
assign n_33227 = n_33215 ^ n_33211;
assign n_33228 = n_33216 ^ n_31225;
assign n_33229 = n_33217 ^ x33;
assign n_33230 = n_33218 ^ n_33217;
assign n_33231 = n_33219 ^ n_31188;
assign n_33232 = n_31871 & ~n_33220;
assign n_33233 = n_33220 ^ n_32852;
assign n_33234 = n_32529 & ~n_33221;
assign n_33235 = n_33222 ^ n_31449;
assign n_33236 = n_33223 ^ n_33214;
assign n_33237 = n_33224 ^ n_33222;
assign n_33238 = n_33223 & ~n_33226;
assign n_33239 = ~n_33227 & n_33225;
assign n_33240 = n_33227 ^ n_32709;
assign n_33241 = n_33218 ^ n_33229;
assign n_33242 = n_33229 & ~n_33230;
assign n_33243 = n_33231 ^ n_33228;
assign n_33244 = n_33231 ^ n_33216;
assign n_33245 = n_33232 ^ n_32519;
assign n_33246 = n_33234 ^ n_32341;
assign n_33247 = n_33210 & ~n_33236;
assign n_33248 = n_33236 ^ n_33210;
assign n_33249 = n_33237 & n_33235;
assign n_33250 = n_33237 ^ n_31449;
assign n_33251 = n_33238 ^ x349;
assign n_33252 = n_33239 ^ n_32709;
assign n_33253 = ~n_32087 & n_33240;
assign n_33254 = ~n_33212 & ~n_33241;
assign n_33255 = n_33241 ^ n_33212;
assign n_33256 = n_33242 ^ x33;
assign n_33257 = n_33243 ^ x32;
assign n_33258 = n_33228 & n_33244;
assign n_33259 = n_33245 ^ n_31491;
assign n_33260 = n_33246 ^ n_32552;
assign n_33261 = n_33248 ^ n_32729;
assign n_33262 = n_33249 ^ n_31449;
assign n_33263 = n_33250 ^ x348;
assign n_33264 = n_33250 ^ n_33251;
assign n_33265 = n_33252 ^ n_33248;
assign n_33266 = n_33253 ^ n_32709;
assign n_33267 = n_33256 ^ x32;
assign n_33268 = n_33243 ^ n_33256;
assign n_33269 = n_33257 ^ n_33256;
assign n_33270 = n_33258 ^ n_31225;
assign n_33271 = n_33260 ^ n_32361;
assign n_33272 = n_33260 & n_32565;
assign n_33273 = n_33245 ^ n_33262;
assign n_33274 = n_33259 ^ n_33262;
assign n_33275 = n_33263 ^ n_33251;
assign n_33276 = ~n_33263 & n_33264;
assign n_33277 = n_33265 & n_33261;
assign n_33278 = n_33265 ^ n_32729;
assign n_33279 = n_33266 ^ n_31271;
assign n_33280 = n_33267 & n_33268;
assign n_33281 = n_33254 & n_33269;
assign n_33282 = n_33269 ^ n_33254;
assign n_33283 = n_33270 ^ n_31271;
assign n_33284 = n_33270 ^ n_33266;
assign n_33285 = n_31898 & ~n_33271;
assign n_33286 = n_32873 ^ n_33271;
assign n_33287 = n_33272 ^ n_32361;
assign n_33288 = n_33259 & n_33273;
assign n_33289 = n_33274 ^ x347;
assign n_33290 = n_33247 & n_33275;
assign n_33291 = n_33275 ^ n_33247;
assign n_33292 = n_33276 ^ x348;
assign n_33293 = n_33277 ^ n_32729;
assign n_33294 = ~n_32111 & n_33278;
assign n_33295 = n_33280 ^ x32;
assign n_33296 = n_33283 ^ n_33266;
assign n_33297 = ~n_33279 & ~n_33284;
assign n_33298 = n_33285 ^ n_32552;
assign n_33299 = n_33287 ^ n_32592;
assign n_33300 = n_33287 ^ n_32380;
assign n_33301 = n_33288 ^ n_31491;
assign n_33302 = n_33291 ^ n_32741;
assign n_33303 = n_33274 ^ n_33292;
assign n_33304 = n_33289 ^ n_33292;
assign n_33305 = n_33293 ^ n_33291;
assign n_33306 = n_33294 ^ n_32729;
assign n_33307 = n_33295 ^ x47;
assign n_33308 = n_33296 ^ x47;
assign n_33309 = n_33295 ^ n_33296;
assign n_33310 = n_33297 ^ n_31271;
assign n_33311 = n_33298 ^ n_31534;
assign n_33312 = n_33299 ^ n_32380;
assign n_33313 = ~n_33299 & n_33300;
assign n_33314 = n_33301 ^ n_33298;
assign n_33315 = n_33289 & ~n_33303;
assign n_33316 = n_33290 & ~n_33304;
assign n_33317 = n_33304 ^ n_33290;
assign n_33318 = n_33305 & n_33302;
assign n_33319 = n_33305 ^ n_32741;
assign n_33320 = n_33306 ^ n_31307;
assign n_33321 = n_33307 ^ n_33296;
assign n_33322 = ~n_33308 & n_33309;
assign n_33323 = n_33310 ^ n_31307;
assign n_33324 = n_33310 ^ n_33306;
assign n_33325 = n_31917 & n_33312;
assign n_33326 = n_32656 ^ n_33313;
assign n_33327 = n_33314 & ~n_33311;
assign n_33328 = n_33314 ^ n_31534;
assign n_33329 = n_33315 ^ x347;
assign n_33330 = n_33317 ^ n_32762;
assign n_33331 = n_33318 ^ n_32741;
assign n_33332 = ~n_32126 & ~n_33319;
assign n_33333 = n_33321 & n_33281;
assign n_33334 = n_33281 ^ n_33321;
assign n_33335 = n_33322 ^ x47;
assign n_33336 = n_33323 ^ n_33306;
assign n_33337 = ~n_33320 & ~n_33324;
assign n_33338 = n_33325 ^ n_32592;
assign n_33339 = ~n_31940 & n_33326;
assign n_33340 = n_32907 ^ n_33326;
assign n_33341 = n_33327 ^ n_31534;
assign n_33342 = n_33328 ^ x346;
assign n_33343 = n_33328 ^ n_33329;
assign n_33344 = n_33331 ^ n_33317;
assign n_33345 = n_33332 ^ n_32741;
assign n_33346 = n_33335 ^ n_33336;
assign n_33347 = n_33336 ^ x46;
assign n_33348 = n_33337 ^ n_31307;
assign n_33349 = n_33338 ^ n_31576;
assign n_33350 = n_33339 ^ n_32618;
assign n_33351 = n_33340 ^ n_32889;
assign n_33352 = n_33341 ^ n_33338;
assign n_33353 = n_33342 ^ n_33329;
assign n_33354 = n_33342 & ~n_33343;
assign n_33355 = n_33344 & ~n_33330;
assign n_33356 = n_33344 ^ n_32762;
assign n_33357 = n_33345 ^ n_31337;
assign n_33358 = n_33346 ^ x46;
assign n_33359 = ~n_33346 & n_33347;
assign n_33360 = n_33348 ^ n_31337;
assign n_33361 = n_33348 ^ n_33345;
assign n_33362 = n_33341 ^ n_33349;
assign n_33363 = n_33350 ^ n_31604;
assign n_33364 = ~n_33349 & n_33352;
assign n_33365 = n_33316 & ~n_33353;
assign n_33366 = n_33353 ^ n_33316;
assign n_33367 = n_33354 ^ x346;
assign n_33368 = n_33355 ^ n_32762;
assign n_33369 = ~n_32146 & ~n_33356;
assign n_33370 = ~n_33333 & n_33358;
assign n_33371 = n_33358 ^ n_33333;
assign n_33372 = n_33359 ^ x46;
assign n_33373 = n_33360 ^ n_33345;
assign n_33374 = n_33357 & ~n_33361;
assign n_33375 = n_33362 ^ x345;
assign n_33376 = n_33364 ^ n_31576;
assign n_33377 = n_33366 ^ n_32780;
assign n_33378 = n_33362 ^ n_33367;
assign n_33379 = n_33368 ^ n_33366;
assign n_33380 = n_33369 ^ n_32762;
assign n_33381 = n_33372 ^ x45;
assign n_33382 = n_33373 ^ x45;
assign n_33383 = n_33372 ^ n_33373;
assign n_33384 = n_33374 ^ n_31337;
assign n_33385 = n_33375 ^ n_33367;
assign n_33386 = n_33376 ^ n_33363;
assign n_33387 = n_33368 ^ n_33377;
assign n_33388 = n_33375 & ~n_33378;
assign n_33389 = n_33377 & n_33379;
assign n_33390 = n_33380 ^ n_31386;
assign n_33391 = n_33381 ^ n_33373;
assign n_33392 = n_33382 & ~n_33383;
assign n_33393 = n_33384 ^ n_33380;
assign n_33394 = n_33365 & ~n_33385;
assign n_33395 = n_33385 ^ n_33365;
assign n_33396 = n_33386 ^ x344;
assign n_33397 = n_32165 & n_33387;
assign n_33398 = n_33388 ^ x345;
assign n_33399 = n_33389 ^ n_32780;
assign n_33400 = n_33384 ^ n_33390;
assign n_33401 = ~n_33370 & ~n_33391;
assign n_33402 = n_33391 ^ n_33370;
assign n_33403 = n_33392 ^ x45;
assign n_33404 = n_33390 & ~n_33393;
assign n_33405 = n_33395 ^ n_32805;
assign n_33406 = n_33397 ^ n_32780;
assign n_33407 = n_33398 ^ n_33396;
assign n_33408 = n_33399 ^ n_33395;
assign n_33409 = n_33400 ^ x44;
assign n_33410 = n_33403 ^ n_33400;
assign n_33411 = n_33404 ^ n_31386;
assign n_33412 = n_33406 ^ n_31428;
assign n_33413 = n_33407 ^ n_33394;
assign n_33414 = ~n_33408 & n_33405;
assign n_33415 = n_33408 ^ n_32805;
assign n_33416 = n_33403 ^ n_33409;
assign n_33417 = n_33409 & ~n_33410;
assign n_33418 = n_33411 ^ n_31428;
assign n_33419 = n_33411 ^ n_33406;
assign n_33420 = n_33413 ^ n_32817;
assign n_33421 = n_33414 ^ n_32805;
assign n_33422 = ~n_32192 & ~n_33415;
assign n_33423 = n_33401 & ~n_33416;
assign n_33424 = n_33416 ^ n_33401;
assign n_33425 = n_33417 ^ x44;
assign n_33426 = n_33418 ^ n_33406;
assign n_33427 = ~n_33412 & n_33419;
assign n_33428 = n_33421 ^ n_33413;
assign n_33429 = n_33421 ^ n_32817;
assign n_33430 = n_33422 ^ n_32805;
assign n_33431 = ~n_32938 & n_33424;
assign n_33432 = n_33424 ^ n_32938;
assign n_33433 = n_33424 ^ n_32930;
assign n_33434 = n_33426 ^ x43;
assign n_33435 = n_33425 ^ n_33426;
assign n_33436 = n_33427 ^ n_31428;
assign n_33437 = ~n_33420 & ~n_33428;
assign n_33438 = n_33429 ^ n_33413;
assign n_33439 = n_33430 ^ n_31475;
assign n_33440 = n_33431 ^ n_32975;
assign n_33441 = ~n_32437 & n_33432;
assign n_33442 = n_33425 ^ n_33434;
assign n_33443 = ~n_33434 & n_33435;
assign n_33444 = n_33436 ^ n_33430;
assign n_33445 = n_33437 ^ n_32817;
assign n_33446 = ~n_32206 & n_33438;
assign n_33447 = n_33436 ^ n_33439;
assign n_33448 = n_33441 ^ n_32938;
assign n_33449 = n_32939 ^ n_33441;
assign n_33450 = n_33423 & n_33442;
assign n_33451 = n_33442 ^ n_33423;
assign n_33452 = n_33443 ^ x43;
assign n_33453 = n_33439 & n_33444;
assign n_33454 = n_33445 ^ n_32841;
assign n_33455 = n_33445 ^ n_32465;
assign n_33456 = n_33446 ^ n_32817;
assign n_33457 = n_33447 ^ x42;
assign n_33458 = n_31896 & n_33448;
assign n_33459 = x263 & n_33449;
assign n_33460 = n_33449 ^ x263;
assign n_33461 = n_33451 ^ n_33431;
assign n_33462 = n_33451 ^ n_33440;
assign n_33463 = n_33452 ^ n_33447;
assign n_33464 = n_33453 ^ n_31475;
assign n_33465 = n_32847 & n_33454;
assign n_33466 = n_33455 ^ n_32841;
assign n_33467 = n_33456 ^ n_31513;
assign n_33468 = n_33452 ^ n_33457;
assign n_33469 = n_33458 ^ n_31923;
assign n_33470 = n_33459 ^ x262;
assign n_33471 = n_33440 & n_33461;
assign n_33472 = n_32453 & n_33462;
assign n_33473 = n_33457 & ~n_33463;
assign n_33474 = n_33464 ^ n_31513;
assign n_33475 = n_33464 ^ n_33456;
assign n_33476 = n_33465 ^ n_32465;
assign n_33477 = n_32225 & n_33466;
assign n_33478 = ~n_33450 & n_33468;
assign n_33479 = n_33468 ^ n_33450;
assign n_33480 = n_33471 ^ n_32975;
assign n_33481 = n_33472 ^ n_32975;
assign n_33482 = n_33473 ^ x42;
assign n_33483 = n_33474 ^ n_33456;
assign n_33484 = n_33467 & n_33475;
assign n_33485 = n_33476 ^ n_32855;
assign n_33486 = n_33476 ^ n_32861;
assign n_33487 = n_33477 ^ n_32841;
assign n_33488 = n_33479 ^ n_33006;
assign n_33489 = n_33480 ^ n_33479;
assign n_33490 = n_33481 ^ n_33458;
assign n_33491 = n_33481 ^ n_33469;
assign n_33492 = n_33482 ^ n_33483;
assign n_33493 = n_33483 ^ x41;
assign n_33494 = n_33484 ^ n_31513;
assign n_33495 = ~n_32861 & ~n_33485;
assign n_33496 = n_32250 & n_33486;
assign n_33497 = n_33487 ^ n_31542;
assign n_33498 = n_33489 & ~n_33488;
assign n_33499 = n_33489 ^ n_33006;
assign n_33500 = ~n_33469 & n_33490;
assign n_33501 = n_33491 ^ n_33459;
assign n_33502 = n_33491 ^ x262;
assign n_33503 = n_33492 ^ x41;
assign n_33504 = n_33492 & ~n_33493;
assign n_33505 = n_33494 ^ n_33487;
assign n_33506 = n_33495 ^ n_32516;
assign n_33507 = n_33496 ^ n_32855;
assign n_33508 = n_33498 ^ n_33006;
assign n_33509 = ~n_32498 & n_33499;
assign n_33510 = n_33500 ^ n_31923;
assign n_33511 = n_33470 & ~n_33501;
assign n_33512 = n_33502 ^ n_33459;
assign n_33513 = ~n_33478 & n_33503;
assign n_33514 = n_33503 ^ n_33478;
assign n_33515 = n_33504 ^ x41;
assign n_33516 = n_33505 ^ n_31542;
assign n_33517 = n_33505 & n_33497;
assign n_33518 = n_33506 ^ n_32880;
assign n_33519 = n_33506 ^ n_32571;
assign n_33520 = n_33507 ^ n_31584;
assign n_33521 = n_33508 ^ n_33042;
assign n_33522 = n_33509 ^ n_33006;
assign n_33523 = n_33511 ^ x262;
assign n_33524 = ~n_33460 & ~n_33512;
assign n_33525 = n_33512 ^ n_33460;
assign n_33526 = n_33514 ^ n_33042;
assign n_33527 = n_33508 ^ n_33514;
assign n_33528 = n_33516 ^ x40;
assign n_33529 = n_33515 ^ n_33516;
assign n_33530 = n_33517 ^ n_31542;
assign n_33531 = n_32886 & ~n_33518;
assign n_33532 = n_33519 ^ n_32880;
assign n_33533 = n_33521 ^ n_33514;
assign n_33534 = n_33522 ^ n_31965;
assign n_33535 = n_33510 ^ n_33522;
assign n_33536 = n_33523 ^ x261;
assign n_33537 = n_33526 & ~n_33527;
assign n_33538 = n_33515 ^ n_33528;
assign n_33539 = n_33528 & ~n_33529;
assign n_33540 = n_33530 ^ n_33520;
assign n_33541 = n_33530 ^ n_33507;
assign n_33542 = n_33531 ^ n_32571;
assign n_33543 = n_32269 & n_33532;
assign n_33544 = ~n_32537 & ~n_33533;
assign n_33545 = n_33510 ^ n_33534;
assign n_33546 = n_33534 & ~n_33535;
assign n_33547 = n_33537 ^ n_33042;
assign n_33548 = n_33513 ^ n_33538;
assign n_33549 = n_33538 & ~n_33513;
assign n_33550 = n_33539 ^ x40;
assign n_33551 = n_33540 ^ x55;
assign n_33552 = ~n_33520 & ~n_33541;
assign n_33553 = n_33542 ^ n_32894;
assign n_33554 = n_33542 ^ n_32900;
assign n_33555 = n_33543 ^ n_32880;
assign n_33556 = n_33544 ^ n_33042;
assign n_33557 = n_33545 ^ x261;
assign n_33558 = n_33523 ^ n_33545;
assign n_33559 = n_33536 ^ n_33545;
assign n_33560 = n_33546 ^ n_31965;
assign n_33561 = n_33548 ^ n_33079;
assign n_33562 = n_33547 ^ n_33548;
assign n_33563 = n_33550 ^ n_33540;
assign n_33564 = n_33552 ^ n_31584;
assign n_33565 = n_32900 & ~n_33553;
assign n_33566 = ~n_32288 & n_33554;
assign n_33567 = n_33555 ^ n_31636;
assign n_33568 = ~n_33557 & n_33558;
assign n_33569 = n_33524 & n_33559;
assign n_33570 = n_33559 ^ n_33524;
assign n_33571 = n_33556 ^ n_33560;
assign n_33572 = n_33560 ^ n_31990;
assign n_33573 = n_33547 ^ n_33561;
assign n_33574 = ~n_33561 & n_33562;
assign n_33575 = n_33563 ^ x55;
assign n_33576 = ~n_33563 & n_33551;
assign n_33577 = n_33564 ^ n_33555;
assign n_33578 = n_33565 ^ n_32623;
assign n_33579 = n_33566 ^ n_32894;
assign n_33580 = n_33564 ^ n_33567;
assign n_33581 = n_33568 ^ x261;
assign n_33582 = n_33571 ^ n_31990;
assign n_33583 = ~n_33571 & ~n_33572;
assign n_33584 = n_32569 & n_33573;
assign n_33585 = n_33574 ^ n_33079;
assign n_33586 = n_33549 ^ n_33575;
assign n_33587 = n_33575 & n_33549;
assign n_33588 = n_33576 ^ x55;
assign n_33589 = ~n_33567 & ~n_33577;
assign n_33590 = n_33578 ^ n_32918;
assign n_33591 = n_33578 ^ n_32924;
assign n_33592 = n_33579 ^ n_31665;
assign n_33593 = n_33580 ^ x54;
assign n_33594 = n_33581 ^ n_33582;
assign n_33595 = n_33582 ^ x260;
assign n_33596 = n_33583 ^ n_31990;
assign n_33597 = n_33584 ^ n_33079;
assign n_33598 = n_33585 ^ n_33586;
assign n_33599 = n_33586 ^ n_33126;
assign n_33600 = n_33588 ^ n_33580;
assign n_33601 = n_33589 ^ n_31636;
assign n_33602 = n_32924 & n_33590;
assign n_33603 = n_32304 & n_33591;
assign n_33604 = n_33594 ^ x260;
assign n_33605 = ~n_33594 & n_33595;
assign n_33606 = n_33596 ^ n_32019;
assign n_33607 = n_33597 ^ n_33596;
assign n_33608 = n_33598 ^ n_33126;
assign n_33609 = ~n_33598 & ~n_33599;
assign n_33610 = n_33600 ^ x54;
assign n_33611 = n_33600 & ~n_33593;
assign n_33612 = n_33601 ^ n_31665;
assign n_33613 = n_33601 ^ n_33579;
assign n_33614 = n_33602 ^ n_32659;
assign n_33615 = n_33603 ^ n_32918;
assign n_33616 = n_33569 & ~n_33604;
assign n_33617 = n_33604 ^ n_33569;
assign n_33618 = n_33605 ^ x260;
assign n_33619 = n_33597 ^ n_33606;
assign n_33620 = n_33606 & n_33607;
assign n_33621 = n_32603 & n_33608;
assign n_33622 = n_33609 ^ n_33126;
assign n_33623 = n_33587 ^ n_33610;
assign n_33624 = ~n_33610 & n_33587;
assign n_33625 = n_33611 ^ x54;
assign n_33626 = n_33612 ^ n_33579;
assign n_33627 = ~n_33592 & n_33613;
assign n_33628 = n_33614 ^ n_32687;
assign n_33629 = n_33614 ^ n_32943;
assign n_33630 = n_33615 ^ n_31697;
assign n_33631 = n_33618 ^ n_33619;
assign n_33632 = n_33619 ^ x259;
assign n_33633 = n_33620 ^ n_32019;
assign n_33634 = n_33621 ^ n_33126;
assign n_33635 = n_33623 ^ n_33163;
assign n_33636 = n_33622 ^ n_33623;
assign n_33637 = n_33625 ^ n_33626;
assign n_33638 = n_33626 ^ x53;
assign n_33639 = n_33627 ^ n_31665;
assign n_33640 = n_33628 ^ n_32943;
assign n_33641 = n_32952 & ~n_33629;
assign n_33642 = n_33631 ^ x259;
assign n_33643 = n_33631 & ~n_33632;
assign n_33644 = n_33634 ^ n_32036;
assign n_33645 = n_33633 ^ n_33634;
assign n_33646 = n_33622 ^ n_33635;
assign n_33647 = ~n_33635 & ~n_33636;
assign n_33648 = n_33637 ^ x53;
assign n_33649 = ~n_33637 & n_33638;
assign n_33650 = n_33639 ^ n_31697;
assign n_33651 = n_33639 ^ n_33615;
assign n_33652 = ~n_32325 & ~n_33640;
assign n_33653 = n_33641 ^ n_32687;
assign n_33654 = ~n_33616 & ~n_33642;
assign n_33655 = n_33642 ^ n_33616;
assign n_33656 = n_33643 ^ x259;
assign n_33657 = n_33633 ^ n_33644;
assign n_33658 = n_33644 & ~n_33645;
assign n_33659 = n_32642 & ~n_33646;
assign n_33660 = n_33460 ^ n_33646;
assign n_33661 = n_33647 ^ n_33163;
assign n_33662 = n_33648 ^ n_33624;
assign n_33663 = ~n_33624 & ~n_33648;
assign n_33664 = n_33649 ^ x53;
assign n_33665 = n_33650 ^ n_33615;
assign n_33666 = n_33630 & ~n_33651;
assign n_33667 = n_33652 ^ n_32943;
assign n_33668 = n_33653 ^ n_32981;
assign n_33669 = n_33653 ^ n_32970;
assign n_33670 = n_33656 ^ x258;
assign n_33671 = n_33657 ^ x258;
assign n_33672 = n_33656 ^ n_33657;
assign n_33673 = n_33658 ^ n_32036;
assign n_33674 = n_33659 ^ n_33163;
assign n_33675 = n_33662 ^ n_33188;
assign n_33676 = n_33661 ^ n_33662;
assign n_33677 = n_33665 ^ x52;
assign n_33678 = n_33664 ^ n_33665;
assign n_33679 = n_33666 ^ n_31697;
assign n_33680 = n_33667 ^ n_31717;
assign n_33681 = ~n_32344 & ~n_33668;
assign n_33682 = n_33668 ^ n_32967;
assign n_33683 = n_32981 & ~n_33669;
assign n_33684 = n_33670 ^ n_33657;
assign n_33685 = n_33671 & ~n_33672;
assign n_33686 = n_33674 ^ n_32058;
assign n_33687 = n_33673 ^ n_33674;
assign n_33688 = n_33661 ^ n_33675;
assign n_33689 = ~n_33675 & n_33676;
assign n_33690 = n_33664 ^ n_33677;
assign n_33691 = ~n_33677 & n_33678;
assign n_33692 = n_33679 ^ n_31717;
assign n_33693 = n_33679 ^ n_33667;
assign n_33694 = n_33681 ^ n_32970;
assign n_33695 = n_33683 ^ n_32714;
assign n_33696 = n_33654 & n_33684;
assign n_33697 = n_33684 ^ n_33654;
assign n_33698 = n_33685 ^ x258;
assign n_33699 = n_33673 ^ n_33686;
assign n_33700 = n_33686 & n_33687;
assign n_33701 = ~n_32685 & n_33688;
assign n_33702 = n_33525 ^ n_33688;
assign n_33703 = n_33689 ^ n_33188;
assign n_33704 = n_33663 ^ n_33690;
assign n_33705 = ~n_33690 & ~n_33663;
assign n_33706 = n_33691 ^ x52;
assign n_33707 = n_33692 ^ n_33667;
assign n_33708 = ~n_33680 & ~n_33693;
assign n_33709 = n_33694 ^ n_31733;
assign n_33710 = n_33695 ^ n_32990;
assign n_33711 = n_33699 ^ x257;
assign n_33712 = n_33698 ^ n_33699;
assign n_33713 = n_33700 ^ n_32058;
assign n_33714 = n_33701 ^ n_33188;
assign n_33715 = n_33704 ^ n_33240;
assign n_33716 = n_33703 ^ n_33704;
assign n_33717 = n_33707 ^ x51;
assign n_33718 = n_33706 ^ n_33707;
assign n_33719 = n_33708 ^ n_31717;
assign n_33720 = n_32734 ^ n_33710;
assign n_33721 = n_33710 & ~n_33001;
assign n_33722 = n_33698 ^ n_33711;
assign n_33723 = n_33711 & ~n_33712;
assign n_33724 = n_33714 ^ n_33713;
assign n_33725 = n_33714 ^ n_32070;
assign n_33726 = n_33703 ^ n_33715;
assign n_33727 = ~n_33715 & ~n_33716;
assign n_33728 = n_33706 ^ n_33717;
assign n_33729 = n_33717 & ~n_33718;
assign n_33730 = n_33719 ^ n_31733;
assign n_33731 = n_33719 ^ n_33694;
assign n_33732 = ~n_32364 & n_33720;
assign n_33733 = n_33033 ^ n_33720;
assign n_33734 = n_33721 ^ n_32734;
assign n_33735 = ~n_33696 & ~n_33722;
assign n_33736 = n_33722 ^ n_33696;
assign n_33737 = n_33723 ^ x257;
assign n_33738 = n_33724 ^ n_32070;
assign n_33739 = ~n_33724 & n_33725;
assign n_33740 = ~n_32709 & n_33726;
assign n_33741 = n_33570 ^ n_33726;
assign n_33742 = n_33727 ^ n_33240;
assign n_33743 = n_33705 ^ n_33728;
assign n_33744 = n_33728 & n_33705;
assign n_33745 = n_33729 ^ x51;
assign n_33746 = n_33730 ^ n_33694;
assign n_33747 = n_33709 & n_33731;
assign n_33748 = n_33732 ^ n_32990;
assign n_33749 = n_33734 ^ n_33023;
assign n_33750 = n_33734 ^ n_32758;
assign n_33751 = n_33737 ^ n_33738;
assign n_33752 = n_33738 ^ x256;
assign n_33753 = n_33739 ^ n_32070;
assign n_33754 = n_33740 ^ n_33240;
assign n_33755 = n_33743 ^ n_33278;
assign n_33756 = n_33742 ^ n_33743;
assign n_33757 = n_33745 ^ n_33746;
assign n_33758 = n_33746 ^ x50;
assign n_33759 = n_33747 ^ n_31733;
assign n_33760 = n_33748 ^ n_31758;
assign n_33761 = n_33038 & n_33749;
assign n_33762 = n_33750 ^ n_33023;
assign n_33763 = n_33751 ^ x256;
assign n_33764 = n_33751 & ~n_33752;
assign n_33765 = n_33754 ^ n_32087;
assign n_33766 = n_33753 ^ n_33754;
assign n_33767 = n_33742 ^ n_33755;
assign n_33768 = ~n_33755 & n_33756;
assign n_33769 = n_33757 ^ x50;
assign n_33770 = ~n_33757 & n_33758;
assign n_33771 = n_33759 ^ n_31758;
assign n_33772 = n_33748 ^ n_33759;
assign n_33773 = n_33761 ^ n_32758;
assign n_33774 = n_32388 & ~n_33762;
assign n_33775 = n_33084 ^ n_33762;
assign n_33776 = ~n_33763 & ~n_33735;
assign n_33777 = n_33735 ^ n_33763;
assign n_33778 = n_33764 ^ x256;
assign n_33779 = n_33753 ^ n_33765;
assign n_33780 = ~n_33765 & n_33766;
assign n_33781 = n_32729 & ~n_33767;
assign n_33782 = n_33617 ^ n_33767;
assign n_33783 = n_33768 ^ n_33278;
assign n_33784 = n_33769 ^ n_33744;
assign n_33785 = n_33744 & n_33769;
assign n_33786 = n_33770 ^ x50;
assign n_33787 = n_33748 ^ n_33771;
assign n_33788 = ~n_33760 & n_33772;
assign n_33789 = n_33773 ^ n_33061;
assign n_33790 = n_33773 ^ n_33076;
assign n_33791 = n_33774 ^ n_33023;
assign n_33792 = n_33779 ^ x271;
assign n_33793 = n_33778 ^ n_33779;
assign n_33794 = n_33780 ^ n_32087;
assign n_33795 = n_33781 ^ n_33278;
assign n_33796 = n_33783 ^ n_33784;
assign n_33797 = n_33784 ^ n_33319;
assign n_33798 = n_33786 ^ n_33787;
assign n_33799 = n_33787 ^ x49;
assign n_33800 = n_33788 ^ n_31758;
assign n_33801 = n_33076 & n_33789;
assign n_33802 = ~n_32408 & n_33790;
assign n_33803 = n_33133 ^ n_33790;
assign n_33804 = n_33791 ^ n_31777;
assign n_33805 = n_33778 ^ n_33792;
assign n_33806 = n_33792 & ~n_33793;
assign n_33807 = n_33795 ^ n_32111;
assign n_33808 = n_33794 ^ n_33795;
assign n_33809 = n_33796 ^ n_33319;
assign n_33810 = n_33796 & n_33797;
assign n_33811 = n_33798 ^ x49;
assign n_33812 = ~n_33798 & n_33799;
assign n_33813 = n_33800 ^ n_33791;
assign n_33814 = n_33800 ^ n_31777;
assign n_33815 = n_33801 ^ n_32777;
assign n_33816 = n_33802 ^ n_33061;
assign n_33817 = n_33805 & n_33776;
assign n_33818 = n_33776 ^ n_33805;
assign n_33819 = n_33806 ^ x271;
assign n_33820 = n_33794 ^ n_33807;
assign n_33821 = ~n_33807 & n_33808;
assign n_33822 = ~n_32741 & n_33809;
assign n_33823 = n_33655 ^ n_33809;
assign n_33824 = n_33810 ^ n_33319;
assign n_33825 = n_33811 ^ n_33785;
assign n_33826 = n_33785 & n_33811;
assign n_33827 = n_33812 ^ x49;
assign n_33828 = ~n_33804 & n_33813;
assign n_33829 = n_33814 ^ n_33791;
assign n_33830 = n_33815 ^ n_33116;
assign n_33831 = n_33815 ^ n_33101;
assign n_33832 = n_33816 ^ n_31791;
assign n_33833 = n_33820 ^ x270;
assign n_33834 = n_33819 ^ n_33820;
assign n_33835 = n_33821 ^ n_32111;
assign n_33836 = n_33822 ^ n_33319;
assign n_33837 = n_33824 ^ n_33825;
assign n_33838 = n_33825 ^ n_33356;
assign n_33839 = n_33828 ^ n_31777;
assign n_33840 = n_33829 ^ x48;
assign n_33841 = n_33829 ^ n_33827;
assign n_33842 = n_32431 & ~n_33830;
assign n_33843 = n_33172 ^ n_33830;
assign n_33844 = n_33116 & n_33831;
assign n_33845 = n_33819 ^ n_33833;
assign n_33846 = n_33833 & ~n_33834;
assign n_33847 = n_33836 ^ n_32126;
assign n_33848 = n_33835 ^ n_33836;
assign n_33849 = n_33837 ^ n_33356;
assign n_33850 = ~n_33837 & n_33838;
assign n_33851 = n_33839 ^ n_33816;
assign n_33852 = n_33839 ^ n_33832;
assign n_33853 = n_33840 ^ n_33827;
assign n_33854 = n_33840 & ~n_33841;
assign n_33855 = n_33842 ^ n_33101;
assign n_33856 = n_33844 ^ n_32798;
assign n_33857 = ~n_33817 & ~n_33845;
assign n_33858 = n_33845 ^ n_33817;
assign n_33859 = n_33846 ^ x270;
assign n_33860 = n_33835 ^ n_33847;
assign n_33861 = n_33847 & ~n_33848;
assign n_33862 = ~n_32762 & ~n_33849;
assign n_33863 = n_33697 ^ n_33849;
assign n_33864 = n_33850 ^ n_33356;
assign n_33865 = n_33832 & ~n_33851;
assign n_33866 = n_33852 ^ x63;
assign n_33867 = ~n_33826 & ~n_33853;
assign n_33868 = n_33853 ^ n_33826;
assign n_33869 = n_33854 ^ x48;
assign n_33870 = n_33855 ^ n_31817;
assign n_33871 = n_33856 ^ n_33168;
assign n_33872 = n_33856 ^ n_33155;
assign n_33873 = n_33860 ^ x269;
assign n_33874 = n_33859 ^ n_33860;
assign n_33875 = n_33861 ^ n_32126;
assign n_33876 = n_33862 ^ n_33356;
assign n_33877 = n_33864 ^ n_33387;
assign n_33878 = n_33865 ^ n_31791;
assign n_33879 = n_33868 ^ n_33387;
assign n_33880 = n_33868 ^ n_33864;
assign n_33881 = n_33869 ^ n_33852;
assign n_33882 = ~n_32457 & ~n_33871;
assign n_33883 = n_33213 ^ n_33871;
assign n_33884 = ~n_33168 & ~n_33872;
assign n_33885 = n_33859 ^ n_33873;
assign n_33886 = ~n_33873 & n_33874;
assign n_33887 = n_33876 ^ n_32146;
assign n_33888 = n_33876 ^ n_33875;
assign n_33889 = n_33868 ^ n_33877;
assign n_33890 = n_33878 ^ n_33855;
assign n_33891 = n_33878 ^ n_31817;
assign n_33892 = n_33879 & n_33880;
assign n_33893 = n_33881 & ~n_33866;
assign n_33894 = n_33881 ^ x63;
assign n_33895 = n_33882 ^ n_33155;
assign n_33896 = n_33884 ^ n_32810;
assign n_33897 = n_33857 & n_33885;
assign n_33898 = n_33885 ^ n_33857;
assign n_33899 = n_33886 ^ x269;
assign n_33900 = n_33887 ^ n_33875;
assign n_33901 = n_33887 & ~n_33888;
assign n_33902 = n_33736 ^ n_33889;
assign n_33903 = n_32780 & ~n_33889;
assign n_33904 = ~n_33870 & n_33890;
assign n_33905 = n_33891 ^ n_33855;
assign n_33906 = n_33892 ^ n_33387;
assign n_33907 = n_33893 ^ x63;
assign n_33908 = n_33894 & n_33867;
assign n_33909 = n_33867 ^ n_33894;
assign n_33910 = n_33895 ^ n_31831;
assign n_33911 = n_33896 ^ n_33207;
assign n_33912 = n_33896 ^ n_33194;
assign n_33913 = n_33899 ^ x268;
assign n_33914 = n_33900 ^ x268;
assign n_33915 = n_33900 ^ n_33899;
assign n_33916 = n_33901 ^ n_32146;
assign n_33917 = n_33903 ^ n_33387;
assign n_33918 = n_33904 ^ n_31817;
assign n_33919 = n_33905 ^ x62;
assign n_33920 = n_33907 ^ n_33905;
assign n_33921 = n_33909 ^ n_33415;
assign n_33922 = n_33909 ^ n_33906;
assign n_33923 = ~n_32481 & n_33911;
assign n_33924 = n_33255 ^ n_33911;
assign n_33925 = ~n_33207 & n_33912;
assign n_33926 = n_33900 ^ n_33913;
assign n_33927 = ~n_33914 & n_33915;
assign n_33928 = n_33916 ^ n_32165;
assign n_33929 = n_33917 ^ n_32165;
assign n_33930 = n_33917 ^ n_33916;
assign n_33931 = n_33918 ^ n_31831;
assign n_33932 = n_33918 ^ n_33895;
assign n_33933 = ~n_33920 & n_33919;
assign n_33934 = n_33920 ^ x62;
assign n_33935 = n_33921 ^ n_33906;
assign n_33936 = ~n_33921 & ~n_33922;
assign n_33937 = n_33923 ^ n_33194;
assign n_33938 = n_33925 ^ n_32834;
assign n_33939 = n_33897 ^ n_33926;
assign n_33940 = n_33926 & n_33897;
assign n_33941 = n_33927 ^ x268;
assign n_33942 = n_33917 ^ n_33928;
assign n_33943 = n_33929 & n_33930;
assign n_33944 = n_33931 ^ n_33895;
assign n_33945 = n_33910 & n_33932;
assign n_33946 = n_33933 ^ x62;
assign n_33947 = n_33934 & ~n_33908;
assign n_33948 = n_33908 ^ n_33934;
assign n_33949 = n_33777 ^ n_33935;
assign n_33950 = n_32805 & ~n_33935;
assign n_33951 = n_33936 ^ n_33415;
assign n_33952 = n_33937 ^ n_31852;
assign n_33953 = n_33938 ^ n_33233;
assign n_33954 = n_33938 ^ n_33220;
assign n_33955 = n_33941 ^ x267;
assign n_33956 = n_33942 ^ x267;
assign n_33957 = n_33942 ^ n_33941;
assign n_33958 = n_33943 ^ n_32165;
assign n_33959 = n_33944 ^ x61;
assign n_33960 = n_33945 ^ n_31831;
assign n_33961 = n_33946 ^ n_33944;
assign n_33962 = n_33948 ^ n_33438;
assign n_33963 = n_33950 ^ n_33415;
assign n_33964 = n_33948 ^ n_33951;
assign n_33965 = n_32519 & n_33953;
assign n_33966 = n_33282 ^ n_33953;
assign n_33967 = ~n_33233 & ~n_33954;
assign n_33968 = n_33942 ^ n_33955;
assign n_33969 = ~n_33956 & n_33957;
assign n_33970 = n_33946 ^ n_33959;
assign n_33971 = n_33960 ^ n_33952;
assign n_33972 = n_33960 ^ n_33937;
assign n_33973 = ~n_33959 & n_33961;
assign n_33974 = n_33962 ^ n_33951;
assign n_33975 = n_33963 ^ n_32192;
assign n_33976 = n_33963 ^ n_33958;
assign n_33977 = n_33962 & n_33964;
assign n_33978 = n_33965 ^ n_33220;
assign n_33979 = n_33967 ^ n_32852;
assign n_33980 = n_33940 & n_33968;
assign n_33981 = n_33968 ^ n_33940;
assign n_33982 = n_33969 ^ x267;
assign n_33983 = ~n_33947 & n_33970;
assign n_33984 = n_33970 ^ n_33947;
assign n_33985 = n_33971 ^ x60;
assign n_33986 = n_33952 & ~n_33972;
assign n_33987 = n_33973 ^ x61;
assign n_33988 = n_33818 ^ n_33974;
assign n_33989 = ~n_32817 & ~n_33974;
assign n_33990 = n_33975 ^ n_33958;
assign n_33991 = n_33975 & n_33976;
assign n_33992 = n_33977 ^ n_33438;
assign n_33993 = n_33978 ^ n_31871;
assign n_33994 = n_33286 ^ n_33979;
assign n_33995 = n_33979 ^ n_33271;
assign n_33996 = n_33984 ^ n_33466;
assign n_33997 = n_33986 ^ n_31852;
assign n_33998 = n_33987 ^ n_33985;
assign n_33999 = n_33987 ^ x60;
assign n_34000 = n_33987 ^ n_33971;
assign n_34001 = n_33989 ^ n_33438;
assign n_34002 = n_33990 ^ x266;
assign n_34003 = n_33990 ^ n_33982;
assign n_34004 = n_33991 ^ n_32192;
assign n_34005 = n_33992 ^ n_33984;
assign n_34006 = ~n_32552 & ~n_33994;
assign n_34007 = n_33334 ^ n_33994;
assign n_34008 = ~n_33286 & n_33995;
assign n_34009 = n_33997 ^ n_33993;
assign n_34010 = n_33997 ^ n_33978;
assign n_34011 = n_33998 & ~n_33983;
assign n_34012 = n_33983 ^ n_33998;
assign n_34013 = n_33999 & ~n_34000;
assign n_34014 = n_34001 ^ n_32206;
assign n_34015 = n_34002 ^ n_33982;
assign n_34016 = n_34002 & ~n_34003;
assign n_34017 = n_34001 ^ n_34004;
assign n_34018 = n_34005 & ~n_33996;
assign n_34019 = n_34005 ^ n_33466;
assign n_34020 = n_34006 ^ n_33271;
assign n_34021 = n_34008 ^ n_32873;
assign n_34022 = n_34009 ^ x59;
assign n_34023 = ~n_33993 & n_34010;
assign n_34024 = n_34012 ^ n_33486;
assign n_34025 = n_34013 ^ x60;
assign n_34026 = n_34014 ^ n_34004;
assign n_34027 = n_33980 & ~n_34015;
assign n_34028 = n_34015 ^ n_33980;
assign n_34029 = n_34016 ^ x266;
assign n_34030 = ~n_34014 & n_34017;
assign n_34031 = n_34018 ^ n_33466;
assign n_34032 = n_33858 ^ n_34019;
assign n_34033 = n_32841 & ~n_34019;
assign n_34034 = n_34020 ^ n_31898;
assign n_34035 = n_34021 ^ n_32889;
assign n_34036 = n_34021 ^ n_33312;
assign n_34037 = n_34023 ^ n_31871;
assign n_34038 = n_34025 ^ n_34022;
assign n_34039 = n_34025 ^ x59;
assign n_34040 = n_34025 ^ n_34009;
assign n_34041 = n_34026 ^ x265;
assign n_34042 = n_34026 ^ n_34029;
assign n_34043 = n_34029 ^ x265;
assign n_34044 = n_34030 ^ n_32206;
assign n_34045 = n_34012 ^ n_34031;
assign n_34046 = n_34024 ^ n_34031;
assign n_34047 = n_34033 ^ n_33466;
assign n_34048 = n_34035 ^ n_33312;
assign n_34049 = ~n_34035 & ~n_34036;
assign n_34050 = n_34037 ^ n_34034;
assign n_34051 = n_34037 ^ n_34020;
assign n_34052 = n_34011 ^ n_34038;
assign n_34053 = ~n_34038 & n_34011;
assign n_34054 = n_34039 & n_34040;
assign n_34055 = n_34041 & ~n_34042;
assign n_34056 = n_34026 ^ n_34043;
assign n_34057 = n_34024 & ~n_34045;
assign n_34058 = n_33898 ^ n_34046;
assign n_34059 = n_32855 & n_34046;
assign n_34060 = n_34047 ^ n_32225;
assign n_34061 = n_34047 ^ n_34044;
assign n_34062 = ~n_32592 & ~n_34048;
assign n_34063 = n_33351 ^ n_34049;
assign n_34064 = n_34050 ^ x58;
assign n_34065 = ~n_34034 & n_34051;
assign n_34066 = n_34052 ^ n_33532;
assign n_34067 = n_34054 ^ x59;
assign n_34068 = n_34055 ^ x265;
assign n_34069 = n_34027 & ~n_34056;
assign n_34070 = n_34056 ^ n_34027;
assign n_34071 = n_34057 ^ n_33486;
assign n_34072 = n_34059 ^ n_33486;
assign n_34073 = n_34060 ^ n_34044;
assign n_34074 = n_34060 & n_34061;
assign n_34075 = n_34062 ^ n_33312;
assign n_34076 = ~n_32618 & ~n_34063;
assign n_34077 = n_33402 ^ n_34063;
assign n_34078 = n_34065 ^ n_31898;
assign n_34079 = n_34067 ^ n_34064;
assign n_34080 = n_34067 ^ n_34050;
assign n_34081 = n_34071 ^ n_33532;
assign n_34082 = n_34052 ^ n_34071;
assign n_34083 = n_34072 ^ n_32250;
assign n_34084 = n_34073 ^ x264;
assign n_34085 = n_34073 ^ n_34068;
assign n_34086 = n_34074 ^ n_32225;
assign n_34087 = n_34075 ^ n_31917;
assign n_34088 = n_34076 ^ n_33326;
assign n_34089 = n_34077 ^ n_33371;
assign n_34090 = n_34075 ^ n_34078;
assign n_34091 = n_34053 & ~n_34079;
assign n_34092 = n_34079 ^ n_34053;
assign n_34093 = ~n_34064 & n_34080;
assign n_34094 = n_34052 ^ n_34081;
assign n_34095 = n_34066 & ~n_34082;
assign n_34096 = n_34084 ^ n_34068;
assign n_34097 = ~n_34084 & n_34085;
assign n_34098 = n_34072 ^ n_34086;
assign n_34099 = n_34083 ^ n_34086;
assign n_34100 = n_34087 ^ n_34078;
assign n_34101 = n_34087 & ~n_34090;
assign n_34102 = n_34092 ^ n_33554;
assign n_34103 = n_34093 ^ x58;
assign n_34104 = n_33939 ^ n_34094;
assign n_34105 = ~n_32880 & n_34094;
assign n_34106 = n_34095 ^ n_33532;
assign n_34107 = ~n_34069 & ~n_34096;
assign n_34108 = n_34096 ^ n_34069;
assign n_34109 = n_34097 ^ x264;
assign n_34110 = n_34083 & ~n_34098;
assign n_34111 = n_34099 ^ x279;
assign n_34112 = n_34100 ^ x57;
assign n_34113 = n_34101 ^ n_31917;
assign n_34114 = n_34103 ^ x57;
assign n_34115 = n_34103 ^ n_34100;
assign n_34116 = n_34105 ^ n_33532;
assign n_34117 = n_34092 ^ n_34106;
assign n_34118 = n_34102 ^ n_34106;
assign n_34119 = n_34099 ^ n_34109;
assign n_34120 = n_34109 ^ x279;
assign n_34121 = n_34110 ^ n_32250;
assign n_34122 = n_34103 ^ n_34112;
assign n_34123 = n_34113 ^ n_31940;
assign n_34124 = n_34114 & ~n_34115;
assign n_34125 = n_34116 ^ n_32269;
assign n_34126 = n_34102 & ~n_34117;
assign n_34127 = ~n_32894 & n_34118;
assign n_34128 = n_33981 ^ n_34118;
assign n_34129 = n_34111 & ~n_34119;
assign n_34130 = n_34099 ^ n_34120;
assign n_34131 = n_34121 ^ n_34116;
assign n_34132 = n_34091 ^ n_34122;
assign n_34133 = n_34122 & n_34091;
assign n_34134 = n_34123 ^ n_34088;
assign n_34135 = n_34124 ^ x57;
assign n_34136 = n_34126 ^ n_33554;
assign n_34137 = n_34127 ^ n_33554;
assign n_34138 = n_34129 ^ x279;
assign n_34139 = n_34107 & n_34130;
assign n_34140 = n_34130 ^ n_34107;
assign n_34141 = ~n_34131 & n_34125;
assign n_34142 = n_34131 ^ n_32269;
assign n_34143 = n_34132 ^ n_33591;
assign n_34144 = n_34134 ^ x56;
assign n_34145 = n_34132 ^ n_34136;
assign n_34146 = n_34137 ^ n_32288;
assign n_34147 = n_34141 ^ n_32269;
assign n_34148 = n_34142 ^ x278;
assign n_34149 = n_34142 ^ n_34138;
assign n_34150 = n_34143 ^ n_34136;
assign n_34151 = n_34135 ^ n_34144;
assign n_34152 = ~n_34143 & n_34145;
assign n_34153 = n_34137 ^ n_34147;
assign n_34154 = n_34147 ^ n_32288;
assign n_34155 = n_34148 ^ n_34138;
assign n_34156 = n_34148 & ~n_34149;
assign n_34157 = n_32918 & ~n_34150;
assign n_34158 = n_34028 ^ n_34150;
assign n_34159 = n_34151 ^ n_34133;
assign n_34160 = n_34152 ^ n_33591;
assign n_34161 = ~n_34146 & ~n_34153;
assign n_34162 = n_34137 ^ n_34154;
assign n_34163 = n_34139 & n_34155;
assign n_34164 = n_34155 ^ n_34139;
assign n_34165 = n_34156 ^ x278;
assign n_34166 = n_34157 ^ n_33591;
assign n_34167 = n_34159 ^ n_33640;
assign n_34168 = n_34160 ^ n_34159;
assign n_34169 = n_34161 ^ n_32288;
assign n_34170 = n_34162 ^ x277;
assign n_34171 = n_34165 ^ n_34162;
assign n_34172 = n_34166 ^ n_32304;
assign n_34173 = n_34168 & n_34167;
assign n_34174 = n_34168 ^ n_33640;
assign n_34175 = n_34166 ^ n_34169;
assign n_34176 = n_34169 ^ n_32304;
assign n_34177 = n_34171 & ~n_34170;
assign n_34178 = n_34171 ^ x277;
assign n_34179 = n_34173 ^ n_33640;
assign n_34180 = n_32943 & n_34174;
assign n_34181 = n_34070 ^ n_34174;
assign n_34182 = n_34172 & n_34175;
assign n_34183 = n_34166 ^ n_34176;
assign n_34184 = n_34177 ^ x277;
assign n_34185 = n_34163 & ~n_34178;
assign n_34186 = n_34178 ^ n_34163;
assign n_34187 = n_34179 ^ n_33668;
assign n_34188 = n_34179 ^ n_32967;
assign n_34189 = n_34180 ^ n_33640;
assign n_34190 = n_34182 ^ n_32304;
assign n_34191 = n_34183 ^ x276;
assign n_34192 = n_34183 ^ n_34184;
assign n_34193 = n_34184 ^ x276;
assign n_34194 = ~n_33682 & ~n_34187;
assign n_34195 = n_34188 ^ n_33668;
assign n_34196 = n_34189 ^ n_32325;
assign n_34197 = n_34190 ^ n_34189;
assign n_34198 = ~n_34191 & n_34192;
assign n_34199 = n_34183 ^ n_34193;
assign n_34200 = n_34194 ^ n_32967;
assign n_34201 = n_32970 & n_34195;
assign n_34202 = n_34108 ^ n_34195;
assign n_34203 = n_34197 & n_34196;
assign n_34204 = n_34197 ^ n_32325;
assign n_34205 = n_34198 ^ x276;
assign n_34206 = ~n_34185 & n_34199;
assign n_34207 = n_34199 ^ n_34185;
assign n_34208 = n_34200 ^ n_33720;
assign n_34209 = n_34200 ^ n_33733;
assign n_34210 = n_34201 ^ n_33668;
assign n_34211 = n_34203 ^ n_32325;
assign n_34212 = n_34204 ^ x275;
assign n_34213 = n_34204 ^ n_34205;
assign n_34214 = ~n_33733 & ~n_34208;
assign n_34215 = ~n_32990 & ~n_34209;
assign n_34216 = n_34209 ^ n_34140;
assign n_34217 = n_34210 ^ n_32344;
assign n_34218 = n_34210 ^ n_34211;
assign n_34219 = n_34211 ^ n_32344;
assign n_34220 = n_34212 ^ n_34205;
assign n_34221 = n_34212 & ~n_34213;
assign n_34222 = n_34214 ^ n_33033;
assign n_34223 = n_34215 ^ n_33720;
assign n_34224 = n_34217 & ~n_34218;
assign n_34225 = n_34210 ^ n_34219;
assign n_34226 = ~n_34206 & n_34220;
assign n_34227 = n_34220 ^ n_34206;
assign n_34228 = n_34221 ^ x275;
assign n_34229 = n_34222 ^ n_33762;
assign n_34230 = n_34222 ^ n_33775;
assign n_34231 = n_34223 ^ n_32364;
assign n_34232 = n_34224 ^ n_32344;
assign n_34233 = n_34225 ^ x274;
assign n_34234 = n_34225 ^ n_34228;
assign n_34235 = n_33775 & ~n_34229;
assign n_34236 = ~n_33023 & ~n_34230;
assign n_34237 = n_34164 ^ n_34230;
assign n_34238 = n_34223 ^ n_34232;
assign n_34239 = n_34231 ^ n_34232;
assign n_34240 = n_34233 ^ n_34228;
assign n_34241 = ~n_34233 & n_34234;
assign n_34242 = n_34235 ^ n_33084;
assign n_34243 = n_34236 ^ n_33762;
assign n_34244 = ~n_34231 & n_34238;
assign n_34245 = n_34239 ^ x273;
assign n_34246 = ~n_34226 & n_34240;
assign n_34247 = n_34240 ^ n_34226;
assign n_34248 = n_34241 ^ x274;
assign n_34249 = n_34242 ^ n_33790;
assign n_34250 = n_34242 ^ n_33803;
assign n_34251 = n_34243 ^ n_32388;
assign n_34252 = n_34244 ^ n_32364;
assign n_34253 = n_34239 ^ n_34248;
assign n_34254 = n_34248 ^ x273;
assign n_34255 = ~n_33803 & n_34249;
assign n_34256 = n_33061 & n_34250;
assign n_34257 = n_34250 ^ n_34186;
assign n_34258 = n_34243 ^ n_34252;
assign n_34259 = n_34252 ^ n_32388;
assign n_34260 = n_34245 & ~n_34253;
assign n_34261 = n_34239 ^ n_34254;
assign n_34262 = n_34255 ^ n_33133;
assign n_34263 = n_34256 ^ n_33790;
assign n_34264 = ~n_34251 & ~n_34258;
assign n_34265 = n_34243 ^ n_34259;
assign n_34266 = n_34260 ^ x273;
assign n_34267 = ~n_34246 & n_34261;
assign n_34268 = n_34261 ^ n_34246;
assign n_34269 = n_34262 ^ n_33830;
assign n_34270 = n_34262 ^ n_33843;
assign n_34271 = n_34263 ^ n_32408;
assign n_34272 = n_34264 ^ n_32388;
assign n_34273 = n_34265 ^ x272;
assign n_34274 = n_34265 ^ n_34266;
assign n_34275 = n_33843 & ~n_34269;
assign n_34276 = ~n_33101 & ~n_34270;
assign n_34277 = n_34270 ^ n_34207;
assign n_34278 = n_34263 ^ n_34272;
assign n_34279 = n_34273 ^ n_34266;
assign n_34280 = n_34273 & ~n_34274;
assign n_34281 = n_34275 ^ n_33172;
assign n_34282 = n_34276 ^ n_33830;
assign n_34283 = ~n_34278 & ~n_34271;
assign n_34284 = n_34278 ^ n_32408;
assign n_34285 = ~n_34267 & ~n_34279;
assign n_34286 = n_34279 ^ n_34267;
assign n_34287 = n_34280 ^ x272;
assign n_34288 = n_34281 ^ n_33871;
assign n_34289 = n_34282 ^ n_32431;
assign n_34290 = n_34283 ^ n_32408;
assign n_34291 = n_34284 ^ x287;
assign n_34292 = n_34284 ^ n_34287;
assign n_34293 = n_34287 ^ x287;
assign n_34294 = ~n_34288 & ~n_33883;
assign n_34295 = n_33213 ^ n_34288;
assign n_34296 = n_34282 ^ n_34290;
assign n_34297 = ~n_34291 & n_34292;
assign n_34298 = n_34284 ^ n_34293;
assign n_34299 = n_34294 ^ n_33213;
assign n_34300 = ~n_33155 & n_34295;
assign n_34301 = n_34295 ^ n_34227;
assign n_34302 = ~n_34296 & ~n_34289;
assign n_34303 = n_34296 ^ n_32431;
assign n_34304 = n_34297 ^ x287;
assign n_34305 = n_34285 & n_34298;
assign n_34306 = n_34298 ^ n_34285;
assign n_34307 = n_34299 ^ n_33911;
assign n_34308 = n_33924 ^ n_34299;
assign n_34309 = n_34300 ^ n_33871;
assign n_34310 = n_34302 ^ n_32431;
assign n_34311 = n_34303 ^ x286;
assign n_34312 = n_34304 ^ n_34303;
assign n_34313 = n_33924 & ~n_34307;
assign n_34314 = ~n_33194 & n_34308;
assign n_34315 = n_34308 ^ n_34247;
assign n_34316 = n_34309 ^ n_32457;
assign n_34317 = n_34309 ^ n_34310;
assign n_34318 = ~n_34312 & n_34311;
assign n_34319 = n_34312 ^ x286;
assign n_34320 = n_34313 ^ n_33255;
assign n_34321 = n_34314 ^ n_33911;
assign n_34322 = n_34316 ^ n_34310;
assign n_34323 = n_34316 & n_34317;
assign n_34324 = n_34318 ^ x286;
assign n_34325 = n_34305 & ~n_34319;
assign n_34326 = n_34319 ^ n_34305;
assign n_34327 = n_34320 ^ n_33282;
assign n_34328 = n_34320 ^ n_33953;
assign n_34329 = n_34321 ^ n_32481;
assign n_34330 = n_34322 ^ x285;
assign n_34331 = n_34323 ^ n_32457;
assign n_34332 = n_34322 ^ n_34324;
assign n_34333 = n_34324 ^ x285;
assign n_34334 = n_34327 ^ n_33953;
assign n_34335 = n_33966 & ~n_34328;
assign n_34336 = n_34321 ^ n_34331;
assign n_34337 = n_34331 ^ n_32481;
assign n_34338 = n_34330 & ~n_34332;
assign n_34339 = n_34322 ^ n_34333;
assign n_34340 = n_33220 & n_34334;
assign n_34341 = n_34268 ^ n_34334;
assign n_34342 = n_34335 ^ n_33282;
assign n_34343 = ~n_34329 & n_34336;
assign n_34344 = n_34321 ^ n_34337;
assign n_34345 = n_34338 ^ x285;
assign n_34346 = n_34325 & ~n_34339;
assign n_34347 = n_34339 ^ n_34325;
assign n_34348 = n_34340 ^ n_33953;
assign n_34349 = n_34342 ^ n_33334;
assign n_34350 = n_34342 ^ n_33994;
assign n_34351 = n_34343 ^ n_32481;
assign n_34352 = n_34344 ^ x284;
assign n_34353 = n_34344 ^ n_34345;
assign n_34354 = ~n_33432 & n_34347;
assign n_34355 = n_34347 ^ n_33432;
assign n_34356 = n_34347 ^ n_33424;
assign n_34357 = n_34348 ^ n_32519;
assign n_34358 = n_34349 ^ n_33994;
assign n_34359 = ~n_34007 & n_34350;
assign n_34360 = n_34348 ^ n_34351;
assign n_34361 = n_34351 ^ n_32519;
assign n_34362 = n_34352 ^ n_34345;
assign n_34363 = n_34352 & ~n_34353;
assign n_34364 = n_34354 ^ n_33462;
assign n_34365 = ~n_32938 & n_34355;
assign n_34366 = n_33271 & ~n_34358;
assign n_34367 = n_34286 ^ n_34358;
assign n_34368 = n_34359 ^ n_33334;
assign n_34369 = n_34357 & n_34360;
assign n_34370 = n_34348 ^ n_34361;
assign n_34371 = n_34346 & ~n_34362;
assign n_34372 = n_34362 ^ n_34346;
assign n_34373 = n_34363 ^ x284;
assign n_34374 = n_34365 ^ n_33432;
assign n_34375 = n_33433 ^ n_34365;
assign n_34376 = n_34366 ^ n_33994;
assign n_34377 = n_34368 ^ n_33371;
assign n_34378 = n_34368 ^ n_34048;
assign n_34379 = n_34369 ^ n_32519;
assign n_34380 = n_34370 ^ x283;
assign n_34381 = n_34372 ^ n_34354;
assign n_34382 = n_34372 ^ n_34364;
assign n_34383 = n_34370 ^ n_34373;
assign n_34384 = ~n_32437 & n_34374;
assign n_34385 = x487 & ~n_34375;
assign n_34386 = n_34375 ^ x487;
assign n_34387 = n_34376 ^ n_32552;
assign n_34388 = n_34377 ^ n_34048;
assign n_34389 = n_34377 & n_34378;
assign n_34390 = n_34379 ^ n_34376;
assign n_34391 = n_34380 ^ n_34373;
assign n_34392 = ~n_34364 & ~n_34381;
assign n_34393 = n_32975 & n_34382;
assign n_34394 = ~n_34380 & n_34383;
assign n_34395 = n_34384 ^ n_32453;
assign n_34396 = n_34385 ^ x486;
assign n_34397 = ~n_33312 & ~n_34388;
assign n_34398 = n_34306 ^ n_34388;
assign n_34399 = n_34089 ^ n_34389;
assign n_34400 = n_34390 ^ n_32552;
assign n_34401 = n_34390 & n_34387;
assign n_34402 = ~n_34371 & ~n_34391;
assign n_34403 = n_34391 ^ n_34371;
assign n_34404 = n_34392 ^ n_33462;
assign n_34405 = n_34393 ^ n_33462;
assign n_34406 = n_34394 ^ x283;
assign n_34407 = n_34397 ^ n_34048;
assign n_34408 = ~n_33326 & ~n_34399;
assign n_34409 = n_34326 ^ n_34399;
assign n_34410 = n_34400 ^ x282;
assign n_34411 = n_34401 ^ n_32552;
assign n_34412 = n_34403 ^ n_33499;
assign n_34413 = n_34404 ^ n_34403;
assign n_34414 = n_34404 ^ n_33499;
assign n_34415 = n_34405 ^ n_34384;
assign n_34416 = n_34405 ^ n_34395;
assign n_34417 = n_34400 ^ n_34406;
assign n_34418 = n_34407 ^ n_32592;
assign n_34419 = n_34408 ^ n_34063;
assign n_34420 = n_34409 ^ n_34388;
assign n_34421 = n_34410 ^ n_34406;
assign n_34422 = n_34407 ^ n_34411;
assign n_34423 = ~n_34412 & n_34413;
assign n_34424 = n_34414 ^ n_34403;
assign n_34425 = n_34395 & ~n_34415;
assign n_34426 = n_34416 ^ n_34385;
assign n_34427 = n_34416 ^ n_34396;
assign n_34428 = n_34410 & ~n_34417;
assign n_34429 = n_34418 ^ n_34411;
assign n_34430 = ~n_34402 & ~n_34421;
assign n_34431 = n_34421 ^ n_34402;
assign n_34432 = n_34418 & ~n_34422;
assign n_34433 = n_34423 ^ n_33499;
assign n_34434 = n_33006 & ~n_34424;
assign n_34435 = n_34425 ^ n_32453;
assign n_34436 = n_34396 & ~n_34426;
assign n_34437 = n_34428 ^ x282;
assign n_34438 = n_34429 ^ x281;
assign n_34439 = n_34431 ^ n_33533;
assign n_34440 = n_34432 ^ n_32592;
assign n_34441 = n_34433 ^ n_34431;
assign n_34442 = n_34434 ^ n_33499;
assign n_34443 = n_34435 ^ n_32498;
assign n_34444 = n_34436 ^ x486;
assign n_34445 = n_34437 ^ n_34429;
assign n_34446 = n_34440 ^ n_32618;
assign n_34447 = ~n_34441 & ~n_34439;
assign n_34448 = n_34441 ^ n_33533;
assign n_34449 = n_34442 ^ n_32498;
assign n_34450 = n_34435 ^ n_34442;
assign n_34451 = n_34443 ^ n_34442;
assign n_34452 = n_34445 & ~n_34438;
assign n_34453 = n_34445 ^ x281;
assign n_34454 = n_34446 ^ n_34419;
assign n_34455 = n_34447 ^ n_33533;
assign n_34456 = n_33042 & ~n_34448;
assign n_34457 = ~n_34449 & ~n_34450;
assign n_34458 = n_34444 ^ n_34451;
assign n_34459 = n_34451 ^ x485;
assign n_34460 = n_34452 ^ x281;
assign n_34461 = n_34430 & n_34453;
assign n_34462 = n_34453 ^ n_34430;
assign n_34463 = n_34454 ^ x280;
assign n_34464 = n_34456 ^ n_33533;
assign n_34465 = n_34457 ^ n_32498;
assign n_34466 = n_34458 ^ x485;
assign n_34467 = n_34458 & ~n_34459;
assign n_34468 = n_34455 ^ n_34462;
assign n_34469 = n_34462 ^ n_33573;
assign n_34470 = n_34460 ^ n_34463;
assign n_34471 = n_34464 ^ n_32537;
assign n_34472 = n_34465 ^ n_34464;
assign n_34473 = n_34467 ^ x485;
assign n_34474 = n_34468 ^ n_33573;
assign n_34475 = n_34468 & n_34469;
assign n_34476 = n_34470 ^ n_34461;
assign n_34477 = ~n_34472 & n_34471;
assign n_34478 = n_34472 ^ n_32537;
assign n_34479 = n_33079 & ~n_34474;
assign n_34480 = n_34475 ^ n_33573;
assign n_34481 = n_34476 ^ n_33608;
assign n_34482 = n_34477 ^ n_32537;
assign n_34483 = n_34478 ^ x484;
assign n_34484 = n_34473 ^ n_34478;
assign n_34485 = n_34479 ^ n_33573;
assign n_34486 = n_34480 ^ n_34476;
assign n_34487 = n_34480 ^ n_34481;
assign n_34488 = n_34473 ^ n_34483;
assign n_34489 = ~n_34483 & n_34484;
assign n_34490 = n_34482 ^ n_34485;
assign n_34491 = n_34485 ^ n_32569;
assign n_34492 = ~n_34481 & n_34486;
assign n_34493 = ~n_33126 & ~n_34487;
assign n_34494 = n_34489 ^ x484;
assign n_34495 = n_34490 ^ n_32569;
assign n_34496 = n_34490 & n_34491;
assign n_34497 = n_34492 ^ n_33608;
assign n_34498 = n_34493 ^ n_33608;
assign n_34499 = n_34494 ^ x483;
assign n_34500 = n_34495 ^ x483;
assign n_34501 = n_34494 ^ n_34495;
assign n_34502 = n_34496 ^ n_32569;
assign n_34503 = n_34497 ^ n_33646;
assign n_34504 = n_34497 ^ n_33660;
assign n_34505 = n_34498 ^ n_32603;
assign n_34506 = n_34499 ^ n_34495;
assign n_34507 = ~n_34500 & n_34501;
assign n_34508 = n_34502 ^ n_34498;
assign n_34509 = ~n_33660 & n_34503;
assign n_34510 = n_33163 & ~n_34504;
assign n_34511 = n_34502 ^ n_34505;
assign n_34512 = n_34507 ^ x483;
assign n_34513 = n_34505 & ~n_34508;
assign n_34514 = n_34509 ^ n_33460;
assign n_34515 = n_34510 ^ n_33646;
assign n_34516 = n_34511 ^ x482;
assign n_34517 = n_34512 ^ n_34511;
assign n_34518 = n_34513 ^ n_32603;
assign n_34519 = n_34514 ^ n_33688;
assign n_34520 = n_34515 ^ n_32642;
assign n_34521 = n_34512 ^ n_34516;
assign n_34522 = n_34516 & ~n_34517;
assign n_34523 = n_34518 ^ n_34515;
assign n_34524 = ~n_34519 & n_33702;
assign n_34525 = n_33525 ^ n_34519;
assign n_34526 = n_34522 ^ x482;
assign n_34527 = n_34523 & ~n_34520;
assign n_34528 = n_34523 ^ n_32642;
assign n_34529 = n_34524 ^ n_33525;
assign n_34530 = n_33188 & n_34525;
assign n_34531 = n_34527 ^ n_32642;
assign n_34532 = n_34528 ^ x481;
assign n_34533 = n_34526 ^ n_34528;
assign n_34534 = n_34529 ^ n_33726;
assign n_34535 = n_34529 ^ n_33741;
assign n_34536 = n_34530 ^ n_33688;
assign n_34537 = n_34526 ^ n_34532;
assign n_34538 = ~n_34532 & n_34533;
assign n_34539 = n_33741 & ~n_34534;
assign n_34540 = ~n_33240 & n_34535;
assign n_34541 = n_34536 ^ n_32685;
assign n_34542 = n_34531 ^ n_34536;
assign n_34543 = ~n_34521 & n_34537;
assign n_34544 = n_34537 ^ n_34521;
assign n_34545 = n_34538 ^ x481;
assign n_34546 = n_34539 ^ n_33570;
assign n_34547 = n_34540 ^ n_33726;
assign n_34548 = n_34531 ^ n_34541;
assign n_34549 = ~n_34541 & ~n_34542;
assign n_34550 = n_34546 ^ n_33767;
assign n_34551 = n_34546 ^ n_33782;
assign n_34552 = n_34547 ^ n_32709;
assign n_34553 = n_34548 ^ x480;
assign n_34554 = n_34545 ^ n_34548;
assign n_34555 = n_34549 ^ n_32685;
assign n_34556 = n_33782 & n_34550;
assign n_34557 = ~n_33278 & n_34551;
assign n_34558 = n_34545 ^ n_34553;
assign n_34559 = ~n_34553 & n_34554;
assign n_34560 = n_34547 ^ n_34555;
assign n_34561 = n_34556 ^ n_33617;
assign n_34562 = n_34557 ^ n_33767;
assign n_34563 = n_34543 & n_34558;
assign n_34564 = n_34558 ^ n_34543;
assign n_34565 = n_34559 ^ x480;
assign n_34566 = n_34560 & ~n_34552;
assign n_34567 = n_34560 ^ n_32709;
assign n_34568 = n_34561 ^ n_33809;
assign n_34569 = n_34562 ^ n_32729;
assign n_34570 = n_34566 ^ n_32709;
assign n_34571 = n_34567 ^ x495;
assign n_34572 = n_34565 ^ n_34567;
assign n_34573 = n_34568 & ~n_33823;
assign n_34574 = n_33655 ^ n_34568;
assign n_34575 = n_34562 ^ n_34570;
assign n_34576 = n_34565 ^ n_34571;
assign n_34577 = n_34571 & ~n_34572;
assign n_34578 = n_34573 ^ n_33655;
assign n_34579 = n_33319 & n_34574;
assign n_34580 = n_34386 ^ n_34574;
assign n_34581 = ~n_34575 & ~n_34569;
assign n_34582 = n_34575 ^ n_32729;
assign n_34583 = ~n_34563 & n_34576;
assign n_34584 = n_34576 ^ n_34563;
assign n_34585 = n_34577 ^ x495;
assign n_34586 = n_34578 ^ n_33849;
assign n_34587 = n_34578 ^ n_33863;
assign n_34588 = n_34579 ^ n_33809;
assign n_34589 = n_34581 ^ n_32729;
assign n_34590 = n_34582 ^ x494;
assign n_34591 = n_34585 ^ n_34582;
assign n_34592 = n_33863 & ~n_34586;
assign n_34593 = n_33356 & ~n_34587;
assign n_34594 = n_34427 ^ n_34587;
assign n_34595 = n_34588 ^ n_32741;
assign n_34596 = n_34589 ^ n_34588;
assign n_34597 = ~n_34591 & n_34590;
assign n_34598 = n_34591 ^ x494;
assign n_34599 = n_34592 ^ n_33697;
assign n_34600 = n_34593 ^ n_33849;
assign n_34601 = n_34589 ^ n_34595;
assign n_34602 = ~n_34595 & ~n_34596;
assign n_34603 = n_34597 ^ x494;
assign n_34604 = ~n_34583 & ~n_34598;
assign n_34605 = n_34598 ^ n_34583;
assign n_34606 = n_34599 ^ n_33889;
assign n_34607 = n_34599 ^ n_33902;
assign n_34608 = n_34600 ^ n_32762;
assign n_34609 = n_34601 ^ x493;
assign n_34610 = n_34602 ^ n_32741;
assign n_34611 = n_34603 ^ n_34601;
assign n_34612 = ~n_33902 & ~n_34606;
assign n_34613 = ~n_33387 & n_34607;
assign n_34614 = n_34466 ^ n_34607;
assign n_34615 = n_34610 ^ n_34600;
assign n_34616 = n_34610 ^ n_32762;
assign n_34617 = n_34611 & ~n_34609;
assign n_34618 = n_34611 ^ x493;
assign n_34619 = n_34612 ^ n_33736;
assign n_34620 = n_34613 ^ n_33889;
assign n_34621 = n_34608 & ~n_34615;
assign n_34622 = n_34616 ^ n_34600;
assign n_34623 = n_34617 ^ x493;
assign n_34624 = n_34604 & n_34618;
assign n_34625 = n_34618 ^ n_34604;
assign n_34626 = n_34619 ^ n_33935;
assign n_34627 = n_34619 ^ n_33777;
assign n_34628 = n_34620 ^ n_32780;
assign n_34629 = n_34621 ^ n_32762;
assign n_34630 = n_34622 ^ x492;
assign n_34631 = n_34623 ^ n_34622;
assign n_34632 = n_34623 ^ x492;
assign n_34633 = n_33949 & n_34626;
assign n_34634 = n_34627 ^ n_33935;
assign n_34635 = n_34629 ^ n_34620;
assign n_34636 = n_34629 ^ n_34628;
assign n_34637 = ~n_34630 & n_34631;
assign n_34638 = n_34632 ^ n_34622;
assign n_34639 = n_34633 ^ n_33777;
assign n_34640 = n_33415 & n_34634;
assign n_34641 = n_34488 ^ n_34634;
assign n_34642 = ~n_34628 & ~n_34635;
assign n_34643 = n_34636 ^ x491;
assign n_34644 = n_34637 ^ x492;
assign n_34645 = ~n_34624 & ~n_34638;
assign n_34646 = n_34638 ^ n_34624;
assign n_34647 = n_34639 ^ n_33974;
assign n_34648 = n_34639 ^ n_33988;
assign n_34649 = n_34640 ^ n_33935;
assign n_34650 = n_34642 ^ n_32780;
assign n_34651 = n_34644 ^ n_34636;
assign n_34652 = n_34644 ^ x491;
assign n_34653 = n_33988 & ~n_34647;
assign n_34654 = ~n_33438 & ~n_34648;
assign n_34655 = n_34506 ^ n_34648;
assign n_34656 = n_34649 ^ n_32805;
assign n_34657 = n_34650 ^ n_34649;
assign n_34658 = n_34643 & ~n_34651;
assign n_34659 = n_34652 ^ n_34636;
assign n_34660 = n_34653 ^ n_33818;
assign n_34661 = n_34654 ^ n_33974;
assign n_34662 = n_34650 ^ n_34656;
assign n_34663 = ~n_34656 & n_34657;
assign n_34664 = n_34658 ^ x491;
assign n_34665 = n_34645 & n_34659;
assign n_34666 = n_34659 ^ n_34645;
assign n_34667 = n_34660 ^ n_34019;
assign n_34668 = n_34660 ^ n_34032;
assign n_34669 = n_34661 ^ n_32817;
assign n_34670 = n_34662 ^ x490;
assign n_34671 = n_34663 ^ n_32805;
assign n_34672 = n_34664 ^ n_34662;
assign n_34673 = ~n_34032 & ~n_34667;
assign n_34674 = ~n_33466 & n_34668;
assign n_34675 = n_34521 ^ n_34668;
assign n_34676 = n_34664 ^ n_34670;
assign n_34677 = n_34661 ^ n_34671;
assign n_34678 = ~n_34670 & n_34672;
assign n_34679 = n_34673 ^ n_33858;
assign n_34680 = n_34674 ^ n_34019;
assign n_34681 = ~n_34665 & n_34676;
assign n_34682 = n_34676 ^ n_34665;
assign n_34683 = n_34677 & n_34669;
assign n_34684 = n_34677 ^ n_32817;
assign n_34685 = n_34678 ^ x490;
assign n_34686 = n_34679 ^ n_34046;
assign n_34687 = n_34679 ^ n_33898;
assign n_34688 = n_34680 ^ n_32841;
assign n_34689 = n_34683 ^ n_32817;
assign n_34690 = n_34684 ^ x489;
assign n_34691 = n_34685 ^ n_34684;
assign n_34692 = n_34685 ^ x489;
assign n_34693 = n_34058 & ~n_34686;
assign n_34694 = n_34687 ^ n_34046;
assign n_34695 = n_34689 ^ n_34680;
assign n_34696 = n_34690 & ~n_34691;
assign n_34697 = n_34692 ^ n_34684;
assign n_34698 = n_34693 ^ n_33898;
assign n_34699 = ~n_33486 & n_34694;
assign n_34700 = n_34544 ^ n_34694;
assign n_34701 = ~n_34695 & ~n_34688;
assign n_34702 = n_34695 ^ n_32841;
assign n_34703 = n_34696 ^ x489;
assign n_34704 = n_34681 & ~n_34697;
assign n_34705 = n_34697 ^ n_34681;
assign n_34706 = n_34698 ^ n_34094;
assign n_34707 = n_34698 ^ n_33939;
assign n_34708 = n_34699 ^ n_34046;
assign n_34709 = n_34701 ^ n_32841;
assign n_34710 = n_34702 ^ x488;
assign n_34711 = n_34703 ^ n_34702;
assign n_34712 = n_34703 ^ x488;
assign n_34713 = n_34104 & ~n_34706;
assign n_34714 = n_34707 ^ n_34094;
assign n_34715 = n_34708 ^ n_32855;
assign n_34716 = n_34709 ^ n_34708;
assign n_34717 = n_34710 & ~n_34711;
assign n_34718 = n_34712 ^ n_34702;
assign n_34719 = n_34713 ^ n_33939;
assign n_34720 = ~n_33532 & n_34714;
assign n_34721 = n_34564 ^ n_34714;
assign n_34722 = n_34709 ^ n_34715;
assign n_34723 = n_34715 & ~n_34716;
assign n_34724 = n_34717 ^ x488;
assign n_34725 = n_34704 & ~n_34718;
assign n_34726 = n_34718 ^ n_34704;
assign n_34727 = n_34719 ^ n_34118;
assign n_34728 = n_34720 ^ n_34094;
assign n_34729 = n_34722 ^ x503;
assign n_34730 = n_34723 ^ n_32855;
assign n_34731 = n_34724 ^ n_34722;
assign n_34732 = ~n_34727 & n_34128;
assign n_34733 = n_33981 ^ n_34727;
assign n_34734 = n_34728 ^ n_32880;
assign n_34735 = n_34724 ^ n_34729;
assign n_34736 = n_34730 ^ n_34728;
assign n_34737 = n_34730 ^ n_32880;
assign n_34738 = n_34729 & ~n_34731;
assign n_34739 = n_34732 ^ n_33981;
assign n_34740 = ~n_33554 & n_34733;
assign n_34741 = n_34584 ^ n_34733;
assign n_34742 = n_34735 & ~n_34725;
assign n_34743 = n_34725 ^ n_34735;
assign n_34744 = ~n_34734 & ~n_34736;
assign n_34745 = n_34737 ^ n_34728;
assign n_34746 = n_34738 ^ x503;
assign n_34747 = n_34739 ^ n_34150;
assign n_34748 = n_34740 ^ n_34118;
assign n_34749 = n_34744 ^ n_32880;
assign n_34750 = n_34745 ^ x502;
assign n_34751 = n_34746 ^ n_34745;
assign n_34752 = n_34747 & n_34158;
assign n_34753 = n_34028 ^ n_34747;
assign n_34754 = n_34748 ^ n_32894;
assign n_34755 = n_34749 ^ n_34748;
assign n_34756 = n_34749 ^ n_32894;
assign n_34757 = n_34751 & ~n_34750;
assign n_34758 = n_34751 ^ x502;
assign n_34759 = n_34752 ^ n_34028;
assign n_34760 = ~n_33591 & n_34753;
assign n_34761 = n_34605 ^ n_34753;
assign n_34762 = ~n_34754 & n_34755;
assign n_34763 = n_34756 ^ n_34748;
assign n_34764 = n_34757 ^ x502;
assign n_34765 = n_34742 & ~n_34758;
assign n_34766 = n_34758 ^ n_34742;
assign n_34767 = n_34759 ^ n_34070;
assign n_34768 = n_34759 ^ n_34174;
assign n_34769 = n_34760 ^ n_34150;
assign n_34770 = n_34762 ^ n_32894;
assign n_34771 = n_34763 ^ x501;
assign n_34772 = n_34764 ^ n_34763;
assign n_34773 = n_34767 ^ n_34174;
assign n_34774 = ~n_34181 & n_34768;
assign n_34775 = n_34769 ^ n_32918;
assign n_34776 = n_34770 ^ n_34769;
assign n_34777 = n_34764 ^ n_34771;
assign n_34778 = n_34771 & ~n_34772;
assign n_34779 = n_33640 & n_34773;
assign n_34780 = n_34625 ^ n_34773;
assign n_34781 = n_34774 ^ n_34070;
assign n_34782 = ~n_34776 & ~n_34775;
assign n_34783 = n_34776 ^ n_32918;
assign n_34784 = ~n_34765 & ~n_34777;
assign n_34785 = n_34777 ^ n_34765;
assign n_34786 = n_34778 ^ x501;
assign n_34787 = n_34779 ^ n_34174;
assign n_34788 = n_34781 ^ n_34108;
assign n_34789 = n_34781 ^ n_34195;
assign n_34790 = n_34782 ^ n_32918;
assign n_34791 = n_34783 ^ x500;
assign n_34792 = n_34786 ^ n_34783;
assign n_34793 = n_34786 ^ x500;
assign n_34794 = n_34787 ^ n_32943;
assign n_34795 = n_34788 ^ n_34195;
assign n_34796 = ~n_34202 & n_34789;
assign n_34797 = n_34790 ^ n_34787;
assign n_34798 = n_34790 ^ n_32943;
assign n_34799 = n_34791 & ~n_34792;
assign n_34800 = n_34793 ^ n_34783;
assign n_34801 = n_33668 & n_34795;
assign n_34802 = n_34646 ^ n_34795;
assign n_34803 = n_34796 ^ n_34108;
assign n_34804 = n_34794 & ~n_34797;
assign n_34805 = n_34798 ^ n_34787;
assign n_34806 = n_34799 ^ x500;
assign n_34807 = n_34784 & ~n_34800;
assign n_34808 = n_34800 ^ n_34784;
assign n_34809 = n_34801 ^ n_34195;
assign n_34810 = n_34803 ^ n_34216;
assign n_34811 = n_34803 ^ n_34209;
assign n_34812 = n_34804 ^ n_32943;
assign n_34813 = n_34805 ^ x499;
assign n_34814 = n_34806 ^ n_34805;
assign n_34815 = n_34809 ^ n_32970;
assign n_34816 = ~n_33720 & ~n_34810;
assign n_34817 = n_34666 ^ n_34810;
assign n_34818 = n_34216 & ~n_34811;
assign n_34819 = n_34812 ^ n_34809;
assign n_34820 = n_34806 ^ n_34813;
assign n_34821 = n_34813 & ~n_34814;
assign n_34822 = n_34812 ^ n_34815;
assign n_34823 = n_34816 ^ n_34209;
assign n_34824 = n_34818 ^ n_34140;
assign n_34825 = n_34815 & ~n_34819;
assign n_34826 = ~n_34807 & n_34820;
assign n_34827 = n_34820 ^ n_34807;
assign n_34828 = n_34821 ^ x499;
assign n_34829 = n_34822 ^ x498;
assign n_34830 = n_34823 ^ n_32990;
assign n_34831 = n_34824 ^ n_34230;
assign n_34832 = n_34825 ^ n_32970;
assign n_34833 = n_34828 ^ n_34822;
assign n_34834 = n_34828 ^ n_34829;
assign n_34835 = n_34164 ^ n_34831;
assign n_34836 = ~n_34831 & n_34237;
assign n_34837 = n_34832 ^ n_34823;
assign n_34838 = n_34829 & ~n_34833;
assign n_34839 = ~n_34826 & ~n_34834;
assign n_34840 = n_34834 ^ n_34826;
assign n_34841 = n_33762 & ~n_34835;
assign n_34842 = n_34682 ^ n_34835;
assign n_34843 = n_34836 ^ n_34164;
assign n_34844 = n_34837 ^ n_32990;
assign n_34845 = n_34837 & n_34830;
assign n_34846 = n_34838 ^ x498;
assign n_34847 = n_34841 ^ n_34230;
assign n_34848 = n_34843 ^ n_34250;
assign n_34849 = n_34843 ^ n_34257;
assign n_34850 = n_34844 ^ x497;
assign n_34851 = n_34845 ^ n_32990;
assign n_34852 = n_34846 ^ n_34844;
assign n_34853 = n_34847 ^ n_33023;
assign n_34854 = n_34257 & n_34848;
assign n_34855 = ~n_33790 & ~n_34849;
assign n_34856 = n_34705 ^ n_34849;
assign n_34857 = n_34851 ^ n_34847;
assign n_34858 = ~n_34852 & n_34850;
assign n_34859 = n_34852 ^ x497;
assign n_34860 = n_34851 ^ n_34853;
assign n_34861 = n_34854 ^ n_34186;
assign n_34862 = n_34855 ^ n_34250;
assign n_34863 = n_34853 & ~n_34857;
assign n_34864 = n_34858 ^ x497;
assign n_34865 = ~n_34839 & n_34859;
assign n_34866 = n_34859 ^ n_34839;
assign n_34867 = n_34860 ^ x496;
assign n_34868 = n_34861 ^ n_34270;
assign n_34869 = n_34861 ^ n_34277;
assign n_34870 = n_34862 ^ n_33061;
assign n_34871 = n_34863 ^ n_33023;
assign n_34872 = n_34864 ^ n_34860;
assign n_34873 = ~n_34355 & ~n_34866;
assign n_34874 = n_34866 ^ n_34355;
assign n_34875 = n_34866 ^ n_34347;
assign n_34876 = n_34277 & n_34868;
assign n_34877 = n_33830 & n_34869;
assign n_34878 = n_34726 ^ n_34869;
assign n_34879 = n_34871 ^ n_34862;
assign n_34880 = n_34871 ^ n_33061;
assign n_34881 = n_34872 ^ x496;
assign n_34882 = n_34872 & ~n_34867;
assign n_34883 = n_34873 ^ n_34382;
assign n_34884 = ~n_33432 & ~n_34874;
assign n_34885 = n_34876 ^ n_34207;
assign n_34886 = n_34877 ^ n_34270;
assign n_34887 = n_34870 & n_34879;
assign n_34888 = n_34880 ^ n_34862;
assign n_34889 = n_34881 ^ n_34865;
assign n_34890 = n_34865 & ~n_34881;
assign n_34891 = n_34882 ^ x496;
assign n_34892 = n_34884 ^ n_34355;
assign n_34893 = n_34356 ^ n_34884;
assign n_34894 = n_34885 ^ n_34295;
assign n_34895 = n_34885 ^ n_34227;
assign n_34896 = n_34886 ^ n_33101;
assign n_34897 = n_34887 ^ n_33061;
assign n_34898 = n_34888 ^ x511;
assign n_34899 = n_34889 ^ n_34883;
assign n_34900 = n_34889 ^ n_34873;
assign n_34901 = n_34891 ^ n_34888;
assign n_34902 = n_34891 ^ x511;
assign n_34903 = ~n_32938 & n_34892;
assign n_34904 = x199 & ~n_34893;
assign n_34905 = n_34893 ^ x199;
assign n_34906 = n_34301 & n_34894;
assign n_34907 = n_34895 ^ n_34295;
assign n_34908 = n_34897 ^ n_34886;
assign n_34909 = n_34897 ^ n_33101;
assign n_34910 = ~n_33462 & ~n_34899;
assign n_34911 = ~n_34883 & n_34900;
assign n_34912 = ~n_34898 & n_34901;
assign n_34913 = n_34902 ^ n_34888;
assign n_34914 = n_34903 ^ n_32975;
assign n_34915 = n_34904 ^ x198;
assign n_34916 = n_34906 ^ n_34227;
assign n_34917 = n_33871 & ~n_34907;
assign n_34918 = n_34743 ^ n_34907;
assign n_34919 = n_34896 & n_34908;
assign n_34920 = n_34909 ^ n_34886;
assign n_34921 = n_34910 ^ n_34382;
assign n_34922 = n_34911 ^ n_34382;
assign n_34923 = n_34912 ^ x511;
assign n_34924 = n_34890 & ~n_34913;
assign n_34925 = n_34913 ^ n_34890;
assign n_34926 = n_34916 ^ n_34308;
assign n_34927 = n_34916 ^ n_34247;
assign n_34928 = n_34917 ^ n_34295;
assign n_34929 = n_34919 ^ n_33101;
assign n_34930 = n_34920 ^ x510;
assign n_34931 = n_34921 ^ n_34903;
assign n_34932 = n_34921 ^ n_34914;
assign n_34933 = n_34923 ^ n_34920;
assign n_34934 = n_34925 ^ n_34424;
assign n_34935 = n_34922 ^ n_34925;
assign n_34936 = ~n_34315 & ~n_34926;
assign n_34937 = n_34927 ^ n_34308;
assign n_34938 = n_34928 ^ n_33155;
assign n_34939 = n_34929 ^ n_34928;
assign n_34940 = n_34929 ^ n_33155;
assign n_34941 = n_34923 ^ n_34930;
assign n_34942 = n_34914 & ~n_34931;
assign n_34943 = n_34932 ^ n_34904;
assign n_34944 = n_34932 ^ n_34915;
assign n_34945 = n_34930 & ~n_34933;
assign n_34946 = n_34922 ^ n_34934;
assign n_34947 = ~n_34934 & ~n_34935;
assign n_34948 = n_34936 ^ n_34247;
assign n_34949 = ~n_33911 & ~n_34937;
assign n_34950 = n_34766 ^ n_34937;
assign n_34951 = ~n_34938 & n_34939;
assign n_34952 = n_34940 ^ n_34928;
assign n_34953 = ~n_34924 & ~n_34941;
assign n_34954 = n_34941 ^ n_34924;
assign n_34955 = n_34942 ^ n_32975;
assign n_34956 = n_34915 & ~n_34943;
assign n_34957 = n_34945 ^ x510;
assign n_34958 = ~n_33499 & ~n_34946;
assign n_34959 = n_34947 ^ n_34424;
assign n_34960 = n_34948 ^ n_34334;
assign n_34961 = n_34341 ^ n_34948;
assign n_34962 = n_34949 ^ n_34308;
assign n_34963 = n_34951 ^ n_33155;
assign n_34964 = n_34952 ^ x509;
assign n_34965 = n_34954 ^ n_34448;
assign n_34966 = n_34956 ^ x198;
assign n_34967 = n_34957 ^ n_34952;
assign n_34968 = n_34958 ^ n_34424;
assign n_34969 = n_34959 ^ n_34954;
assign n_34970 = n_34341 & n_34960;
assign n_34971 = ~n_33953 & ~n_34961;
assign n_34972 = n_34785 ^ n_34961;
assign n_34973 = n_34962 ^ n_33194;
assign n_34974 = n_34963 ^ n_34962;
assign n_34975 = n_34963 ^ n_33194;
assign n_34976 = n_34959 ^ n_34965;
assign n_34977 = ~n_34967 & n_34964;
assign n_34978 = n_34967 ^ x509;
assign n_34979 = n_34968 ^ n_33006;
assign n_34980 = n_34955 ^ n_34968;
assign n_34981 = ~n_34965 & n_34969;
assign n_34982 = n_34970 ^ n_34268;
assign n_34983 = n_34971 ^ n_34334;
assign n_34984 = ~n_34973 & n_34974;
assign n_34985 = n_34975 ^ n_34962;
assign n_34986 = n_33533 & n_34976;
assign n_34987 = n_34977 ^ x509;
assign n_34988 = n_34953 & ~n_34978;
assign n_34989 = n_34978 ^ n_34953;
assign n_34990 = n_34955 ^ n_34979;
assign n_34991 = ~n_34979 & n_34980;
assign n_34992 = n_34981 ^ n_34448;
assign n_34993 = n_34982 ^ n_34286;
assign n_34994 = n_34982 ^ n_34358;
assign n_34995 = n_34983 ^ n_33220;
assign n_34996 = n_34984 ^ n_33194;
assign n_34997 = n_34985 ^ x508;
assign n_34998 = n_34986 ^ n_34448;
assign n_34999 = n_34987 ^ n_34985;
assign n_35000 = n_34987 ^ x508;
assign n_35001 = n_34989 ^ n_34474;
assign n_35002 = n_34966 ^ n_34990;
assign n_35003 = n_34990 ^ x197;
assign n_35004 = n_34991 ^ n_33006;
assign n_35005 = n_34992 ^ n_34989;
assign n_35006 = n_34992 ^ n_34474;
assign n_35007 = n_34993 ^ n_34358;
assign n_35008 = ~n_34367 & n_34994;
assign n_35009 = n_34996 ^ n_34983;
assign n_35010 = n_34998 ^ n_33042;
assign n_35011 = n_34997 & ~n_34999;
assign n_35012 = n_35000 ^ n_34985;
assign n_35013 = n_35002 ^ x197;
assign n_35014 = n_35002 & ~n_35003;
assign n_35015 = n_35004 ^ n_34998;
assign n_35016 = n_35001 & ~n_35005;
assign n_35017 = n_35006 ^ n_34989;
assign n_35018 = n_33994 & ~n_35007;
assign n_35019 = n_34808 ^ n_35007;
assign n_35020 = n_35008 ^ n_34286;
assign n_35021 = n_35009 & n_34995;
assign n_35022 = n_35009 ^ n_33220;
assign n_35023 = n_35004 ^ n_35010;
assign n_35024 = n_35011 ^ x508;
assign n_35025 = n_34988 & ~n_35012;
assign n_35026 = n_35012 ^ n_34988;
assign n_35027 = n_35014 ^ x197;
assign n_35028 = ~n_35010 & n_35015;
assign n_35029 = n_35016 ^ n_34474;
assign n_35030 = ~n_33573 & ~n_35017;
assign n_35031 = n_35018 ^ n_34358;
assign n_35032 = n_34398 ^ n_35020;
assign n_35033 = n_35020 ^ n_34388;
assign n_35034 = n_34306 ^ n_35020;
assign n_35035 = n_35021 ^ n_33220;
assign n_35036 = n_35022 ^ x507;
assign n_35037 = n_35023 ^ x196;
assign n_35038 = n_35024 ^ n_35022;
assign n_35039 = n_35024 ^ x507;
assign n_35040 = n_35026 ^ n_34487;
assign n_35041 = n_35027 ^ n_35023;
assign n_35042 = n_35027 ^ x196;
assign n_35043 = n_35028 ^ n_33042;
assign n_35044 = n_35029 ^ n_35026;
assign n_35045 = n_35030 ^ n_34474;
assign n_35046 = n_35031 ^ n_33271;
assign n_35047 = n_34048 & ~n_35032;
assign n_35048 = ~n_35033 & ~n_35034;
assign n_35049 = n_35031 ^ n_35035;
assign n_35050 = ~n_35036 & n_35038;
assign n_35051 = n_35039 ^ n_35022;
assign n_35052 = n_35029 ^ n_35040;
assign n_35053 = ~n_35037 & n_35041;
assign n_35054 = n_35042 ^ n_35023;
assign n_35055 = n_35043 ^ n_33079;
assign n_35056 = n_35040 & ~n_35044;
assign n_35057 = n_35045 ^ n_33079;
assign n_35058 = n_35043 ^ n_35045;
assign n_35059 = n_35046 ^ n_35035;
assign n_35060 = n_35047 ^ n_34388;
assign n_35061 = n_34420 ^ n_35048;
assign n_35062 = ~n_35046 & n_35049;
assign n_35063 = n_35050 ^ x507;
assign n_35064 = n_35051 & n_35025;
assign n_35065 = n_35025 ^ n_35051;
assign n_35066 = ~n_33608 & ~n_35052;
assign n_35067 = n_35053 ^ x196;
assign n_35068 = ~n_35013 & ~n_35054;
assign n_35069 = n_35054 ^ n_35013;
assign n_35070 = n_35055 ^ n_35045;
assign n_35071 = n_35056 ^ n_34487;
assign n_35072 = ~n_35057 & n_35058;
assign n_35073 = n_35059 ^ x506;
assign n_35074 = n_35060 ^ n_33312;
assign n_35075 = n_34063 & ~n_35061;
assign n_35076 = n_34840 ^ n_35061;
assign n_35077 = n_35062 ^ n_33271;
assign n_35078 = n_35063 ^ n_35059;
assign n_35079 = n_35065 ^ n_34504;
assign n_35080 = n_35066 ^ n_34487;
assign n_35081 = n_35070 ^ x195;
assign n_35082 = n_35067 ^ n_35070;
assign n_35083 = n_35071 ^ n_35065;
assign n_35084 = n_35072 ^ n_33079;
assign n_35085 = n_35063 ^ n_35073;
assign n_35086 = n_35075 ^ n_34399;
assign n_35087 = n_35076 ^ n_34827;
assign n_35088 = n_35077 ^ n_35060;
assign n_35089 = ~n_35073 & n_35078;
assign n_35090 = n_35080 ^ n_33126;
assign n_35091 = n_35067 ^ n_35081;
assign n_35092 = ~n_35081 & n_35082;
assign n_35093 = n_35083 & ~n_35079;
assign n_35094 = n_35083 ^ n_34504;
assign n_35095 = n_35084 ^ n_35080;
assign n_35096 = n_35085 & n_35064;
assign n_35097 = n_35064 ^ n_35085;
assign n_35098 = n_35088 ^ n_33312;
assign n_35099 = n_35088 & n_35074;
assign n_35100 = n_35089 ^ x506;
assign n_35101 = n_35084 ^ n_35090;
assign n_35102 = ~n_35068 & n_35091;
assign n_35103 = n_35091 ^ n_35068;
assign n_35104 = n_35092 ^ x195;
assign n_35105 = n_35093 ^ n_34504;
assign n_35106 = n_33646 & n_35094;
assign n_35107 = n_35090 & n_35095;
assign n_35108 = n_35097 ^ n_34525;
assign n_35109 = n_35098 ^ x505;
assign n_35110 = n_35099 ^ n_33312;
assign n_35111 = n_35098 ^ n_35100;
assign n_35112 = n_35101 ^ x194;
assign n_35113 = n_35104 ^ n_35101;
assign n_35114 = n_35105 ^ n_35097;
assign n_35115 = n_35106 ^ n_34504;
assign n_35116 = n_35107 ^ n_33126;
assign n_35117 = n_35105 ^ n_35108;
assign n_35118 = n_35109 ^ n_35100;
assign n_35119 = n_35110 ^ n_33326;
assign n_35120 = n_35109 & ~n_35111;
assign n_35121 = n_35104 ^ n_35112;
assign n_35122 = n_35112 & ~n_35113;
assign n_35123 = n_35108 & n_35114;
assign n_35124 = n_35115 ^ n_33163;
assign n_35125 = n_35116 ^ n_35115;
assign n_35126 = ~n_33688 & ~n_35117;
assign n_35127 = n_35096 & ~n_35118;
assign n_35128 = n_35118 ^ n_35096;
assign n_35129 = n_35119 ^ n_35086;
assign n_35130 = n_35120 ^ x505;
assign n_35131 = ~n_35102 & n_35121;
assign n_35132 = n_35121 ^ n_35102;
assign n_35133 = n_35122 ^ x194;
assign n_35134 = n_35123 ^ n_34525;
assign n_35135 = ~n_35125 & ~n_35124;
assign n_35136 = n_35125 ^ n_33163;
assign n_35137 = n_35126 ^ n_34525;
assign n_35138 = n_35128 ^ n_34535;
assign n_35139 = n_35129 ^ x504;
assign n_35140 = n_35134 ^ n_35128;
assign n_35141 = n_35135 ^ n_33163;
assign n_35142 = n_35136 ^ x193;
assign n_35143 = n_35133 ^ n_35136;
assign n_35144 = n_35137 ^ n_33188;
assign n_35145 = n_35130 ^ n_35139;
assign n_35146 = n_35140 & ~n_35138;
assign n_35147 = n_35140 ^ n_34535;
assign n_35148 = n_35141 ^ n_35137;
assign n_35149 = n_35133 ^ n_35142;
assign n_35150 = n_35142 & ~n_35143;
assign n_35151 = n_35141 ^ n_35144;
assign n_35152 = n_35145 ^ n_35127;
assign n_35153 = n_35146 ^ n_34535;
assign n_35154 = ~n_33726 & ~n_35147;
assign n_35155 = n_35144 & ~n_35148;
assign n_35156 = n_35131 & n_35149;
assign n_35157 = n_35149 ^ n_35131;
assign n_35158 = n_35150 ^ x193;
assign n_35159 = n_35151 ^ x192;
assign n_35160 = n_35152 ^ n_34551;
assign n_35161 = n_35153 ^ n_35152;
assign n_35162 = n_35154 ^ n_34535;
assign n_35163 = n_35155 ^ n_33188;
assign n_35164 = n_35158 ^ n_35151;
assign n_35165 = n_35158 ^ x192;
assign n_35166 = n_35153 ^ n_35160;
assign n_35167 = n_35160 & ~n_35161;
assign n_35168 = n_35162 ^ n_33240;
assign n_35169 = n_35163 ^ n_35162;
assign n_35170 = n_35159 & ~n_35164;
assign n_35171 = n_35165 ^ n_35151;
assign n_35172 = n_33767 & n_35166;
assign n_35173 = n_35167 ^ n_34551;
assign n_35174 = n_35163 ^ n_35168;
assign n_35175 = ~n_35168 & ~n_35169;
assign n_35176 = n_35170 ^ x192;
assign n_35177 = n_35156 & n_35171;
assign n_35178 = n_35171 ^ n_35156;
assign n_35179 = n_35172 ^ n_34551;
assign n_35180 = n_35173 ^ n_34574;
assign n_35181 = n_35173 ^ n_34580;
assign n_35182 = n_35174 ^ x207;
assign n_35183 = n_35175 ^ n_33240;
assign n_35184 = n_35176 ^ n_35174;
assign n_35185 = n_35179 ^ n_33278;
assign n_35186 = n_34580 & ~n_35180;
assign n_35187 = ~n_33809 & n_35181;
assign n_35188 = n_35176 ^ n_35182;
assign n_35189 = n_35183 ^ n_35179;
assign n_35190 = ~n_35182 & n_35184;
assign n_35191 = n_35186 ^ n_34386;
assign n_35192 = n_35187 ^ n_34574;
assign n_35193 = ~n_35177 & n_35188;
assign n_35194 = n_35188 ^ n_35177;
assign n_35195 = n_35189 & ~n_35185;
assign n_35196 = n_35189 ^ n_33278;
assign n_35197 = n_35190 ^ x207;
assign n_35198 = n_35191 ^ n_34587;
assign n_35199 = n_35191 ^ n_34594;
assign n_35200 = n_35192 ^ n_33319;
assign n_35201 = n_35195 ^ n_33278;
assign n_35202 = n_35196 ^ x206;
assign n_35203 = n_35197 ^ n_35196;
assign n_35204 = n_34594 & n_35198;
assign n_35205 = n_33849 & n_35199;
assign n_35206 = n_35201 ^ n_35192;
assign n_35207 = n_35201 ^ n_33319;
assign n_35208 = ~n_35203 & n_35202;
assign n_35209 = n_35203 ^ x206;
assign n_35210 = n_35204 ^ n_34427;
assign n_35211 = n_35205 ^ n_34587;
assign n_35212 = n_35200 & n_35206;
assign n_35213 = n_35207 ^ n_35192;
assign n_35214 = n_35208 ^ x206;
assign n_35215 = n_35193 & ~n_35209;
assign n_35216 = n_35209 ^ n_35193;
assign n_35217 = n_35210 ^ n_34607;
assign n_35218 = n_35211 ^ n_33356;
assign n_35219 = n_35212 ^ n_33319;
assign n_35220 = n_35213 ^ x205;
assign n_35221 = n_35214 ^ n_35213;
assign n_35222 = n_35217 & n_34614;
assign n_35223 = n_34466 ^ n_35217;
assign n_35224 = n_35219 ^ n_35211;
assign n_35225 = n_35219 ^ n_35218;
assign n_35226 = n_35214 ^ n_35220;
assign n_35227 = ~n_35220 & n_35221;
assign n_35228 = n_35222 ^ n_34466;
assign n_35229 = n_33889 & ~n_35223;
assign n_35230 = ~n_35218 & n_35224;
assign n_35231 = n_35225 ^ x204;
assign n_35232 = ~n_35215 & ~n_35226;
assign n_35233 = n_35226 ^ n_35215;
assign n_35234 = n_35227 ^ x205;
assign n_35235 = n_35228 ^ n_34634;
assign n_35236 = n_35228 ^ n_34488;
assign n_35237 = n_35229 ^ n_34607;
assign n_35238 = n_35230 ^ n_33356;
assign n_35239 = n_35234 ^ n_35225;
assign n_35240 = n_35234 ^ x204;
assign n_35241 = n_34641 & ~n_35235;
assign n_35242 = n_35236 ^ n_34634;
assign n_35243 = n_35237 ^ n_33387;
assign n_35244 = n_35238 ^ n_35237;
assign n_35245 = n_35238 ^ n_33387;
assign n_35246 = ~n_35231 & n_35239;
assign n_35247 = n_35240 ^ n_35225;
assign n_35248 = n_35241 ^ n_34488;
assign n_35249 = n_33935 & n_35242;
assign n_35250 = ~n_35243 & ~n_35244;
assign n_35251 = n_35245 ^ n_35237;
assign n_35252 = n_35246 ^ x204;
assign n_35253 = n_35232 & ~n_35247;
assign n_35254 = n_35247 ^ n_35232;
assign n_35255 = n_35248 ^ n_34648;
assign n_35256 = n_35248 ^ n_34655;
assign n_35257 = n_35249 ^ n_34634;
assign n_35258 = n_35250 ^ n_33387;
assign n_35259 = n_35251 ^ x203;
assign n_35260 = n_35252 ^ n_35251;
assign n_35261 = n_35252 ^ x203;
assign n_35262 = ~n_34655 & n_35255;
assign n_35263 = n_33974 & ~n_35256;
assign n_35264 = n_35257 ^ n_33415;
assign n_35265 = n_35258 ^ n_35257;
assign n_35266 = ~n_35259 & n_35260;
assign n_35267 = n_35261 ^ n_35251;
assign n_35268 = n_35262 ^ n_34506;
assign n_35269 = n_35263 ^ n_34648;
assign n_35270 = n_35258 ^ n_35264;
assign n_35271 = n_35264 & n_35265;
assign n_35272 = n_35266 ^ x203;
assign n_35273 = n_35253 & ~n_35267;
assign n_35274 = n_35267 ^ n_35253;
assign n_35275 = n_35268 ^ n_34668;
assign n_35276 = n_35268 ^ n_34675;
assign n_35277 = n_35269 ^ n_33438;
assign n_35278 = n_35270 ^ x202;
assign n_35279 = n_35271 ^ n_33415;
assign n_35280 = n_35272 ^ n_35270;
assign n_35281 = n_35272 ^ x202;
assign n_35282 = n_34675 & ~n_35275;
assign n_35283 = n_34019 & n_35276;
assign n_35284 = n_35276 ^ n_34905;
assign n_35285 = n_35279 ^ n_35269;
assign n_35286 = n_35279 ^ n_35277;
assign n_35287 = ~n_35278 & n_35280;
assign n_35288 = n_35281 ^ n_35270;
assign n_35289 = n_35282 ^ n_34521;
assign n_35290 = n_35283 ^ n_34668;
assign n_35291 = n_35277 & n_35285;
assign n_35292 = n_35286 ^ x201;
assign n_35293 = n_35287 ^ x202;
assign n_35294 = n_35273 & ~n_35288;
assign n_35295 = n_35288 ^ n_35273;
assign n_35296 = n_35289 ^ n_34694;
assign n_35297 = n_35289 ^ n_34700;
assign n_35298 = n_35290 ^ n_33466;
assign n_35299 = n_35291 ^ n_33438;
assign n_35300 = n_35293 ^ n_35286;
assign n_35301 = n_35293 ^ x201;
assign n_35302 = ~n_34700 & ~n_35296;
assign n_35303 = ~n_34046 & ~n_35297;
assign n_35304 = n_35297 ^ n_34944;
assign n_35305 = n_35299 ^ n_35290;
assign n_35306 = n_35299 ^ n_35298;
assign n_35307 = n_35292 & ~n_35300;
assign n_35308 = n_35301 ^ n_35286;
assign n_35309 = n_35302 ^ n_34544;
assign n_35310 = n_35303 ^ n_34694;
assign n_35311 = ~n_35298 & n_35305;
assign n_35312 = n_35306 ^ x200;
assign n_35313 = n_35307 ^ x201;
assign n_35314 = ~n_35294 & ~n_35308;
assign n_35315 = n_35308 ^ n_35294;
assign n_35316 = n_35309 ^ n_34714;
assign n_35317 = n_35309 ^ n_34721;
assign n_35318 = n_35310 ^ n_33486;
assign n_35319 = n_35311 ^ n_33466;
assign n_35320 = n_35313 ^ n_35306;
assign n_35321 = n_34721 & n_35316;
assign n_35322 = ~n_34094 & ~n_35317;
assign n_35323 = n_35013 ^ n_35317;
assign n_35324 = n_35319 ^ n_35310;
assign n_35325 = n_35319 ^ n_33486;
assign n_35326 = ~n_35320 & n_35312;
assign n_35327 = n_35320 ^ x200;
assign n_35328 = n_35321 ^ n_34564;
assign n_35329 = n_35322 ^ n_34714;
assign n_35330 = ~n_35318 & n_35324;
assign n_35331 = n_35325 ^ n_35310;
assign n_35332 = n_35326 ^ x200;
assign n_35333 = ~n_35314 & n_35327;
assign n_35334 = n_35327 ^ n_35314;
assign n_35335 = n_35328 ^ n_34733;
assign n_35336 = n_35329 ^ n_33532;
assign n_35337 = n_35330 ^ n_33486;
assign n_35338 = n_35331 ^ x215;
assign n_35339 = n_35332 ^ n_35331;
assign n_35340 = ~n_35335 & n_34741;
assign n_35341 = n_34584 ^ n_35335;
assign n_35342 = n_35337 ^ n_35329;
assign n_35343 = n_35337 ^ n_35336;
assign n_35344 = ~n_35339 & n_35338;
assign n_35345 = n_35339 ^ x215;
assign n_35346 = n_35340 ^ n_34584;
assign n_35347 = ~n_34118 & n_35341;
assign n_35348 = n_35069 ^ n_35341;
assign n_35349 = ~n_35336 & n_35342;
assign n_35350 = n_35343 ^ x214;
assign n_35351 = n_35344 ^ x215;
assign n_35352 = ~n_35333 & ~n_35345;
assign n_35353 = n_35345 ^ n_35333;
assign n_35354 = n_35346 ^ n_34753;
assign n_35355 = n_35346 ^ n_34761;
assign n_35356 = n_35347 ^ n_34733;
assign n_35357 = n_35349 ^ n_33532;
assign n_35358 = n_35351 ^ n_35343;
assign n_35359 = n_35351 ^ n_35350;
assign n_35360 = n_34761 & ~n_35354;
assign n_35361 = n_34150 & n_35355;
assign n_35362 = n_35103 ^ n_35355;
assign n_35363 = n_35356 ^ n_33554;
assign n_35364 = n_35357 ^ n_35356;
assign n_35365 = n_35357 ^ n_33554;
assign n_35366 = n_35350 & ~n_35358;
assign n_35367 = ~n_35352 & n_35359;
assign n_35368 = n_35359 ^ n_35352;
assign n_35369 = n_35360 ^ n_34605;
assign n_35370 = n_35361 ^ n_34753;
assign n_35371 = ~n_35363 & n_35364;
assign n_35372 = n_35365 ^ n_35356;
assign n_35373 = n_35366 ^ x214;
assign n_35374 = n_34874 & ~n_35368;
assign n_35375 = n_35368 ^ n_34874;
assign n_35376 = n_35369 ^ n_34773;
assign n_35377 = n_35370 ^ n_33591;
assign n_35378 = n_35371 ^ n_33554;
assign n_35379 = n_35372 ^ x213;
assign n_35380 = n_35373 ^ n_35372;
assign n_35381 = n_35373 ^ x213;
assign n_35382 = n_35374 ^ n_34899;
assign n_35383 = ~n_34355 & n_35375;
assign n_35384 = ~n_35376 & n_34780;
assign n_35385 = n_34625 ^ n_35376;
assign n_35386 = n_35378 ^ n_35370;
assign n_35387 = n_35378 ^ n_35377;
assign n_35388 = n_35379 & ~n_35380;
assign n_35389 = n_35381 ^ n_35372;
assign n_35390 = n_35383 ^ n_34874;
assign n_35391 = n_34875 ^ n_35383;
assign n_35392 = n_35384 ^ n_34625;
assign n_35393 = ~n_34174 & n_35385;
assign n_35394 = n_35132 ^ n_35385;
assign n_35395 = ~n_35377 & n_35386;
assign n_35396 = n_35387 ^ x212;
assign n_35397 = n_35388 ^ x213;
assign n_35398 = n_35367 & n_35389;
assign n_35399 = n_35389 ^ n_35367;
assign n_35400 = ~n_33432 & ~n_35390;
assign n_35401 = x423 & n_35391;
assign n_35402 = n_35391 ^ x423;
assign n_35403 = n_35392 ^ n_34795;
assign n_35404 = n_35392 ^ n_34802;
assign n_35405 = n_35393 ^ n_34773;
assign n_35406 = n_35395 ^ n_33591;
assign n_35407 = n_35397 ^ n_35387;
assign n_35408 = n_35399 ^ n_35374;
assign n_35409 = n_35399 ^ n_35382;
assign n_35410 = n_35400 ^ n_33462;
assign n_35411 = n_35401 ^ x422;
assign n_35412 = ~n_34802 & ~n_35403;
assign n_35413 = ~n_34195 & ~n_35404;
assign n_35414 = n_35157 ^ n_35404;
assign n_35415 = n_35405 ^ n_33640;
assign n_35416 = n_35406 ^ n_35405;
assign n_35417 = ~n_35407 & n_35396;
assign n_35418 = n_35407 ^ x212;
assign n_35419 = n_35382 & ~n_35408;
assign n_35420 = ~n_34382 & ~n_35409;
assign n_35421 = n_35412 ^ n_34646;
assign n_35422 = n_35413 ^ n_34795;
assign n_35423 = n_35406 ^ n_35415;
assign n_35424 = n_35415 & n_35416;
assign n_35425 = n_35417 ^ x212;
assign n_35426 = n_35418 & n_35398;
assign n_35427 = n_35398 ^ n_35418;
assign n_35428 = n_35419 ^ n_34899;
assign n_35429 = n_35420 ^ n_34899;
assign n_35430 = n_35421 ^ n_34810;
assign n_35431 = n_35422 ^ n_33668;
assign n_35432 = n_35423 ^ x211;
assign n_35433 = n_35424 ^ n_33640;
assign n_35434 = n_35425 ^ n_35423;
assign n_35435 = n_35427 ^ n_34946;
assign n_35436 = n_35428 ^ n_35427;
assign n_35437 = n_35429 ^ n_35400;
assign n_35438 = ~n_35430 & n_34817;
assign n_35439 = n_34666 ^ n_35430;
assign n_35440 = n_35425 ^ n_35432;
assign n_35441 = n_35433 ^ n_35422;
assign n_35442 = ~n_35432 & n_35434;
assign n_35443 = ~n_35436 & n_35435;
assign n_35444 = n_35436 ^ n_34946;
assign n_35445 = n_35437 & ~n_35410;
assign n_35446 = n_35437 ^ n_33462;
assign n_35447 = n_35438 ^ n_34666;
assign n_35448 = n_34209 & ~n_35439;
assign n_35449 = n_35178 ^ n_35439;
assign n_35450 = ~n_35440 & n_35426;
assign n_35451 = n_35426 ^ n_35440;
assign n_35452 = ~n_35441 & n_35431;
assign n_35453 = n_35441 ^ n_33668;
assign n_35454 = n_35442 ^ x211;
assign n_35455 = n_35443 ^ n_34946;
assign n_35456 = n_34424 & ~n_35444;
assign n_35457 = n_35445 ^ n_33462;
assign n_35458 = n_35446 ^ n_35401;
assign n_35459 = n_35446 ^ n_35411;
assign n_35460 = n_35447 ^ n_34842;
assign n_35461 = n_35447 ^ n_34835;
assign n_35462 = n_35448 ^ n_34810;
assign n_35463 = n_35451 ^ n_34976;
assign n_35464 = n_35452 ^ n_33668;
assign n_35465 = n_35453 ^ x210;
assign n_35466 = n_35454 ^ n_35453;
assign n_35467 = n_35455 ^ n_35451;
assign n_35468 = n_35455 ^ n_34976;
assign n_35469 = n_35456 ^ n_34946;
assign n_35470 = n_35411 & ~n_35458;
assign n_35471 = n_35402 & n_35459;
assign n_35472 = n_35459 ^ n_35402;
assign n_35473 = n_34230 & ~n_35460;
assign n_35474 = n_35194 ^ n_35460;
assign n_35475 = n_34842 & ~n_35461;
assign n_35476 = n_35462 ^ n_33720;
assign n_35477 = n_35464 ^ n_35462;
assign n_35478 = ~n_35466 & n_35465;
assign n_35479 = n_35466 ^ x210;
assign n_35480 = n_35463 & n_35467;
assign n_35481 = n_35468 ^ n_35451;
assign n_35482 = n_35469 ^ n_33499;
assign n_35483 = n_35457 ^ n_35469;
assign n_35484 = n_35470 ^ x422;
assign n_35485 = n_35473 ^ n_34835;
assign n_35486 = n_35475 ^ n_34682;
assign n_35487 = n_35464 ^ n_35476;
assign n_35488 = n_35476 & n_35477;
assign n_35489 = n_35478 ^ x210;
assign n_35490 = n_35450 & n_35479;
assign n_35491 = n_35479 ^ n_35450;
assign n_35492 = n_35480 ^ n_34976;
assign n_35493 = n_34448 & ~n_35481;
assign n_35494 = n_35457 ^ n_35482;
assign n_35495 = n_35482 & ~n_35483;
assign n_35496 = n_35484 ^ x421;
assign n_35497 = n_35485 ^ n_33762;
assign n_35498 = n_35486 ^ n_34849;
assign n_35499 = n_35487 ^ x209;
assign n_35500 = n_35488 ^ n_33720;
assign n_35501 = n_35489 ^ n_35487;
assign n_35502 = n_35491 ^ n_35017;
assign n_35503 = n_35492 ^ n_35491;
assign n_35504 = n_35493 ^ n_34976;
assign n_35505 = n_35484 ^ n_35494;
assign n_35506 = n_35495 ^ n_33499;
assign n_35507 = n_34705 ^ n_35498;
assign n_35508 = ~n_35498 & n_34856;
assign n_35509 = n_35489 ^ n_35499;
assign n_35510 = n_35485 ^ n_35500;
assign n_35511 = n_35499 & ~n_35501;
assign n_35512 = n_35492 ^ n_35502;
assign n_35513 = n_35502 & n_35503;
assign n_35514 = n_35504 ^ n_33533;
assign n_35515 = n_35505 & n_35496;
assign n_35516 = n_35505 ^ x421;
assign n_35517 = n_35506 ^ n_35504;
assign n_35518 = ~n_34250 & ~n_35507;
assign n_35519 = n_35216 ^ n_35507;
assign n_35520 = n_35508 ^ n_34705;
assign n_35521 = n_35509 & n_35490;
assign n_35522 = n_35490 ^ n_35509;
assign n_35523 = ~n_35510 & ~n_35497;
assign n_35524 = n_35510 ^ n_33762;
assign n_35525 = n_35511 ^ x209;
assign n_35526 = n_34474 & n_35512;
assign n_35527 = n_35513 ^ n_35017;
assign n_35528 = n_35506 ^ n_35514;
assign n_35529 = n_35515 ^ x421;
assign n_35530 = n_35471 & ~n_35516;
assign n_35531 = n_35516 ^ n_35471;
assign n_35532 = n_35514 & n_35517;
assign n_35533 = n_35518 ^ n_34849;
assign n_35534 = n_35520 ^ n_34726;
assign n_35535 = n_35520 ^ n_34869;
assign n_35536 = n_35522 ^ n_35052;
assign n_35537 = n_35523 ^ n_33762;
assign n_35538 = n_35524 ^ x208;
assign n_35539 = n_35525 ^ n_35524;
assign n_35540 = n_35526 ^ n_35017;
assign n_35541 = n_35527 ^ n_35522;
assign n_35542 = n_35528 ^ x420;
assign n_35543 = n_35529 ^ n_35528;
assign n_35544 = n_35532 ^ n_33533;
assign n_35545 = n_35533 ^ n_33790;
assign n_35546 = n_35534 ^ n_34869;
assign n_35547 = ~n_34878 & n_35535;
assign n_35548 = n_35527 ^ n_35536;
assign n_35549 = n_35537 ^ n_33790;
assign n_35550 = n_35537 ^ n_35533;
assign n_35551 = n_35525 ^ n_35538;
assign n_35552 = n_35538 & ~n_35539;
assign n_35553 = n_35536 & ~n_35541;
assign n_35554 = n_35529 ^ n_35542;
assign n_35555 = ~n_35542 & n_35543;
assign n_35556 = n_35544 ^ n_33573;
assign n_35557 = n_35540 ^ n_35544;
assign n_35558 = n_34270 & n_35546;
assign n_35559 = n_35233 ^ n_35546;
assign n_35560 = n_35547 ^ n_34726;
assign n_35561 = n_34487 & ~n_35548;
assign n_35562 = n_35549 ^ n_35533;
assign n_35563 = n_35545 & n_35550;
assign n_35564 = n_35551 & n_35521;
assign n_35565 = n_35521 ^ n_35551;
assign n_35566 = n_35552 ^ x208;
assign n_35567 = n_35553 ^ n_35052;
assign n_35568 = n_35530 & ~n_35554;
assign n_35569 = n_35554 ^ n_35530;
assign n_35570 = n_35555 ^ x420;
assign n_35571 = n_35540 ^ n_35556;
assign n_35572 = ~n_35556 & n_35557;
assign n_35573 = n_35558 ^ n_34869;
assign n_35574 = n_35560 ^ n_34918;
assign n_35575 = n_35560 ^ n_34907;
assign n_35576 = n_35561 ^ n_35052;
assign n_35577 = n_35562 ^ x223;
assign n_35578 = n_35563 ^ n_33790;
assign n_35579 = n_35565 ^ n_35094;
assign n_35580 = n_35566 ^ n_35562;
assign n_35581 = n_35566 ^ x223;
assign n_35582 = n_35567 ^ n_35565;
assign n_35583 = n_35570 ^ x419;
assign n_35584 = n_35571 ^ n_35570;
assign n_35585 = n_35572 ^ n_33573;
assign n_35586 = n_35573 ^ n_33830;
assign n_35587 = ~n_34295 & n_35574;
assign n_35588 = n_35254 ^ n_35574;
assign n_35589 = ~n_34918 & ~n_35575;
assign n_35590 = n_35576 ^ n_33608;
assign n_35591 = n_35578 ^ n_33830;
assign n_35592 = n_35578 ^ n_35573;
assign n_35593 = n_35567 ^ n_35579;
assign n_35594 = n_35577 & ~n_35580;
assign n_35595 = n_35581 ^ n_35562;
assign n_35596 = ~n_35579 & ~n_35582;
assign n_35597 = n_35571 ^ n_35583;
assign n_35598 = n_35583 & ~n_35584;
assign n_35599 = n_35585 ^ n_35576;
assign n_35600 = n_35585 ^ n_33608;
assign n_35601 = n_35587 ^ n_34907;
assign n_35602 = n_35589 ^ n_34743;
assign n_35603 = n_35591 ^ n_35573;
assign n_35604 = n_35586 & n_35592;
assign n_35605 = n_34504 & n_35593;
assign n_35606 = n_35594 ^ x223;
assign n_35607 = ~n_35595 & ~n_35564;
assign n_35608 = n_35564 ^ n_35595;
assign n_35609 = n_35596 ^ n_35094;
assign n_35610 = n_35597 & n_35568;
assign n_35611 = n_35568 ^ n_35597;
assign n_35612 = n_35598 ^ x419;
assign n_35613 = n_35590 & ~n_35599;
assign n_35614 = n_35600 ^ n_35576;
assign n_35615 = n_35601 ^ n_33871;
assign n_35616 = n_35602 ^ n_34937;
assign n_35617 = n_35603 ^ x222;
assign n_35618 = n_35604 ^ n_33830;
assign n_35619 = n_35605 ^ n_35094;
assign n_35620 = n_35606 ^ n_35603;
assign n_35621 = n_35608 ^ n_35117;
assign n_35622 = n_35609 ^ n_35608;
assign n_35623 = n_35609 ^ n_35117;
assign n_35624 = n_35613 ^ n_33608;
assign n_35625 = n_35614 ^ x418;
assign n_35626 = n_35612 ^ n_35614;
assign n_35627 = n_34766 ^ n_35616;
assign n_35628 = n_35616 & ~n_34950;
assign n_35629 = n_35606 ^ n_35617;
assign n_35630 = n_35618 ^ n_35615;
assign n_35631 = n_35618 ^ n_35601;
assign n_35632 = n_35619 ^ n_33646;
assign n_35633 = ~n_35617 & n_35620;
assign n_35634 = ~n_35621 & ~n_35622;
assign n_35635 = n_35623 ^ n_35608;
assign n_35636 = n_35624 ^ n_35619;
assign n_35637 = n_35612 ^ n_35625;
assign n_35638 = ~n_35625 & n_35626;
assign n_35639 = ~n_34308 & ~n_35627;
assign n_35640 = n_35274 ^ n_35627;
assign n_35641 = n_35628 ^ n_34766;
assign n_35642 = n_35629 & n_35607;
assign n_35643 = n_35607 ^ n_35629;
assign n_35644 = n_35630 ^ x221;
assign n_35645 = ~n_35615 & n_35631;
assign n_35646 = n_35624 ^ n_35632;
assign n_35647 = n_35633 ^ x222;
assign n_35648 = n_35634 ^ n_35117;
assign n_35649 = ~n_34525 & ~n_35635;
assign n_35650 = n_35632 & n_35636;
assign n_35651 = ~n_35610 & n_35637;
assign n_35652 = n_35637 ^ n_35610;
assign n_35653 = n_35638 ^ x418;
assign n_35654 = n_35639 ^ n_34937;
assign n_35655 = n_35641 ^ n_34972;
assign n_35656 = n_35641 ^ n_34961;
assign n_35657 = n_35643 ^ n_35147;
assign n_35658 = n_35645 ^ n_33871;
assign n_35659 = n_35646 ^ x417;
assign n_35660 = n_35647 ^ x221;
assign n_35661 = n_35647 ^ n_35630;
assign n_35662 = n_35648 ^ n_35643;
assign n_35663 = n_35649 ^ n_35117;
assign n_35664 = n_35650 ^ n_33646;
assign n_35665 = n_35653 ^ n_35646;
assign n_35666 = n_35654 ^ n_33911;
assign n_35667 = ~n_34334 & ~n_35655;
assign n_35668 = n_35295 ^ n_35655;
assign n_35669 = ~n_34972 & n_35656;
assign n_35670 = n_35648 ^ n_35657;
assign n_35671 = n_35658 ^ n_33911;
assign n_35672 = n_35658 ^ n_35654;
assign n_35673 = n_35653 ^ n_35659;
assign n_35674 = n_35660 ^ n_35630;
assign n_35675 = ~n_35644 & n_35661;
assign n_35676 = ~n_35657 & n_35662;
assign n_35677 = n_35663 ^ n_33688;
assign n_35678 = n_35664 ^ n_35663;
assign n_35679 = ~n_35659 & n_35665;
assign n_35680 = n_35667 ^ n_34961;
assign n_35681 = n_35669 ^ n_34785;
assign n_35682 = ~n_34535 & n_35670;
assign n_35683 = n_35671 ^ n_35654;
assign n_35684 = n_35666 & n_35672;
assign n_35685 = ~n_35651 & ~n_35673;
assign n_35686 = n_35673 ^ n_35651;
assign n_35687 = n_35642 ^ n_35674;
assign n_35688 = ~n_35674 & ~n_35642;
assign n_35689 = n_35675 ^ x221;
assign n_35690 = n_35676 ^ n_35147;
assign n_35691 = n_35664 ^ n_35677;
assign n_35692 = n_35677 & n_35678;
assign n_35693 = n_35679 ^ x417;
assign n_35694 = n_35680 ^ n_33953;
assign n_35695 = n_35019 ^ n_35681;
assign n_35696 = n_35681 ^ n_35007;
assign n_35697 = n_35682 ^ n_35147;
assign n_35698 = n_35683 ^ x220;
assign n_35699 = n_35684 ^ n_33911;
assign n_35700 = n_35687 ^ n_35166;
assign n_35701 = n_35689 ^ n_35683;
assign n_35702 = n_35690 ^ n_35687;
assign n_35703 = n_35691 ^ x416;
assign n_35704 = n_35692 ^ n_33688;
assign n_35705 = n_35693 ^ n_35691;
assign n_35706 = n_35693 ^ x416;
assign n_35707 = n_34358 & n_35695;
assign n_35708 = n_35315 ^ n_35695;
assign n_35709 = n_35019 & n_35696;
assign n_35710 = n_35697 ^ n_33726;
assign n_35711 = n_35689 ^ n_35698;
assign n_35712 = n_35680 ^ n_35699;
assign n_35713 = n_35690 ^ n_35700;
assign n_35714 = n_35698 & ~n_35701;
assign n_35715 = ~n_35700 & ~n_35702;
assign n_35716 = n_35704 ^ n_35697;
assign n_35717 = n_35703 & ~n_35705;
assign n_35718 = n_35706 ^ n_35691;
assign n_35719 = n_35707 ^ n_35007;
assign n_35720 = n_35709 ^ n_34808;
assign n_35721 = n_35704 ^ n_35710;
assign n_35722 = n_35711 ^ n_35688;
assign n_35723 = n_35688 & n_35711;
assign n_35724 = n_35712 ^ n_33953;
assign n_35725 = ~n_35712 & n_35694;
assign n_35726 = ~n_34551 & n_35713;
assign n_35727 = n_35714 ^ x220;
assign n_35728 = n_35715 ^ n_35166;
assign n_35729 = n_35710 & ~n_35716;
assign n_35730 = n_35717 ^ x416;
assign n_35731 = ~n_35685 & ~n_35718;
assign n_35732 = n_35718 ^ n_35685;
assign n_35733 = n_35719 ^ n_33994;
assign n_35734 = n_35720 ^ n_34827;
assign n_35735 = n_35720 ^ n_35032;
assign n_35736 = n_35721 ^ x431;
assign n_35737 = n_35722 ^ n_35181;
assign n_35738 = n_35724 ^ x219;
assign n_35739 = n_35725 ^ n_33953;
assign n_35740 = n_35726 ^ n_35166;
assign n_35741 = n_35727 ^ x219;
assign n_35742 = n_35727 ^ n_35724;
assign n_35743 = n_35728 ^ n_35181;
assign n_35744 = n_35728 ^ n_35722;
assign n_35745 = n_35729 ^ n_33726;
assign n_35746 = n_35730 ^ n_35721;
assign n_35747 = n_35730 ^ x431;
assign n_35748 = n_35734 ^ n_35032;
assign n_35749 = ~n_35734 & ~n_35735;
assign n_35750 = n_35739 ^ n_35719;
assign n_35751 = n_35740 ^ n_33767;
assign n_35752 = n_35741 ^ n_35724;
assign n_35753 = ~n_35738 & n_35742;
assign n_35754 = n_35743 ^ n_35722;
assign n_35755 = ~n_35737 & n_35744;
assign n_35756 = n_35745 ^ n_35740;
assign n_35757 = n_35745 ^ n_33767;
assign n_35758 = ~n_35736 & n_35746;
assign n_35759 = n_35747 ^ n_35721;
assign n_35760 = n_34388 & n_35748;
assign n_35761 = n_35087 ^ n_35749;
assign n_35762 = n_35750 ^ n_33994;
assign n_35763 = ~n_35750 & ~n_35733;
assign n_35764 = n_35723 ^ n_35752;
assign n_35765 = ~n_35752 & n_35723;
assign n_35766 = n_35753 ^ x219;
assign n_35767 = ~n_34574 & ~n_35754;
assign n_35768 = n_35755 ^ n_35181;
assign n_35769 = n_35751 & n_35756;
assign n_35770 = n_35757 ^ n_35740;
assign n_35771 = n_35758 ^ x431;
assign n_35772 = n_35731 & n_35759;
assign n_35773 = n_35759 ^ n_35731;
assign n_35774 = n_35760 ^ n_35032;
assign n_35775 = n_34399 & ~n_35761;
assign n_35776 = n_35353 ^ n_35761;
assign n_35777 = n_35762 ^ x218;
assign n_35778 = n_35763 ^ n_33994;
assign n_35779 = n_35764 ^ n_35199;
assign n_35780 = n_35766 ^ x218;
assign n_35781 = n_35762 ^ n_35766;
assign n_35782 = n_35767 ^ n_35181;
assign n_35783 = n_35768 ^ n_35764;
assign n_35784 = n_35769 ^ n_33767;
assign n_35785 = n_35770 ^ x430;
assign n_35786 = n_35771 ^ n_35770;
assign n_35787 = n_35771 ^ x430;
assign n_35788 = n_35774 ^ n_34048;
assign n_35789 = n_35775 ^ n_35061;
assign n_35790 = n_35776 ^ n_35334;
assign n_35791 = n_35777 ^ n_35766;
assign n_35792 = n_35778 ^ n_34048;
assign n_35793 = n_35774 ^ n_35778;
assign n_35794 = n_35768 ^ n_35779;
assign n_35795 = n_35780 & ~n_35781;
assign n_35796 = n_35782 ^ n_33809;
assign n_35797 = n_35779 & ~n_35783;
assign n_35798 = n_35784 ^ n_35782;
assign n_35799 = ~n_35785 & n_35786;
assign n_35800 = n_35787 ^ n_35770;
assign n_35801 = n_35789 ^ n_34063;
assign n_35802 = n_35791 ^ n_35765;
assign n_35803 = ~n_35765 & ~n_35791;
assign n_35804 = n_35774 ^ n_35792;
assign n_35805 = ~n_35788 & n_35793;
assign n_35806 = n_34587 & n_35794;
assign n_35807 = n_35795 ^ x218;
assign n_35808 = n_35784 ^ n_35796;
assign n_35809 = n_35797 ^ n_35199;
assign n_35810 = ~n_35796 & ~n_35798;
assign n_35811 = n_35799 ^ x430;
assign n_35812 = ~n_35772 & ~n_35800;
assign n_35813 = n_35800 ^ n_35772;
assign n_35814 = n_35802 ^ n_35223;
assign n_35815 = n_35804 ^ x217;
assign n_35816 = n_35805 ^ n_34048;
assign n_35817 = n_35806 ^ n_35199;
assign n_35818 = n_35807 ^ n_35804;
assign n_35819 = n_35808 ^ x429;
assign n_35820 = n_35809 ^ n_35802;
assign n_35821 = n_35810 ^ n_33809;
assign n_35822 = n_35811 ^ n_35808;
assign n_35823 = n_35811 ^ x429;
assign n_35824 = n_35809 ^ n_35814;
assign n_35825 = n_35807 ^ n_35815;
assign n_35826 = n_35816 ^ n_35801;
assign n_35827 = n_35817 ^ n_33849;
assign n_35828 = ~n_35815 & n_35818;
assign n_35829 = ~n_35814 & ~n_35820;
assign n_35830 = n_35821 ^ n_35817;
assign n_35831 = ~n_35819 & n_35822;
assign n_35832 = n_35823 ^ n_35808;
assign n_35833 = ~n_34607 & ~n_35824;
assign n_35834 = n_35803 ^ n_35825;
assign n_35835 = ~n_35825 & ~n_35803;
assign n_35836 = n_35821 ^ n_35827;
assign n_35837 = n_35828 ^ x217;
assign n_35838 = n_35829 ^ n_35223;
assign n_35839 = n_35827 & n_35830;
assign n_35840 = n_35831 ^ x429;
assign n_35841 = n_35812 & ~n_35832;
assign n_35842 = n_35833 ^ n_35223;
assign n_35843 = n_35834 ^ n_35242;
assign n_35844 = n_35836 ^ x428;
assign n_35845 = n_35837 ^ x216;
assign n_35846 = n_35838 ^ n_35834;
assign n_35847 = n_35839 ^ n_33849;
assign n_35848 = n_35840 ^ n_35836;
assign n_35849 = n_35842 ^ n_33889;
assign n_35850 = n_35838 ^ n_35843;
assign n_35851 = n_35840 ^ n_35844;
assign n_35852 = n_35845 ^ n_35826;
assign n_35853 = ~n_35843 & ~n_35846;
assign n_35854 = n_35847 ^ n_33889;
assign n_35855 = n_35847 ^ n_35842;
assign n_35856 = ~n_35844 & n_35848;
assign n_35857 = ~n_34634 & n_35850;
assign n_35858 = n_35841 & ~n_35851;
assign n_35859 = n_35851 ^ n_35841;
assign n_35860 = n_35852 ^ n_35835;
assign n_35861 = n_35853 ^ n_35242;
assign n_35862 = n_35854 ^ n_35842;
assign n_35863 = ~n_35849 & n_35855;
assign n_35864 = n_35856 ^ x428;
assign n_35865 = n_35857 ^ n_35242;
assign n_35866 = ~n_35375 & ~n_35859;
assign n_35867 = n_35859 ^ n_35368;
assign n_35868 = n_35860 ^ n_35256;
assign n_35869 = n_35861 ^ n_35256;
assign n_35870 = n_35861 ^ n_35860;
assign n_35871 = n_35862 ^ x427;
assign n_35872 = n_35863 ^ n_33889;
assign n_35873 = n_35864 ^ n_35862;
assign n_35874 = n_35865 ^ n_33935;
assign n_35875 = n_35866 ^ n_35409;
assign n_35876 = n_35867 ^ n_34874;
assign n_35877 = n_35869 ^ n_35860;
assign n_35878 = n_35868 & n_35870;
assign n_35879 = n_35864 ^ n_35871;
assign n_35880 = n_35872 ^ n_35865;
assign n_35881 = n_35872 ^ n_33935;
assign n_35882 = ~n_35871 & n_35873;
assign n_35883 = n_34874 & ~n_35876;
assign n_35884 = n_34648 & n_35877;
assign n_35885 = n_35878 ^ n_35256;
assign n_35886 = n_35879 ^ n_35858;
assign n_35887 = ~n_35858 & n_35879;
assign n_35888 = n_35874 & ~n_35880;
assign n_35889 = n_35881 ^ n_35865;
assign n_35890 = n_35882 ^ x427;
assign n_35891 = n_35883 ^ n_35368;
assign n_35892 = n_35884 ^ n_35256;
assign n_35893 = n_35885 ^ n_35284;
assign n_35894 = n_35885 ^ n_35276;
assign n_35895 = n_35886 ^ n_35875;
assign n_35896 = n_35886 ^ n_35866;
assign n_35897 = n_35888 ^ n_33935;
assign n_35898 = n_35889 ^ x426;
assign n_35899 = n_35890 ^ n_35889;
assign n_35900 = n_35891 ^ n_34874;
assign n_35901 = n_35891 ^ n_34866;
assign n_35902 = n_35892 ^ n_33974;
assign n_35903 = ~n_34668 & ~n_35893;
assign n_35904 = n_35284 & n_35894;
assign n_35905 = n_34899 & ~n_35895;
assign n_35906 = n_35875 & ~n_35896;
assign n_35907 = n_35897 ^ n_35892;
assign n_35908 = n_35890 ^ n_35898;
assign n_35909 = n_35898 & ~n_35899;
assign n_35910 = ~n_34355 & n_35900;
assign n_35911 = x135 & ~n_35901;
assign n_35912 = n_35901 ^ x135;
assign n_35913 = n_35897 ^ n_35902;
assign n_35914 = n_35903 ^ n_35276;
assign n_35915 = n_35904 ^ n_34905;
assign n_35916 = n_35905 ^ n_35409;
assign n_35917 = n_35906 ^ n_35409;
assign n_35918 = ~n_35902 & n_35907;
assign n_35919 = ~n_35887 & n_35908;
assign n_35920 = n_35908 ^ n_35887;
assign n_35921 = n_35909 ^ x426;
assign n_35922 = n_35910 ^ n_34382;
assign n_35923 = n_35911 ^ x134;
assign n_35924 = n_35913 ^ x425;
assign n_35925 = n_35914 ^ n_34019;
assign n_35926 = n_35915 ^ n_35304;
assign n_35927 = n_35915 ^ n_35297;
assign n_35928 = n_35916 ^ n_35910;
assign n_35929 = n_35918 ^ n_33974;
assign n_35930 = n_35920 ^ n_35444;
assign n_35931 = n_35917 ^ n_35920;
assign n_35932 = n_35921 ^ n_35913;
assign n_35933 = n_35921 ^ n_35924;
assign n_35934 = ~n_34694 & n_35926;
assign n_35935 = n_35304 & n_35927;
assign n_35936 = n_35928 ^ n_34382;
assign n_35937 = n_35928 & ~n_35922;
assign n_35938 = n_35929 ^ n_35925;
assign n_35939 = n_35929 ^ n_35914;
assign n_35940 = n_35917 ^ n_35930;
assign n_35941 = ~n_35930 & n_35931;
assign n_35942 = ~n_35924 & n_35932;
assign n_35943 = n_35919 & ~n_35933;
assign n_35944 = n_35933 ^ n_35919;
assign n_35945 = n_35934 ^ n_35297;
assign n_35946 = n_35935 ^ n_34944;
assign n_35947 = n_35936 ^ n_35923;
assign n_35948 = n_35936 ^ n_35911;
assign n_35949 = n_35937 ^ n_34382;
assign n_35950 = n_35938 ^ x424;
assign n_35951 = n_35925 & ~n_35939;
assign n_35952 = n_34946 & n_35940;
assign n_35953 = n_35941 ^ n_35444;
assign n_35954 = n_35942 ^ x425;
assign n_35955 = n_35944 ^ n_35481;
assign n_35956 = n_35945 ^ n_34046;
assign n_35957 = n_35946 ^ n_35323;
assign n_35958 = n_35946 ^ n_35317;
assign n_35959 = n_35923 & ~n_35948;
assign n_35960 = n_35951 ^ n_34019;
assign n_35961 = n_35952 ^ n_35444;
assign n_35962 = n_35953 ^ n_35944;
assign n_35963 = n_35954 ^ n_35938;
assign n_35964 = n_35954 ^ n_35950;
assign n_35965 = n_35953 ^ n_35955;
assign n_35966 = ~n_34714 & ~n_35957;
assign n_35967 = n_35323 & ~n_35958;
assign n_35968 = n_35959 ^ x134;
assign n_35969 = n_35960 ^ n_34046;
assign n_35970 = n_35960 ^ n_35945;
assign n_35971 = n_35961 ^ n_34424;
assign n_35972 = n_35949 ^ n_35961;
assign n_35973 = ~n_35955 & n_35962;
assign n_35974 = n_35950 & ~n_35963;
assign n_35975 = n_35943 & n_35964;
assign n_35976 = n_35964 ^ n_35943;
assign n_35977 = ~n_34976 & n_35965;
assign n_35978 = n_35966 ^ n_35317;
assign n_35979 = n_35967 ^ n_35013;
assign n_35980 = n_35968 ^ x133;
assign n_35981 = n_35969 ^ n_35945;
assign n_35982 = n_35956 & n_35970;
assign n_35983 = n_35949 ^ n_35971;
assign n_35984 = ~n_35971 & ~n_35972;
assign n_35985 = n_35973 ^ n_35481;
assign n_35986 = n_35974 ^ x424;
assign n_35987 = n_35976 ^ n_35512;
assign n_35988 = n_35977 ^ n_35481;
assign n_35989 = n_35978 ^ n_34094;
assign n_35990 = n_35979 ^ n_35341;
assign n_35991 = n_35981 ^ x439;
assign n_35992 = n_35982 ^ n_34046;
assign n_35993 = n_35968 ^ n_35983;
assign n_35994 = n_35984 ^ n_34424;
assign n_35995 = n_35985 ^ n_35976;
assign n_35996 = n_35985 ^ n_35512;
assign n_35997 = n_35986 ^ n_35981;
assign n_35998 = n_35988 ^ n_34448;
assign n_35999 = n_35069 ^ n_35990;
assign n_36000 = n_35990 & ~n_35348;
assign n_36001 = n_35992 ^ n_35978;
assign n_36002 = ~n_35993 & n_35980;
assign n_36003 = n_35993 ^ x133;
assign n_36004 = n_35994 ^ n_35988;
assign n_36005 = ~n_35987 & ~n_35995;
assign n_36006 = n_35996 ^ n_35976;
assign n_36007 = ~n_35997 & n_35991;
assign n_36008 = n_35997 ^ x439;
assign n_36009 = n_35994 ^ n_35998;
assign n_36010 = ~n_34733 & n_35999;
assign n_36011 = n_36000 ^ n_35069;
assign n_36012 = n_36001 ^ n_34094;
assign n_36013 = ~n_36001 & n_35989;
assign n_36014 = n_36002 ^ x133;
assign n_36015 = n_35947 & n_36003;
assign n_36016 = n_36003 ^ n_35947;
assign n_36017 = ~n_35998 & n_36004;
assign n_36018 = n_36005 ^ n_35512;
assign n_36019 = n_35017 & n_36006;
assign n_36020 = n_36007 ^ x439;
assign n_36021 = n_35975 & n_36008;
assign n_36022 = n_36008 ^ n_35975;
assign n_36023 = n_36009 ^ x132;
assign n_36024 = n_36010 ^ n_35341;
assign n_36025 = n_36011 ^ n_35355;
assign n_36026 = n_35362 ^ n_36011;
assign n_36027 = n_36012 ^ x438;
assign n_36028 = n_36013 ^ n_34094;
assign n_36029 = n_36014 ^ n_36009;
assign n_36030 = n_36017 ^ n_34448;
assign n_36031 = n_36018 ^ n_35548;
assign n_36032 = n_36019 ^ n_35512;
assign n_36033 = n_36020 ^ n_36012;
assign n_36034 = n_36018 ^ n_36022;
assign n_36035 = n_36014 ^ n_36023;
assign n_36036 = n_36024 ^ n_34118;
assign n_36037 = ~n_35362 & n_36025;
assign n_36038 = ~n_34753 & n_36026;
assign n_36039 = n_36020 ^ n_36027;
assign n_36040 = n_36028 ^ n_36024;
assign n_36041 = ~n_36023 & n_36029;
assign n_36042 = n_36032 ^ n_36030;
assign n_36043 = n_36032 ^ n_34474;
assign n_36044 = ~n_36027 & n_36033;
assign n_36045 = n_36034 & ~n_36031;
assign n_36046 = n_36034 ^ n_35548;
assign n_36047 = n_36015 & ~n_36035;
assign n_36048 = n_36035 ^ n_36015;
assign n_36049 = n_36028 ^ n_36036;
assign n_36050 = n_36037 ^ n_35103;
assign n_36051 = n_36038 ^ n_35355;
assign n_36052 = n_36039 ^ n_36021;
assign n_36053 = n_36021 & ~n_36039;
assign n_36054 = ~n_36036 & n_36040;
assign n_36055 = n_36041 ^ x132;
assign n_36056 = n_36042 ^ n_34474;
assign n_36057 = ~n_36042 & n_36043;
assign n_36058 = n_36044 ^ x438;
assign n_36059 = n_36045 ^ n_35548;
assign n_36060 = n_35052 & n_36046;
assign n_36061 = n_36049 ^ x437;
assign n_36062 = n_36050 ^ n_35385;
assign n_36063 = n_35394 ^ n_36050;
assign n_36064 = n_36051 ^ n_34150;
assign n_36065 = n_36052 ^ n_35593;
assign n_36066 = n_36054 ^ n_34118;
assign n_36067 = n_36056 ^ x131;
assign n_36068 = n_36055 ^ n_36056;
assign n_36069 = n_36057 ^ n_34474;
assign n_36070 = n_36058 ^ x437;
assign n_36071 = n_36049 ^ n_36058;
assign n_36072 = n_36059 ^ n_36052;
assign n_36073 = n_36059 ^ n_35593;
assign n_36074 = n_36060 ^ n_35548;
assign n_36075 = n_36061 ^ n_36058;
assign n_36076 = n_35394 & n_36062;
assign n_36077 = ~n_34773 & ~n_36063;
assign n_36078 = n_36051 ^ n_36066;
assign n_36079 = n_36064 ^ n_36066;
assign n_36080 = n_36055 ^ n_36067;
assign n_36081 = n_36067 & ~n_36068;
assign n_36082 = n_36070 & ~n_36071;
assign n_36083 = n_36065 & n_36072;
assign n_36084 = n_36073 ^ n_36052;
assign n_36085 = n_36074 ^ n_34487;
assign n_36086 = n_36069 ^ n_36074;
assign n_36087 = n_36053 ^ n_36075;
assign n_36088 = n_36075 & n_36053;
assign n_36089 = n_36076 ^ n_35132;
assign n_36090 = n_36077 ^ n_35385;
assign n_36091 = n_36064 & n_36078;
assign n_36092 = n_36079 ^ x436;
assign n_36093 = n_36047 & n_36080;
assign n_36094 = n_36080 ^ n_36047;
assign n_36095 = n_36081 ^ x131;
assign n_36096 = n_36082 ^ x437;
assign n_36097 = n_36083 ^ n_35593;
assign n_36098 = ~n_35094 & ~n_36084;
assign n_36099 = n_35912 ^ n_36084;
assign n_36100 = n_36069 ^ n_36085;
assign n_36101 = ~n_36085 & n_36086;
assign n_36102 = n_36087 ^ n_35635;
assign n_36103 = n_36089 ^ n_35414;
assign n_36104 = n_36089 ^ n_35404;
assign n_36105 = n_36090 ^ n_34174;
assign n_36106 = n_36091 ^ n_34150;
assign n_36107 = n_36095 ^ x130;
assign n_36108 = n_36079 ^ n_36096;
assign n_36109 = n_36092 ^ n_36096;
assign n_36110 = n_36097 ^ n_35635;
assign n_36111 = n_36097 ^ n_36087;
assign n_36112 = n_36098 ^ n_35593;
assign n_36113 = n_36100 ^ n_36095;
assign n_36114 = n_36100 ^ x130;
assign n_36115 = n_36101 ^ n_34487;
assign n_36116 = n_36103 ^ n_35402;
assign n_36117 = ~n_34795 & n_36103;
assign n_36118 = n_35414 & n_36104;
assign n_36119 = n_36090 ^ n_36106;
assign n_36120 = n_36105 ^ n_36106;
assign n_36121 = ~n_36092 & n_36108;
assign n_36122 = n_36109 & ~n_36088;
assign n_36123 = n_36088 ^ n_36109;
assign n_36124 = n_36110 ^ n_36087;
assign n_36125 = n_36102 & n_36111;
assign n_36126 = n_36112 ^ n_34504;
assign n_36127 = n_36107 & n_36113;
assign n_36128 = n_36114 ^ n_36095;
assign n_36129 = n_36112 ^ n_36115;
assign n_36130 = n_36117 ^ n_35404;
assign n_36131 = n_36118 ^ n_35157;
assign n_36132 = ~n_36105 & ~n_36119;
assign n_36133 = n_36120 ^ x435;
assign n_36134 = n_36121 ^ x436;
assign n_36135 = n_36123 ^ n_35670;
assign n_36136 = n_35947 ^ n_36124;
assign n_36137 = n_35117 & n_36124;
assign n_36138 = n_36125 ^ n_35635;
assign n_36139 = n_36127 ^ x130;
assign n_36140 = n_36093 & ~n_36128;
assign n_36141 = n_36128 ^ n_36093;
assign n_36142 = ~n_36129 & n_36126;
assign n_36143 = n_36129 ^ n_34504;
assign n_36144 = n_36130 ^ n_34195;
assign n_36145 = n_36131 ^ n_35439;
assign n_36146 = n_36132 ^ n_34174;
assign n_36147 = n_36120 ^ n_36134;
assign n_36148 = n_36134 ^ x435;
assign n_36149 = n_36137 ^ n_35635;
assign n_36150 = n_36138 ^ n_36123;
assign n_36151 = n_36142 ^ n_34504;
assign n_36152 = n_36143 ^ x129;
assign n_36153 = n_36139 ^ n_36143;
assign n_36154 = ~n_36145 & n_35449;
assign n_36155 = n_36145 ^ n_35178;
assign n_36156 = n_36130 ^ n_36146;
assign n_36157 = n_36144 ^ n_36146;
assign n_36158 = ~n_36133 & n_36147;
assign n_36159 = n_36120 ^ n_36148;
assign n_36160 = n_36149 ^ n_34525;
assign n_36161 = ~n_36150 & ~n_36135;
assign n_36162 = n_36150 ^ n_35670;
assign n_36163 = n_36151 ^ n_36149;
assign n_36164 = n_36139 ^ n_36152;
assign n_36165 = n_36152 & ~n_36153;
assign n_36166 = n_36154 ^ n_35178;
assign n_36167 = n_34810 & ~n_36155;
assign n_36168 = n_35472 ^ n_36155;
assign n_36169 = n_36144 & ~n_36156;
assign n_36170 = n_36157 ^ x434;
assign n_36171 = n_36158 ^ x435;
assign n_36172 = ~n_36159 & ~n_36122;
assign n_36173 = n_36122 ^ n_36159;
assign n_36174 = n_36161 ^ n_35670;
assign n_36175 = n_35147 & n_36162;
assign n_36176 = n_36016 ^ n_36162;
assign n_36177 = n_36163 & n_36160;
assign n_36178 = n_36163 ^ n_34525;
assign n_36179 = n_36140 & n_36164;
assign n_36180 = n_36164 ^ n_36140;
assign n_36181 = n_36165 ^ x129;
assign n_36182 = n_36166 ^ n_35460;
assign n_36183 = n_35474 ^ n_36166;
assign n_36184 = n_36167 ^ n_35439;
assign n_36185 = n_36169 ^ n_34195;
assign n_36186 = n_36157 ^ n_36171;
assign n_36187 = n_36170 ^ n_36171;
assign n_36188 = n_36173 ^ n_35713;
assign n_36189 = n_36173 ^ n_36174;
assign n_36190 = n_36175 ^ n_35670;
assign n_36191 = n_36177 ^ n_34525;
assign n_36192 = n_36178 ^ x128;
assign n_36193 = n_36181 ^ n_36178;
assign n_36194 = n_35474 & ~n_36182;
assign n_36195 = n_34835 & ~n_36183;
assign n_36196 = n_35531 ^ n_36183;
assign n_36197 = n_36184 ^ n_34209;
assign n_36198 = n_36185 ^ n_36184;
assign n_36199 = ~n_36170 & n_36186;
assign n_36200 = ~n_36187 & n_36172;
assign n_36201 = n_36172 ^ n_36187;
assign n_36202 = n_36188 ^ n_36174;
assign n_36203 = ~n_36188 & n_36189;
assign n_36204 = n_36190 ^ n_34535;
assign n_36205 = n_36190 ^ n_36191;
assign n_36206 = n_36191 ^ n_34535;
assign n_36207 = n_36181 ^ n_36192;
assign n_36208 = n_36192 & ~n_36193;
assign n_36209 = n_36194 ^ n_35194;
assign n_36210 = n_36195 ^ n_35460;
assign n_36211 = ~n_36198 & ~n_36197;
assign n_36212 = n_36198 ^ n_34209;
assign n_36213 = n_36199 ^ x434;
assign n_36214 = n_36201 ^ n_35754;
assign n_36215 = ~n_35166 & ~n_36202;
assign n_36216 = n_36048 ^ n_36202;
assign n_36217 = n_36203 ^ n_35713;
assign n_36218 = ~n_36204 & n_36205;
assign n_36219 = n_36190 ^ n_36206;
assign n_36220 = ~n_36179 & ~n_36207;
assign n_36221 = n_36207 ^ n_36179;
assign n_36222 = n_36208 ^ x128;
assign n_36223 = n_36209 ^ n_35507;
assign n_36224 = n_35519 ^ n_36209;
assign n_36225 = n_36210 ^ n_34230;
assign n_36226 = n_36211 ^ n_34209;
assign n_36227 = n_36212 ^ x433;
assign n_36228 = n_36212 ^ n_36213;
assign n_36229 = n_36215 ^ n_35713;
assign n_36230 = n_36201 ^ n_36217;
assign n_36231 = n_36217 ^ n_35754;
assign n_36232 = n_36218 ^ n_34535;
assign n_36233 = n_36219 ^ x143;
assign n_36234 = n_36219 ^ n_36222;
assign n_36235 = n_36222 ^ x143;
assign n_36236 = n_35519 & ~n_36223;
assign n_36237 = n_34849 & ~n_36224;
assign n_36238 = n_35569 ^ n_36224;
assign n_36239 = n_36210 ^ n_36226;
assign n_36240 = n_36225 ^ n_36226;
assign n_36241 = n_36227 ^ n_36213;
assign n_36242 = n_36227 & ~n_36228;
assign n_36243 = n_36229 ^ n_34551;
assign n_36244 = ~n_36214 & ~n_36230;
assign n_36245 = n_36201 ^ n_36231;
assign n_36246 = n_36232 ^ n_36229;
assign n_36247 = n_36233 & ~n_36234;
assign n_36248 = n_36219 ^ n_36235;
assign n_36249 = n_36236 ^ n_35216;
assign n_36250 = n_36237 ^ n_35507;
assign n_36251 = ~n_36225 & n_36239;
assign n_36252 = n_36240 ^ x432;
assign n_36253 = n_36241 & n_36200;
assign n_36254 = n_36200 ^ n_36241;
assign n_36255 = n_36242 ^ x433;
assign n_36256 = n_36244 ^ n_35754;
assign n_36257 = ~n_35181 & ~n_36245;
assign n_36258 = n_36094 ^ n_36245;
assign n_36259 = n_36246 & ~n_36243;
assign n_36260 = n_36246 ^ n_34551;
assign n_36261 = n_36247 ^ x143;
assign n_36262 = n_36248 & ~n_36220;
assign n_36263 = n_36220 ^ n_36248;
assign n_36264 = n_35559 ^ n_36249;
assign n_36265 = n_36249 ^ n_35546;
assign n_36266 = n_36250 ^ n_34250;
assign n_36267 = n_36251 ^ n_34230;
assign n_36268 = n_36254 ^ n_35794;
assign n_36269 = n_36240 ^ n_36255;
assign n_36270 = n_36255 ^ x432;
assign n_36271 = n_36254 ^ n_36256;
assign n_36272 = n_36256 ^ n_35794;
assign n_36273 = n_36257 ^ n_35754;
assign n_36274 = n_36259 ^ n_34551;
assign n_36275 = n_36260 ^ x142;
assign n_36276 = n_36260 ^ n_36261;
assign n_36277 = n_36261 ^ x142;
assign n_36278 = ~n_34869 & n_36264;
assign n_36279 = n_35611 ^ n_36264;
assign n_36280 = ~n_35559 & n_36265;
assign n_36281 = n_36267 ^ n_36250;
assign n_36282 = ~n_36252 & n_36269;
assign n_36283 = n_36240 ^ n_36270;
assign n_36284 = ~n_36268 & ~n_36271;
assign n_36285 = n_36254 ^ n_36272;
assign n_36286 = n_36273 ^ n_34574;
assign n_36287 = n_36274 ^ n_36273;
assign n_36288 = n_36275 & ~n_36276;
assign n_36289 = n_36260 ^ n_36277;
assign n_36290 = n_36278 ^ n_35546;
assign n_36291 = n_36280 ^ n_35233;
assign n_36292 = n_36281 & n_36266;
assign n_36293 = n_36281 ^ n_34250;
assign n_36294 = n_36282 ^ x432;
assign n_36295 = ~n_36283 & n_36253;
assign n_36296 = n_36253 ^ n_36283;
assign n_36297 = n_36284 ^ n_35794;
assign n_36298 = ~n_35199 & n_36285;
assign n_36299 = n_36141 ^ n_36285;
assign n_36300 = ~n_36287 & n_36286;
assign n_36301 = n_36287 ^ n_34574;
assign n_36302 = n_36288 ^ x142;
assign n_36303 = ~n_36262 & ~n_36289;
assign n_36304 = n_36289 ^ n_36262;
assign n_36305 = n_36290 ^ n_34270;
assign n_36306 = n_36291 ^ n_35254;
assign n_36307 = n_36291 ^ n_35574;
assign n_36308 = n_36292 ^ n_34250;
assign n_36309 = n_36293 ^ x447;
assign n_36310 = n_36294 ^ n_36293;
assign n_36311 = n_36296 ^ n_35824;
assign n_36312 = n_36296 ^ n_36297;
assign n_36313 = n_36298 ^ n_35794;
assign n_36314 = n_36300 ^ n_34574;
assign n_36315 = n_36301 ^ x141;
assign n_36316 = n_36301 ^ n_36302;
assign n_36317 = n_36306 ^ n_35574;
assign n_36318 = n_35588 & n_36307;
assign n_36319 = n_36290 ^ n_36308;
assign n_36320 = n_36305 ^ n_36308;
assign n_36321 = ~n_36310 & n_36309;
assign n_36322 = n_36310 ^ x447;
assign n_36323 = n_36311 ^ n_36297;
assign n_36324 = ~n_36311 & ~n_36312;
assign n_36325 = n_36313 ^ n_34587;
assign n_36326 = n_36313 ^ n_36314;
assign n_36327 = n_36315 ^ n_36302;
assign n_36328 = ~n_36315 & n_36316;
assign n_36329 = n_34907 & ~n_36317;
assign n_36330 = n_35652 ^ n_36317;
assign n_36331 = n_36318 ^ n_35254;
assign n_36332 = n_36305 & n_36319;
assign n_36333 = n_36320 ^ x446;
assign n_36334 = n_36321 ^ x447;
assign n_36335 = n_36322 & n_36295;
assign n_36336 = n_36295 ^ n_36322;
assign n_36337 = n_35223 & ~n_36323;
assign n_36338 = n_36180 ^ n_36323;
assign n_36339 = n_36324 ^ n_35824;
assign n_36340 = n_36325 ^ n_36314;
assign n_36341 = n_36325 & n_36326;
assign n_36342 = n_36303 & n_36327;
assign n_36343 = n_36327 ^ n_36303;
assign n_36344 = n_36328 ^ x141;
assign n_36345 = n_36329 ^ n_35574;
assign n_36346 = n_36331 ^ n_35640;
assign n_36347 = n_36331 ^ n_35627;
assign n_36348 = n_36332 ^ n_34270;
assign n_36349 = n_36320 ^ n_36334;
assign n_36350 = n_36334 ^ x446;
assign n_36351 = n_36336 ^ n_35850;
assign n_36352 = n_36337 ^ n_35824;
assign n_36353 = n_36336 ^ n_36339;
assign n_36354 = n_36339 ^ n_35850;
assign n_36355 = n_36341 ^ n_34587;
assign n_36356 = n_36344 ^ n_36340;
assign n_36357 = n_36344 ^ x140;
assign n_36358 = n_36345 ^ n_34295;
assign n_36359 = n_34937 & ~n_36346;
assign n_36360 = n_35686 ^ n_36346;
assign n_36361 = ~n_35640 & n_36347;
assign n_36362 = n_36348 ^ n_36345;
assign n_36363 = ~n_36333 & n_36349;
assign n_36364 = n_36320 ^ n_36350;
assign n_36365 = n_36352 ^ n_34607;
assign n_36366 = ~n_36351 & ~n_36353;
assign n_36367 = n_36336 ^ n_36354;
assign n_36368 = n_36352 ^ n_36355;
assign n_36369 = n_36355 ^ n_34607;
assign n_36370 = n_36356 ^ x140;
assign n_36371 = n_36356 & n_36357;
assign n_36372 = n_36359 ^ n_35627;
assign n_36373 = n_36361 ^ n_35274;
assign n_36374 = ~n_36362 & ~n_36358;
assign n_36375 = n_36362 ^ n_34295;
assign n_36376 = n_36363 ^ x446;
assign n_36377 = n_36364 & ~n_36335;
assign n_36378 = n_36335 ^ n_36364;
assign n_36379 = n_36366 ^ n_35850;
assign n_36380 = ~n_35242 & n_36367;
assign n_36381 = n_36221 ^ n_36367;
assign n_36382 = n_36365 & n_36368;
assign n_36383 = n_36352 ^ n_36369;
assign n_36384 = n_36342 & n_36370;
assign n_36385 = n_36370 ^ n_36342;
assign n_36386 = n_36371 ^ x140;
assign n_36387 = n_36372 ^ n_34308;
assign n_36388 = n_36373 ^ n_35295;
assign n_36389 = n_36373 ^ n_35655;
assign n_36390 = n_36374 ^ n_34295;
assign n_36391 = n_36375 ^ x445;
assign n_36392 = n_36375 ^ n_36376;
assign n_36393 = n_36376 ^ x445;
assign n_36394 = n_36378 ^ n_35877;
assign n_36395 = n_36378 ^ n_36379;
assign n_36396 = n_36380 ^ n_35850;
assign n_36397 = n_36382 ^ n_34607;
assign n_36398 = n_36383 ^ x139;
assign n_36399 = n_36386 ^ n_36383;
assign n_36400 = n_36388 ^ n_35655;
assign n_36401 = ~n_35668 & n_36389;
assign n_36402 = n_36390 ^ n_36372;
assign n_36403 = ~n_36391 & n_36392;
assign n_36404 = n_36375 ^ n_36393;
assign n_36405 = n_36394 ^ n_36379;
assign n_36406 = ~n_36394 & n_36395;
assign n_36407 = n_36396 ^ n_34634;
assign n_36408 = n_36397 ^ n_36396;
assign n_36409 = ~n_36399 & n_36398;
assign n_36410 = n_36399 ^ x139;
assign n_36411 = n_34961 & ~n_36400;
assign n_36412 = n_35732 ^ n_36400;
assign n_36413 = n_36401 ^ n_35295;
assign n_36414 = ~n_36402 & n_36387;
assign n_36415 = n_36402 ^ n_34308;
assign n_36416 = n_36403 ^ x445;
assign n_36417 = n_36404 & n_36377;
assign n_36418 = n_36377 ^ n_36404;
assign n_36419 = n_35256 & ~n_36405;
assign n_36420 = n_36263 ^ n_36405;
assign n_36421 = n_36406 ^ n_35877;
assign n_36422 = n_36408 & ~n_36407;
assign n_36423 = n_36408 ^ n_34634;
assign n_36424 = n_36409 ^ x139;
assign n_36425 = n_36384 & ~n_36410;
assign n_36426 = n_36410 ^ n_36384;
assign n_36427 = n_36411 ^ n_35655;
assign n_36428 = n_36413 ^ n_35315;
assign n_36429 = n_36413 ^ n_35695;
assign n_36430 = n_36414 ^ n_34308;
assign n_36431 = n_36415 ^ x444;
assign n_36432 = n_36415 ^ n_36416;
assign n_36433 = n_36418 ^ n_35893;
assign n_36434 = n_36419 ^ n_35877;
assign n_36435 = n_36418 ^ n_36421;
assign n_36436 = n_36421 ^ n_35893;
assign n_36437 = n_36422 ^ n_34634;
assign n_36438 = n_36423 ^ x138;
assign n_36439 = n_36424 ^ n_36423;
assign n_36440 = n_36427 ^ n_34334;
assign n_36441 = n_36428 ^ n_35695;
assign n_36442 = n_35708 & ~n_36429;
assign n_36443 = n_36430 ^ n_36427;
assign n_36444 = n_36431 ^ n_36416;
assign n_36445 = ~n_36431 & n_36432;
assign n_36446 = n_36434 ^ n_34648;
assign n_36447 = ~n_36433 & ~n_36435;
assign n_36448 = n_36418 ^ n_36436;
assign n_36449 = n_36434 ^ n_36437;
assign n_36450 = n_36437 ^ n_34648;
assign n_36451 = ~n_36439 & n_36438;
assign n_36452 = n_36439 ^ x138;
assign n_36453 = n_36430 ^ n_36440;
assign n_36454 = n_35007 & n_36441;
assign n_36455 = n_35773 ^ n_36441;
assign n_36456 = n_36442 ^ n_35315;
assign n_36457 = n_36440 & ~n_36443;
assign n_36458 = n_36444 & n_36417;
assign n_36459 = n_36417 ^ n_36444;
assign n_36460 = n_36445 ^ x444;
assign n_36461 = n_36447 ^ n_35893;
assign n_36462 = ~n_35276 & ~n_36448;
assign n_36463 = n_36304 ^ n_36448;
assign n_36464 = n_36446 & n_36449;
assign n_36465 = n_36434 ^ n_36450;
assign n_36466 = n_36451 ^ x138;
assign n_36467 = n_36425 & ~n_36452;
assign n_36468 = n_36452 ^ n_36425;
assign n_36469 = n_36453 ^ x443;
assign n_36470 = n_36454 ^ n_35695;
assign n_36471 = n_36456 ^ n_35748;
assign n_36472 = n_36456 ^ n_35334;
assign n_36473 = n_36457 ^ n_34334;
assign n_36474 = n_36459 ^ n_35926;
assign n_36475 = n_36453 ^ n_36460;
assign n_36476 = n_36461 ^ n_36459;
assign n_36477 = n_36462 ^ n_35893;
assign n_36478 = n_36464 ^ n_34648;
assign n_36479 = n_36465 ^ x137;
assign n_36480 = n_36466 ^ n_36465;
assign n_36481 = n_36469 ^ n_36460;
assign n_36482 = n_36470 ^ n_34358;
assign n_36483 = n_36471 ^ n_35334;
assign n_36484 = ~n_36471 & n_36472;
assign n_36485 = n_36473 ^ n_34358;
assign n_36486 = n_36473 ^ n_36470;
assign n_36487 = ~n_36469 & n_36475;
assign n_36488 = n_36476 & n_36474;
assign n_36489 = n_36476 ^ n_35926;
assign n_36490 = n_36477 ^ n_34668;
assign n_36491 = n_36477 ^ n_36478;
assign n_36492 = n_36478 ^ n_34668;
assign n_36493 = n_36480 & ~n_36479;
assign n_36494 = n_36480 ^ x137;
assign n_36495 = ~n_36481 & ~n_36458;
assign n_36496 = n_36458 ^ n_36481;
assign n_36497 = n_35032 & n_36483;
assign n_36498 = n_35790 ^ n_36484;
assign n_36499 = n_36485 ^ n_36470;
assign n_36500 = n_36482 & n_36486;
assign n_36501 = n_36487 ^ x443;
assign n_36502 = n_36488 ^ n_35926;
assign n_36503 = n_35297 & ~n_36489;
assign n_36504 = n_36343 ^ n_36489;
assign n_36505 = n_36490 & n_36491;
assign n_36506 = n_36477 ^ n_36492;
assign n_36507 = n_36493 ^ x137;
assign n_36508 = n_36467 & n_36494;
assign n_36509 = n_36494 ^ n_36467;
assign n_36510 = n_36496 ^ n_35957;
assign n_36511 = n_36497 ^ n_35748;
assign n_36512 = n_35061 & ~n_36498;
assign n_36513 = n_36498 ^ n_35812;
assign n_36514 = n_36499 ^ x442;
assign n_36515 = n_36500 ^ n_34358;
assign n_36516 = n_36501 ^ n_36499;
assign n_36517 = n_36502 ^ n_36496;
assign n_36518 = n_36503 ^ n_35926;
assign n_36519 = n_36505 ^ n_34668;
assign n_36520 = n_36506 ^ x136;
assign n_36521 = n_36507 ^ n_36506;
assign n_36522 = n_36511 ^ n_34388;
assign n_36523 = n_36512 ^ n_35761;
assign n_36524 = n_36513 ^ n_35832;
assign n_36525 = n_36515 ^ n_36511;
assign n_36526 = n_36516 & ~n_36514;
assign n_36527 = n_36516 ^ x442;
assign n_36528 = n_36517 & n_36510;
assign n_36529 = n_36517 ^ n_35957;
assign n_36530 = n_36518 ^ n_34694;
assign n_36531 = n_36518 ^ n_36519;
assign n_36532 = n_36519 ^ n_34694;
assign n_36533 = ~n_36521 & n_36520;
assign n_36534 = n_36521 ^ x136;
assign n_36535 = n_36524 ^ n_35813;
assign n_36536 = n_36525 ^ n_34388;
assign n_36537 = ~n_36525 & n_36522;
assign n_36538 = n_36526 ^ x442;
assign n_36539 = ~n_36527 & n_36495;
assign n_36540 = n_36495 ^ n_36527;
assign n_36541 = n_36528 ^ n_35957;
assign n_36542 = n_35317 & n_36529;
assign n_36543 = n_36385 ^ n_36529;
assign n_36544 = ~n_36530 & n_36531;
assign n_36545 = n_36518 ^ n_36532;
assign n_36546 = n_36533 ^ x136;
assign n_36547 = ~n_36508 & n_36534;
assign n_36548 = n_36534 ^ n_36508;
assign n_36549 = n_36536 ^ x441;
assign n_36550 = n_36537 ^ n_34388;
assign n_36551 = n_36538 ^ n_36536;
assign n_36552 = n_36540 ^ n_35999;
assign n_36553 = n_36541 ^ n_36540;
assign n_36554 = n_36542 ^ n_35957;
assign n_36555 = n_36544 ^ n_34694;
assign n_36556 = n_36545 ^ x151;
assign n_36557 = n_36545 ^ n_36546;
assign n_36558 = n_36546 ^ x151;
assign n_36559 = n_36550 ^ n_34399;
assign n_36560 = ~n_36551 & n_36549;
assign n_36561 = n_36551 ^ x441;
assign n_36562 = n_36553 & n_36552;
assign n_36563 = n_36553 ^ n_35999;
assign n_36564 = n_36554 ^ n_34714;
assign n_36565 = n_36555 ^ n_36554;
assign n_36566 = n_36556 & ~n_36557;
assign n_36567 = n_36545 ^ n_36558;
assign n_36568 = n_36559 ^ n_36523;
assign n_36569 = n_36560 ^ x441;
assign n_36570 = ~n_36561 & ~n_36539;
assign n_36571 = n_36539 ^ n_36561;
assign n_36572 = n_36562 ^ n_35999;
assign n_36573 = ~n_35341 & ~n_36563;
assign n_36574 = n_36426 ^ n_36563;
assign n_36575 = ~n_36565 & n_36564;
assign n_36576 = n_36565 ^ n_34714;
assign n_36577 = n_36566 ^ x151;
assign n_36578 = ~n_36547 & ~n_36567;
assign n_36579 = n_36567 ^ n_36547;
assign n_36580 = n_36569 ^ n_36568;
assign n_36581 = n_36571 ^ n_36026;
assign n_36582 = n_36571 ^ n_36572;
assign n_36583 = n_36572 ^ n_36026;
assign n_36584 = n_36573 ^ n_35999;
assign n_36585 = n_36575 ^ n_34714;
assign n_36586 = n_36576 ^ x150;
assign n_36587 = n_36577 ^ n_36576;
assign n_36588 = n_36580 ^ x440;
assign n_36589 = n_36581 & ~n_36582;
assign n_36590 = n_36571 ^ n_36583;
assign n_36591 = n_36584 ^ n_34733;
assign n_36592 = n_36584 ^ n_36585;
assign n_36593 = n_36585 ^ n_34733;
assign n_36594 = n_36587 & ~n_36586;
assign n_36595 = n_36587 ^ x150;
assign n_36596 = n_36588 ^ n_36570;
assign n_36597 = n_36589 ^ n_36026;
assign n_36598 = ~n_35355 & n_36590;
assign n_36599 = n_36468 ^ n_36590;
assign n_36600 = ~n_36591 & n_36592;
assign n_36601 = n_36584 ^ n_36593;
assign n_36602 = n_36594 ^ x150;
assign n_36603 = n_36578 & n_36595;
assign n_36604 = n_36595 ^ n_36578;
assign n_36605 = n_36596 ^ n_36063;
assign n_36606 = n_36596 ^ n_36597;
assign n_36607 = n_36597 ^ n_36063;
assign n_36608 = n_36598 ^ n_36026;
assign n_36609 = n_36600 ^ n_34733;
assign n_36610 = n_36601 ^ x149;
assign n_36611 = n_36602 ^ n_36601;
assign n_36612 = n_36605 & n_36606;
assign n_36613 = n_36596 ^ n_36607;
assign n_36614 = n_36608 ^ n_34753;
assign n_36615 = n_36608 ^ n_36609;
assign n_36616 = n_36609 ^ n_34753;
assign n_36617 = ~n_36611 & n_36610;
assign n_36618 = n_36611 ^ x149;
assign n_36619 = n_36612 ^ n_36063;
assign n_36620 = ~n_35385 & n_36613;
assign n_36621 = n_36509 ^ n_36613;
assign n_36622 = ~n_36614 & n_36615;
assign n_36623 = n_36608 ^ n_36616;
assign n_36624 = n_36617 ^ x149;
assign n_36625 = ~n_36603 & n_36618;
assign n_36626 = n_36618 ^ n_36603;
assign n_36627 = n_36619 ^ n_36103;
assign n_36628 = n_36116 ^ n_36619;
assign n_36629 = n_36620 ^ n_36063;
assign n_36630 = n_36622 ^ n_34753;
assign n_36631 = n_36623 ^ x148;
assign n_36632 = n_36624 ^ n_36623;
assign n_36633 = n_36116 & n_36627;
assign n_36634 = n_35404 & ~n_36628;
assign n_36635 = n_36548 ^ n_36628;
assign n_36636 = n_36629 ^ n_34773;
assign n_36637 = n_36629 ^ n_36630;
assign n_36638 = n_36630 ^ n_34773;
assign n_36639 = ~n_36632 & n_36631;
assign n_36640 = n_36632 ^ x148;
assign n_36641 = n_36633 ^ n_35402;
assign n_36642 = n_36634 ^ n_36103;
assign n_36643 = n_36636 & ~n_36637;
assign n_36644 = n_36629 ^ n_36638;
assign n_36645 = n_36639 ^ x148;
assign n_36646 = n_36625 & n_36640;
assign n_36647 = n_36640 ^ n_36625;
assign n_36648 = n_36641 ^ n_36155;
assign n_36649 = n_36643 ^ n_34773;
assign n_36650 = n_36644 ^ x147;
assign n_36651 = n_36645 ^ n_36644;
assign n_36652 = n_36648 & n_36168;
assign n_36653 = n_36648 ^ n_35472;
assign n_36654 = n_36649 ^ n_34795;
assign n_36655 = n_36649 ^ n_36642;
assign n_36656 = n_36651 & ~n_36650;
assign n_36657 = n_36651 ^ x147;
assign n_36658 = n_36652 ^ n_35472;
assign n_36659 = n_35439 & n_36653;
assign n_36660 = n_36579 ^ n_36653;
assign n_36661 = n_36654 ^ n_36642;
assign n_36662 = n_36654 & n_36655;
assign n_36663 = n_36656 ^ x147;
assign n_36664 = ~n_36646 & n_36657;
assign n_36665 = n_36657 ^ n_36646;
assign n_36666 = n_36658 ^ n_36183;
assign n_36667 = n_36659 ^ n_36155;
assign n_36668 = n_36661 ^ x146;
assign n_36669 = n_36662 ^ n_34795;
assign n_36670 = n_36663 ^ n_36661;
assign n_36671 = n_35531 ^ n_36666;
assign n_36672 = ~n_36666 & ~n_36196;
assign n_36673 = n_36667 ^ n_34810;
assign n_36674 = n_36667 ^ n_36669;
assign n_36675 = n_36669 ^ n_34810;
assign n_36676 = ~n_36670 & n_36668;
assign n_36677 = n_36670 ^ x146;
assign n_36678 = n_35460 & n_36671;
assign n_36679 = n_36604 ^ n_36671;
assign n_36680 = n_36672 ^ n_35531;
assign n_36681 = ~n_36673 & ~n_36674;
assign n_36682 = n_36667 ^ n_36675;
assign n_36683 = n_36676 ^ x146;
assign n_36684 = ~n_36664 & n_36677;
assign n_36685 = n_36677 ^ n_36664;
assign n_36686 = n_36678 ^ n_36183;
assign n_36687 = n_36680 ^ n_35569;
assign n_36688 = n_36680 ^ n_36224;
assign n_36689 = n_36681 ^ n_34810;
assign n_36690 = n_36682 ^ x145;
assign n_36691 = n_36683 ^ n_36682;
assign n_36692 = n_36686 ^ n_34835;
assign n_36693 = n_36687 ^ n_36224;
assign n_36694 = ~n_36238 & n_36688;
assign n_36695 = n_36686 ^ n_36689;
assign n_36696 = n_36689 ^ n_34835;
assign n_36697 = ~n_36691 & n_36690;
assign n_36698 = n_36691 ^ x145;
assign n_36699 = n_35507 & ~n_36693;
assign n_36700 = n_36626 ^ n_36693;
assign n_36701 = n_36694 ^ n_35569;
assign n_36702 = ~n_36692 & n_36695;
assign n_36703 = n_36686 ^ n_36696;
assign n_36704 = n_36697 ^ x145;
assign n_36705 = ~n_36684 & ~n_36698;
assign n_36706 = n_36698 ^ n_36684;
assign n_36707 = n_36699 ^ n_36224;
assign n_36708 = n_36701 ^ n_35611;
assign n_36709 = n_36701 ^ n_36264;
assign n_36710 = n_36702 ^ n_34835;
assign n_36711 = n_36703 ^ x144;
assign n_36712 = n_36704 ^ n_36703;
assign n_36713 = n_36707 ^ n_34849;
assign n_36714 = n_36708 ^ n_36264;
assign n_36715 = ~n_36279 & ~n_36709;
assign n_36716 = n_36710 ^ n_34849;
assign n_36717 = n_36710 ^ n_36707;
assign n_36718 = n_36712 & ~n_36711;
assign n_36719 = n_36712 ^ x144;
assign n_36720 = ~n_35546 & ~n_36714;
assign n_36721 = n_36647 ^ n_36714;
assign n_36722 = n_36715 ^ n_35611;
assign n_36723 = n_36716 ^ n_36707;
assign n_36724 = ~n_36713 & n_36717;
assign n_36725 = n_36718 ^ x144;
assign n_36726 = ~n_36705 & ~n_36719;
assign n_36727 = n_36719 ^ n_36705;
assign n_36728 = n_36720 ^ n_36264;
assign n_36729 = n_36722 ^ n_36317;
assign n_36730 = n_36723 ^ x159;
assign n_36731 = n_36724 ^ n_34849;
assign n_36732 = n_36723 ^ n_36725;
assign n_36733 = n_36725 ^ x159;
assign n_36734 = n_36728 ^ n_34869;
assign n_36735 = n_35652 ^ n_36729;
assign n_36736 = ~n_36729 & n_36330;
assign n_36737 = n_36731 ^ n_36728;
assign n_36738 = ~n_36730 & n_36732;
assign n_36739 = n_36723 ^ n_36733;
assign n_36740 = ~n_35574 & ~n_36735;
assign n_36741 = n_36665 ^ n_36735;
assign n_36742 = n_36736 ^ n_35652;
assign n_36743 = n_36737 ^ n_34869;
assign n_36744 = ~n_36737 & ~n_36734;
assign n_36745 = n_36738 ^ x159;
assign n_36746 = ~n_36726 & n_36739;
assign n_36747 = n_36739 ^ n_36726;
assign n_36748 = n_36740 ^ n_36317;
assign n_36749 = n_36742 ^ n_36346;
assign n_36750 = n_36743 ^ x158;
assign n_36751 = n_36744 ^ n_34869;
assign n_36752 = n_36745 ^ n_36743;
assign n_36753 = n_36748 ^ n_34907;
assign n_36754 = n_36749 ^ n_35686;
assign n_36755 = ~n_36749 & n_36360;
assign n_36756 = n_36751 ^ n_34907;
assign n_36757 = n_36751 ^ n_36748;
assign n_36758 = n_36752 & ~n_36750;
assign n_36759 = n_36752 ^ x158;
assign n_36760 = n_35627 & ~n_36754;
assign n_36761 = n_36685 ^ n_36754;
assign n_36762 = n_36755 ^ n_35686;
assign n_36763 = n_36756 ^ n_36748;
assign n_36764 = ~n_36753 & ~n_36757;
assign n_36765 = n_36758 ^ x158;
assign n_36766 = n_36746 & n_36759;
assign n_36767 = n_36759 ^ n_36746;
assign n_36768 = n_36760 ^ n_36346;
assign n_36769 = n_36762 ^ n_36400;
assign n_36770 = n_36763 ^ x157;
assign n_36771 = n_36764 ^ n_34907;
assign n_36772 = n_36765 ^ n_36763;
assign n_36773 = n_36768 ^ n_34937;
assign n_36774 = n_36769 ^ n_35732;
assign n_36775 = ~n_36769 & ~n_36412;
assign n_36776 = n_36771 ^ n_34937;
assign n_36777 = n_36771 ^ n_36768;
assign n_36778 = ~n_36772 & n_36770;
assign n_36779 = n_36772 ^ x157;
assign n_36780 = n_35655 & n_36774;
assign n_36781 = n_36706 ^ n_36774;
assign n_36782 = n_36775 ^ n_35732;
assign n_36783 = n_36776 ^ n_36768;
assign n_36784 = ~n_36773 & n_36777;
assign n_36785 = n_36778 ^ x157;
assign n_36786 = n_36766 & ~n_36779;
assign n_36787 = n_36779 ^ n_36766;
assign n_36788 = n_36780 ^ n_36400;
assign n_36789 = n_36782 ^ n_36441;
assign n_36790 = n_36783 ^ x156;
assign n_36791 = n_36784 ^ n_34937;
assign n_36792 = n_36785 ^ n_36783;
assign n_36793 = n_35876 & n_36787;
assign n_36794 = n_36787 ^ n_35876;
assign n_36795 = n_36787 ^ n_35859;
assign n_36796 = n_36788 ^ n_34961;
assign n_36797 = n_36789 ^ n_35773;
assign n_36798 = ~n_36789 & n_36455;
assign n_36799 = n_36791 ^ n_34961;
assign n_36800 = n_36791 ^ n_36788;
assign n_36801 = n_36792 & ~n_36790;
assign n_36802 = n_36792 ^ x156;
assign n_36803 = n_36793 ^ n_35895;
assign n_36804 = ~n_35375 & ~n_36794;
assign y7 = ~n_36794;
assign n_36805 = ~n_35695 & n_36797;
assign n_36806 = n_36727 ^ n_36797;
assign n_36807 = n_36798 ^ n_35773;
assign n_36808 = n_36799 ^ n_36788;
assign n_36809 = ~n_36796 & n_36800;
assign n_36810 = n_36801 ^ x156;
assign n_36811 = ~n_36786 & ~n_36802;
assign n_36812 = n_36802 ^ n_36786;
assign n_36813 = n_36804 ^ n_35876;
assign n_36814 = n_36804 ^ n_35867;
assign n_36815 = n_36805 ^ n_36441;
assign n_36816 = n_36807 ^ n_36483;
assign n_36817 = n_36807 ^ n_35813;
assign n_36818 = n_36808 ^ x155;
assign n_36819 = n_36809 ^ n_34961;
assign n_36820 = n_36810 ^ n_36808;
assign n_36821 = n_36812 ^ n_36793;
assign n_36822 = n_34874 & ~n_36813;
assign n_36823 = x359 & ~n_36814;
assign n_36824 = n_36814 ^ x359;
assign n_36825 = n_36815 ^ n_35007;
assign n_36826 = n_36816 ^ n_35813;
assign n_36827 = ~n_36816 & ~n_36817;
assign n_36828 = n_36819 ^ n_35007;
assign n_36829 = n_36819 ^ n_36815;
assign n_36830 = n_36820 & ~n_36818;
assign n_36831 = n_36820 ^ x155;
assign n_36832 = ~n_36821 & n_36803;
assign n_36833 = n_36821 ^ n_35895;
assign n_36834 = n_36822 ^ n_34899;
assign n_36835 = n_36823 ^ x358;
assign n_36836 = ~n_35748 & ~n_36826;
assign n_36837 = n_36747 ^ n_36826;
assign n_36838 = n_36535 ^ n_36827;
assign n_36839 = n_36828 ^ n_36815;
assign n_36840 = n_36825 & ~n_36829;
assign n_36841 = n_36830 ^ x155;
assign n_36842 = ~n_36811 & n_36831;
assign n_36843 = n_36831 ^ n_36811;
assign n_36844 = n_36832 ^ n_35895;
assign n_36845 = n_36794 & n_36833;
assign n_36846 = n_36833 ^ n_36794;
assign n_36847 = n_35409 & ~n_36833;
assign n_36848 = n_36836 ^ n_36483;
assign n_36849 = n_35761 & n_36838;
assign n_36850 = n_36839 ^ x154;
assign n_36851 = n_36840 ^ n_35007;
assign n_36852 = n_36841 ^ n_36839;
assign n_36853 = n_36844 ^ n_36843;
assign n_36854 = n_36844 ^ n_35940;
assign y6 = n_36846;
assign n_36855 = n_36847 ^ n_35895;
assign n_36856 = n_36848 ^ n_35032;
assign n_36857 = n_36849 ^ n_36498;
assign n_36858 = n_36851 ^ n_35032;
assign n_36859 = n_36851 ^ n_36848;
assign n_36860 = ~n_36852 & n_36850;
assign n_36861 = n_36852 ^ x154;
assign n_36862 = n_36853 ^ n_35940;
assign n_36863 = ~n_36853 & ~n_36854;
assign n_36864 = n_36855 ^ n_36834;
assign n_36865 = n_36855 ^ n_36822;
assign n_36866 = n_36858 ^ n_36848;
assign n_36867 = n_36856 & ~n_36859;
assign n_36868 = n_36860 ^ x154;
assign n_36869 = n_36842 & ~n_36861;
assign n_36870 = n_36861 ^ n_36842;
assign n_36871 = n_36845 & ~n_36862;
assign n_36872 = n_36862 ^ n_36845;
assign n_36873 = n_35444 & n_36862;
assign n_36874 = n_36863 ^ n_35940;
assign n_36875 = n_36864 ^ n_36823;
assign n_36876 = n_36834 & n_36865;
assign n_36877 = n_36866 ^ x153;
assign n_36878 = n_36867 ^ n_35032;
assign n_36879 = n_36868 ^ n_36866;
assign n_36880 = n_36870 ^ n_35965;
assign y5 = ~n_36872;
assign n_36881 = n_36873 ^ n_35940;
assign n_36882 = n_36870 ^ n_36874;
assign n_36883 = n_36874 ^ n_35965;
assign n_36884 = n_36875 & n_36835;
assign n_36885 = n_36875 ^ x358;
assign n_36886 = n_36876 ^ n_34899;
assign n_36887 = n_36878 ^ n_35061;
assign n_36888 = ~n_36879 & n_36877;
assign n_36889 = n_36879 ^ x153;
assign n_36890 = n_36881 ^ n_34946;
assign n_36891 = ~n_36880 & n_36882;
assign n_36892 = n_36870 ^ n_36883;
assign n_36893 = n_36884 ^ x358;
assign n_36894 = ~n_36824 & ~n_36885;
assign n_36895 = n_36885 ^ n_36824;
assign n_36896 = n_36886 ^ n_34946;
assign n_36897 = n_36886 ^ n_36881;
assign n_36898 = n_36887 ^ n_36857;
assign n_36899 = n_36888 ^ x153;
assign n_36900 = n_36869 & ~n_36889;
assign n_36901 = n_36889 ^ n_36869;
assign n_36902 = n_36891 ^ n_35965;
assign n_36903 = n_36871 & n_36892;
assign n_36904 = n_36892 ^ n_36871;
assign n_36905 = n_35481 & ~n_36892;
assign n_36906 = n_36893 ^ x357;
assign n_36907 = n_36896 ^ n_36881;
assign n_36908 = n_36890 & ~n_36897;
assign n_36909 = n_36899 ^ n_36898;
assign n_36910 = n_36901 ^ n_36006;
assign n_36911 = n_36901 ^ n_36902;
assign n_36912 = n_36902 ^ n_36006;
assign y4 = n_36904;
assign n_36913 = n_36905 ^ n_35965;
assign n_36914 = n_36893 ^ n_36907;
assign n_36915 = n_36908 ^ n_34946;
assign n_36916 = n_36909 ^ x152;
assign n_36917 = ~n_36910 & n_36911;
assign n_36918 = n_36901 ^ n_36912;
assign n_36919 = ~n_36914 & n_36906;
assign n_36920 = n_36914 ^ x357;
assign n_36921 = n_36915 ^ n_34976;
assign n_36922 = n_36913 ^ n_36915;
assign n_36923 = n_36916 ^ n_36900;
assign n_36924 = n_36917 ^ n_36006;
assign n_36925 = n_36903 & n_36918;
assign n_36926 = n_36918 ^ n_36903;
assign n_36927 = ~n_35512 & ~n_36918;
assign n_36928 = n_36919 ^ x357;
assign n_36929 = ~n_36894 & ~n_36920;
assign n_36930 = n_36920 ^ n_36894;
assign n_36931 = n_36913 ^ n_36921;
assign n_36932 = ~n_36921 & ~n_36922;
assign n_36933 = n_36923 ^ n_36046;
assign n_36934 = n_36923 ^ n_36924;
assign n_36935 = n_36924 ^ n_36046;
assign y3 = n_36926;
assign n_36936 = n_36927 ^ n_36006;
assign n_36937 = n_36928 ^ x356;
assign n_36938 = n_36928 ^ n_36931;
assign n_36939 = n_36932 ^ n_34976;
assign n_36940 = n_36933 & ~n_36934;
assign n_36941 = n_36923 ^ n_36935;
assign n_36942 = n_36936 ^ n_35017;
assign n_36943 = n_36938 & n_36937;
assign n_36944 = n_36938 ^ x356;
assign n_36945 = n_36939 ^ n_35017;
assign n_36946 = n_36939 ^ n_36936;
assign n_36947 = n_36940 ^ n_36046;
assign n_36948 = n_36925 & ~n_36941;
assign n_36949 = n_36941 ^ n_36925;
assign n_36950 = n_35548 & n_36941;
assign n_36951 = n_36943 ^ x356;
assign n_36952 = ~n_36929 & ~n_36944;
assign n_36953 = n_36944 ^ n_36929;
assign n_36954 = n_36945 ^ n_36936;
assign n_36955 = n_36942 & n_36946;
assign n_36956 = n_36947 ^ n_36084;
assign y2 = ~n_36949;
assign n_36957 = n_36950 ^ n_36046;
assign n_36958 = n_36951 ^ x355;
assign n_36959 = n_36951 ^ n_36954;
assign n_36960 = n_36955 ^ n_35017;
assign n_36961 = n_36956 & ~n_36099;
assign n_36962 = n_36956 ^ n_35912;
assign n_36963 = n_36959 & n_36958;
assign n_36964 = n_36959 ^ x355;
assign n_36965 = n_36960 ^ n_35052;
assign n_36966 = n_36957 ^ n_36960;
assign n_36967 = n_36961 ^ n_35912;
assign n_36968 = n_36948 & n_36962;
assign n_36969 = n_36962 ^ n_36948;
assign n_36970 = ~n_35593 & ~n_36962;
assign n_36971 = n_36963 ^ x355;
assign n_36972 = ~n_36952 & n_36964;
assign n_36973 = n_36964 ^ n_36952;
assign n_36974 = n_36957 ^ n_36965;
assign n_36975 = n_36965 & ~n_36966;
assign n_36976 = n_36136 ^ n_36967;
assign n_36977 = n_36967 ^ n_35947;
assign y1 = n_36969;
assign n_36978 = n_36970 ^ n_36084;
assign n_36979 = n_36971 ^ n_36974;
assign n_36980 = n_36974 ^ x354;
assign n_36981 = n_36975 ^ n_35052;
assign n_36982 = n_36976 ^ n_36968;
assign n_36983 = n_36968 & ~n_36976;
assign n_36984 = n_35635 & n_36976;
assign n_36985 = n_36136 & ~n_36977;
assign n_36986 = n_36978 ^ n_35094;
assign n_36987 = n_36979 ^ x354;
assign n_36988 = ~n_36979 & n_36980;
assign n_36989 = n_36981 ^ n_35094;
assign n_36990 = n_36981 ^ n_36978;
assign y0 = ~n_36982;
assign n_36991 = n_36984 ^ n_36124;
assign n_36992 = n_36985 ^ n_36124;
assign n_36993 = n_36972 & ~n_36987;
assign n_36994 = n_36987 ^ n_36972;
assign n_36995 = n_36988 ^ x354;
assign n_36996 = n_36989 ^ n_36978;
assign n_36997 = n_36986 & n_36990;
assign n_36998 = n_36992 ^ n_36162;
assign n_36999 = n_36995 ^ n_36996;
assign n_37000 = n_36996 ^ x353;
assign n_37001 = n_36997 ^ n_35094;
assign n_37002 = ~n_36998 & ~n_36176;
assign n_37003 = n_36998 ^ n_36016;
assign n_37004 = n_36999 ^ x353;
assign n_37005 = ~n_36999 & n_37000;
assign n_37006 = n_37001 ^ n_35117;
assign n_37007 = n_36991 ^ n_37001;
assign n_37008 = n_37002 ^ n_36016;
assign n_37009 = ~n_37003 & ~n_36983;
assign n_37010 = n_36983 ^ n_37003;
assign n_37011 = ~n_35670 & ~n_37003;
assign n_37012 = ~n_36993 & n_37004;
assign n_37013 = n_37004 ^ n_36993;
assign n_37014 = n_37005 ^ x353;
assign n_37015 = n_36991 ^ n_37006;
assign n_37016 = ~n_37006 & n_37007;
assign n_37017 = n_37008 ^ n_36202;
assign y15 = ~n_37010;
assign n_37018 = n_37011 ^ n_36162;
assign n_37019 = n_37014 ^ x352;
assign n_37020 = n_37014 ^ n_37015;
assign n_37021 = n_37016 ^ n_35117;
assign n_37022 = ~n_37017 & ~n_36216;
assign n_37023 = n_37017 ^ n_36048;
assign n_37024 = n_37018 ^ n_35147;
assign n_37025 = n_37020 & n_37019;
assign n_37026 = n_37020 ^ x352;
assign n_37027 = n_37021 ^ n_35147;
assign n_37028 = n_37021 ^ n_37018;
assign n_37029 = n_37022 ^ n_36048;
assign n_37030 = n_37009 & n_37023;
assign n_37031 = n_37023 ^ n_37009;
assign n_37032 = ~n_35713 & n_37023;
assign n_37033 = n_37025 ^ x352;
assign n_37034 = ~n_37026 & n_37012;
assign n_37035 = n_37012 ^ n_37026;
assign n_37036 = n_37027 ^ n_37018;
assign n_37037 = n_37024 & ~n_37028;
assign n_37038 = n_37029 ^ n_36245;
assign n_37039 = n_36094 ^ n_37029;
assign y14 = ~n_37031;
assign n_37040 = n_37032 ^ n_36202;
assign n_37041 = n_37033 ^ n_37036;
assign n_37042 = n_37036 ^ x367;
assign n_37043 = n_37037 ^ n_35147;
assign n_37044 = n_36258 & n_37038;
assign n_37045 = n_37039 ^ n_36245;
assign n_37046 = n_37040 ^ n_35166;
assign n_37047 = n_37041 ^ x367;
assign n_37048 = ~n_37041 & n_37042;
assign n_37049 = n_37043 ^ n_35166;
assign n_37050 = n_37043 ^ n_37040;
assign n_37051 = n_37044 ^ n_36094;
assign n_37052 = ~n_37030 & ~n_37045;
assign n_37053 = n_37045 ^ n_37030;
assign n_37054 = n_35754 & n_37045;
assign n_37055 = n_36824 ^ n_37045;
assign n_37056 = n_37034 & n_37047;
assign n_37057 = n_37047 ^ n_37034;
assign n_37058 = n_37048 ^ x367;
assign n_37059 = n_37049 ^ n_37040;
assign n_37060 = n_37046 & n_37050;
assign n_37061 = n_37051 ^ n_36285;
assign y13 = n_37053;
assign n_37062 = n_37054 ^ n_36245;
assign n_37063 = n_37058 ^ n_37059;
assign n_37064 = n_37059 ^ x366;
assign n_37065 = n_37060 ^ n_35166;
assign n_37066 = n_37061 & n_36299;
assign n_37067 = n_37061 ^ n_36141;
assign n_37068 = n_37062 ^ n_35181;
assign n_37069 = n_37063 ^ x366;
assign n_37070 = ~n_37063 & n_37064;
assign n_37071 = n_37065 ^ n_35181;
assign n_37072 = n_37065 ^ n_37062;
assign n_37073 = n_37066 ^ n_36141;
assign n_37074 = n_37052 & n_37067;
assign n_37075 = n_37067 ^ n_37052;
assign n_37076 = ~n_35794 & ~n_37067;
assign n_37077 = n_36895 ^ n_37067;
assign n_37078 = ~n_37056 & ~n_37069;
assign n_37079 = n_37069 ^ n_37056;
assign n_37080 = n_37070 ^ x366;
assign n_37081 = n_37071 ^ n_37062;
assign n_37082 = n_37068 & ~n_37072;
assign n_37083 = n_37073 ^ n_36323;
assign n_37084 = n_36180 ^ n_37073;
assign y12 = n_37075;
assign n_37085 = n_37076 ^ n_36285;
assign n_37086 = n_37080 ^ n_37081;
assign n_37087 = n_37081 ^ x365;
assign n_37088 = n_37082 ^ n_35181;
assign n_37089 = n_36338 & n_37083;
assign n_37090 = n_37084 ^ n_36323;
assign n_37091 = n_37085 ^ n_35199;
assign n_37092 = n_37086 ^ x365;
assign n_37093 = n_37086 & ~n_37087;
assign n_37094 = n_37088 ^ n_35199;
assign n_37095 = n_37088 ^ n_37085;
assign n_37096 = n_37089 ^ n_36180;
assign n_37097 = n_37074 & ~n_37090;
assign n_37098 = n_37090 ^ n_37074;
assign n_37099 = n_35824 & n_37090;
assign n_37100 = n_36930 ^ n_37090;
assign n_37101 = ~n_37078 & ~n_37092;
assign n_37102 = n_37092 ^ n_37078;
assign n_37103 = n_37093 ^ x365;
assign n_37104 = n_37094 ^ n_37085;
assign n_37105 = ~n_37091 & n_37095;
assign n_37106 = n_37096 ^ n_36367;
assign y11 = ~n_37098;
assign n_37107 = n_37099 ^ n_36323;
assign n_37108 = n_37103 ^ n_37104;
assign n_37109 = n_37104 ^ x364;
assign n_37110 = n_37105 ^ n_35199;
assign n_37111 = n_37106 & n_36381;
assign n_37112 = n_37106 ^ n_36221;
assign n_37113 = n_37107 ^ n_35223;
assign n_37114 = n_37108 ^ x364;
assign n_37115 = ~n_37108 & n_37109;
assign n_37116 = n_37110 ^ n_35223;
assign n_37117 = n_37110 ^ n_37107;
assign n_37118 = n_37111 ^ n_36221;
assign n_37119 = ~n_37097 & ~n_37112;
assign n_37120 = n_37112 ^ n_37097;
assign n_37121 = ~n_35850 & ~n_37112;
assign n_37122 = n_36953 ^ n_37112;
assign n_37123 = n_37101 & n_37114;
assign n_37124 = n_37114 ^ n_37101;
assign n_37125 = n_37115 ^ x364;
assign n_37126 = n_37116 ^ n_37107;
assign n_37127 = ~n_37113 & ~n_37117;
assign n_37128 = n_37118 ^ n_36405;
assign y10 = ~n_37120;
assign n_37129 = n_37121 ^ n_36367;
assign n_37130 = n_37125 ^ n_37126;
assign n_37131 = n_37126 ^ x363;
assign n_37132 = n_37127 ^ n_35223;
assign n_37133 = n_37128 & ~n_36420;
assign n_37134 = n_37128 ^ n_36263;
assign n_37135 = n_37129 ^ n_35242;
assign n_37136 = n_37130 ^ x363;
assign n_37137 = ~n_37130 & n_37131;
assign n_37138 = n_37132 ^ n_35242;
assign n_37139 = n_37132 ^ n_37129;
assign n_37140 = n_37133 ^ n_36263;
assign n_37141 = ~n_37119 & n_37134;
assign n_37142 = n_37134 ^ n_37119;
assign n_37143 = ~n_35877 & ~n_37134;
assign n_37144 = n_36973 ^ n_37134;
assign n_37145 = ~n_37123 & ~n_37136;
assign n_37146 = n_37136 ^ n_37123;
assign n_37147 = n_37137 ^ x363;
assign n_37148 = n_37138 ^ n_37129;
assign n_37149 = ~n_37135 & ~n_37139;
assign n_37150 = n_37140 ^ n_36448;
assign y9 = ~n_37142;
assign n_37151 = n_37143 ^ n_36405;
assign n_37152 = n_37147 ^ n_37148;
assign n_37153 = n_37148 ^ x362;
assign n_37154 = n_37149 ^ n_35242;
assign n_37155 = n_37150 ^ n_36304;
assign n_37156 = n_37150 & ~n_36463;
assign n_37157 = n_37151 ^ n_35256;
assign n_37158 = n_37152 ^ x362;
assign n_37159 = n_37152 & ~n_37153;
assign n_37160 = n_37154 ^ n_35256;
assign n_37161 = n_37154 ^ n_37151;
assign n_37162 = n_37155 ^ n_37141;
assign n_37163 = n_37141 & n_37155;
assign n_37164 = n_35893 & ~n_37155;
assign n_37165 = n_36994 ^ n_37155;
assign n_37166 = n_37156 ^ n_36304;
assign n_37167 = n_37158 & n_37145;
assign n_37168 = n_37145 ^ n_37158;
assign n_37169 = n_37159 ^ x362;
assign n_37170 = n_37160 ^ n_37151;
assign n_37171 = ~n_37157 & ~n_37161;
assign y8 = n_37162;
assign n_37172 = n_37164 ^ n_36448;
assign n_37173 = n_36343 ^ n_37166;
assign n_37174 = n_36504 ^ n_37166;
assign n_37175 = n_37169 ^ n_37170;
assign n_37176 = n_37170 ^ x361;
assign n_37177 = n_37171 ^ n_35256;
assign n_37178 = n_37172 ^ n_35276;
assign n_37179 = ~n_36504 & ~n_37173;
assign n_37180 = ~n_37163 & ~n_37174;
assign n_37181 = n_37174 ^ n_37163;
assign n_37182 = ~n_35926 & ~n_37174;
assign n_37183 = n_37013 ^ n_37174;
assign n_37184 = n_37175 ^ x361;
assign n_37185 = ~n_37175 & n_37176;
assign n_37186 = n_37177 ^ n_35276;
assign n_37187 = n_37177 ^ n_37172;
assign n_37188 = n_37179 ^ n_36489;
assign y23 = ~n_37181;
assign n_37189 = n_37182 ^ n_36489;
assign n_37190 = n_37167 & ~n_37184;
assign n_37191 = n_37184 ^ n_37167;
assign n_37192 = n_37185 ^ x361;
assign n_37193 = n_37186 ^ n_37172;
assign n_37194 = n_37178 & n_37187;
assign n_37195 = n_37188 ^ n_36529;
assign n_37196 = n_36385 ^ n_37188;
assign n_37197 = n_37189 ^ n_35297;
assign n_37198 = n_37192 ^ n_37193;
assign n_37199 = n_37193 ^ x360;
assign n_37200 = n_37194 ^ n_35276;
assign n_37201 = n_36543 & n_37195;
assign n_37202 = n_37196 ^ n_36529;
assign n_37203 = n_37198 ^ x360;
assign n_37204 = ~n_37198 & n_37199;
assign n_37205 = n_37200 ^ n_35297;
assign n_37206 = n_37200 ^ n_37189;
assign n_37207 = n_37201 ^ n_36385;
assign n_37208 = ~n_37180 & n_37202;
assign n_37209 = n_37202 ^ n_37180;
assign n_37210 = n_35957 & ~n_37202;
assign n_37211 = n_37035 ^ n_37202;
assign n_37212 = n_37190 & ~n_37203;
assign n_37213 = n_37203 ^ n_37190;
assign n_37214 = n_37204 ^ x360;
assign n_37215 = n_37205 ^ n_37189;
assign n_37216 = ~n_37197 & ~n_37206;
assign n_37217 = n_37207 ^ n_36563;
assign y22 = ~n_37209;
assign n_37218 = n_37210 ^ n_36529;
assign n_37219 = n_37214 ^ x375;
assign n_37220 = n_37215 ^ x375;
assign n_37221 = n_37214 ^ n_37215;
assign n_37222 = n_37216 ^ n_35297;
assign n_37223 = n_37217 & n_36574;
assign n_37224 = n_37217 ^ n_36426;
assign n_37225 = n_37218 ^ n_35317;
assign n_37226 = n_37219 ^ n_37215;
assign n_37227 = n_37220 & ~n_37221;
assign n_37228 = n_37222 ^ n_37218;
assign n_37229 = n_37223 ^ n_36426;
assign n_37230 = ~n_37208 & n_37224;
assign n_37231 = n_37224 ^ n_37208;
assign n_37232 = ~n_35999 & n_37224;
assign n_37233 = n_37057 ^ n_37224;
assign n_37234 = ~n_37212 & n_37226;
assign n_37235 = n_37226 ^ n_37212;
assign n_37236 = n_37227 ^ x375;
assign n_37237 = n_37228 ^ n_35317;
assign n_37238 = ~n_37228 & n_37225;
assign n_37239 = n_37229 ^ n_36590;
assign y21 = n_37231;
assign n_37240 = n_37232 ^ n_36563;
assign n_37241 = n_37236 ^ n_37237;
assign n_37242 = n_37237 ^ x374;
assign n_37243 = n_37238 ^ n_35317;
assign n_37244 = n_37239 & ~n_36599;
assign n_37245 = n_37239 ^ n_36468;
assign n_37246 = n_37240 ^ n_35341;
assign n_37247 = n_37241 ^ x374;
assign n_37248 = ~n_37241 & n_37242;
assign n_37249 = n_37243 ^ n_35341;
assign n_37250 = n_37243 ^ n_37240;
assign n_37251 = n_37244 ^ n_36468;
assign n_37252 = ~n_37230 & ~n_37245;
assign n_37253 = n_37245 ^ n_37230;
assign n_37254 = ~n_36026 & n_37245;
assign n_37255 = n_37079 ^ n_37245;
assign n_37256 = ~n_37234 & ~n_37247;
assign n_37257 = n_37247 ^ n_37234;
assign n_37258 = n_37248 ^ x374;
assign n_37259 = n_37249 ^ n_37240;
assign n_37260 = n_37246 & n_37250;
assign n_37261 = n_37251 ^ n_36613;
assign y20 = n_37253;
assign n_37262 = n_37254 ^ n_36590;
assign n_37263 = n_37258 ^ n_37259;
assign n_37264 = n_37259 ^ x373;
assign n_37265 = n_37260 ^ n_35341;
assign n_37266 = n_37261 & n_36621;
assign n_37267 = n_37261 ^ n_36509;
assign n_37268 = n_37262 ^ n_35355;
assign n_37269 = n_37263 ^ x373;
assign n_37270 = ~n_37263 & n_37264;
assign n_37271 = n_37265 ^ n_35355;
assign n_37272 = n_37265 ^ n_37262;
assign n_37273 = n_37266 ^ n_36509;
assign n_37274 = n_37252 & n_37267;
assign n_37275 = n_37267 ^ n_37252;
assign n_37276 = n_37102 ^ n_37267;
assign n_37277 = n_36063 & ~n_37267;
assign n_37278 = ~n_37256 & n_37269;
assign n_37279 = n_37269 ^ n_37256;
assign n_37280 = n_37270 ^ x373;
assign n_37281 = n_37271 ^ n_37262;
assign n_37282 = ~n_37268 & n_37272;
assign n_37283 = n_37273 ^ n_36628;
assign y19 = n_37275;
assign n_37284 = n_37277 ^ n_36613;
assign n_37285 = n_37280 ^ n_37281;
assign n_37286 = n_37281 ^ x372;
assign n_37287 = n_37282 ^ n_35355;
assign n_37288 = n_37283 & ~n_36635;
assign n_37289 = n_37283 ^ n_36548;
assign n_37290 = n_37284 ^ n_35385;
assign n_37291 = n_37285 ^ x372;
assign n_37292 = ~n_37285 & n_37286;
assign n_37293 = n_37287 ^ n_37284;
assign n_37294 = n_37287 ^ n_35385;
assign n_37295 = n_37288 ^ n_36548;
assign n_37296 = n_37274 & n_37289;
assign n_37297 = n_37289 ^ n_37274;
assign n_37298 = ~n_36103 & ~n_37289;
assign n_37299 = n_37124 ^ n_37289;
assign n_37300 = n_37278 ^ n_37291;
assign n_37301 = ~n_37291 & ~n_37278;
assign n_37302 = n_37292 ^ x372;
assign n_37303 = ~n_37290 & n_37293;
assign n_37304 = n_37294 ^ n_37284;
assign n_37305 = n_37295 ^ n_36653;
assign n_37306 = n_36660 ^ n_37295;
assign y18 = n_37297;
assign n_37307 = n_37298 ^ n_36628;
assign n_37308 = n_37303 ^ n_35385;
assign n_37309 = n_37304 ^ x371;
assign n_37310 = n_37302 ^ n_37304;
assign n_37311 = n_36660 & ~n_37305;
assign n_37312 = ~n_37296 & n_37306;
assign n_37313 = n_37306 ^ n_37296;
assign n_37314 = n_37146 ^ n_37306;
assign n_37315 = n_36155 & n_37306;
assign n_37316 = n_37307 ^ n_35404;
assign n_37317 = n_37308 ^ n_37307;
assign n_37318 = n_37308 ^ n_35404;
assign n_37319 = n_37302 ^ n_37309;
assign n_37320 = n_37309 & ~n_37310;
assign n_37321 = n_37311 ^ n_36579;
assign y17 = n_37313;
assign n_37322 = n_37315 ^ n_36653;
assign n_37323 = ~n_37316 & ~n_37317;
assign n_37324 = n_37318 ^ n_37307;
assign n_37325 = n_37301 & ~n_37319;
assign n_37326 = n_37319 ^ n_37301;
assign n_37327 = n_37320 ^ x371;
assign n_37328 = n_36679 ^ n_37321;
assign n_37329 = n_37321 ^ n_36671;
assign n_37330 = n_37322 ^ n_35439;
assign n_37331 = n_37323 ^ n_35404;
assign n_37332 = n_37324 ^ x370;
assign n_37333 = n_37327 ^ n_37324;
assign n_37334 = n_37327 ^ x370;
assign n_37335 = n_37328 ^ n_37312;
assign n_37336 = ~n_37312 & ~n_37328;
assign n_37337 = n_37168 ^ n_37328;
assign n_37338 = n_36183 & n_37328;
assign n_37339 = n_36679 & ~n_37329;
assign n_37340 = n_37322 ^ n_37331;
assign n_37341 = n_37332 & ~n_37333;
assign n_37342 = n_37334 ^ n_37324;
assign y16 = n_37335;
assign n_37343 = n_37338 ^ n_36671;
assign n_37344 = n_37339 ^ n_36604;
assign n_37345 = ~n_37340 & n_37330;
assign n_37346 = n_37340 ^ n_35439;
assign n_37347 = n_37341 ^ x370;
assign n_37348 = n_37325 & ~n_37342;
assign n_37349 = n_37342 ^ n_37325;
assign n_37350 = n_37343 ^ n_35460;
assign n_37351 = n_37344 ^ n_36626;
assign n_37352 = n_37344 ^ n_36700;
assign n_37353 = n_37345 ^ n_35439;
assign n_37354 = n_37346 ^ x369;
assign n_37355 = n_37347 ^ n_37346;
assign n_37356 = ~n_36700 & ~n_37351;
assign n_37357 = ~n_37336 & ~n_37352;
assign n_37358 = n_37352 ^ n_37336;
assign n_37359 = n_37191 ^ n_37352;
assign n_37360 = n_36224 & ~n_37352;
assign n_37361 = n_37343 ^ n_37353;
assign n_37362 = n_37350 ^ n_37353;
assign n_37363 = ~n_37355 & n_37354;
assign n_37364 = n_37355 ^ x369;
assign n_37365 = n_37356 ^ n_36693;
assign y31 = ~n_37358;
assign n_37366 = n_37360 ^ n_36693;
assign n_37367 = n_37350 & ~n_37361;
assign n_37368 = n_37362 ^ x368;
assign n_37369 = n_37363 ^ x369;
assign n_37370 = n_37364 & ~n_37348;
assign n_37371 = n_37348 ^ n_37364;
assign n_37372 = n_37365 ^ n_36714;
assign n_37373 = n_37367 ^ n_35460;
assign n_37374 = n_37362 ^ n_37369;
assign n_37375 = n_37368 ^ n_37369;
assign n_37376 = n_36794 & ~n_37371;
assign n_37377 = n_37371 ^ n_36787;
assign n_37378 = ~n_37372 & n_36721;
assign n_37379 = n_37372 ^ n_36647;
assign n_37380 = n_37373 ^ n_35507;
assign n_37381 = n_37373 ^ n_37366;
assign n_37382 = n_37368 & ~n_37374;
assign n_37383 = n_37375 & n_37370;
assign n_37384 = n_37370 ^ n_37375;
assign n_37385 = n_37377 ^ n_35876;
assign n_37386 = n_37378 ^ n_36647;
assign n_37387 = ~n_37379 & n_37357;
assign n_37388 = n_37357 ^ n_37379;
assign n_37389 = n_37213 ^ n_37379;
assign n_37390 = ~n_36264 & ~n_37379;
assign n_37391 = n_37380 ^ n_37366;
assign n_37392 = n_37380 & n_37381;
assign n_37393 = n_37382 ^ x368;
assign n_37394 = n_37384 ^ n_36833;
assign n_37395 = n_37384 ^ n_37376;
assign n_37396 = n_35876 & n_37385;
assign y103 = ~n_37385;
assign n_37397 = n_37386 ^ n_36735;
assign y30 = n_37388;
assign n_37398 = n_37390 ^ n_36714;
assign n_37399 = n_37391 ^ x383;
assign n_37400 = n_37392 ^ n_35507;
assign n_37401 = n_37391 ^ n_37393;
assign n_37402 = n_37393 ^ x383;
assign n_37403 = n_37394 ^ n_37376;
assign n_37404 = n_37394 & ~n_37395;
assign n_37405 = n_37396 ^ n_36794;
assign n_37406 = n_37396 ^ n_36795;
assign n_37407 = ~n_37397 & n_36741;
assign n_37408 = n_37397 ^ n_36665;
assign n_37409 = n_37398 ^ n_35546;
assign n_37410 = n_37400 ^ n_37398;
assign n_37411 = ~n_37399 & n_37401;
assign n_37412 = n_37391 ^ n_37402;
assign n_37413 = n_35895 & ~n_37403;
assign y102 = ~n_37403;
assign n_37414 = n_37404 ^ n_36833;
assign n_37415 = ~n_35375 & ~n_37405;
assign n_37416 = x71 & n_37406;
assign n_37417 = n_37406 ^ x71;
assign n_37418 = n_37407 ^ n_36665;
assign n_37419 = n_37387 & ~n_37408;
assign n_37420 = n_37408 ^ n_37387;
assign n_37421 = n_36317 & ~n_37408;
assign n_37422 = n_37235 ^ n_37408;
assign n_37423 = n_37410 & n_37409;
assign n_37424 = n_37410 ^ n_35546;
assign n_37425 = n_37411 ^ x383;
assign n_37426 = n_37412 & ~n_37383;
assign n_37427 = n_37383 ^ n_37412;
assign n_37428 = n_37413 ^ n_36833;
assign n_37429 = n_37415 ^ n_35409;
assign n_37430 = n_37418 ^ n_36754;
assign y29 = n_37420;
assign n_37431 = n_37421 ^ n_36735;
assign n_37432 = n_37423 ^ n_35546;
assign n_37433 = n_37425 ^ n_37424;
assign n_37434 = n_37425 ^ x382;
assign n_37435 = n_37414 ^ n_37427;
assign n_37436 = n_37427 ^ n_36862;
assign n_37437 = n_37428 ^ n_37415;
assign n_37438 = ~n_37430 & ~n_36761;
assign n_37439 = n_37430 ^ n_36685;
assign n_37440 = n_37431 ^ n_35574;
assign n_37441 = n_37431 ^ n_37432;
assign n_37442 = n_37433 ^ x382;
assign n_37443 = ~n_37433 & n_37434;
assign n_37444 = n_37435 ^ n_36862;
assign n_37445 = ~n_37435 & ~n_37436;
assign n_37446 = n_37437 & n_37429;
assign n_37447 = n_37437 ^ n_35409;
assign n_37448 = n_37438 ^ n_36685;
assign n_37449 = ~n_37419 & ~n_37439;
assign n_37450 = n_37439 ^ n_37419;
assign n_37451 = n_37257 ^ n_37439;
assign n_37452 = n_36346 & n_37439;
assign n_37453 = n_37440 ^ n_37432;
assign n_37454 = n_37440 & ~n_37441;
assign n_37455 = n_37442 & ~n_37426;
assign n_37456 = n_37426 ^ n_37442;
assign n_37457 = n_37443 ^ x382;
assign n_37458 = ~n_35940 & n_37444;
assign n_37459 = ~n_37403 & n_37444;
assign n_37460 = n_37444 ^ n_37403;
assign n_37461 = n_37445 ^ n_36862;
assign n_37462 = n_37446 ^ n_35409;
assign n_37463 = n_37447 ^ x70;
assign n_37464 = n_37447 ^ n_37416;
assign n_37465 = n_37448 ^ n_36774;
assign n_37466 = n_36706 ^ n_37448;
assign y28 = n_37450;
assign n_37467 = n_37452 ^ n_36754;
assign n_37468 = n_37453 ^ x381;
assign n_37469 = n_37454 ^ n_35574;
assign n_37470 = n_37456 ^ n_36892;
assign n_37471 = n_37453 ^ n_37457;
assign n_37472 = n_37458 ^ n_36862;
assign y101 = n_37460;
assign n_37473 = n_37456 ^ n_37461;
assign n_37474 = n_37462 ^ n_35444;
assign n_37475 = n_37463 ^ n_37416;
assign n_37476 = ~n_37463 & n_37464;
assign n_37477 = n_36781 & ~n_37465;
assign n_37478 = n_37466 ^ n_36774;
assign n_37479 = n_37467 ^ n_35627;
assign n_37480 = n_37468 ^ n_37457;
assign n_37481 = n_37467 ^ n_37469;
assign n_37482 = n_37470 ^ n_37461;
assign n_37483 = ~n_37468 & n_37471;
assign n_37484 = n_37472 ^ n_35444;
assign n_37485 = n_37472 ^ n_37462;
assign n_37486 = ~n_37470 & ~n_37473;
assign n_37487 = n_37472 ^ n_37474;
assign n_37488 = ~n_37417 & n_37475;
assign n_37489 = n_37475 ^ n_37417;
assign n_37490 = n_37476 ^ x70;
assign n_37491 = n_37477 ^ n_36706;
assign n_37492 = n_37449 & ~n_37478;
assign n_37493 = n_37478 ^ n_37449;
assign n_37494 = n_36400 & n_37478;
assign n_37495 = n_37279 ^ n_37478;
assign n_37496 = n_37479 ^ n_37469;
assign n_37497 = n_37480 & ~n_37455;
assign n_37498 = n_37455 ^ n_37480;
assign n_37499 = ~n_37479 & ~n_37481;
assign n_37500 = ~n_35965 & ~n_37482;
assign n_37501 = n_37482 & ~n_37459;
assign n_37502 = n_37459 ^ n_37482;
assign n_37503 = n_37483 ^ x381;
assign n_37504 = n_37484 & ~n_37485;
assign n_37505 = n_37486 ^ n_36892;
assign n_37506 = n_37487 ^ x69;
assign n_37507 = n_37487 ^ n_37490;
assign n_37508 = n_36727 ^ n_37491;
assign n_37509 = n_36806 ^ n_37491;
assign y27 = ~n_37493;
assign n_37510 = n_37494 ^ n_36774;
assign n_37511 = n_37496 ^ x380;
assign n_37512 = n_37499 ^ n_35627;
assign n_37513 = n_37500 ^ n_36892;
assign y100 = ~n_37502;
assign n_37514 = n_37496 ^ n_37503;
assign n_37515 = n_37503 ^ x380;
assign n_37516 = n_37504 ^ n_35444;
assign n_37517 = n_37505 ^ n_37498;
assign n_37518 = n_37505 ^ n_36918;
assign n_37519 = n_37506 ^ n_37490;
assign n_37520 = n_37506 & ~n_37507;
assign n_37521 = ~n_36806 & n_37508;
assign n_37522 = ~n_37492 & ~n_37509;
assign n_37523 = n_37509 ^ n_37492;
assign n_37524 = n_37300 ^ n_37509;
assign n_37525 = ~n_36441 & ~n_37509;
assign n_37526 = n_37510 ^ n_35655;
assign n_37527 = n_37512 ^ n_37510;
assign n_37528 = n_37511 & ~n_37514;
assign n_37529 = n_37496 ^ n_37515;
assign n_37530 = n_37516 ^ n_35481;
assign n_37531 = n_37516 ^ n_37513;
assign n_37532 = n_37517 ^ n_36918;
assign n_37533 = ~n_37517 & n_37518;
assign n_37534 = ~n_37488 & n_37519;
assign n_37535 = n_37519 ^ n_37488;
assign n_37536 = n_37520 ^ x69;
assign n_37537 = n_37521 ^ n_36797;
assign y26 = ~n_37523;
assign n_37538 = n_37525 ^ n_36797;
assign n_37539 = ~n_37527 & n_37526;
assign n_37540 = n_37527 ^ n_35655;
assign n_37541 = n_37528 ^ x380;
assign n_37542 = n_37497 & ~n_37529;
assign n_37543 = n_37529 ^ n_37497;
assign n_37544 = n_37530 ^ n_37513;
assign n_37545 = n_37530 & n_37531;
assign n_37546 = ~n_36006 & ~n_37532;
assign n_37547 = ~n_37532 & ~n_37501;
assign n_37548 = n_37501 ^ n_37532;
assign n_37549 = n_37533 ^ n_36918;
assign n_37550 = n_37537 ^ n_36826;
assign n_37551 = n_36837 ^ n_37537;
assign n_37552 = n_37538 ^ n_35695;
assign n_37553 = n_37539 ^ n_35655;
assign n_37554 = n_37540 ^ x379;
assign n_37555 = n_37541 ^ n_37540;
assign n_37556 = n_37543 ^ n_36941;
assign n_37557 = n_37536 ^ n_37544;
assign n_37558 = n_37544 ^ x68;
assign n_37559 = n_37545 ^ n_35481;
assign n_37560 = n_37546 ^ n_36918;
assign y99 = ~n_37548;
assign n_37561 = n_37543 ^ n_37549;
assign n_37562 = n_37549 ^ n_36941;
assign n_37563 = n_36837 & n_37550;
assign n_37564 = n_37522 & n_37551;
assign n_37565 = n_37551 ^ n_37522;
assign n_37566 = ~n_36483 & n_37551;
assign n_37567 = n_37553 ^ n_35695;
assign n_37568 = n_37553 ^ n_37538;
assign n_37569 = ~n_37555 & n_37554;
assign n_37570 = n_37555 ^ x379;
assign n_37571 = n_37557 ^ x68;
assign n_37572 = n_37557 & ~n_37558;
assign n_37573 = n_37559 ^ n_35512;
assign n_37574 = n_37560 ^ n_35512;
assign n_37575 = n_37560 ^ n_37559;
assign n_37576 = ~n_37556 & ~n_37561;
assign n_37577 = n_37543 ^ n_37562;
assign n_37578 = n_37563 ^ n_36747;
assign y25 = ~n_37565;
assign n_37579 = n_37566 ^ n_36826;
assign n_37580 = n_37567 ^ n_37538;
assign n_37581 = ~n_37552 & ~n_37568;
assign n_37582 = n_37569 ^ x379;
assign n_37583 = ~n_37570 & n_37542;
assign n_37584 = n_37542 ^ n_37570;
assign n_37585 = ~n_37534 & n_37571;
assign n_37586 = n_37571 ^ n_37534;
assign n_37587 = n_37572 ^ x68;
assign n_37588 = n_37560 ^ n_37573;
assign n_37589 = n_37574 & n_37575;
assign n_37590 = n_37576 ^ n_36941;
assign n_37591 = ~n_36046 & n_37577;
assign n_37592 = n_37577 & n_37547;
assign n_37593 = n_37547 ^ n_37577;
assign n_37594 = n_37578 ^ n_36767;
assign n_37595 = n_37579 ^ n_35748;
assign n_37596 = n_37580 ^ x378;
assign n_37597 = n_37581 ^ n_35695;
assign n_37598 = n_37580 ^ n_37582;
assign n_37599 = n_37584 ^ n_36962;
assign n_37600 = n_37587 ^ x67;
assign n_37601 = n_37588 ^ n_37587;
assign n_37602 = n_37589 ^ n_35512;
assign n_37603 = n_37584 ^ n_37590;
assign n_37604 = n_37591 ^ n_36941;
assign y98 = ~n_37593;
assign n_37605 = n_37594 ^ n_36838;
assign n_37606 = n_37596 ^ n_37582;
assign n_37607 = n_37597 ^ n_35748;
assign n_37608 = n_37597 ^ n_37579;
assign n_37609 = ~n_37596 & n_37598;
assign n_37610 = n_37599 ^ n_37590;
assign n_37611 = ~n_37601 & n_37600;
assign n_37612 = n_37601 ^ x67;
assign n_37613 = n_37602 ^ n_35548;
assign n_37614 = n_37599 & n_37603;
assign n_37615 = n_37604 ^ n_35548;
assign n_37616 = n_37604 ^ n_37602;
assign n_37617 = n_37605 ^ n_37564;
assign n_37618 = n_36498 & ~n_37605;
assign n_37619 = n_37349 ^ n_37605;
assign n_37620 = n_37606 & n_37583;
assign n_37621 = n_37583 ^ n_37606;
assign n_37622 = n_37607 ^ n_37579;
assign n_37623 = n_37595 & ~n_37608;
assign n_37624 = n_37609 ^ x378;
assign n_37625 = n_36084 & n_37610;
assign n_37626 = n_37610 & n_37592;
assign n_37627 = n_37592 ^ n_37610;
assign n_37628 = n_37611 ^ x67;
assign n_37629 = n_37585 & ~n_37612;
assign n_37630 = n_37612 ^ n_37585;
assign n_37631 = n_37604 ^ n_37613;
assign n_37632 = n_37614 ^ n_36962;
assign n_37633 = n_37615 & n_37616;
assign y24 = ~n_37617;
assign n_37634 = n_37618 ^ n_36838;
assign n_37635 = n_37619 ^ n_37326;
assign n_37636 = n_37621 ^ n_36976;
assign n_37637 = n_37622 ^ x377;
assign n_37638 = n_37623 ^ n_35748;
assign n_37639 = n_37624 ^ n_37622;
assign n_37640 = n_37625 ^ n_36962;
assign y97 = ~n_37627;
assign n_37641 = n_37631 ^ x66;
assign n_37642 = n_37631 ^ n_37628;
assign n_37643 = n_37621 ^ n_37632;
assign n_37644 = n_37633 ^ n_35548;
assign n_37645 = n_37636 ^ n_37632;
assign n_37646 = n_37638 ^ n_35761;
assign n_37647 = n_37639 & ~n_37637;
assign n_37648 = n_37639 ^ x377;
assign n_37649 = n_37640 ^ n_35593;
assign n_37650 = n_37641 ^ n_37628;
assign n_37651 = ~n_37641 & n_37642;
assign n_37652 = n_37636 & n_37643;
assign n_37653 = n_37640 ^ n_37644;
assign n_37654 = n_37644 ^ n_35593;
assign n_37655 = ~n_36124 & ~n_37645;
assign n_37656 = n_37626 ^ n_37645;
assign n_37657 = n_37645 & ~n_37626;
assign n_37658 = n_37646 ^ n_37634;
assign n_37659 = n_37647 ^ x377;
assign n_37660 = ~n_37648 & ~n_37620;
assign n_37661 = n_37620 ^ n_37648;
assign n_37662 = n_37629 & n_37650;
assign n_37663 = n_37650 ^ n_37629;
assign n_37664 = n_37651 ^ x66;
assign n_37665 = n_37652 ^ n_36976;
assign n_37666 = n_37649 & n_37653;
assign n_37667 = n_37640 ^ n_37654;
assign n_37668 = n_37655 ^ n_36976;
assign y96 = ~n_37656;
assign n_37669 = n_37659 ^ n_37658;
assign n_37670 = n_37661 ^ n_37003;
assign n_37671 = n_37664 ^ x65;
assign n_37672 = n_37665 ^ n_37661;
assign n_37673 = n_37666 ^ n_35593;
assign n_37674 = n_37667 ^ x65;
assign n_37675 = n_37667 ^ n_37664;
assign n_37676 = n_37668 ^ n_35635;
assign n_37677 = n_37669 ^ x376;
assign n_37678 = n_37667 ^ n_37671;
assign n_37679 = n_37672 & n_37670;
assign n_37680 = n_37672 ^ n_37003;
assign n_37681 = n_37668 ^ n_37673;
assign n_37682 = n_37673 ^ n_35635;
assign n_37683 = n_37674 & ~n_37675;
assign n_37684 = n_37677 ^ n_37660;
assign n_37685 = ~n_37662 & n_37678;
assign n_37686 = n_37678 ^ n_37662;
assign n_37687 = n_37679 ^ n_37003;
assign n_37688 = ~n_36162 & n_37680;
assign n_37689 = ~n_37680 & n_37657;
assign n_37690 = n_37657 ^ n_37680;
assign n_37691 = n_37676 & n_37681;
assign n_37692 = n_37668 ^ n_37682;
assign n_37693 = n_37683 ^ x65;
assign n_37694 = n_37684 ^ n_37023;
assign n_37695 = n_37684 ^ n_37687;
assign n_37696 = n_37687 ^ n_37023;
assign n_37697 = n_37688 ^ n_37003;
assign y111 = ~n_37690;
assign n_37698 = n_37691 ^ n_35635;
assign n_37699 = n_37692 ^ x64;
assign n_37700 = n_37692 ^ n_37693;
assign n_37701 = ~n_37694 & ~n_37695;
assign n_37702 = n_37684 ^ n_37696;
assign n_37703 = n_37697 ^ n_35670;
assign n_37704 = n_37697 ^ n_37698;
assign n_37705 = n_37698 ^ n_35670;
assign n_37706 = n_37699 ^ n_37693;
assign n_37707 = ~n_37699 & n_37700;
assign n_37708 = n_37701 ^ n_37023;
assign n_37709 = n_36202 & n_37702;
assign n_37710 = ~n_37702 & n_37689;
assign n_37711 = n_37689 ^ n_37702;
assign n_37712 = n_37703 & n_37704;
assign n_37713 = n_37697 ^ n_37705;
assign n_37714 = ~n_37685 & n_37706;
assign n_37715 = n_37706 ^ n_37685;
assign n_37716 = n_37707 ^ x64;
assign n_37717 = n_37708 ^ n_37045;
assign n_37718 = n_37708 ^ n_36824;
assign n_37719 = n_37709 ^ n_37023;
assign y110 = ~n_37711;
assign n_37720 = n_37712 ^ n_35670;
assign n_37721 = n_37713 ^ x79;
assign n_37722 = n_37716 ^ n_37713;
assign n_37723 = ~n_37055 & ~n_37717;
assign n_37724 = n_37718 ^ n_37045;
assign n_37725 = n_37719 ^ n_35713;
assign n_37726 = n_37719 ^ n_37720;
assign n_37727 = ~n_37722 & n_37721;
assign n_37728 = n_37722 ^ x79;
assign n_37729 = n_37723 ^ n_36824;
assign n_37730 = n_36245 & ~n_37724;
assign n_37731 = ~n_37724 & ~n_37710;
assign n_37732 = n_37710 ^ n_37724;
assign n_37733 = n_37725 ^ n_37720;
assign n_37734 = ~n_37725 & n_37726;
assign n_37735 = n_37727 ^ x79;
assign n_37736 = ~n_37714 & n_37728;
assign n_37737 = n_37728 ^ n_37714;
assign n_37738 = n_37729 ^ n_37067;
assign n_37739 = n_37730 ^ n_37045;
assign y109 = ~n_37732;
assign n_37740 = n_37733 ^ x78;
assign n_37741 = n_37734 ^ n_35713;
assign n_37742 = n_37733 ^ n_37735;
assign n_37743 = n_37735 ^ x78;
assign n_37744 = ~n_37738 & n_37077;
assign n_37745 = n_37738 ^ n_36895;
assign n_37746 = n_37739 ^ n_35754;
assign n_37747 = n_37739 ^ n_37741;
assign n_37748 = n_37741 ^ n_35754;
assign n_37749 = n_37740 & ~n_37742;
assign n_37750 = n_37733 ^ n_37743;
assign n_37751 = n_37744 ^ n_36895;
assign n_37752 = ~n_36285 & ~n_37745;
assign n_37753 = n_37745 & ~n_37731;
assign n_37754 = n_37731 ^ n_37745;
assign n_37755 = n_37746 & n_37747;
assign n_37756 = n_37739 ^ n_37748;
assign n_37757 = n_37749 ^ x78;
assign n_37758 = ~n_37736 & ~n_37750;
assign n_37759 = n_37750 ^ n_37736;
assign n_37760 = n_36930 ^ n_37751;
assign n_37761 = n_37100 ^ n_37751;
assign n_37762 = n_37752 ^ n_37067;
assign y108 = ~n_37754;
assign n_37763 = n_37755 ^ n_35754;
assign n_37764 = n_37756 ^ x77;
assign n_37765 = n_37756 ^ n_37757;
assign n_37766 = n_37757 ^ x77;
assign n_37767 = n_37100 & n_37760;
assign n_37768 = n_36323 & ~n_37761;
assign n_37769 = ~n_37761 & ~n_37753;
assign n_37770 = n_37753 ^ n_37761;
assign n_37771 = n_37762 ^ n_35794;
assign n_37772 = n_37763 ^ n_37762;
assign n_37773 = ~n_37764 & n_37765;
assign n_37774 = n_37756 ^ n_37766;
assign n_37775 = n_37767 ^ n_37090;
assign n_37776 = n_37768 ^ n_37090;
assign y107 = ~n_37770;
assign n_37777 = n_37772 & n_37771;
assign n_37778 = n_37772 ^ n_35794;
assign n_37779 = n_37773 ^ x77;
assign n_37780 = ~n_37758 & ~n_37774;
assign n_37781 = n_37774 ^ n_37758;
assign n_37782 = n_37775 ^ n_37112;
assign n_37783 = n_36953 ^ n_37775;
assign n_37784 = n_37776 ^ n_35824;
assign n_37785 = n_37777 ^ n_35794;
assign n_37786 = n_37778 ^ x76;
assign n_37787 = n_37779 ^ n_37778;
assign n_37788 = n_37122 & n_37782;
assign n_37789 = n_37783 ^ n_37112;
assign n_37790 = n_37776 ^ n_37785;
assign n_37791 = n_37785 ^ n_35824;
assign n_37792 = ~n_37787 & n_37786;
assign n_37793 = n_37787 ^ x76;
assign n_37794 = n_37788 ^ n_36953;
assign n_37795 = ~n_36367 & n_37789;
assign n_37796 = ~n_37789 & ~n_37769;
assign n_37797 = n_37769 ^ n_37789;
assign n_37798 = n_37784 & n_37790;
assign n_37799 = n_37776 ^ n_37791;
assign n_37800 = n_37792 ^ x76;
assign n_37801 = n_37780 & n_37793;
assign n_37802 = n_37793 ^ n_37780;
assign n_37803 = n_37794 ^ n_37134;
assign n_37804 = n_37795 ^ n_37112;
assign y106 = n_37797;
assign n_37805 = n_37798 ^ n_35824;
assign n_37806 = n_37799 ^ x75;
assign n_37807 = n_37800 ^ n_37799;
assign n_37808 = ~n_37803 & n_37144;
assign n_37809 = n_37803 ^ n_36973;
assign n_37810 = n_37804 ^ n_35850;
assign n_37811 = n_37804 ^ n_37805;
assign n_37812 = n_37805 ^ n_35850;
assign n_37813 = n_37807 & ~n_37806;
assign n_37814 = n_37807 ^ x75;
assign n_37815 = n_37808 ^ n_36973;
assign n_37816 = n_36405 & ~n_37809;
assign n_37817 = ~n_37809 & ~n_37796;
assign n_37818 = n_37796 ^ n_37809;
assign n_37819 = n_37810 & n_37811;
assign n_37820 = n_37804 ^ n_37812;
assign n_37821 = n_37813 ^ x75;
assign n_37822 = ~n_37801 & n_37814;
assign n_37823 = n_37814 ^ n_37801;
assign n_37824 = n_36994 ^ n_37815;
assign n_37825 = n_37165 ^ n_37815;
assign n_37826 = n_37816 ^ n_37134;
assign y105 = ~n_37818;
assign n_37827 = n_37819 ^ n_35850;
assign n_37828 = n_37820 ^ x74;
assign n_37829 = n_37821 ^ n_37820;
assign n_37830 = n_37165 & ~n_37824;
assign n_37831 = n_36448 & ~n_37825;
assign n_37832 = n_37825 ^ n_37417;
assign n_37833 = n_37817 ^ n_37825;
assign n_37834 = n_37825 & ~n_37817;
assign n_37835 = n_37826 ^ n_35877;
assign n_37836 = n_37826 ^ n_37827;
assign n_37837 = ~n_37829 & n_37828;
assign n_37838 = n_37829 ^ x74;
assign n_37839 = n_37830 ^ n_37155;
assign n_37840 = n_37831 ^ n_37155;
assign y104 = ~n_37833;
assign n_37841 = n_37835 ^ n_37827;
assign n_37842 = n_37835 & ~n_37836;
assign n_37843 = n_37837 ^ x74;
assign n_37844 = ~n_37822 & n_37838;
assign n_37845 = n_37838 ^ n_37822;
assign n_37846 = n_37839 ^ n_37174;
assign n_37847 = n_37840 ^ n_35893;
assign n_37848 = n_37841 ^ x73;
assign n_37849 = n_37842 ^ n_35877;
assign n_37850 = n_37841 ^ n_37843;
assign n_37851 = n_37843 ^ x73;
assign n_37852 = ~n_37846 & ~n_37183;
assign n_37853 = n_37846 ^ n_37013;
assign n_37854 = n_37840 ^ n_37849;
assign n_37855 = n_37847 ^ n_37849;
assign n_37856 = ~n_37848 & n_37850;
assign n_37857 = n_37841 ^ n_37851;
assign n_37858 = n_37852 ^ n_37013;
assign n_37859 = n_36489 & n_37853;
assign n_37860 = n_37489 ^ n_37853;
assign n_37861 = ~n_37853 & n_37834;
assign n_37862 = n_37834 ^ n_37853;
assign n_37863 = ~n_37847 & ~n_37854;
assign n_37864 = n_37855 ^ x72;
assign n_37865 = n_37856 ^ x73;
assign n_37866 = ~n_37844 & n_37857;
assign n_37867 = n_37857 ^ n_37844;
assign n_37868 = n_37035 ^ n_37858;
assign n_37869 = n_37211 ^ n_37858;
assign n_37870 = n_37859 ^ n_37174;
assign y119 = ~n_37862;
assign n_37871 = n_37863 ^ n_35893;
assign n_37872 = n_37865 ^ n_37855;
assign n_37873 = ~n_37211 & ~n_37868;
assign n_37874 = ~n_36529 & ~n_37869;
assign n_37875 = n_37535 ^ n_37869;
assign n_37876 = ~n_37869 & ~n_37861;
assign n_37877 = n_37861 ^ n_37869;
assign n_37878 = n_37870 ^ n_35926;
assign n_37879 = n_37870 ^ n_37871;
assign n_37880 = n_37871 ^ n_35926;
assign n_37881 = ~n_37872 & n_37864;
assign n_37882 = n_37872 ^ x72;
assign n_37883 = n_37873 ^ n_37202;
assign n_37884 = n_37874 ^ n_37202;
assign y118 = ~n_37877;
assign n_37885 = n_37878 & n_37879;
assign n_37886 = n_37870 ^ n_37880;
assign n_37887 = n_37881 ^ x72;
assign n_37888 = n_37866 & ~n_37882;
assign n_37889 = n_37882 ^ n_37866;
assign n_37890 = n_37883 ^ n_37224;
assign n_37891 = n_37884 ^ n_35957;
assign n_37892 = n_37885 ^ n_35926;
assign n_37893 = n_37886 ^ x87;
assign n_37894 = n_37886 ^ n_37887;
assign n_37895 = n_37890 & ~n_37233;
assign n_37896 = n_37890 ^ n_37057;
assign n_37897 = n_37884 ^ n_37892;
assign n_37898 = n_37891 ^ n_37892;
assign n_37899 = n_37893 ^ n_37887;
assign n_37900 = n_37893 & ~n_37894;
assign n_37901 = n_37895 ^ n_37057;
assign n_37902 = n_36563 & n_37896;
assign n_37903 = n_37586 ^ n_37896;
assign n_37904 = ~n_37896 & ~n_37876;
assign n_37905 = n_37876 ^ n_37896;
assign n_37906 = ~n_37891 & ~n_37897;
assign n_37907 = n_37898 ^ x86;
assign n_37908 = n_37888 & ~n_37899;
assign n_37909 = n_37899 ^ n_37888;
assign n_37910 = n_37900 ^ x87;
assign n_37911 = n_37901 ^ n_37245;
assign n_37912 = n_37902 ^ n_37224;
assign y117 = n_37905;
assign n_37913 = n_37906 ^ n_35957;
assign n_37914 = n_37898 ^ n_37910;
assign n_37915 = n_37907 ^ n_37910;
assign n_37916 = n_37911 & n_37255;
assign n_37917 = n_37911 ^ n_37079;
assign n_37918 = n_37912 ^ n_35999;
assign n_37919 = n_37913 ^ n_37912;
assign n_37920 = n_37913 ^ n_35999;
assign n_37921 = n_37907 & ~n_37914;
assign n_37922 = n_37908 & ~n_37915;
assign n_37923 = n_37915 ^ n_37908;
assign n_37924 = n_37916 ^ n_37079;
assign n_37925 = ~n_36590 & ~n_37917;
assign n_37926 = n_37630 ^ n_37917;
assign n_37927 = n_37917 & n_37904;
assign n_37928 = n_37904 ^ n_37917;
assign n_37929 = ~n_37918 & ~n_37919;
assign n_37930 = n_37920 ^ n_37912;
assign n_37931 = n_37921 ^ x86;
assign n_37932 = ~n_37385 & n_37923;
assign n_37933 = n_37923 ^ n_37385;
assign n_37934 = n_37924 ^ n_37267;
assign n_37935 = n_37102 ^ n_37924;
assign n_37936 = n_37925 ^ n_37245;
assign y116 = n_37928;
assign n_37937 = n_37929 ^ n_35999;
assign n_37938 = n_37930 ^ x85;
assign n_37939 = n_37931 ^ n_37930;
assign n_37940 = n_37932 ^ n_37403;
assign n_37941 = n_36794 & n_37933;
assign y71 = ~n_37933;
assign n_37942 = n_37276 & n_37934;
assign n_37943 = n_37935 ^ n_37267;
assign n_37944 = n_37936 ^ n_36026;
assign n_37945 = n_37936 ^ n_37937;
assign n_37946 = n_37937 ^ n_36026;
assign n_37947 = n_37931 ^ n_37938;
assign n_37948 = ~n_37938 & n_37939;
assign n_37949 = n_37941 ^ n_37385;
assign n_37950 = n_37941 ^ n_37377;
assign n_37951 = n_37942 ^ n_37102;
assign n_37952 = ~n_36613 & n_37943;
assign n_37953 = n_37663 ^ n_37943;
assign n_37954 = n_37943 & ~n_37927;
assign n_37955 = n_37927 ^ n_37943;
assign n_37956 = ~n_37944 & n_37945;
assign n_37957 = n_37936 ^ n_37946;
assign n_37958 = n_37922 & n_37947;
assign n_37959 = n_37947 ^ n_37922;
assign n_37960 = n_37948 ^ x85;
assign n_37961 = n_35876 & n_37949;
assign n_37962 = x295 & n_37950;
assign n_37963 = n_37950 ^ x295;
assign n_37964 = n_37951 ^ n_37289;
assign n_37965 = n_37952 ^ n_37267;
assign y115 = n_37955;
assign n_37966 = n_37956 ^ n_36026;
assign n_37967 = n_37957 ^ x84;
assign n_37968 = n_37959 ^ n_37932;
assign n_37969 = n_37959 ^ n_37940;
assign n_37970 = n_37960 ^ n_37957;
assign n_37971 = n_37961 ^ n_35895;
assign n_37972 = n_37962 ^ x294;
assign n_37973 = ~n_37964 & n_37299;
assign n_37974 = n_37964 ^ n_37124;
assign n_37975 = n_37965 ^ n_36063;
assign n_37976 = n_37965 ^ n_37966;
assign n_37977 = n_37940 & n_37968;
assign n_37978 = n_36833 & n_37969;
assign y70 = n_37969;
assign n_37979 = ~n_37970 & n_37967;
assign n_37980 = n_37970 ^ x84;
assign n_37981 = n_37973 ^ n_37124;
assign n_37982 = n_36628 & ~n_37974;
assign n_37983 = n_37686 ^ n_37974;
assign n_37984 = ~n_37974 & n_37954;
assign n_37985 = n_37954 ^ n_37974;
assign n_37986 = n_37975 ^ n_37966;
assign n_37987 = ~n_37975 & ~n_37976;
assign n_37988 = n_37977 ^ n_37403;
assign n_37989 = n_37978 ^ n_37403;
assign n_37990 = n_37979 ^ x84;
assign n_37991 = n_37980 & ~n_37958;
assign n_37992 = n_37958 ^ n_37980;
assign n_37993 = n_37981 ^ n_37306;
assign n_37994 = n_37314 ^ n_37981;
assign n_37995 = n_37982 ^ n_37289;
assign y114 = n_37985;
assign n_37996 = n_37986 ^ x83;
assign n_37997 = n_37987 ^ n_36063;
assign n_37998 = n_37989 ^ n_37961;
assign n_37999 = n_37989 ^ n_37971;
assign n_38000 = n_37986 ^ n_37990;
assign n_38001 = n_37990 ^ x83;
assign n_38002 = n_37992 ^ n_37444;
assign n_38003 = n_37988 ^ n_37992;
assign n_38004 = n_37314 & n_37993;
assign n_38005 = ~n_36653 & ~n_37994;
assign n_38006 = n_37715 ^ n_37994;
assign n_38007 = n_37994 & ~n_37984;
assign n_38008 = n_37984 ^ n_37994;
assign n_38009 = n_37995 ^ n_36103;
assign n_38010 = n_37997 ^ n_37995;
assign n_38011 = n_37971 & n_37998;
assign n_38012 = n_37999 ^ n_37962;
assign n_38013 = n_37999 ^ n_37972;
assign n_38014 = n_37996 & ~n_38000;
assign n_38015 = n_37986 ^ n_38001;
assign n_38016 = n_37988 ^ n_38002;
assign n_38017 = n_38002 & n_38003;
assign n_38018 = n_38004 ^ n_37146;
assign n_38019 = n_38005 ^ n_37306;
assign y113 = ~n_38008;
assign n_38020 = n_38010 & n_38009;
assign n_38021 = n_38010 ^ n_36103;
assign n_38022 = n_38011 ^ n_35895;
assign n_38023 = n_37972 & n_38012;
assign n_38024 = n_37963 & ~n_38013;
assign n_38025 = n_38013 ^ n_37963;
assign n_38026 = n_38014 ^ x83;
assign n_38027 = ~n_38015 & ~n_37991;
assign n_38028 = n_37991 ^ n_38015;
assign n_38029 = ~n_36862 & ~n_38016;
assign n_38030 = ~n_38016 & n_37969;
assign n_38031 = n_37969 ^ n_38016;
assign n_38032 = n_38017 ^ n_37444;
assign n_38033 = n_37168 ^ n_38018;
assign n_38034 = n_37337 ^ n_38018;
assign n_38035 = n_38019 ^ n_36155;
assign n_38036 = n_38020 ^ n_36103;
assign n_38037 = n_38021 ^ x82;
assign n_38038 = n_38023 ^ x294;
assign n_38039 = n_38026 ^ n_38021;
assign n_38040 = n_38028 ^ n_37482;
assign n_38041 = n_38029 ^ n_37444;
assign y69 = n_38031;
assign n_38042 = n_38028 ^ n_38032;
assign n_38043 = n_38032 ^ n_37482;
assign n_38044 = n_37337 & ~n_38033;
assign n_38045 = ~n_36671 & n_38034;
assign n_38046 = n_37737 ^ n_38034;
assign n_38047 = n_38007 ^ n_38034;
assign n_38048 = ~n_38034 & n_38007;
assign n_38049 = n_38019 ^ n_38036;
assign n_38050 = n_38036 ^ n_36155;
assign n_38051 = ~n_38039 & n_38037;
assign n_38052 = n_38039 ^ x82;
assign n_38053 = n_38041 ^ n_35940;
assign n_38054 = n_38022 ^ n_38041;
assign n_38055 = ~n_38040 & ~n_38042;
assign n_38056 = n_38028 ^ n_38043;
assign n_38057 = n_38044 ^ n_37328;
assign n_38058 = n_38045 ^ n_37328;
assign y112 = ~n_38047;
assign n_38059 = n_38035 & n_38049;
assign n_38060 = n_38019 ^ n_38050;
assign n_38061 = n_38051 ^ x82;
assign n_38062 = n_38052 & ~n_38027;
assign n_38063 = n_38027 ^ n_38052;
assign n_38064 = n_38022 ^ n_38053;
assign n_38065 = ~n_38053 & ~n_38054;
assign n_38066 = n_38055 ^ n_37482;
assign n_38067 = n_36892 & ~n_38056;
assign n_38068 = ~n_38056 & n_38030;
assign n_38069 = n_38030 ^ n_38056;
assign n_38070 = n_38057 ^ n_37352;
assign n_38071 = n_37359 ^ n_38057;
assign n_38072 = n_38058 ^ n_36183;
assign n_38073 = n_38059 ^ n_36155;
assign n_38074 = n_38060 ^ x81;
assign n_38075 = n_38060 ^ n_38061;
assign n_38076 = n_38063 ^ n_37532;
assign n_38077 = n_38038 ^ n_38064;
assign n_38078 = n_38064 ^ x293;
assign n_38079 = n_38065 ^ n_35940;
assign n_38080 = n_38063 ^ n_38066;
assign n_38081 = n_38067 ^ n_37482;
assign y68 = n_38069;
assign n_38082 = n_37359 & n_38070;
assign n_38083 = n_36693 & n_38071;
assign n_38084 = n_37759 ^ n_38071;
assign n_38085 = ~n_38071 & n_38048;
assign n_38086 = n_38048 ^ n_38071;
assign n_38087 = n_38058 ^ n_38073;
assign n_38088 = n_38072 ^ n_38073;
assign n_38089 = n_38074 ^ n_38061;
assign n_38090 = ~n_38074 & n_38075;
assign n_38091 = n_38076 ^ n_38066;
assign n_38092 = n_38077 ^ x293;
assign n_38093 = n_38077 & ~n_38078;
assign n_38094 = n_38079 ^ n_35965;
assign n_38095 = ~n_38076 & n_38080;
assign n_38096 = n_38081 ^ n_35965;
assign n_38097 = n_38079 ^ n_38081;
assign n_38098 = n_38082 ^ n_37191;
assign n_38099 = n_38083 ^ n_37352;
assign y127 = ~n_38086;
assign n_38100 = n_38072 & ~n_38087;
assign n_38101 = n_38088 ^ x80;
assign n_38102 = n_38089 & ~n_38062;
assign n_38103 = n_38062 ^ n_38089;
assign n_38104 = n_38090 ^ x81;
assign n_38105 = n_36918 & n_38091;
assign n_38106 = n_38091 & n_38068;
assign n_38107 = n_38068 ^ n_38091;
assign n_38108 = ~n_38092 & n_38024;
assign n_38109 = n_38024 ^ n_38092;
assign n_38110 = n_38093 ^ x293;
assign n_38111 = n_38094 ^ n_38081;
assign n_38112 = n_38095 ^ n_37532;
assign n_38113 = n_38096 & ~n_38097;
assign n_38114 = n_37213 ^ n_38098;
assign n_38115 = n_37389 ^ n_38098;
assign n_38116 = n_38099 ^ n_36224;
assign n_38117 = n_38100 ^ n_36183;
assign n_38118 = n_38104 ^ n_38088;
assign n_38119 = n_38105 ^ n_37532;
assign y67 = ~n_38107;
assign n_38120 = n_38110 ^ x292;
assign n_38121 = n_38111 ^ x292;
assign n_38122 = n_38110 ^ n_38111;
assign n_38123 = n_38112 ^ n_38103;
assign n_38124 = n_38112 ^ n_37577;
assign n_38125 = n_38113 ^ n_35965;
assign n_38126 = n_37389 & ~n_38114;
assign n_38127 = n_36714 & ~n_38115;
assign n_38128 = n_37781 ^ n_38115;
assign n_38129 = n_38115 & n_38085;
assign n_38130 = n_38085 ^ n_38115;
assign n_38131 = n_38099 ^ n_38117;
assign n_38132 = n_38117 ^ n_36224;
assign n_38133 = ~n_38118 & n_38101;
assign n_38134 = n_38118 ^ x80;
assign n_38135 = n_38119 ^ n_36006;
assign n_38136 = n_38120 ^ n_38111;
assign n_38137 = ~n_38121 & n_38122;
assign n_38138 = n_38123 ^ n_37577;
assign n_38139 = ~n_38123 & ~n_38124;
assign n_38140 = n_38119 ^ n_38125;
assign n_38141 = n_38125 ^ n_36006;
assign n_38142 = n_38126 ^ n_37379;
assign n_38143 = n_38127 ^ n_37379;
assign y126 = n_38130;
assign n_38144 = ~n_38116 & n_38131;
assign n_38145 = n_38099 ^ n_38132;
assign n_38146 = n_38133 ^ x80;
assign n_38147 = n_38102 & ~n_38134;
assign n_38148 = n_38134 ^ n_38102;
assign n_38149 = n_38108 & ~n_38136;
assign n_38150 = n_38136 ^ n_38108;
assign n_38151 = n_38137 ^ x292;
assign n_38152 = ~n_36941 & n_38138;
assign n_38153 = n_38138 & n_38106;
assign n_38154 = n_38106 ^ n_38138;
assign n_38155 = n_38139 ^ n_37577;
assign n_38156 = n_38135 & ~n_38140;
assign n_38157 = n_38119 ^ n_38141;
assign n_38158 = n_38142 ^ n_37408;
assign n_38159 = n_38143 ^ n_36264;
assign n_38160 = n_38144 ^ n_36224;
assign n_38161 = n_38145 ^ x95;
assign n_38162 = n_38145 ^ n_38146;
assign n_38163 = n_38146 ^ x95;
assign n_38164 = n_38148 ^ n_37610;
assign n_38165 = n_38151 ^ x291;
assign n_38166 = n_38152 ^ n_37577;
assign y66 = ~n_38154;
assign n_38167 = n_38155 ^ n_38148;
assign n_38168 = n_38156 ^ n_36006;
assign n_38169 = n_38157 ^ x291;
assign n_38170 = n_38151 ^ n_38157;
assign n_38171 = ~n_38158 & ~n_37422;
assign n_38172 = n_38158 ^ n_37235;
assign n_38173 = n_38143 ^ n_38160;
assign n_38174 = n_38160 ^ n_36264;
assign n_38175 = ~n_38161 & n_38162;
assign n_38176 = n_38145 ^ n_38163;
assign n_38177 = n_38165 ^ n_38157;
assign n_38178 = n_38166 ^ n_36046;
assign n_38179 = n_38167 & ~n_38164;
assign n_38180 = n_38167 ^ n_37610;
assign n_38181 = n_38168 ^ n_38166;
assign n_38182 = ~n_38169 & n_38170;
assign n_38183 = n_38171 ^ n_37235;
assign n_38184 = n_36735 & n_38172;
assign n_38185 = n_37802 ^ n_38172;
assign n_38186 = ~n_38172 & n_38129;
assign n_38187 = n_38129 ^ n_38172;
assign n_38188 = n_38159 & n_38173;
assign n_38189 = n_38143 ^ n_38174;
assign n_38190 = n_38175 ^ x95;
assign n_38191 = ~n_38147 & ~n_38176;
assign n_38192 = n_38176 ^ n_38147;
assign n_38193 = ~n_38149 & n_38177;
assign n_38194 = n_38177 ^ n_38149;
assign n_38195 = n_38179 ^ n_37610;
assign n_38196 = n_36962 & ~n_38180;
assign n_38197 = ~n_38180 & n_38153;
assign n_38198 = n_38153 ^ n_38180;
assign n_38199 = n_38181 & ~n_38178;
assign n_38200 = n_38181 ^ n_36046;
assign n_38201 = n_38182 ^ x291;
assign n_38202 = n_38183 ^ n_37439;
assign n_38203 = n_37257 ^ n_38183;
assign n_38204 = n_38184 ^ n_37408;
assign y125 = ~n_38187;
assign n_38205 = n_38188 ^ n_36264;
assign n_38206 = n_38189 ^ x94;
assign n_38207 = n_38189 ^ n_38190;
assign n_38208 = n_38192 ^ n_37645;
assign n_38209 = n_38192 ^ n_38195;
assign n_38210 = n_38196 ^ n_37610;
assign y65 = n_38198;
assign n_38211 = n_38199 ^ n_36046;
assign n_38212 = n_38200 ^ x290;
assign n_38213 = n_38200 ^ n_38201;
assign n_38214 = n_38201 ^ x290;
assign n_38215 = n_37451 & ~n_38202;
assign n_38216 = n_38203 ^ n_37439;
assign n_38217 = n_38204 ^ n_36317;
assign n_38218 = n_38204 ^ n_38205;
assign n_38219 = n_38205 ^ n_36317;
assign n_38220 = n_38206 ^ n_38190;
assign n_38221 = n_38206 & ~n_38207;
assign n_38222 = n_38208 ^ n_38195;
assign n_38223 = n_38208 & n_38209;
assign n_38224 = n_38210 ^ n_36084;
assign n_38225 = n_38211 ^ n_38210;
assign n_38226 = n_38212 & ~n_38213;
assign n_38227 = n_38200 ^ n_38214;
assign n_38228 = n_38215 ^ n_37257;
assign n_38229 = n_36754 & n_38216;
assign n_38230 = n_37823 ^ n_38216;
assign n_38231 = ~n_38216 & n_38186;
assign n_38232 = n_38186 ^ n_38216;
assign n_38233 = ~n_38217 & ~n_38218;
assign n_38234 = n_38204 ^ n_38219;
assign n_38235 = ~n_38220 & ~n_38191;
assign n_38236 = n_38191 ^ n_38220;
assign n_38237 = n_38221 ^ x94;
assign n_38238 = ~n_36976 & n_38222;
assign n_38239 = n_38197 ^ n_38222;
assign n_38240 = n_38222 & n_38197;
assign n_38241 = n_38223 ^ n_37645;
assign n_38242 = n_38225 & n_38224;
assign n_38243 = n_38225 ^ n_36084;
assign n_38244 = n_38226 ^ x290;
assign n_38245 = n_38227 & ~n_38193;
assign n_38246 = n_38193 ^ n_38227;
assign n_38247 = n_38228 ^ n_37478;
assign n_38248 = n_38228 ^ n_37279;
assign n_38249 = n_38228 ^ n_37495;
assign n_38250 = n_38229 ^ n_37439;
assign y124 = ~n_38232;
assign n_38251 = n_38233 ^ n_36317;
assign n_38252 = n_38234 ^ x93;
assign n_38253 = n_38236 ^ n_37680;
assign n_38254 = n_38234 ^ n_38237;
assign n_38255 = n_38238 ^ n_37645;
assign y64 = ~n_38239;
assign n_38256 = n_38236 ^ n_38241;
assign n_38257 = n_38241 ^ n_37680;
assign n_38258 = n_38242 ^ n_36084;
assign n_38259 = n_38243 ^ x289;
assign n_38260 = n_38243 ^ n_38244;
assign n_38261 = n_38247 & ~n_38248;
assign n_38262 = ~n_36774 & n_38249;
assign n_38263 = n_37845 ^ n_38249;
assign n_38264 = n_38249 & ~n_38231;
assign n_38265 = n_38231 ^ n_38249;
assign n_38266 = n_38250 ^ n_36346;
assign n_38267 = n_38250 ^ n_38251;
assign n_38268 = n_38251 ^ n_36346;
assign n_38269 = n_38252 ^ n_38237;
assign n_38270 = n_38252 & ~n_38254;
assign n_38271 = n_38255 ^ n_36124;
assign n_38272 = n_38253 & n_38256;
assign n_38273 = n_38236 ^ n_38257;
assign n_38274 = n_38255 ^ n_38258;
assign n_38275 = n_38259 ^ n_38244;
assign n_38276 = ~n_38259 & n_38260;
assign n_38277 = n_38261 ^ n_37478;
assign n_38278 = n_38262 ^ n_37478;
assign y123 = n_38265;
assign n_38279 = n_38266 & ~n_38267;
assign n_38280 = n_38250 ^ n_38268;
assign n_38281 = n_38269 & ~n_38235;
assign n_38282 = n_38235 ^ n_38269;
assign n_38283 = n_38270 ^ x93;
assign n_38284 = n_38271 ^ n_38258;
assign n_38285 = n_38272 ^ n_37680;
assign n_38286 = n_37003 & ~n_38273;
assign n_38287 = n_38273 & ~n_38240;
assign n_38288 = n_38240 ^ n_38273;
assign n_38289 = n_38271 & n_38274;
assign n_38290 = n_38245 & ~n_38275;
assign n_38291 = n_38275 ^ n_38245;
assign n_38292 = n_38276 ^ x289;
assign n_38293 = n_38277 ^ n_37509;
assign n_38294 = n_37300 ^ n_38277;
assign n_38295 = n_38278 ^ n_36400;
assign n_38296 = n_38279 ^ n_36346;
assign n_38297 = n_38280 ^ x92;
assign n_38298 = n_38282 ^ n_37702;
assign n_38299 = n_38283 ^ n_38280;
assign n_38300 = n_38284 ^ x288;
assign n_38301 = n_38282 ^ n_38285;
assign n_38302 = n_38286 ^ n_37680;
assign y79 = ~n_38288;
assign n_38303 = n_38289 ^ n_36124;
assign n_38304 = n_38284 ^ n_38292;
assign n_38305 = ~n_37524 & n_38293;
assign n_38306 = n_38294 ^ n_37509;
assign n_38307 = n_38278 ^ n_38296;
assign n_38308 = n_38296 ^ n_36400;
assign n_38309 = n_38298 ^ n_38285;
assign n_38310 = ~n_38299 & n_38297;
assign n_38311 = n_38299 ^ x92;
assign n_38312 = n_38300 ^ n_38292;
assign n_38313 = n_38298 & ~n_38301;
assign n_38314 = n_38302 ^ n_36162;
assign n_38315 = n_38302 ^ n_38303;
assign n_38316 = n_38300 & ~n_38304;
assign n_38317 = n_38305 ^ n_37300;
assign n_38318 = ~n_36797 & ~n_38306;
assign n_38319 = n_37867 ^ n_38306;
assign n_38320 = n_38306 & ~n_38264;
assign n_38321 = n_38264 ^ n_38306;
assign n_38322 = n_38295 & ~n_38307;
assign n_38323 = n_38278 ^ n_38308;
assign n_38324 = ~n_37023 & n_38309;
assign n_38325 = ~n_38309 & n_38287;
assign n_38326 = n_38287 ^ n_38309;
assign n_38327 = n_38310 ^ x92;
assign n_38328 = ~n_38281 & ~n_38311;
assign n_38329 = n_38311 ^ n_38281;
assign n_38330 = ~n_38290 & ~n_38312;
assign n_38331 = n_38312 ^ n_38290;
assign n_38332 = n_38313 ^ n_37702;
assign n_38333 = n_38314 ^ n_38303;
assign n_38334 = ~n_38314 & n_38315;
assign n_38335 = n_38316 ^ x288;
assign n_38336 = n_38317 ^ n_37326;
assign n_38337 = n_38317 ^ n_37551;
assign n_38338 = n_38318 ^ n_37509;
assign y122 = ~n_38321;
assign n_38339 = n_38322 ^ n_36400;
assign n_38340 = n_38323 ^ x91;
assign n_38341 = n_38324 ^ n_37702;
assign y78 = ~n_38326;
assign n_38342 = n_38323 ^ n_38327;
assign n_38343 = n_38327 ^ x91;
assign n_38344 = n_38329 ^ n_37724;
assign n_38345 = n_38329 ^ n_38332;
assign n_38346 = n_38333 ^ x303;
assign n_38347 = n_38334 ^ n_36162;
assign n_38348 = n_38335 ^ n_38333;
assign n_38349 = n_38336 ^ n_37551;
assign n_38350 = ~n_38336 & ~n_38337;
assign n_38351 = n_38338 ^ n_36441;
assign n_38352 = n_38339 ^ n_38338;
assign n_38353 = n_38341 ^ n_36202;
assign n_38354 = n_38340 & ~n_38342;
assign n_38355 = n_38323 ^ n_38343;
assign n_38356 = n_38344 ^ n_38332;
assign n_38357 = ~n_38344 & ~n_38345;
assign n_38358 = n_38347 ^ n_36202;
assign n_38359 = n_38347 ^ n_38341;
assign n_38360 = ~n_38348 & n_38346;
assign n_38361 = n_38348 ^ x303;
assign n_38362 = n_36826 & ~n_38349;
assign n_38363 = n_38349 & n_38320;
assign n_38364 = n_38320 ^ n_38349;
assign n_38365 = n_37635 ^ n_38350;
assign n_38366 = n_38352 & n_38351;
assign n_38367 = n_38352 ^ n_36441;
assign n_38368 = n_38347 ^ n_38353;
assign n_38369 = n_38354 ^ x91;
assign n_38370 = ~n_38328 & n_38355;
assign n_38371 = n_38355 ^ n_38328;
assign n_38372 = ~n_37045 & ~n_38356;
assign n_38373 = ~n_38356 & ~n_38325;
assign n_38374 = n_38325 ^ n_38356;
assign n_38375 = n_38357 ^ n_37724;
assign n_38376 = ~n_38358 & n_38359;
assign n_38377 = n_38360 ^ x303;
assign n_38378 = n_38330 & ~n_38361;
assign n_38379 = n_38361 ^ n_38330;
assign n_38380 = n_38362 ^ n_37551;
assign y121 = n_38364;
assign n_38381 = ~n_36838 & ~n_38365;
assign n_38382 = n_37909 ^ n_38365;
assign n_38383 = n_38363 ^ n_38365;
assign n_38384 = n_38366 ^ n_36441;
assign n_38385 = n_38367 ^ x90;
assign n_38386 = n_38368 ^ x302;
assign n_38387 = n_38367 ^ n_38369;
assign n_38388 = n_38369 ^ x90;
assign n_38389 = n_38371 ^ n_37745;
assign n_38390 = n_38372 ^ n_37724;
assign y77 = ~n_38374;
assign n_38391 = n_38371 ^ n_38375;
assign n_38392 = n_38375 ^ n_37745;
assign n_38393 = n_38376 ^ n_36202;
assign n_38394 = n_38368 ^ n_38377;
assign n_38395 = n_38380 ^ n_36483;
assign n_38396 = n_38381 ^ n_37605;
assign n_38397 = n_38382 ^ n_37889;
assign y120 = n_38383;
assign n_38398 = n_38380 ^ n_38384;
assign n_38399 = n_38386 ^ n_38377;
assign n_38400 = n_38385 & ~n_38387;
assign n_38401 = n_38367 ^ n_38388;
assign n_38402 = n_38390 ^ n_36245;
assign n_38403 = ~n_38389 & n_38391;
assign n_38404 = n_38371 ^ n_38392;
assign n_38405 = n_38390 ^ n_38393;
assign n_38406 = ~n_38386 & n_38394;
assign n_38407 = n_38395 ^ n_38384;
assign n_38408 = ~n_38395 & n_38398;
assign n_38409 = n_38378 & n_38399;
assign n_38410 = n_38399 ^ n_38378;
assign n_38411 = n_38400 ^ x90;
assign n_38412 = ~n_38370 & ~n_38401;
assign n_38413 = n_38401 ^ n_38370;
assign n_38414 = n_38402 ^ n_38393;
assign n_38415 = n_38403 ^ n_37745;
assign n_38416 = n_37067 & n_38404;
assign n_38417 = n_38404 & n_38373;
assign n_38418 = n_38373 ^ n_38404;
assign n_38419 = ~n_38402 & n_38405;
assign n_38420 = n_38406 ^ x302;
assign n_38421 = n_38407 ^ x89;
assign n_38422 = n_38408 ^ n_36483;
assign n_38423 = n_38407 ^ n_38411;
assign n_38424 = n_38413 ^ n_37761;
assign n_38425 = n_38414 ^ x301;
assign n_38426 = n_38415 ^ n_38413;
assign n_38427 = n_38416 ^ n_37745;
assign y76 = ~n_38418;
assign n_38428 = n_38419 ^ n_36245;
assign n_38429 = n_38420 ^ n_38414;
assign n_38430 = n_38421 ^ n_38411;
assign n_38431 = n_38422 ^ n_36498;
assign n_38432 = n_38421 & ~n_38423;
assign n_38433 = n_38426 & ~n_38424;
assign n_38434 = n_38426 ^ n_37761;
assign n_38435 = n_38427 ^ n_36285;
assign n_38436 = n_38427 ^ n_38428;
assign n_38437 = n_38428 ^ n_36285;
assign n_38438 = n_38429 & ~n_38425;
assign n_38439 = n_38429 ^ x301;
assign n_38440 = ~n_38412 & n_38430;
assign n_38441 = n_38430 ^ n_38412;
assign n_38442 = n_38431 ^ n_38396;
assign n_38443 = n_38432 ^ x89;
assign n_38444 = n_38433 ^ n_37761;
assign n_38445 = ~n_37090 & n_38434;
assign n_38446 = n_38434 & n_38417;
assign n_38447 = n_38417 ^ n_38434;
assign n_38448 = n_38435 & n_38436;
assign n_38449 = n_38427 ^ n_38437;
assign n_38450 = n_38438 ^ x301;
assign n_38451 = ~n_38409 & ~n_38439;
assign n_38452 = n_38439 ^ n_38409;
assign n_38453 = n_38441 ^ n_37789;
assign n_38454 = n_38442 ^ x88;
assign n_38455 = n_38441 ^ n_38444;
assign n_38456 = n_38444 ^ n_37789;
assign n_38457 = n_38445 ^ n_37761;
assign y75 = ~n_38447;
assign n_38458 = n_38448 ^ n_36285;
assign n_38459 = n_38449 ^ x300;
assign n_38460 = n_38449 ^ n_38450;
assign n_38461 = n_38443 ^ n_38454;
assign n_38462 = n_38453 & n_38455;
assign n_38463 = n_38441 ^ n_38456;
assign n_38464 = n_38457 ^ n_36323;
assign n_38465 = n_38457 ^ n_38458;
assign n_38466 = n_38459 ^ n_38450;
assign n_38467 = n_38459 & ~n_38460;
assign n_38468 = n_38461 ^ n_38440;
assign n_38469 = n_38462 ^ n_37789;
assign n_38470 = n_37112 & ~n_38463;
assign n_38471 = n_38463 & ~n_38446;
assign n_38472 = n_38446 ^ n_38463;
assign n_38473 = n_38464 ^ n_38458;
assign n_38474 = ~n_38464 & ~n_38465;
assign n_38475 = n_38451 & n_38466;
assign n_38476 = n_38466 ^ n_38451;
assign n_38477 = n_38467 ^ x300;
assign n_38478 = n_38468 ^ n_37809;
assign n_38479 = n_38468 ^ n_38469;
assign n_38480 = n_38469 ^ n_37809;
assign n_38481 = n_38470 ^ n_37789;
assign y74 = ~n_38472;
assign n_38482 = n_38473 ^ x299;
assign n_38483 = n_38474 ^ n_36323;
assign n_38484 = ~n_37933 & n_38476;
assign n_38485 = n_38476 ^ n_37933;
assign n_38486 = n_38477 ^ n_38473;
assign n_38487 = n_38478 & n_38479;
assign n_38488 = n_38468 ^ n_38480;
assign n_38489 = n_38481 ^ n_36367;
assign n_38490 = n_38481 ^ n_38483;
assign n_38491 = n_38483 ^ n_36367;
assign n_38492 = n_38484 ^ n_37969;
assign y39 = n_38485;
assign n_38493 = ~n_38486 & n_38482;
assign n_38494 = n_38486 ^ x299;
assign n_38495 = n_38487 ^ n_37809;
assign n_38496 = n_37134 & n_38488;
assign n_38497 = n_38488 & ~n_38471;
assign n_38498 = n_38471 ^ n_38488;
assign n_38499 = ~n_38489 & ~n_38490;
assign n_38500 = n_38481 ^ n_38491;
assign n_38501 = n_38493 ^ x299;
assign n_38502 = ~n_38475 & ~n_38494;
assign n_38503 = n_38494 ^ n_38475;
assign n_38504 = n_38495 ^ n_37832;
assign n_38505 = n_38495 ^ n_37825;
assign n_38506 = n_38496 ^ n_37809;
assign y73 = n_38498;
assign n_38507 = n_38499 ^ n_36367;
assign n_38508 = n_38500 ^ x298;
assign n_38509 = n_38500 ^ n_38501;
assign n_38510 = n_38501 ^ x298;
assign n_38511 = n_38503 ^ n_38484;
assign n_38512 = n_38503 ^ n_38492;
assign n_38513 = n_37155 & n_38504;
assign n_38514 = n_38497 ^ n_38504;
assign n_38515 = n_38504 & n_38497;
assign n_38516 = ~n_37832 & ~n_38505;
assign n_38517 = n_38506 ^ n_36405;
assign n_38518 = n_38507 ^ n_38506;
assign n_38519 = ~n_38508 & n_38509;
assign n_38520 = n_38500 ^ n_38510;
assign n_38521 = ~n_38492 & n_38511;
assign n_38522 = ~n_38485 & n_38512;
assign n_38523 = n_38512 ^ n_38485;
assign n_38524 = n_38513 ^ n_37825;
assign y72 = ~n_38514;
assign n_38525 = n_38516 ^ n_37417;
assign n_38526 = ~n_38518 & ~n_38517;
assign n_38527 = n_38518 ^ n_36405;
assign n_38528 = n_38519 ^ x298;
assign n_38529 = ~n_38502 & ~n_38520;
assign n_38530 = n_38520 ^ n_38502;
assign n_38531 = n_38521 ^ n_37969;
assign y38 = ~n_38523;
assign n_38532 = n_38524 ^ n_36448;
assign n_38533 = n_37860 ^ n_38525;
assign n_38534 = n_38525 ^ n_37853;
assign n_38535 = n_38526 ^ n_36405;
assign n_38536 = n_38527 ^ x297;
assign n_38537 = n_38527 ^ n_38528;
assign n_38538 = n_38528 ^ x297;
assign n_38539 = n_38530 ^ n_38016;
assign n_38540 = n_38530 ^ n_38531;
assign n_38541 = n_38531 ^ n_38016;
assign n_38542 = n_37174 & ~n_38533;
assign n_38543 = n_38533 & ~n_38515;
assign n_38544 = n_38515 ^ n_38533;
assign n_38545 = ~n_37860 & ~n_38534;
assign n_38546 = n_38535 ^ n_36448;
assign n_38547 = n_38524 ^ n_38535;
assign n_38548 = n_38536 & ~n_38537;
assign n_38549 = n_38527 ^ n_38538;
assign n_38550 = n_38539 & n_38540;
assign n_38551 = n_38530 ^ n_38541;
assign n_38552 = n_38542 ^ n_37853;
assign y87 = ~n_38544;
assign n_38553 = n_38545 ^ n_37489;
assign n_38554 = n_38524 ^ n_38546;
assign n_38555 = ~n_38532 & n_38547;
assign n_38556 = n_38548 ^ x297;
assign n_38557 = ~n_38529 & ~n_38549;
assign n_38558 = n_38549 ^ n_38529;
assign n_38559 = n_38550 ^ n_38016;
assign n_38560 = ~n_38551 & n_38522;
assign n_38561 = n_38522 ^ n_38551;
assign n_38562 = n_38552 ^ n_36489;
assign n_38563 = n_38553 ^ n_37535;
assign n_38564 = n_38553 ^ n_37869;
assign n_38565 = n_38554 ^ x296;
assign n_38566 = n_38555 ^ n_36448;
assign n_38567 = n_38554 ^ n_38556;
assign n_38568 = n_38558 ^ n_38056;
assign n_38569 = n_38559 ^ n_38558;
assign y37 = ~n_38561;
assign n_38570 = n_38563 ^ n_37869;
assign n_38571 = ~n_37875 & ~n_38564;
assign n_38572 = n_38565 ^ n_38556;
assign n_38573 = n_38552 ^ n_38566;
assign n_38574 = ~n_38565 & n_38567;
assign n_38575 = n_38569 & ~n_38568;
assign n_38576 = n_38569 ^ n_38056;
assign n_38577 = n_37202 & n_38570;
assign n_38578 = n_38570 & ~n_38543;
assign n_38579 = n_38543 ^ n_38570;
assign n_38580 = n_38571 ^ n_37535;
assign n_38581 = n_38557 & n_38572;
assign n_38582 = n_38572 ^ n_38557;
assign n_38583 = n_38573 ^ n_36489;
assign n_38584 = ~n_38573 & n_38562;
assign n_38585 = n_38574 ^ x296;
assign n_38586 = n_38575 ^ n_38056;
assign n_38587 = ~n_38560 & n_38576;
assign n_38588 = n_38576 ^ n_38560;
assign n_38589 = n_38577 ^ n_37869;
assign y86 = n_38579;
assign n_38590 = n_38580 ^ n_37896;
assign n_38591 = n_38582 ^ n_38091;
assign n_38592 = n_38583 ^ x311;
assign n_38593 = n_38584 ^ n_36489;
assign n_38594 = n_38585 ^ n_38583;
assign n_38595 = n_38586 ^ n_38582;
assign y36 = n_38588;
assign n_38596 = n_38589 ^ n_36529;
assign n_38597 = n_38590 ^ n_37586;
assign n_38598 = ~n_38590 & ~n_37903;
assign n_38599 = n_38593 ^ n_38589;
assign n_38600 = ~n_38594 & n_38592;
assign n_38601 = n_38594 ^ x311;
assign n_38602 = n_38595 & n_38591;
assign n_38603 = n_38595 ^ n_38091;
assign n_38604 = ~n_37224 & ~n_38597;
assign n_38605 = n_38597 & ~n_38578;
assign n_38606 = n_38578 ^ n_38597;
assign n_38607 = n_38598 ^ n_37586;
assign n_38608 = n_38599 ^ n_36529;
assign n_38609 = n_38599 & n_38596;
assign n_38610 = n_38600 ^ x311;
assign n_38611 = ~n_38581 & n_38601;
assign n_38612 = n_38601 ^ n_38581;
assign n_38613 = n_38602 ^ n_38091;
assign n_38614 = ~n_38587 & n_38603;
assign n_38615 = n_38603 ^ n_38587;
assign n_38616 = n_38604 ^ n_37896;
assign y85 = ~n_38606;
assign n_38617 = n_38607 ^ n_37917;
assign n_38618 = n_37926 ^ n_38607;
assign n_38619 = n_38608 ^ x310;
assign n_38620 = n_38609 ^ n_36529;
assign n_38621 = n_38610 ^ n_38608;
assign n_38622 = n_38612 ^ n_38138;
assign n_38623 = n_38612 ^ n_38613;
assign n_38624 = n_38613 ^ n_38138;
assign y35 = ~n_38615;
assign n_38625 = n_38616 ^ n_36563;
assign n_38626 = n_37926 & ~n_38617;
assign n_38627 = ~n_37245 & ~n_38618;
assign n_38628 = ~n_38618 & ~n_38605;
assign n_38629 = n_38605 ^ n_38618;
assign n_38630 = n_38620 ^ n_36563;
assign n_38631 = n_38620 ^ n_38616;
assign n_38632 = n_38621 ^ x310;
assign n_38633 = ~n_38621 & n_38619;
assign n_38634 = n_38622 & ~n_38623;
assign n_38635 = n_38612 ^ n_38624;
assign n_38636 = n_38626 ^ n_37630;
assign n_38637 = n_38627 ^ n_37917;
assign y84 = ~n_38629;
assign n_38638 = n_38630 ^ n_38616;
assign n_38639 = n_38625 & n_38631;
assign n_38640 = n_38632 ^ n_38611;
assign n_38641 = ~n_38611 & ~n_38632;
assign n_38642 = n_38633 ^ x310;
assign n_38643 = n_38634 ^ n_38138;
assign n_38644 = n_38614 & ~n_38635;
assign n_38645 = n_38635 ^ n_38614;
assign n_38646 = n_37663 ^ n_38636;
assign n_38647 = n_37953 ^ n_38636;
assign n_38648 = n_38637 ^ n_36590;
assign n_38649 = n_38638 ^ x309;
assign n_38650 = n_38639 ^ n_36563;
assign n_38651 = n_38640 ^ n_38180;
assign n_38652 = n_38642 ^ n_38638;
assign n_38653 = n_38640 ^ n_38643;
assign y34 = ~n_38645;
assign n_38654 = n_37953 & n_38646;
assign n_38655 = n_37267 & ~n_38647;
assign n_38656 = ~n_38647 & n_38628;
assign n_38657 = n_38628 ^ n_38647;
assign n_38658 = n_38637 ^ n_38650;
assign n_38659 = n_38648 ^ n_38650;
assign n_38660 = n_38651 ^ n_38643;
assign n_38661 = n_38652 ^ x309;
assign n_38662 = n_38652 & ~n_38649;
assign n_38663 = ~n_38651 & ~n_38653;
assign n_38664 = n_38654 ^ n_37943;
assign n_38665 = n_38655 ^ n_37943;
assign y83 = n_38657;
assign n_38666 = n_38648 & n_38658;
assign n_38667 = n_38659 ^ x308;
assign n_38668 = n_38644 & n_38660;
assign n_38669 = n_38660 ^ n_38644;
assign n_38670 = n_38661 ^ n_38641;
assign n_38671 = n_38641 & n_38661;
assign n_38672 = n_38662 ^ x309;
assign n_38673 = n_38663 ^ n_38180;
assign n_38674 = n_38664 ^ n_37974;
assign n_38675 = n_38665 ^ n_36613;
assign n_38676 = n_38666 ^ n_36590;
assign y33 = n_38669;
assign n_38677 = n_38670 ^ n_38222;
assign n_38678 = n_38672 ^ n_38659;
assign n_38679 = n_38673 ^ n_38670;
assign n_38680 = n_38674 & ~n_37983;
assign n_38681 = n_38674 ^ n_37686;
assign n_38682 = n_38665 ^ n_38676;
assign n_38683 = n_38675 ^ n_38676;
assign n_38684 = ~n_38678 & n_38667;
assign n_38685 = n_38678 ^ x308;
assign n_38686 = n_38679 ^ n_38222;
assign n_38687 = n_38679 & n_38677;
assign n_38688 = n_38680 ^ n_37686;
assign n_38689 = n_37289 & ~n_38681;
assign n_38690 = n_38681 ^ n_37963;
assign n_38691 = ~n_38681 & n_38656;
assign n_38692 = n_38656 ^ n_38681;
assign n_38693 = ~n_38675 & n_38682;
assign n_38694 = n_38683 ^ x307;
assign n_38695 = n_38684 ^ x308;
assign n_38696 = ~n_38671 & n_38685;
assign n_38697 = n_38685 ^ n_38671;
assign n_38698 = n_38686 ^ n_38668;
assign n_38699 = ~n_38668 & ~n_38686;
assign n_38700 = n_38687 ^ n_38222;
assign n_38701 = n_38006 ^ n_38688;
assign n_38702 = n_38688 ^ n_37994;
assign n_38703 = n_37715 ^ n_38688;
assign n_38704 = n_38689 ^ n_37974;
assign y82 = n_38692;
assign n_38705 = n_38693 ^ n_36613;
assign n_38706 = n_38683 ^ n_38695;
assign n_38707 = n_38694 ^ n_38695;
assign n_38708 = n_38697 ^ n_38273;
assign y32 = ~n_38698;
assign n_38709 = n_38697 ^ n_38700;
assign n_38710 = ~n_37306 & n_38701;
assign n_38711 = n_38025 ^ n_38701;
assign n_38712 = ~n_38701 & ~n_38691;
assign n_38713 = n_38691 ^ n_38701;
assign n_38714 = ~n_38702 & n_38703;
assign n_38715 = n_38704 ^ n_36628;
assign n_38716 = n_38704 ^ n_38705;
assign n_38717 = n_38705 ^ n_36628;
assign n_38718 = n_38694 & ~n_38706;
assign n_38719 = n_38696 & n_38707;
assign n_38720 = n_38707 ^ n_38696;
assign n_38721 = n_38708 ^ n_38700;
assign n_38722 = ~n_38708 & ~n_38709;
assign n_38723 = n_38710 ^ n_37994;
assign y81 = n_38713;
assign n_38724 = n_38714 ^ n_37994;
assign n_38725 = ~n_38715 & ~n_38716;
assign n_38726 = n_38704 ^ n_38717;
assign n_38727 = n_38718 ^ x307;
assign n_38728 = n_38720 ^ n_38309;
assign n_38729 = n_38699 & ~n_38721;
assign n_38730 = n_38721 ^ n_38699;
assign n_38731 = n_38722 ^ n_38273;
assign n_38732 = n_38723 ^ n_36653;
assign n_38733 = n_38724 ^ n_38034;
assign n_38734 = n_38725 ^ n_36628;
assign n_38735 = n_38726 ^ x306;
assign n_38736 = n_38727 ^ n_38726;
assign y47 = n_38730;
assign n_38737 = n_38731 ^ n_38720;
assign n_38738 = n_38733 ^ n_37737;
assign n_38739 = n_38733 & n_38046;
assign n_38740 = n_38734 ^ n_36653;
assign n_38741 = n_38723 ^ n_38734;
assign n_38742 = ~n_38736 & n_38735;
assign n_38743 = n_38736 ^ x306;
assign n_38744 = ~n_38737 & ~n_38728;
assign n_38745 = n_38737 ^ n_38309;
assign n_38746 = ~n_37328 & ~n_38738;
assign n_38747 = n_38109 ^ n_38738;
assign n_38748 = n_38712 ^ n_38738;
assign n_38749 = ~n_38738 & ~n_38712;
assign n_38750 = n_38739 ^ n_37737;
assign n_38751 = n_38723 ^ n_38740;
assign n_38752 = n_38732 & n_38741;
assign n_38753 = n_38742 ^ x306;
assign n_38754 = n_38719 & n_38743;
assign n_38755 = n_38743 ^ n_38719;
assign n_38756 = n_38744 ^ n_38309;
assign n_38757 = n_38729 & n_38745;
assign n_38758 = n_38745 ^ n_38729;
assign n_38759 = n_38746 ^ n_38034;
assign y80 = ~n_38748;
assign n_38760 = n_38084 ^ n_38750;
assign n_38761 = n_38750 ^ n_38071;
assign n_38762 = n_37759 ^ n_38750;
assign n_38763 = n_38751 ^ x305;
assign n_38764 = n_38752 ^ n_36653;
assign n_38765 = n_38751 ^ n_38753;
assign n_38766 = n_38753 ^ x305;
assign n_38767 = n_38755 ^ n_38356;
assign n_38768 = n_38755 ^ n_38756;
assign n_38769 = n_38756 ^ n_38356;
assign y46 = ~n_38758;
assign n_38770 = n_38759 ^ n_36671;
assign n_38771 = n_37352 & n_38760;
assign n_38772 = n_38150 ^ n_38760;
assign n_38773 = ~n_38760 & ~n_38749;
assign n_38774 = n_38749 ^ n_38760;
assign n_38775 = n_38761 & ~n_38762;
assign n_38776 = n_38764 ^ n_36671;
assign n_38777 = n_38764 ^ n_38759;
assign n_38778 = n_38763 & ~n_38765;
assign n_38779 = n_38751 ^ n_38766;
assign n_38780 = n_38767 & n_38768;
assign n_38781 = n_38755 ^ n_38769;
assign n_38782 = n_38771 ^ n_38071;
assign y95 = n_38774;
assign n_38783 = n_38775 ^ n_38071;
assign n_38784 = n_38776 ^ n_38759;
assign n_38785 = ~n_38770 & n_38777;
assign n_38786 = n_38778 ^ x305;
assign n_38787 = n_38754 & n_38779;
assign n_38788 = n_38779 ^ n_38754;
assign n_38789 = n_38780 ^ n_38356;
assign n_38790 = ~n_38757 & ~n_38781;
assign n_38791 = n_38781 ^ n_38757;
assign n_38792 = n_38782 ^ n_36693;
assign n_38793 = n_38783 ^ n_37781;
assign n_38794 = n_38783 ^ n_38115;
assign n_38795 = n_38784 ^ x304;
assign n_38796 = n_38785 ^ n_36671;
assign n_38797 = n_38786 ^ n_38784;
assign n_38798 = n_38788 ^ n_38404;
assign n_38799 = n_38789 ^ n_38788;
assign y45 = n_38791;
assign n_38800 = n_38793 ^ n_38115;
assign n_38801 = n_38128 & n_38794;
assign n_38802 = n_38792 ^ n_38796;
assign n_38803 = n_38796 ^ n_36693;
assign n_38804 = n_38782 ^ n_38796;
assign n_38805 = ~n_38797 & n_38795;
assign n_38806 = n_38797 ^ x304;
assign n_38807 = ~n_38799 & ~n_38798;
assign n_38808 = n_38799 ^ n_38404;
assign n_38809 = n_37379 & n_38800;
assign n_38810 = n_38194 ^ n_38800;
assign n_38811 = ~n_38800 & n_38773;
assign n_38812 = n_38773 ^ n_38800;
assign n_38813 = n_38801 ^ n_37781;
assign n_38814 = n_38802 ^ x319;
assign n_38815 = ~n_38803 & n_38804;
assign n_38816 = n_38805 ^ x304;
assign n_38817 = ~n_38787 & ~n_38806;
assign n_38818 = n_38806 ^ n_38787;
assign n_38819 = n_38807 ^ n_38404;
assign n_38820 = ~n_38790 & n_38808;
assign n_38821 = n_38808 ^ n_38790;
assign n_38822 = n_38809 ^ n_38115;
assign y94 = ~n_38812;
assign n_38823 = n_38813 ^ n_37802;
assign n_38824 = n_38813 ^ n_38172;
assign n_38825 = n_38815 ^ n_36693;
assign n_38826 = n_38816 ^ n_38802;
assign n_38827 = n_38818 ^ n_38434;
assign n_38828 = n_38818 ^ n_38819;
assign n_38829 = n_38819 ^ n_38434;
assign y44 = n_38821;
assign n_38830 = n_38822 ^ n_36714;
assign n_38831 = n_38823 ^ n_38172;
assign n_38832 = ~n_38185 & n_38824;
assign n_38833 = n_38825 ^ n_36714;
assign n_38834 = n_38822 ^ n_38825;
assign n_38835 = n_38826 & ~n_38814;
assign n_38836 = n_38826 ^ x319;
assign n_38837 = n_38827 & ~n_38828;
assign n_38838 = n_38818 ^ n_38829;
assign n_38839 = n_37408 & n_38831;
assign n_38840 = n_38246 ^ n_38831;
assign n_38841 = ~n_38831 & n_38811;
assign n_38842 = n_38811 ^ n_38831;
assign n_38843 = n_38832 ^ n_37802;
assign n_38844 = n_38822 ^ n_38833;
assign n_38845 = ~n_38830 & n_38834;
assign n_38846 = n_38835 ^ x319;
assign n_38847 = n_38817 & n_38836;
assign n_38848 = n_38836 ^ n_38817;
assign n_38849 = n_38837 ^ n_38434;
assign n_38850 = ~n_38820 & ~n_38838;
assign n_38851 = n_38838 ^ n_38820;
assign n_38852 = n_38839 ^ n_38172;
assign y93 = ~n_38842;
assign n_38853 = n_38843 ^ n_38216;
assign n_38854 = n_38844 ^ x318;
assign n_38855 = n_38845 ^ n_36714;
assign n_38856 = n_38846 ^ n_38844;
assign n_38857 = n_38848 ^ n_38463;
assign n_38858 = n_38849 ^ n_38848;
assign y43 = n_38851;
assign n_38859 = n_38852 ^ n_36735;
assign n_38860 = n_37823 ^ n_38853;
assign n_38861 = n_38853 & ~n_38230;
assign n_38862 = n_38855 ^ n_36735;
assign n_38863 = n_38855 ^ n_38852;
assign n_38864 = n_38856 ^ x318;
assign n_38865 = n_38856 & ~n_38854;
assign n_38866 = ~n_38858 & ~n_38857;
assign n_38867 = n_38858 ^ n_38463;
assign n_38868 = ~n_37439 & n_38860;
assign n_38869 = n_38291 ^ n_38860;
assign n_38870 = n_38860 & ~n_38841;
assign n_38871 = n_38841 ^ n_38860;
assign n_38872 = n_38861 ^ n_37823;
assign n_38873 = n_38862 ^ n_38852;
assign n_38874 = n_38859 & ~n_38863;
assign n_38875 = n_38864 ^ n_38847;
assign n_38876 = n_38847 & n_38864;
assign n_38877 = n_38865 ^ x318;
assign n_38878 = n_38866 ^ n_38463;
assign n_38879 = ~n_38850 & ~n_38867;
assign n_38880 = n_38867 ^ n_38850;
assign n_38881 = n_38868 ^ n_38216;
assign y92 = n_38871;
assign n_38882 = n_38872 ^ n_38249;
assign n_38883 = n_38873 ^ x317;
assign n_38884 = n_38874 ^ n_36735;
assign n_38885 = n_38875 ^ n_38488;
assign n_38886 = n_38877 ^ x317;
assign n_38887 = n_38877 ^ n_38873;
assign n_38888 = n_38875 ^ n_38878;
assign n_38889 = n_38878 ^ n_38488;
assign y42 = ~n_38880;
assign n_38890 = n_38881 ^ n_36754;
assign n_38891 = n_37845 ^ n_38882;
assign n_38892 = n_38882 & n_38263;
assign n_38893 = n_38884 ^ n_36754;
assign n_38894 = n_38884 ^ n_38881;
assign n_38895 = n_38886 ^ n_38873;
assign n_38896 = n_38883 & ~n_38887;
assign n_38897 = n_38885 & n_38888;
assign n_38898 = n_38875 ^ n_38889;
assign n_38899 = ~n_37478 & ~n_38891;
assign n_38900 = n_38331 ^ n_38891;
assign n_38901 = ~n_38891 & n_38870;
assign n_38902 = n_38870 ^ n_38891;
assign n_38903 = n_38892 ^ n_37845;
assign n_38904 = n_38893 ^ n_38881;
assign n_38905 = n_38890 & ~n_38894;
assign n_38906 = n_38895 ^ n_38876;
assign n_38907 = ~n_38876 & n_38895;
assign n_38908 = n_38896 ^ x317;
assign n_38909 = n_38897 ^ n_38488;
assign n_38910 = ~n_38879 & n_38898;
assign n_38911 = n_38898 ^ n_38879;
assign n_38912 = n_38899 ^ n_38249;
assign y91 = n_38902;
assign n_38913 = n_38903 ^ n_38319;
assign n_38914 = n_38903 ^ n_38306;
assign n_38915 = n_38904 ^ x316;
assign n_38916 = n_38905 ^ n_36754;
assign n_38917 = n_38906 ^ n_38504;
assign n_38918 = n_38908 ^ n_38904;
assign n_38919 = n_38908 ^ x316;
assign n_38920 = n_38909 ^ n_38504;
assign n_38921 = n_38909 ^ n_38906;
assign y41 = ~n_38911;
assign n_38922 = n_38912 ^ n_36774;
assign n_38923 = n_37509 & n_38913;
assign n_38924 = n_38379 ^ n_38913;
assign n_38925 = ~n_38913 & ~n_38901;
assign n_38926 = n_38901 ^ n_38913;
assign n_38927 = n_38319 & n_38914;
assign n_38928 = n_38916 ^ n_36774;
assign n_38929 = n_38916 ^ n_38912;
assign n_38930 = n_38915 & ~n_38918;
assign n_38931 = n_38919 ^ n_38904;
assign n_38932 = n_38920 ^ n_38906;
assign n_38933 = n_38917 & ~n_38921;
assign n_38934 = n_38923 ^ n_38306;
assign y90 = n_38926;
assign n_38935 = n_38927 ^ n_37867;
assign n_38936 = n_38928 ^ n_38912;
assign n_38937 = ~n_38922 & ~n_38929;
assign n_38938 = n_38930 ^ x316;
assign n_38939 = ~n_38907 & ~n_38931;
assign n_38940 = n_38931 ^ n_38907;
assign n_38941 = n_38932 ^ n_38910;
assign n_38942 = ~n_38910 & n_38932;
assign n_38943 = n_38933 ^ n_38504;
assign n_38944 = n_38934 ^ n_36797;
assign n_38945 = n_38935 ^ n_38349;
assign n_38946 = n_38935 ^ n_37889;
assign n_38947 = n_38936 ^ x315;
assign n_38948 = n_38937 ^ n_36774;
assign n_38949 = n_38938 ^ n_38936;
assign n_38950 = n_38940 ^ n_38533;
assign y40 = n_38941;
assign n_38951 = n_38943 ^ n_38940;
assign n_38952 = n_38945 ^ n_37889;
assign n_38953 = ~n_38945 & n_38946;
assign n_38954 = n_38948 ^ n_36797;
assign n_38955 = n_38948 ^ n_38934;
assign n_38956 = n_38949 & ~n_38947;
assign n_38957 = n_38949 ^ x315;
assign n_38958 = n_38943 ^ n_38950;
assign n_38959 = ~n_38950 & ~n_38951;
assign n_38960 = ~n_37551 & ~n_38952;
assign n_38961 = n_38410 ^ n_38952;
assign n_38962 = n_38952 & n_38925;
assign n_38963 = n_38925 ^ n_38952;
assign n_38964 = n_38397 ^ n_38953;
assign n_38965 = n_38954 ^ n_38934;
assign n_38966 = n_38944 & ~n_38955;
assign n_38967 = n_38956 ^ x315;
assign n_38968 = ~n_38939 & ~n_38957;
assign n_38969 = n_38957 ^ n_38939;
assign n_38970 = n_38942 & ~n_38958;
assign n_38971 = n_38958 ^ n_38942;
assign n_38972 = n_38959 ^ n_38533;
assign n_38973 = n_38960 ^ n_38349;
assign y89 = n_38963;
assign n_38974 = n_37605 & ~n_38964;
assign n_38975 = n_38452 ^ n_38964;
assign n_38976 = n_38962 ^ n_38964;
assign n_38977 = n_38965 ^ x314;
assign n_38978 = n_38966 ^ n_36797;
assign n_38979 = n_38967 ^ n_38965;
assign n_38980 = n_38969 ^ n_38570;
assign y55 = n_38971;
assign n_38981 = n_38972 ^ n_38969;
assign n_38982 = n_38973 ^ n_36826;
assign n_38983 = n_38974 ^ n_38365;
assign y88 = ~n_38976;
assign n_38984 = n_38978 ^ n_36826;
assign n_38985 = n_38978 ^ n_38973;
assign n_38986 = n_38979 & ~n_38977;
assign n_38987 = n_38979 ^ x314;
assign n_38988 = n_38972 ^ n_38980;
assign n_38989 = ~n_38980 & ~n_38981;
assign n_38990 = n_38984 ^ n_38973;
assign n_38991 = ~n_38982 & ~n_38985;
assign n_38992 = n_38986 ^ x314;
assign n_38993 = ~n_38968 & n_38987;
assign n_38994 = n_38987 ^ n_38968;
assign n_38995 = ~n_38970 & ~n_38988;
assign n_38996 = n_38988 ^ n_38970;
assign n_38997 = n_38989 ^ n_38570;
assign n_38998 = n_38990 ^ x313;
assign n_38999 = n_38991 ^ n_36826;
assign n_39000 = n_38992 ^ n_38990;
assign n_39001 = n_38994 ^ n_38597;
assign y54 = n_38996;
assign n_39002 = n_38997 ^ n_38994;
assign n_39003 = n_38999 ^ n_38983;
assign n_39004 = n_39000 ^ x313;
assign n_39005 = ~n_39000 & n_38998;
assign n_39006 = n_39002 & n_39001;
assign n_39007 = n_39002 ^ n_38597;
assign n_39008 = n_39003 ^ n_36838;
assign n_39009 = n_39004 ^ n_38993;
assign n_39010 = n_38993 & ~n_39004;
assign n_39011 = n_39005 ^ x313;
assign n_39012 = n_39006 ^ n_38597;
assign n_39013 = ~n_38995 & n_39007;
assign n_39014 = n_39007 ^ n_38995;
assign n_39015 = n_39008 ^ x312;
assign n_39016 = n_39009 ^ n_38618;
assign n_39017 = n_39012 ^ n_39009;
assign y53 = n_39014;
assign n_39018 = n_39011 ^ n_39015;
assign n_39019 = n_39012 ^ n_39016;
assign n_39020 = n_39016 & ~n_39017;
assign n_39021 = n_39018 ^ n_39010;
assign n_39022 = n_39013 & ~n_39019;
assign n_39023 = n_39019 ^ n_39013;
assign n_39024 = n_39020 ^ n_38618;
assign n_39025 = n_39021 ^ n_38647;
assign y52 = n_39023;
assign n_39026 = n_39024 ^ n_39021;
assign n_39027 = ~n_39026 & n_39025;
assign n_39028 = n_39026 ^ n_38647;
assign n_39029 = n_39027 ^ n_38647;
assign n_39030 = n_39028 & ~n_39022;
assign n_39031 = n_39022 ^ n_39028;
assign n_39032 = n_39029 ^ n_38681;
assign n_39033 = n_39029 ^ n_38690;
assign y51 = ~n_39031;
assign n_39034 = ~n_38690 & ~n_39032;
assign n_39035 = n_39030 & ~n_39033;
assign n_39036 = n_39033 ^ n_39030;
assign n_39037 = n_39034 ^ n_37963;
assign y50 = ~n_39036;
assign n_39038 = n_39037 ^ n_38701;
assign n_39039 = ~n_39038 & n_38711;
assign n_39040 = n_39038 ^ n_38025;
assign n_39041 = n_39039 ^ n_38025;
assign n_39042 = n_39040 & ~n_39035;
assign n_39043 = n_39035 ^ n_39040;
assign n_39044 = n_39041 ^ n_38738;
assign y49 = n_39043;
assign n_39045 = n_39044 ^ n_38109;
assign n_39046 = n_39044 & ~n_38747;
assign n_39047 = n_39045 ^ n_39042;
assign n_39048 = n_39042 & ~n_39045;
assign n_39049 = n_39046 ^ n_38109;
assign y48 = n_39047;
assign n_39050 = n_39049 ^ n_38760;
assign n_39051 = ~n_39050 & n_38772;
assign n_39052 = n_39050 ^ n_38150;
assign n_39053 = n_39051 ^ n_38150;
assign n_39054 = n_39048 & n_39052;
assign n_39055 = n_39052 ^ n_39048;
assign n_39056 = n_39053 ^ n_38800;
assign n_39057 = n_38194 ^ n_39053;
assign y63 = ~n_39055;
assign n_39058 = ~n_38810 & ~n_39056;
assign n_39059 = n_39057 ^ n_38800;
assign n_39060 = n_39058 ^ n_38194;
assign n_39061 = n_39054 & ~n_39059;
assign n_39062 = n_39059 ^ n_39054;
assign n_39063 = n_39060 ^ n_38831;
assign n_39064 = n_38246 ^ n_39060;
assign y62 = n_39062;
assign n_39065 = n_38840 & n_39063;
assign n_39066 = n_39064 ^ n_38831;
assign n_39067 = n_39065 ^ n_38246;
assign n_39068 = n_39061 & ~n_39066;
assign n_39069 = n_39066 ^ n_39061;
assign n_39070 = n_39067 ^ n_38860;
assign y61 = n_39069;
assign n_39071 = ~n_39070 & n_38869;
assign n_39072 = n_39070 ^ n_38291;
assign n_39073 = n_39071 ^ n_38291;
assign n_39074 = n_39068 & n_39072;
assign n_39075 = n_39072 ^ n_39068;
assign n_39076 = n_39073 ^ n_38891;
assign y60 = ~n_39075;
assign n_39077 = n_39076 & ~n_38900;
assign n_39078 = n_39076 ^ n_38331;
assign n_39079 = n_39077 ^ n_38331;
assign n_39080 = ~n_39074 & n_39078;
assign n_39081 = n_39078 ^ n_39074;
assign n_39082 = n_38379 ^ n_39079;
assign n_39083 = n_38924 ^ n_39079;
assign y59 = ~n_39081;
assign n_39084 = ~n_38924 & n_39082;
assign n_39085 = ~n_39080 & ~n_39083;
assign n_39086 = n_39083 ^ n_39080;
assign n_39087 = n_39084 ^ n_38913;
assign y58 = ~n_39086;
assign n_39088 = n_39087 ^ n_38952;
assign n_39089 = n_39088 & ~n_38961;
assign n_39090 = n_39088 ^ n_38410;
assign n_39091 = n_39089 ^ n_38410;
assign n_39092 = n_39085 & ~n_39090;
assign n_39093 = n_39090 ^ n_39085;
assign n_39094 = n_39091 ^ n_38975;
assign y57 = n_39093;
assign n_39095 = n_39094 ^ n_39092;
assign y56 = ~n_39095;
endmodule